LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L8_1_WROM IS
  PORT (
    weight : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
    address : IN unsigned(weightsbitsAddress(8)-1 DOWNTO 0));
END L8_1_WROM;

ARCHITECTURE RTL OF L8_1_WROM IS

  TYPE ROM_mem IS ARRAY (0 TO 65535) OF STD_LOGIC_VECTOR(8 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem := (0=>"101001000",
  1=>"010010101",
  2=>"011001000",
  3=>"100010111",
  4=>"110101001",
  5=>"011011101",
  6=>"111001011",
  7=>"110100100",
  8=>"010000000",
  9=>"101110000",
  10=>"011100000",
  11=>"001010110",
  12=>"101001111",
  13=>"001000011",
  14=>"111101000",
  15=>"000101001",
  16=>"000100110",
  17=>"100010010",
  18=>"011101111",
  19=>"000000111",
  20=>"011110001",
  21=>"000110100",
  22=>"100100010",
  23=>"000011001",
  24=>"001000101",
  25=>"011111001",
  26=>"000111000",
  27=>"011110100",
  28=>"110110111",
  29=>"110001001",
  30=>"011000010",
  31=>"000101011",
  32=>"001000101",
  33=>"000011000",
  34=>"100111111",
  35=>"111110000",
  36=>"110100001",
  37=>"011001001",
  38=>"110111001",
  39=>"111011010",
  40=>"011010011",
  41=>"001111100",
  42=>"111011101",
  43=>"000100011",
  44=>"001101001",
  45=>"101011110",
  46=>"111001110",
  47=>"110100111",
  48=>"101000000",
  49=>"001100001",
  50=>"000000000",
  51=>"110000011",
  52=>"001000110",
  53=>"111010100",
  54=>"101010010",
  55=>"101010000",
  56=>"110111111",
  57=>"001000001",
  58=>"101100001",
  59=>"101111110",
  60=>"101111101",
  61=>"100100100",
  62=>"001000001",
  63=>"001000111",
  64=>"111111101",
  65=>"011110101",
  66=>"111110010",
  67=>"100101010",
  68=>"000110010",
  69=>"100101110",
  70=>"101010000",
  71=>"110011100",
  72=>"000110010",
  73=>"000011010",
  74=>"100111101",
  75=>"110101000",
  76=>"001101011",
  77=>"101011001",
  78=>"001111010",
  79=>"000111010",
  80=>"011101111",
  81=>"100000001",
  82=>"000111100",
  83=>"001010011",
  84=>"000111110",
  85=>"100101010",
  86=>"101111000",
  87=>"111010001",
  88=>"001011100",
  89=>"001011101",
  90=>"101011011",
  91=>"001010101",
  92=>"010101010",
  93=>"001101001",
  94=>"001010011",
  95=>"001001010",
  96=>"010000110",
  97=>"101111111",
  98=>"110101001",
  99=>"010000000",
  100=>"110001100",
  101=>"100100101",
  102=>"101111001",
  103=>"110011100",
  104=>"000101010",
  105=>"010111101",
  106=>"001000000",
  107=>"010011001",
  108=>"001010111",
  109=>"001110010",
  110=>"100110001",
  111=>"000111001",
  112=>"010100010",
  113=>"100011111",
  114=>"001000100",
  115=>"000011011",
  116=>"100001100",
  117=>"010100010",
  118=>"101110011",
  119=>"101101000",
  120=>"110000010",
  121=>"101010011",
  122=>"011010100",
  123=>"000100010",
  124=>"011010001",
  125=>"000000001",
  126=>"000011100",
  127=>"101101111",
  128=>"101101110",
  129=>"011001010",
  130=>"001101111",
  131=>"011101001",
  132=>"011000101",
  133=>"010011011",
  134=>"011110011",
  135=>"011101001",
  136=>"110101011",
  137=>"010110100",
  138=>"101111001",
  139=>"010010000",
  140=>"011011000",
  141=>"101000010",
  142=>"101100000",
  143=>"011010000",
  144=>"111001000",
  145=>"111110110",
  146=>"011010110",
  147=>"010010111",
  148=>"100111100",
  149=>"100001100",
  150=>"110101101",
  151=>"101101110",
  152=>"111011011",
  153=>"010110110",
  154=>"111011111",
  155=>"111100111",
  156=>"101110110",
  157=>"111011010",
  158=>"110001000",
  159=>"110010001",
  160=>"001000101",
  161=>"101001001",
  162=>"001111101",
  163=>"001101111",
  164=>"110111010",
  165=>"100011000",
  166=>"000100001",
  167=>"011000010",
  168=>"100011000",
  169=>"111010101",
  170=>"011011110",
  171=>"000110100",
  172=>"101000010",
  173=>"000101100",
  174=>"001111101",
  175=>"110111110",
  176=>"111100010",
  177=>"111011100",
  178=>"010110000",
  179=>"011000000",
  180=>"000000011",
  181=>"000010101",
  182=>"001000111",
  183=>"010100111",
  184=>"000001100",
  185=>"101001100",
  186=>"001011000",
  187=>"111011101",
  188=>"110000101",
  189=>"100110101",
  190=>"110101101",
  191=>"110111010",
  192=>"110011011",
  193=>"001000101",
  194=>"000011000",
  195=>"010000101",
  196=>"100011000",
  197=>"110100110",
  198=>"110000101",
  199=>"101110100",
  200=>"110111101",
  201=>"000001100",
  202=>"001010000",
  203=>"101110001",
  204=>"100101101",
  205=>"110101010",
  206=>"101111010",
  207=>"011010110",
  208=>"100001001",
  209=>"000110010",
  210=>"010110011",
  211=>"010101010",
  212=>"100000010",
  213=>"101001000",
  214=>"110010100",
  215=>"111100011",
  216=>"100101100",
  217=>"110001011",
  218=>"011101101",
  219=>"101110110",
  220=>"101001000",
  221=>"011100101",
  222=>"011010001",
  223=>"000111000",
  224=>"101010101",
  225=>"001111101",
  226=>"101100010",
  227=>"110011010",
  228=>"101010101",
  229=>"011111101",
  230=>"000000001",
  231=>"010001010",
  232=>"010010110",
  233=>"110111111",
  234=>"101101110",
  235=>"111110010",
  236=>"011001110",
  237=>"010000010",
  238=>"100111001",
  239=>"101110101",
  240=>"000101110",
  241=>"010111000",
  242=>"110110000",
  243=>"001111000",
  244=>"111011010",
  245=>"110010101",
  246=>"110010010",
  247=>"011110110",
  248=>"000001111",
  249=>"100001000",
  250=>"110011101",
  251=>"010011010",
  252=>"001011001",
  253=>"010011010",
  254=>"001011100",
  255=>"110101011",
  256=>"110111111",
  257=>"100011011",
  258=>"100001111",
  259=>"000000010",
  260=>"011101000",
  261=>"000101101",
  262=>"111101010",
  263=>"101101101",
  264=>"100000001",
  265=>"000011111",
  266=>"100100110",
  267=>"011101110",
  268=>"100000000",
  269=>"000000010",
  270=>"110011110",
  271=>"011001100",
  272=>"001011101",
  273=>"111101100",
  274=>"111101111",
  275=>"010010000",
  276=>"110111111",
  277=>"101001001",
  278=>"111100110",
  279=>"110110011",
  280=>"100001000",
  281=>"000000110",
  282=>"000101101",
  283=>"000111001",
  284=>"010011111",
  285=>"000110100",
  286=>"110111010",
  287=>"100001001",
  288=>"100001100",
  289=>"101001111",
  290=>"010010101",
  291=>"101101110",
  292=>"000100001",
  293=>"110110101",
  294=>"000100110",
  295=>"000110011",
  296=>"001100010",
  297=>"011100000",
  298=>"110001101",
  299=>"100011001",
  300=>"000110010",
  301=>"100011000",
  302=>"101101010",
  303=>"111000101",
  304=>"111011011",
  305=>"011110010",
  306=>"111100111",
  307=>"101100000",
  308=>"001111001",
  309=>"110100000",
  310=>"110111001",
  311=>"100101011",
  312=>"000111001",
  313=>"000101111",
  314=>"010010000",
  315=>"010001001",
  316=>"000010000",
  317=>"001101100",
  318=>"010110110",
  319=>"100001100",
  320=>"101001001",
  321=>"001101111",
  322=>"111000010",
  323=>"001000001",
  324=>"111110001",
  325=>"100100001",
  326=>"001100010",
  327=>"101010011",
  328=>"010111001",
  329=>"111000000",
  330=>"000000000",
  331=>"000011111",
  332=>"001111001",
  333=>"111110111",
  334=>"111000000",
  335=>"010101110",
  336=>"001000001",
  337=>"111011101",
  338=>"001111100",
  339=>"001110101",
  340=>"010001111",
  341=>"001110101",
  342=>"110101100",
  343=>"101000110",
  344=>"101010101",
  345=>"101101100",
  346=>"010110001",
  347=>"001001010",
  348=>"110010001",
  349=>"001011000",
  350=>"101101001",
  351=>"111110010",
  352=>"101101111",
  353=>"111010100",
  354=>"111001100",
  355=>"100111111",
  356=>"101100101",
  357=>"100110101",
  358=>"011011111",
  359=>"000001001",
  360=>"100110000",
  361=>"110010100",
  362=>"111000101",
  363=>"010010011",
  364=>"101110010",
  365=>"000100000",
  366=>"101011101",
  367=>"000000011",
  368=>"101110100",
  369=>"111001111",
  370=>"011100110",
  371=>"010000110",
  372=>"110010101",
  373=>"100000011",
  374=>"110111010",
  375=>"101100011",
  376=>"101001111",
  377=>"111010101",
  378=>"110100100",
  379=>"100111111",
  380=>"111001110",
  381=>"111100001",
  382=>"001111001",
  383=>"101111000",
  384=>"111110011",
  385=>"110000000",
  386=>"000101011",
  387=>"010010100",
  388=>"000001010",
  389=>"010010101",
  390=>"111110011",
  391=>"110001001",
  392=>"000010011",
  393=>"110001110",
  394=>"101100000",
  395=>"110111011",
  396=>"001010001",
  397=>"110111011",
  398=>"110011111",
  399=>"010001101",
  400=>"001001111",
  401=>"000010000",
  402=>"011111011",
  403=>"011100100",
  404=>"110000100",
  405=>"010001000",
  406=>"010111111",
  407=>"011000011",
  408=>"110100010",
  409=>"101000111",
  410=>"011110101",
  411=>"010101001",
  412=>"001101101",
  413=>"110100101",
  414=>"110001000",
  415=>"001000100",
  416=>"001101001",
  417=>"011011011",
  418=>"001010000",
  419=>"001100001",
  420=>"011101010",
  421=>"000101111",
  422=>"100110101",
  423=>"010110110",
  424=>"100100000",
  425=>"000111110",
  426=>"110010000",
  427=>"001010011",
  428=>"000100011",
  429=>"110111101",
  430=>"110100110",
  431=>"000110101",
  432=>"111100001",
  433=>"010001100",
  434=>"101100000",
  435=>"101110000",
  436=>"100000001",
  437=>"000101000",
  438=>"110100010",
  439=>"001011000",
  440=>"111001110",
  441=>"000000110",
  442=>"000001110",
  443=>"101011101",
  444=>"011000111",
  445=>"100110011",
  446=>"110001110",
  447=>"111110000",
  448=>"100001010",
  449=>"111001110",
  450=>"010101010",
  451=>"001111000",
  452=>"111101100",
  453=>"011100110",
  454=>"011100111",
  455=>"010101111",
  456=>"010010110",
  457=>"101011100",
  458=>"011100010",
  459=>"100101111",
  460=>"100101101",
  461=>"101001000",
  462=>"101010101",
  463=>"100011111",
  464=>"111001010",
  465=>"000010110",
  466=>"001110000",
  467=>"001110101",
  468=>"101101110",
  469=>"010111110",
  470=>"101101111",
  471=>"001100101",
  472=>"010101101",
  473=>"010000101",
  474=>"110010010",
  475=>"100100001",
  476=>"011111011",
  477=>"110001011",
  478=>"001101010",
  479=>"011001000",
  480=>"000000110",
  481=>"000000100",
  482=>"100010110",
  483=>"011001010",
  484=>"000010111",
  485=>"011101100",
  486=>"010000000",
  487=>"010010100",
  488=>"000101110",
  489=>"110010111",
  490=>"110111100",
  491=>"011011010",
  492=>"000001101",
  493=>"110001110",
  494=>"011100010",
  495=>"001110110",
  496=>"000000110",
  497=>"100010100",
  498=>"000001001",
  499=>"001100000",
  500=>"010111110",
  501=>"101001100",
  502=>"010001111",
  503=>"100010111",
  504=>"010111001",
  505=>"011000000",
  506=>"000000111",
  507=>"101000000",
  508=>"010010100",
  509=>"110000111",
  510=>"000110101",
  511=>"010011111",
  512=>"000101110",
  513=>"011111111",
  514=>"011111100",
  515=>"100001000",
  516=>"010000111",
  517=>"111001010",
  518=>"001001110",
  519=>"100010000",
  520=>"000011001",
  521=>"111110100",
  522=>"100111011",
  523=>"001001001",
  524=>"000011111",
  525=>"101000011",
  526=>"000100011",
  527=>"101010011",
  528=>"001100100",
  529=>"111101111",
  530=>"101101100",
  531=>"111100011",
  532=>"001100111",
  533=>"000010100",
  534=>"100110100",
  535=>"011100010",
  536=>"100000011",
  537=>"010000110",
  538=>"111110100",
  539=>"010010101",
  540=>"001110110",
  541=>"000011001",
  542=>"000101111",
  543=>"001010101",
  544=>"000110100",
  545=>"101111101",
  546=>"101001101",
  547=>"000101010",
  548=>"111110011",
  549=>"000000101",
  550=>"101001000",
  551=>"000010010",
  552=>"000001001",
  553=>"000110101",
  554=>"011111101",
  555=>"111101101",
  556=>"010001111",
  557=>"101011001",
  558=>"000101000",
  559=>"011000010",
  560=>"010001010",
  561=>"111010011",
  562=>"001001101",
  563=>"011100100",
  564=>"000100100",
  565=>"011110001",
  566=>"101101011",
  567=>"000111011",
  568=>"011011000",
  569=>"011001001",
  570=>"101111011",
  571=>"100010001",
  572=>"100000001",
  573=>"101101001",
  574=>"101101111",
  575=>"110110000",
  576=>"111001110",
  577=>"110011001",
  578=>"110010111",
  579=>"110101001",
  580=>"010000110",
  581=>"110101011",
  582=>"000010000",
  583=>"111111110",
  584=>"111101011",
  585=>"001100011",
  586=>"000101010",
  587=>"100101100",
  588=>"000000100",
  589=>"111111001",
  590=>"111011011",
  591=>"001000000",
  592=>"011110111",
  593=>"110111010",
  594=>"001000010",
  595=>"010100011",
  596=>"000001010",
  597=>"110000001",
  598=>"000100110",
  599=>"000101001",
  600=>"011100110",
  601=>"011101010",
  602=>"001110110",
  603=>"011010111",
  604=>"000000001",
  605=>"100101101",
  606=>"111001011",
  607=>"100110101",
  608=>"001000000",
  609=>"010110101",
  610=>"000101100",
  611=>"000111101",
  612=>"101011101",
  613=>"001110011",
  614=>"110111011",
  615=>"111100011",
  616=>"010101101",
  617=>"000111011",
  618=>"111010001",
  619=>"001011000",
  620=>"000100000",
  621=>"001101100",
  622=>"001011101",
  623=>"101110000",
  624=>"001100110",
  625=>"000100001",
  626=>"000111111",
  627=>"111000011",
  628=>"000010100",
  629=>"110101101",
  630=>"010111101",
  631=>"101101111",
  632=>"001001101",
  633=>"000111001",
  634=>"001000110",
  635=>"110010101",
  636=>"110000001",
  637=>"100000001",
  638=>"000111111",
  639=>"011001011",
  640=>"010001011",
  641=>"100000000",
  642=>"001100011",
  643=>"111100101",
  644=>"110100101",
  645=>"011001110",
  646=>"000000100",
  647=>"001011011",
  648=>"101001011",
  649=>"000010010",
  650=>"011111100",
  651=>"111110101",
  652=>"101000111",
  653=>"111001000",
  654=>"000010000",
  655=>"110100000",
  656=>"011011010",
  657=>"100101000",
  658=>"111100110",
  659=>"101001110",
  660=>"111101110",
  661=>"101111011",
  662=>"101001000",
  663=>"101100110",
  664=>"000110110",
  665=>"100111101",
  666=>"001010000",
  667=>"001110110",
  668=>"000110101",
  669=>"001101111",
  670=>"010010000",
  671=>"101000000",
  672=>"010000101",
  673=>"110011101",
  674=>"110000101",
  675=>"000011110",
  676=>"100100011",
  677=>"100100001",
  678=>"001001010",
  679=>"000000110",
  680=>"110110101",
  681=>"010110001",
  682=>"110110100",
  683=>"110011001",
  684=>"100101101",
  685=>"011100010",
  686=>"000100101",
  687=>"110010011",
  688=>"101010001",
  689=>"101111110",
  690=>"100100101",
  691=>"100001110",
  692=>"011100011",
  693=>"010011101",
  694=>"110100011",
  695=>"010010011",
  696=>"011000001",
  697=>"011100001",
  698=>"111010100",
  699=>"011101001",
  700=>"111101000",
  701=>"000000100",
  702=>"110111111",
  703=>"000010110",
  704=>"100101110",
  705=>"000000100",
  706=>"001111011",
  707=>"011011100",
  708=>"011100011",
  709=>"000000000",
  710=>"001101010",
  711=>"100010100",
  712=>"000110000",
  713=>"001101100",
  714=>"010111110",
  715=>"101010010",
  716=>"110011111",
  717=>"100001000",
  718=>"111110100",
  719=>"111101001",
  720=>"000011110",
  721=>"001001001",
  722=>"101101011",
  723=>"110110010",
  724=>"000110101",
  725=>"010101111",
  726=>"101111100",
  727=>"001000000",
  728=>"111110011",
  729=>"100001001",
  730=>"100100110",
  731=>"000001011",
  732=>"000010100",
  733=>"011101101",
  734=>"011001110",
  735=>"011001011",
  736=>"000011110",
  737=>"000011000",
  738=>"001011110",
  739=>"111110101",
  740=>"100111100",
  741=>"101101100",
  742=>"001100110",
  743=>"110111100",
  744=>"001100000",
  745=>"101000000",
  746=>"110010101",
  747=>"110011000",
  748=>"000100011",
  749=>"110011110",
  750=>"110000110",
  751=>"011010111",
  752=>"000010000",
  753=>"011001000",
  754=>"101111011",
  755=>"010000110",
  756=>"110101101",
  757=>"000011000",
  758=>"010111111",
  759=>"000000011",
  760=>"001011001",
  761=>"011110110",
  762=>"001000100",
  763=>"101010000",
  764=>"011001111",
  765=>"010000001",
  766=>"000101101",
  767=>"010001001",
  768=>"100110011",
  769=>"100010000",
  770=>"011000001",
  771=>"011111001",
  772=>"010101110",
  773=>"110000111",
  774=>"010110111",
  775=>"011100011",
  776=>"110110011",
  777=>"100000101",
  778=>"111100111",
  779=>"110101000",
  780=>"010110001",
  781=>"010101110",
  782=>"101000111",
  783=>"110001001",
  784=>"100100001",
  785=>"110111100",
  786=>"010100000",
  787=>"110001111",
  788=>"000111111",
  789=>"000000101",
  790=>"001101011",
  791=>"110010011",
  792=>"100010010",
  793=>"101110100",
  794=>"001001010",
  795=>"000011010",
  796=>"100010100",
  797=>"101010010",
  798=>"011101000",
  799=>"100110110",
  800=>"010011110",
  801=>"110000100",
  802=>"111000001",
  803=>"111100010",
  804=>"101001001",
  805=>"100111111",
  806=>"001111111",
  807=>"010111001",
  808=>"010101100",
  809=>"110100100",
  810=>"011111111",
  811=>"011001110",
  812=>"011000000",
  813=>"100011011",
  814=>"100110110",
  815=>"000110010",
  816=>"100101101",
  817=>"111100011",
  818=>"111110101",
  819=>"111001010",
  820=>"010110110",
  821=>"010111100",
  822=>"001100000",
  823=>"110110010",
  824=>"011010110",
  825=>"000111010",
  826=>"101001111",
  827=>"101000110",
  828=>"000001100",
  829=>"101111010",
  830=>"000000100",
  831=>"001101100",
  832=>"000111011",
  833=>"011000100",
  834=>"101000010",
  835=>"001101111",
  836=>"100000111",
  837=>"101001011",
  838=>"011101010",
  839=>"101101011",
  840=>"001100111",
  841=>"011000110",
  842=>"110111001",
  843=>"000001100",
  844=>"000100010",
  845=>"111001000",
  846=>"110111110",
  847=>"111001000",
  848=>"111101111",
  849=>"011000100",
  850=>"000000100",
  851=>"000011011",
  852=>"111110011",
  853=>"111010010",
  854=>"000111111",
  855=>"010101110",
  856=>"001100101",
  857=>"101111000",
  858=>"001111100",
  859=>"000000000",
  860=>"110001100",
  861=>"011111111",
  862=>"001100110",
  863=>"000110101",
  864=>"001111100",
  865=>"110000011",
  866=>"010010000",
  867=>"000101100",
  868=>"010100110",
  869=>"110111001",
  870=>"100010011",
  871=>"101011100",
  872=>"111010000",
  873=>"001100011",
  874=>"110010011",
  875=>"010011011",
  876=>"101000101",
  877=>"110000111",
  878=>"011010001",
  879=>"001101100",
  880=>"111110100",
  881=>"011101100",
  882=>"001010000",
  883=>"010111000",
  884=>"001100000",
  885=>"111110011",
  886=>"010001011",
  887=>"000110100",
  888=>"000100110",
  889=>"010011010",
  890=>"000110111",
  891=>"001000100",
  892=>"001110100",
  893=>"100001001",
  894=>"000100111",
  895=>"001110100",
  896=>"000101000",
  897=>"101011001",
  898=>"100010101",
  899=>"100111001",
  900=>"100101000",
  901=>"111101010",
  902=>"000010011",
  903=>"010010010",
  904=>"000100110",
  905=>"001001001",
  906=>"010010010",
  907=>"000000110",
  908=>"100111111",
  909=>"110001100",
  910=>"010001001",
  911=>"101010010",
  912=>"100000110",
  913=>"001111011",
  914=>"100111100",
  915=>"100001010",
  916=>"001000001",
  917=>"110111011",
  918=>"001100000",
  919=>"110110001",
  920=>"100011011",
  921=>"010001111",
  922=>"000101001",
  923=>"011001011",
  924=>"111010111",
  925=>"001110010",
  926=>"011110001",
  927=>"011011100",
  928=>"111000000",
  929=>"111000110",
  930=>"000111011",
  931=>"101000101",
  932=>"010010110",
  933=>"010010101",
  934=>"110111111",
  935=>"010100000",
  936=>"001111101",
  937=>"110111000",
  938=>"101100000",
  939=>"111100110",
  940=>"000000011",
  941=>"000111111",
  942=>"110001011",
  943=>"000011001",
  944=>"111100000",
  945=>"101100001",
  946=>"101111000",
  947=>"111111111",
  948=>"111110010",
  949=>"111100001",
  950=>"000111111",
  951=>"000011011",
  952=>"100001110",
  953=>"000101000",
  954=>"110100110",
  955=>"010000000",
  956=>"000101000",
  957=>"000100110",
  958=>"010110110",
  959=>"101010101",
  960=>"010010001",
  961=>"101010110",
  962=>"100000111",
  963=>"000101111",
  964=>"000001110",
  965=>"000111110",
  966=>"111011010",
  967=>"101000000",
  968=>"001100101",
  969=>"000000000",
  970=>"011110101",
  971=>"111011111",
  972=>"110101011",
  973=>"010001011",
  974=>"111001101",
  975=>"100001101",
  976=>"000110000",
  977=>"000111100",
  978=>"001110111",
  979=>"000001000",
  980=>"001101101",
  981=>"101111111",
  982=>"100011110",
  983=>"000001101",
  984=>"101110011",
  985=>"010101001",
  986=>"111001100",
  987=>"100000010",
  988=>"000000010",
  989=>"001110001",
  990=>"011001110",
  991=>"010101001",
  992=>"011111000",
  993=>"000100111",
  994=>"010111110",
  995=>"000100101",
  996=>"000110010",
  997=>"111010111",
  998=>"001110011",
  999=>"001101001",
  1000=>"110100100",
  1001=>"010001101",
  1002=>"000100000",
  1003=>"100001110",
  1004=>"010000101",
  1005=>"111011100",
  1006=>"011000110",
  1007=>"001000101",
  1008=>"000111100",
  1009=>"110010111",
  1010=>"111011111",
  1011=>"010010010",
  1012=>"001001101",
  1013=>"111110011",
  1014=>"111000100",
  1015=>"111110010",
  1016=>"100100011",
  1017=>"001010000",
  1018=>"000100001",
  1019=>"101001110",
  1020=>"100110011",
  1021=>"110100101",
  1022=>"111011011",
  1023=>"101001010",
  1024=>"110010000",
  1025=>"101010001",
  1026=>"101100100",
  1027=>"011001110",
  1028=>"001100011",
  1029=>"110011011",
  1030=>"011100111",
  1031=>"001101101",
  1032=>"100101010",
  1033=>"110101011",
  1034=>"100111001",
  1035=>"111010010",
  1036=>"001101110",
  1037=>"011101010",
  1038=>"110010111",
  1039=>"110100110",
  1040=>"101111110",
  1041=>"011001000",
  1042=>"110110010",
  1043=>"000000000",
  1044=>"011001011",
  1045=>"001101110",
  1046=>"010011000",
  1047=>"101100111",
  1048=>"000101100",
  1049=>"111001100",
  1050=>"010111000",
  1051=>"000000001",
  1052=>"011001111",
  1053=>"010100010",
  1054=>"010110000",
  1055=>"111011010",
  1056=>"011001011",
  1057=>"000000001",
  1058=>"100111000",
  1059=>"001001111",
  1060=>"111000100",
  1061=>"011001011",
  1062=>"110111100",
  1063=>"001011110",
  1064=>"010111011",
  1065=>"001111000",
  1066=>"100011001",
  1067=>"100100010",
  1068=>"100100001",
  1069=>"101001100",
  1070=>"000001101",
  1071=>"000000111",
  1072=>"101110110",
  1073=>"000100000",
  1074=>"000001011",
  1075=>"101101110",
  1076=>"000101000",
  1077=>"111111011",
  1078=>"101001110",
  1079=>"001111010",
  1080=>"010001111",
  1081=>"010000011",
  1082=>"000011110",
  1083=>"101001000",
  1084=>"000100001",
  1085=>"101001010",
  1086=>"001010001",
  1087=>"000010111",
  1088=>"110010111",
  1089=>"000000010",
  1090=>"100001011",
  1091=>"100100110",
  1092=>"011100001",
  1093=>"000110001",
  1094=>"111111100",
  1095=>"101101101",
  1096=>"010111010",
  1097=>"111111010",
  1098=>"011001000",
  1099=>"101101001",
  1100=>"000100010",
  1101=>"111100001",
  1102=>"010110000",
  1103=>"010011110",
  1104=>"111111000",
  1105=>"110000111",
  1106=>"110001001",
  1107=>"010010011",
  1108=>"000011100",
  1109=>"111101000",
  1110=>"110110111",
  1111=>"101001000",
  1112=>"001110101",
  1113=>"101101000",
  1114=>"101110000",
  1115=>"101010101",
  1116=>"111101101",
  1117=>"000101000",
  1118=>"011100100",
  1119=>"110001001",
  1120=>"100101011",
  1121=>"101010001",
  1122=>"011011100",
  1123=>"001001000",
  1124=>"100000111",
  1125=>"010100110",
  1126=>"000101000",
  1127=>"110110101",
  1128=>"010011011",
  1129=>"100100001",
  1130=>"010001010",
  1131=>"110010000",
  1132=>"011101000",
  1133=>"111011001",
  1134=>"101010000",
  1135=>"001110000",
  1136=>"101010000",
  1137=>"011111111",
  1138=>"001100011",
  1139=>"101110101",
  1140=>"001011110",
  1141=>"100100101",
  1142=>"101111111",
  1143=>"101100011",
  1144=>"110000001",
  1145=>"010110010",
  1146=>"101001100",
  1147=>"100001100",
  1148=>"000010110",
  1149=>"101101100",
  1150=>"100100000",
  1151=>"100011101",
  1152=>"000000000",
  1153=>"111101000",
  1154=>"101001001",
  1155=>"001111101",
  1156=>"000001000",
  1157=>"001011101",
  1158=>"111011101",
  1159=>"001100010",
  1160=>"111001110",
  1161=>"101000111",
  1162=>"100000000",
  1163=>"100111000",
  1164=>"011101001",
  1165=>"000101111",
  1166=>"101011011",
  1167=>"001001011",
  1168=>"110111000",
  1169=>"111000011",
  1170=>"101101111",
  1171=>"010011111",
  1172=>"010101110",
  1173=>"101101010",
  1174=>"000011011",
  1175=>"110001100",
  1176=>"010010000",
  1177=>"100011010",
  1178=>"000101000",
  1179=>"010100111",
  1180=>"011111111",
  1181=>"111100110",
  1182=>"011010101",
  1183=>"100001111",
  1184=>"110000110",
  1185=>"100000110",
  1186=>"110000101",
  1187=>"111000010",
  1188=>"100000001",
  1189=>"001000110",
  1190=>"001101101",
  1191=>"011110011",
  1192=>"000010110",
  1193=>"111010011",
  1194=>"101111011",
  1195=>"010101100",
  1196=>"000001011",
  1197=>"000111101",
  1198=>"000011110",
  1199=>"011011011",
  1200=>"111000001",
  1201=>"011100001",
  1202=>"010011100",
  1203=>"001101110",
  1204=>"000010011",
  1205=>"010101001",
  1206=>"100111100",
  1207=>"101000001",
  1208=>"111011111",
  1209=>"011010000",
  1210=>"011001100",
  1211=>"111110011",
  1212=>"101011000",
  1213=>"000101010",
  1214=>"011010100",
  1215=>"111101010",
  1216=>"110001010",
  1217=>"001001101",
  1218=>"000001010",
  1219=>"000101110",
  1220=>"111111100",
  1221=>"010111111",
  1222=>"011101101",
  1223=>"110101101",
  1224=>"001011100",
  1225=>"110000101",
  1226=>"110010011",
  1227=>"000111110",
  1228=>"010101110",
  1229=>"100010111",
  1230=>"101101100",
  1231=>"000101100",
  1232=>"111111101",
  1233=>"101101010",
  1234=>"111001010",
  1235=>"110100001",
  1236=>"000101111",
  1237=>"000000100",
  1238=>"100101010",
  1239=>"000110010",
  1240=>"100100100",
  1241=>"010001000",
  1242=>"000001010",
  1243=>"110110000",
  1244=>"001111011",
  1245=>"101001100",
  1246=>"001100000",
  1247=>"001011100",
  1248=>"101000000",
  1249=>"111000011",
  1250=>"101010101",
  1251=>"100100101",
  1252=>"000100111",
  1253=>"010110100",
  1254=>"000001000",
  1255=>"011001010",
  1256=>"000101111",
  1257=>"000000110",
  1258=>"010100000",
  1259=>"001010000",
  1260=>"111001110",
  1261=>"101011111",
  1262=>"110000000",
  1263=>"011100010",
  1264=>"000100100",
  1265=>"101101100",
  1266=>"110001100",
  1267=>"111000111",
  1268=>"011000010",
  1269=>"001000001",
  1270=>"001011001",
  1271=>"111000011",
  1272=>"001101000",
  1273=>"111110101",
  1274=>"011100101",
  1275=>"001101001",
  1276=>"101101011",
  1277=>"001010000",
  1278=>"011000010",
  1279=>"101111101",
  1280=>"011101000",
  1281=>"001001111",
  1282=>"111010001",
  1283=>"110110110",
  1284=>"011100000",
  1285=>"000101010",
  1286=>"011011110",
  1287=>"111111101",
  1288=>"010011101",
  1289=>"110001100",
  1290=>"111000100",
  1291=>"000000110",
  1292=>"011101100",
  1293=>"110110011",
  1294=>"110010000",
  1295=>"110011011",
  1296=>"110000001",
  1297=>"111000110",
  1298=>"110011011",
  1299=>"100100000",
  1300=>"000001010",
  1301=>"001100100",
  1302=>"000000101",
  1303=>"001100010",
  1304=>"011100010",
  1305=>"110001010",
  1306=>"101010111",
  1307=>"101001001",
  1308=>"001011111",
  1309=>"100110100",
  1310=>"111011010",
  1311=>"000101111",
  1312=>"001001101",
  1313=>"011111000",
  1314=>"100000101",
  1315=>"000111010",
  1316=>"100010001",
  1317=>"111000010",
  1318=>"101001110",
  1319=>"110010001",
  1320=>"000001100",
  1321=>"111010000",
  1322=>"000100100",
  1323=>"010011101",
  1324=>"010011011",
  1325=>"011101001",
  1326=>"000111011",
  1327=>"001001110",
  1328=>"100000100",
  1329=>"111000101",
  1330=>"000111001",
  1331=>"111101100",
  1332=>"101110101",
  1333=>"111011100",
  1334=>"011011100",
  1335=>"101101000",
  1336=>"111101111",
  1337=>"001011010",
  1338=>"000011011",
  1339=>"001110111",
  1340=>"111001011",
  1341=>"110011111",
  1342=>"000110100",
  1343=>"111011111",
  1344=>"100010001",
  1345=>"001110010",
  1346=>"100110100",
  1347=>"011101001",
  1348=>"001011010",
  1349=>"111010111",
  1350=>"000001001",
  1351=>"100111100",
  1352=>"011111110",
  1353=>"001010110",
  1354=>"111010110",
  1355=>"000100111",
  1356=>"101010101",
  1357=>"001011111",
  1358=>"100110001",
  1359=>"101110010",
  1360=>"111111101",
  1361=>"000000101",
  1362=>"000100110",
  1363=>"100110000",
  1364=>"010111101",
  1365=>"011010110",
  1366=>"000100101",
  1367=>"100101000",
  1368=>"100111011",
  1369=>"100011000",
  1370=>"000001001",
  1371=>"110100001",
  1372=>"101101001",
  1373=>"010111001",
  1374=>"100100101",
  1375=>"001000110",
  1376=>"101001011",
  1377=>"111110010",
  1378=>"000100011",
  1379=>"000001101",
  1380=>"000001011",
  1381=>"010011100",
  1382=>"001111101",
  1383=>"010010011",
  1384=>"010110101",
  1385=>"110101110",
  1386=>"010010101",
  1387=>"101100100",
  1388=>"101111101",
  1389=>"010001001",
  1390=>"011010101",
  1391=>"101001010",
  1392=>"000111011",
  1393=>"000010011",
  1394=>"000100110",
  1395=>"000101100",
  1396=>"000000110",
  1397=>"011000001",
  1398=>"110000001",
  1399=>"111010001",
  1400=>"111110101",
  1401=>"000100000",
  1402=>"110011101",
  1403=>"000000110",
  1404=>"000100000",
  1405=>"111111001",
  1406=>"000011001",
  1407=>"101000111",
  1408=>"111101101",
  1409=>"000101101",
  1410=>"001000101",
  1411=>"011001100",
  1412=>"100100000",
  1413=>"111000010",
  1414=>"010110110",
  1415=>"111001100",
  1416=>"111001001",
  1417=>"000010111",
  1418=>"011101010",
  1419=>"011010101",
  1420=>"001000101",
  1421=>"100101110",
  1422=>"100101000",
  1423=>"100100111",
  1424=>"111111000",
  1425=>"001011100",
  1426=>"010000101",
  1427=>"011010011",
  1428=>"010000011",
  1429=>"000010111",
  1430=>"111101000",
  1431=>"111011000",
  1432=>"111010100",
  1433=>"111010000",
  1434=>"111000101",
  1435=>"100111100",
  1436=>"110010101",
  1437=>"100100000",
  1438=>"010011010",
  1439=>"110010001",
  1440=>"110100101",
  1441=>"100011110",
  1442=>"011000111",
  1443=>"100101110",
  1444=>"000101001",
  1445=>"110111100",
  1446=>"110110101",
  1447=>"100100011",
  1448=>"110111011",
  1449=>"101001000",
  1450=>"001011000",
  1451=>"000010011",
  1452=>"011101000",
  1453=>"010000001",
  1454=>"000010111",
  1455=>"100001011",
  1456=>"000001000",
  1457=>"111111011",
  1458=>"000110100",
  1459=>"010001100",
  1460=>"101111010",
  1461=>"110001010",
  1462=>"110000110",
  1463=>"001111111",
  1464=>"111111111",
  1465=>"111001110",
  1466=>"001010010",
  1467=>"001010101",
  1468=>"010010001",
  1469=>"100101110",
  1470=>"111101101",
  1471=>"100111011",
  1472=>"100010011",
  1473=>"100101111",
  1474=>"100100001",
  1475=>"111101111",
  1476=>"010000001",
  1477=>"000001010",
  1478=>"010000001",
  1479=>"101100011",
  1480=>"100110111",
  1481=>"100111101",
  1482=>"101000000",
  1483=>"100010101",
  1484=>"101010111",
  1485=>"110001010",
  1486=>"000111110",
  1487=>"101110001",
  1488=>"001011110",
  1489=>"001100001",
  1490=>"010111000",
  1491=>"001001011",
  1492=>"101111110",
  1493=>"110011100",
  1494=>"000010000",
  1495=>"001110011",
  1496=>"100110100",
  1497=>"111111011",
  1498=>"111111111",
  1499=>"111011101",
  1500=>"000011011",
  1501=>"110111101",
  1502=>"100110001",
  1503=>"011110001",
  1504=>"100110001",
  1505=>"101010100",
  1506=>"110011011",
  1507=>"001001110",
  1508=>"101111011",
  1509=>"101100101",
  1510=>"111010110",
  1511=>"100001110",
  1512=>"100000001",
  1513=>"011110110",
  1514=>"010101100",
  1515=>"000000011",
  1516=>"011100101",
  1517=>"000100011",
  1518=>"110101011",
  1519=>"001101111",
  1520=>"101110000",
  1521=>"000001001",
  1522=>"100101011",
  1523=>"101010001",
  1524=>"010100100",
  1525=>"110111011",
  1526=>"011111011",
  1527=>"100110100",
  1528=>"101011111",
  1529=>"000000111",
  1530=>"011000011",
  1531=>"110101111",
  1532=>"100010110",
  1533=>"100111110",
  1534=>"011110011",
  1535=>"110011001",
  1536=>"110111100",
  1537=>"101100100",
  1538=>"111000101",
  1539=>"111101000",
  1540=>"000110001",
  1541=>"100101111",
  1542=>"000111110",
  1543=>"100000000",
  1544=>"101011000",
  1545=>"110110100",
  1546=>"101110111",
  1547=>"010000001",
  1548=>"010011010",
  1549=>"001111111",
  1550=>"101001101",
  1551=>"100110110",
  1552=>"011100110",
  1553=>"100001010",
  1554=>"011101110",
  1555=>"110001100",
  1556=>"010011101",
  1557=>"010111010",
  1558=>"100111101",
  1559=>"101101111",
  1560=>"000010111",
  1561=>"101000000",
  1562=>"010010101",
  1563=>"100110100",
  1564=>"110110111",
  1565=>"101100101",
  1566=>"000111110",
  1567=>"010111111",
  1568=>"101011011",
  1569=>"011010000",
  1570=>"101100110",
  1571=>"111000111",
  1572=>"011100101",
  1573=>"010000000",
  1574=>"100011000",
  1575=>"011001100",
  1576=>"010110010",
  1577=>"111001011",
  1578=>"001001011",
  1579=>"100001001",
  1580=>"111101000",
  1581=>"011111101",
  1582=>"101101100",
  1583=>"111100011",
  1584=>"100001101",
  1585=>"111100000",
  1586=>"110101110",
  1587=>"101111101",
  1588=>"000011010",
  1589=>"001011011",
  1590=>"001000011",
  1591=>"000010010",
  1592=>"011010011",
  1593=>"101011001",
  1594=>"100001010",
  1595=>"111111100",
  1596=>"011011100",
  1597=>"000001111",
  1598=>"000110111",
  1599=>"110111010",
  1600=>"111010001",
  1601=>"110100100",
  1602=>"110101010",
  1603=>"100000100",
  1604=>"111011101",
  1605=>"010111101",
  1606=>"001000100",
  1607=>"001110111",
  1608=>"001011000",
  1609=>"011000110",
  1610=>"101001100",
  1611=>"000101110",
  1612=>"101000101",
  1613=>"001101001",
  1614=>"011101110",
  1615=>"011110011",
  1616=>"101011100",
  1617=>"010110010",
  1618=>"100111100",
  1619=>"101010001",
  1620=>"110101011",
  1621=>"010111111",
  1622=>"101010110",
  1623=>"010011010",
  1624=>"001101000",
  1625=>"010010011",
  1626=>"011011110",
  1627=>"101100001",
  1628=>"001111100",
  1629=>"001011101",
  1630=>"001111110",
  1631=>"000110100",
  1632=>"000000000",
  1633=>"000100100",
  1634=>"001000101",
  1635=>"010000011",
  1636=>"100000101",
  1637=>"000000100",
  1638=>"111100100",
  1639=>"100000100",
  1640=>"001000011",
  1641=>"010111000",
  1642=>"111010000",
  1643=>"001100001",
  1644=>"100010101",
  1645=>"011001100",
  1646=>"101011100",
  1647=>"011001111",
  1648=>"001000110",
  1649=>"010111111",
  1650=>"111101001",
  1651=>"011111111",
  1652=>"000100011",
  1653=>"111100111",
  1654=>"101111011",
  1655=>"000101101",
  1656=>"101100010",
  1657=>"110010010",
  1658=>"101001010",
  1659=>"011001101",
  1660=>"010000000",
  1661=>"001001110",
  1662=>"111011111",
  1663=>"010100001",
  1664=>"010011000",
  1665=>"010110011",
  1666=>"111100101",
  1667=>"001111000",
  1668=>"101111000",
  1669=>"011011000",
  1670=>"001001001",
  1671=>"111000110",
  1672=>"100111001",
  1673=>"001110111",
  1674=>"111110100",
  1675=>"000000010",
  1676=>"000100101",
  1677=>"100010110",
  1678=>"010101100",
  1679=>"010100101",
  1680=>"011010010",
  1681=>"010011101",
  1682=>"000010001",
  1683=>"101011110",
  1684=>"001001000",
  1685=>"101101010",
  1686=>"011011110",
  1687=>"110110111",
  1688=>"000110110",
  1689=>"011101100",
  1690=>"100011000",
  1691=>"000000000",
  1692=>"011100101",
  1693=>"111100101",
  1694=>"010100001",
  1695=>"011111010",
  1696=>"100100110",
  1697=>"110001100",
  1698=>"000100100",
  1699=>"101101110",
  1700=>"101111101",
  1701=>"111001110",
  1702=>"000001110",
  1703=>"111100101",
  1704=>"010100110",
  1705=>"100001111",
  1706=>"101110001",
  1707=>"110011011",
  1708=>"111101100",
  1709=>"010011100",
  1710=>"011001011",
  1711=>"101110000",
  1712=>"000110111",
  1713=>"010111110",
  1714=>"001011110",
  1715=>"101101001",
  1716=>"111100110",
  1717=>"110110110",
  1718=>"001101001",
  1719=>"111100101",
  1720=>"110111010",
  1721=>"010011110",
  1722=>"110001101",
  1723=>"001101001",
  1724=>"100001101",
  1725=>"000011011",
  1726=>"011000011",
  1727=>"101110001",
  1728=>"110111100",
  1729=>"010011011",
  1730=>"101011011",
  1731=>"011111100",
  1732=>"011101111",
  1733=>"111001010",
  1734=>"010111101",
  1735=>"001101010",
  1736=>"000110011",
  1737=>"110011001",
  1738=>"001101100",
  1739=>"000111001",
  1740=>"010101100",
  1741=>"111101110",
  1742=>"110001010",
  1743=>"011011001",
  1744=>"000110000",
  1745=>"000010010",
  1746=>"000010010",
  1747=>"001100011",
  1748=>"000100110",
  1749=>"010110000",
  1750=>"110110111",
  1751=>"100010001",
  1752=>"001101111",
  1753=>"010011001",
  1754=>"011110011",
  1755=>"100010100",
  1756=>"100000001",
  1757=>"011001001",
  1758=>"010111111",
  1759=>"111011100",
  1760=>"100110111",
  1761=>"011110010",
  1762=>"011101111",
  1763=>"001001111",
  1764=>"101010110",
  1765=>"110000011",
  1766=>"100001010",
  1767=>"011110011",
  1768=>"010010010",
  1769=>"110010101",
  1770=>"111110111",
  1771=>"111111011",
  1772=>"101001011",
  1773=>"011111000",
  1774=>"111111111",
  1775=>"010111010",
  1776=>"110001100",
  1777=>"011111010",
  1778=>"000100011",
  1779=>"101100111",
  1780=>"101100111",
  1781=>"000101101",
  1782=>"100101011",
  1783=>"010000100",
  1784=>"110100111",
  1785=>"001000010",
  1786=>"100111110",
  1787=>"101001001",
  1788=>"100011010",
  1789=>"000100100",
  1790=>"101011101",
  1791=>"010101011",
  1792=>"010011111",
  1793=>"000000101",
  1794=>"111100011",
  1795=>"000101010",
  1796=>"110010011",
  1797=>"111001101",
  1798=>"101110111",
  1799=>"001010000",
  1800=>"110101110",
  1801=>"010001001",
  1802=>"010000110",
  1803=>"011010100",
  1804=>"011101000",
  1805=>"011110011",
  1806=>"110110001",
  1807=>"110011010",
  1808=>"111011101",
  1809=>"011101100",
  1810=>"010110010",
  1811=>"011000111",
  1812=>"100001000",
  1813=>"000101010",
  1814=>"000001100",
  1815=>"111100011",
  1816=>"001101001",
  1817=>"011011010",
  1818=>"000010011",
  1819=>"111011000",
  1820=>"111110111",
  1821=>"001010110",
  1822=>"101110000",
  1823=>"101010110",
  1824=>"100111101",
  1825=>"111110000",
  1826=>"010100110",
  1827=>"001001001",
  1828=>"110100000",
  1829=>"011100111",
  1830=>"110011110",
  1831=>"100011100",
  1832=>"010000100",
  1833=>"000101010",
  1834=>"110111110",
  1835=>"111110000",
  1836=>"010011010",
  1837=>"011110001",
  1838=>"101000010",
  1839=>"010100100",
  1840=>"011100110",
  1841=>"001000100",
  1842=>"001011001",
  1843=>"010000000",
  1844=>"011010110",
  1845=>"011001010",
  1846=>"111101111",
  1847=>"101100100",
  1848=>"000001011",
  1849=>"101011011",
  1850=>"110000001",
  1851=>"101000111",
  1852=>"001011011",
  1853=>"110001000",
  1854=>"101000111",
  1855=>"001101011",
  1856=>"011101100",
  1857=>"110001010",
  1858=>"111011111",
  1859=>"100000110",
  1860=>"011011100",
  1861=>"001010001",
  1862=>"000111101",
  1863=>"101011011",
  1864=>"111101001",
  1865=>"010010000",
  1866=>"100101010",
  1867=>"110011011",
  1868=>"000110100",
  1869=>"001000110",
  1870=>"100110101",
  1871=>"011011100",
  1872=>"101110001",
  1873=>"000100000",
  1874=>"010001000",
  1875=>"011001000",
  1876=>"111001010",
  1877=>"100100000",
  1878=>"001110001",
  1879=>"010011101",
  1880=>"011101100",
  1881=>"011001111",
  1882=>"100111110",
  1883=>"101010001",
  1884=>"111111111",
  1885=>"001000001",
  1886=>"111000110",
  1887=>"111111010",
  1888=>"001000101",
  1889=>"011001100",
  1890=>"000001010",
  1891=>"101111110",
  1892=>"010111111",
  1893=>"110101011",
  1894=>"110001000",
  1895=>"001001101",
  1896=>"010110000",
  1897=>"100101111",
  1898=>"010110110",
  1899=>"011111011",
  1900=>"010101100",
  1901=>"100000001",
  1902=>"111010011",
  1903=>"010101111",
  1904=>"100100011",
  1905=>"001011011",
  1906=>"100001001",
  1907=>"001100010",
  1908=>"011000010",
  1909=>"000011011",
  1910=>"010011111",
  1911=>"100001001",
  1912=>"001011101",
  1913=>"000000111",
  1914=>"100001000",
  1915=>"100101001",
  1916=>"010101000",
  1917=>"110000110",
  1918=>"011110100",
  1919=>"111011010",
  1920=>"011000110",
  1921=>"110001010",
  1922=>"010101011",
  1923=>"011010000",
  1924=>"010110101",
  1925=>"101111000",
  1926=>"001111011",
  1927=>"110100011",
  1928=>"110101100",
  1929=>"111110111",
  1930=>"111011001",
  1931=>"001001001",
  1932=>"000111000",
  1933=>"010011110",
  1934=>"010100101",
  1935=>"001001100",
  1936=>"000101101",
  1937=>"100001101",
  1938=>"111000001",
  1939=>"011101100",
  1940=>"111111010",
  1941=>"110100011",
  1942=>"101001010",
  1943=>"010011101",
  1944=>"100111011",
  1945=>"100001000",
  1946=>"011011000",
  1947=>"001111111",
  1948=>"100011101",
  1949=>"000000010",
  1950=>"000001010",
  1951=>"110110110",
  1952=>"011110001",
  1953=>"111111010",
  1954=>"110011100",
  1955=>"111001100",
  1956=>"010000111",
  1957=>"111111110",
  1958=>"101101101",
  1959=>"001000010",
  1960=>"100010011",
  1961=>"111100100",
  1962=>"000101110",
  1963=>"001111101",
  1964=>"111100101",
  1965=>"111110010",
  1966=>"000100010",
  1967=>"011110011",
  1968=>"101000011",
  1969=>"001111000",
  1970=>"000110101",
  1971=>"110001011",
  1972=>"001010110",
  1973=>"110001110",
  1974=>"000000111",
  1975=>"011000001",
  1976=>"100110110",
  1977=>"100111001",
  1978=>"101011101",
  1979=>"111101000",
  1980=>"000111111",
  1981=>"010000010",
  1982=>"000010001",
  1983=>"100000111",
  1984=>"100110101",
  1985=>"001010010",
  1986=>"111010100",
  1987=>"101100010",
  1988=>"000110001",
  1989=>"111111010",
  1990=>"101000110",
  1991=>"011000000",
  1992=>"000001011",
  1993=>"100010010",
  1994=>"010000001",
  1995=>"111100011",
  1996=>"110101111",
  1997=>"000010101",
  1998=>"101100101",
  1999=>"001101111",
  2000=>"111000111",
  2001=>"110011001",
  2002=>"101000011",
  2003=>"110000110",
  2004=>"011000000",
  2005=>"101101100",
  2006=>"000101110",
  2007=>"000100100",
  2008=>"010011010",
  2009=>"000001001",
  2010=>"000101100",
  2011=>"110011101",
  2012=>"100101010",
  2013=>"111101010",
  2014=>"011110010",
  2015=>"110011101",
  2016=>"010101010",
  2017=>"011111000",
  2018=>"010000111",
  2019=>"001100111",
  2020=>"100110110",
  2021=>"000110001",
  2022=>"000101110",
  2023=>"011100000",
  2024=>"101100001",
  2025=>"101011011",
  2026=>"101110100",
  2027=>"011000000",
  2028=>"101110101",
  2029=>"000001111",
  2030=>"010110100",
  2031=>"000011111",
  2032=>"101110000",
  2033=>"100100110",
  2034=>"000001111",
  2035=>"011100101",
  2036=>"100100100",
  2037=>"101111010",
  2038=>"000111010",
  2039=>"000000110",
  2040=>"001101000",
  2041=>"110011000",
  2042=>"001001000",
  2043=>"111101101",
  2044=>"011100001",
  2045=>"010000000",
  2046=>"010000111",
  2047=>"111010111",
  2048=>"100101101",
  2049=>"110101101",
  2050=>"101010010",
  2051=>"101000010",
  2052=>"011101011",
  2053=>"100110101",
  2054=>"101010010",
  2055=>"000001001",
  2056=>"000000011",
  2057=>"000000110",
  2058=>"000010000",
  2059=>"100011001",
  2060=>"111000001",
  2061=>"100000011",
  2062=>"001110111",
  2063=>"000000010",
  2064=>"000001100",
  2065=>"111111101",
  2066=>"000010111",
  2067=>"111000111",
  2068=>"110100001",
  2069=>"010010111",
  2070=>"001001111",
  2071=>"011000111",
  2072=>"101100111",
  2073=>"111110011",
  2074=>"111101100",
  2075=>"111000110",
  2076=>"110111000",
  2077=>"110010100",
  2078=>"010100101",
  2079=>"110010001",
  2080=>"110011000",
  2081=>"010110101",
  2082=>"010110011",
  2083=>"110010011",
  2084=>"010010101",
  2085=>"110010101",
  2086=>"111101010",
  2087=>"100101111",
  2088=>"110010000",
  2089=>"110110111",
  2090=>"100010100",
  2091=>"011100100",
  2092=>"010000110",
  2093=>"111111111",
  2094=>"111011010",
  2095=>"100111000",
  2096=>"011011001",
  2097=>"011111001",
  2098=>"100111000",
  2099=>"100100111",
  2100=>"000100011",
  2101=>"010000001",
  2102=>"000001110",
  2103=>"110110111",
  2104=>"100111100",
  2105=>"000001010",
  2106=>"000001110",
  2107=>"000101001",
  2108=>"011010011",
  2109=>"000001011",
  2110=>"111010100",
  2111=>"110010000",
  2112=>"010110011",
  2113=>"001110000",
  2114=>"111100010",
  2115=>"111101000",
  2116=>"110110110",
  2117=>"100011110",
  2118=>"010111100",
  2119=>"000011100",
  2120=>"110110011",
  2121=>"010010011",
  2122=>"010111100",
  2123=>"001010010",
  2124=>"011100000",
  2125=>"111101110",
  2126=>"011101001",
  2127=>"000010000",
  2128=>"111011010",
  2129=>"111101000",
  2130=>"010111001",
  2131=>"010110111",
  2132=>"001011010",
  2133=>"110110000",
  2134=>"011010010",
  2135=>"001011011",
  2136=>"000011111",
  2137=>"100011111",
  2138=>"100111100",
  2139=>"100000001",
  2140=>"011010110",
  2141=>"110000100",
  2142=>"001010001",
  2143=>"110101001",
  2144=>"001101010",
  2145=>"000011001",
  2146=>"001001011",
  2147=>"000100010",
  2148=>"011110000",
  2149=>"100000000",
  2150=>"010111110",
  2151=>"001101010",
  2152=>"101110101",
  2153=>"100011101",
  2154=>"000101011",
  2155=>"011111001",
  2156=>"001111010",
  2157=>"011111000",
  2158=>"101101010",
  2159=>"101011010",
  2160=>"110000000",
  2161=>"110110101",
  2162=>"010111010",
  2163=>"011111000",
  2164=>"101011110",
  2165=>"111001110",
  2166=>"111011111",
  2167=>"110100110",
  2168=>"100011100",
  2169=>"101110111",
  2170=>"110101000",
  2171=>"111011110",
  2172=>"010100001",
  2173=>"101110100",
  2174=>"011001000",
  2175=>"000001000",
  2176=>"010000000",
  2177=>"011100111",
  2178=>"001101001",
  2179=>"011001111",
  2180=>"000101000",
  2181=>"001101110",
  2182=>"100011010",
  2183=>"010100010",
  2184=>"100110111",
  2185=>"000001110",
  2186=>"111000011",
  2187=>"000010101",
  2188=>"110001111",
  2189=>"110011110",
  2190=>"111010111",
  2191=>"100110001",
  2192=>"101111110",
  2193=>"101100100",
  2194=>"101101011",
  2195=>"011001000",
  2196=>"010010011",
  2197=>"110100000",
  2198=>"011101110",
  2199=>"010000010",
  2200=>"001000011",
  2201=>"000001000",
  2202=>"001010110",
  2203=>"010010110",
  2204=>"011000111",
  2205=>"001101000",
  2206=>"000011010",
  2207=>"110110000",
  2208=>"010100100",
  2209=>"110101100",
  2210=>"111010000",
  2211=>"000110101",
  2212=>"000111101",
  2213=>"001000000",
  2214=>"001110011",
  2215=>"000000001",
  2216=>"010101111",
  2217=>"010101011",
  2218=>"010001010",
  2219=>"001100011",
  2220=>"110110100",
  2221=>"010100000",
  2222=>"100100010",
  2223=>"111101010",
  2224=>"001000011",
  2225=>"011000001",
  2226=>"010000001",
  2227=>"100001100",
  2228=>"001001010",
  2229=>"011011000",
  2230=>"000010101",
  2231=>"000100100",
  2232=>"111100100",
  2233=>"000110101",
  2234=>"011001000",
  2235=>"111110000",
  2236=>"101111001",
  2237=>"001010111",
  2238=>"001011000",
  2239=>"011110010",
  2240=>"010101000",
  2241=>"100010001",
  2242=>"000110101",
  2243=>"110111000",
  2244=>"001001110",
  2245=>"101001101",
  2246=>"110111110",
  2247=>"101000111",
  2248=>"111001110",
  2249=>"100000011",
  2250=>"110000011",
  2251=>"101110010",
  2252=>"101001100",
  2253=>"101001110",
  2254=>"001010100",
  2255=>"111100110",
  2256=>"111100110",
  2257=>"000110110",
  2258=>"100100101",
  2259=>"110000001",
  2260=>"011101111",
  2261=>"101100101",
  2262=>"111011101",
  2263=>"101001101",
  2264=>"100010010",
  2265=>"000110001",
  2266=>"111110100",
  2267=>"001010001",
  2268=>"011110001",
  2269=>"010001101",
  2270=>"000001000",
  2271=>"111000001",
  2272=>"000010001",
  2273=>"101001111",
  2274=>"100000111",
  2275=>"010110011",
  2276=>"111110101",
  2277=>"001111110",
  2278=>"001010010",
  2279=>"110010000",
  2280=>"010000100",
  2281=>"000111001",
  2282=>"111000001",
  2283=>"000100000",
  2284=>"101011000",
  2285=>"000101000",
  2286=>"111010100",
  2287=>"011100011",
  2288=>"111010001",
  2289=>"010000111",
  2290=>"100001001",
  2291=>"000011110",
  2292=>"101010110",
  2293=>"111111111",
  2294=>"000000100",
  2295=>"000110001",
  2296=>"011100111",
  2297=>"001001010",
  2298=>"101110100",
  2299=>"000011100",
  2300=>"000001101",
  2301=>"101001110",
  2302=>"011001100",
  2303=>"001001101",
  2304=>"100110011",
  2305=>"111001001",
  2306=>"001111111",
  2307=>"100010001",
  2308=>"101101011",
  2309=>"100001011",
  2310=>"001110001",
  2311=>"010011001",
  2312=>"110110100",
  2313=>"101000000",
  2314=>"001101010",
  2315=>"111110000",
  2316=>"000011011",
  2317=>"100001000",
  2318=>"101001110",
  2319=>"000000000",
  2320=>"111111101",
  2321=>"001110010",
  2322=>"110010000",
  2323=>"010110101",
  2324=>"001110101",
  2325=>"111011111",
  2326=>"101011111",
  2327=>"001001011",
  2328=>"010011111",
  2329=>"111000011",
  2330=>"100011101",
  2331=>"001001000",
  2332=>"010101100",
  2333=>"111100011",
  2334=>"101110111",
  2335=>"000000001",
  2336=>"010001100",
  2337=>"000100100",
  2338=>"010110001",
  2339=>"101001111",
  2340=>"111010011",
  2341=>"000010010",
  2342=>"111010111",
  2343=>"011101000",
  2344=>"110011101",
  2345=>"010001100",
  2346=>"000111100",
  2347=>"101010001",
  2348=>"010111101",
  2349=>"100101000",
  2350=>"110000111",
  2351=>"111110110",
  2352=>"111101101",
  2353=>"100100001",
  2354=>"110001101",
  2355=>"000110000",
  2356=>"000001001",
  2357=>"001101111",
  2358=>"110010111",
  2359=>"111001100",
  2360=>"010011111",
  2361=>"011000010",
  2362=>"011001111",
  2363=>"100111011",
  2364=>"111101001",
  2365=>"101110111",
  2366=>"010001100",
  2367=>"100100010",
  2368=>"101111110",
  2369=>"110011010",
  2370=>"110000111",
  2371=>"100000000",
  2372=>"101001111",
  2373=>"010011000",
  2374=>"110111111",
  2375=>"001000001",
  2376=>"010110110",
  2377=>"100000011",
  2378=>"011111110",
  2379=>"010110011",
  2380=>"100111101",
  2381=>"011010110",
  2382=>"101000000",
  2383=>"001011111",
  2384=>"001010010",
  2385=>"011010010",
  2386=>"101110010",
  2387=>"001110101",
  2388=>"001110000",
  2389=>"001111111",
  2390=>"111100000",
  2391=>"100101111",
  2392=>"001000111",
  2393=>"100010111",
  2394=>"101101000",
  2395=>"010110011",
  2396=>"111011111",
  2397=>"011111110",
  2398=>"100101111",
  2399=>"000111001",
  2400=>"001010000",
  2401=>"001010000",
  2402=>"000101111",
  2403=>"101001110",
  2404=>"011011011",
  2405=>"001101110",
  2406=>"001100101",
  2407=>"111000111",
  2408=>"111000010",
  2409=>"000011111",
  2410=>"010101000",
  2411=>"001011001",
  2412=>"001000000",
  2413=>"011011001",
  2414=>"011010010",
  2415=>"010111101",
  2416=>"111100100",
  2417=>"011001011",
  2418=>"000000101",
  2419=>"011101101",
  2420=>"000110010",
  2421=>"010110000",
  2422=>"110100000",
  2423=>"101111100",
  2424=>"110011111",
  2425=>"111001000",
  2426=>"110111100",
  2427=>"101010000",
  2428=>"001000001",
  2429=>"110101001",
  2430=>"111001011",
  2431=>"000011110",
  2432=>"101010110",
  2433=>"001100101",
  2434=>"101111100",
  2435=>"000110010",
  2436=>"000110011",
  2437=>"000001100",
  2438=>"001111010",
  2439=>"000111101",
  2440=>"000010010",
  2441=>"110000110",
  2442=>"101111000",
  2443=>"100011011",
  2444=>"111010000",
  2445=>"100110111",
  2446=>"000010110",
  2447=>"111010110",
  2448=>"011011101",
  2449=>"001001010",
  2450=>"100110001",
  2451=>"000000011",
  2452=>"100001100",
  2453=>"001100101",
  2454=>"001001010",
  2455=>"101010000",
  2456=>"101010011",
  2457=>"001100101",
  2458=>"101001111",
  2459=>"110010100",
  2460=>"001011111",
  2461=>"001100101",
  2462=>"000010001",
  2463=>"101000101",
  2464=>"101110000",
  2465=>"100000010",
  2466=>"101011010",
  2467=>"111000001",
  2468=>"011011011",
  2469=>"110110000",
  2470=>"010000000",
  2471=>"011011000",
  2472=>"010101111",
  2473=>"011101100",
  2474=>"111000111",
  2475=>"111010001",
  2476=>"111011001",
  2477=>"000100011",
  2478=>"011011111",
  2479=>"000000100",
  2480=>"001001110",
  2481=>"001001000",
  2482=>"110010010",
  2483=>"111110010",
  2484=>"100101101",
  2485=>"001111100",
  2486=>"000000111",
  2487=>"011101011",
  2488=>"111010001",
  2489=>"001000100",
  2490=>"000101110",
  2491=>"010001001",
  2492=>"000001000",
  2493=>"101100000",
  2494=>"011001010",
  2495=>"011101010",
  2496=>"110000101",
  2497=>"100101110",
  2498=>"111001110",
  2499=>"001111000",
  2500=>"100111110",
  2501=>"111101110",
  2502=>"001001001",
  2503=>"010000000",
  2504=>"110111100",
  2505=>"111101110",
  2506=>"010010101",
  2507=>"111001000",
  2508=>"011001101",
  2509=>"010110010",
  2510=>"000000010",
  2511=>"101000101",
  2512=>"110010101",
  2513=>"100000001",
  2514=>"100001111",
  2515=>"111101100",
  2516=>"110111011",
  2517=>"010001100",
  2518=>"011101101",
  2519=>"111011001",
  2520=>"001000000",
  2521=>"000100001",
  2522=>"001111111",
  2523=>"100010001",
  2524=>"010100011",
  2525=>"001001001",
  2526=>"010001010",
  2527=>"010000110",
  2528=>"100011110",
  2529=>"000101000",
  2530=>"101110001",
  2531=>"011000101",
  2532=>"001011010",
  2533=>"011010001",
  2534=>"101000000",
  2535=>"000101101",
  2536=>"010010001",
  2537=>"000010101",
  2538=>"000000101",
  2539=>"011000000",
  2540=>"110100100",
  2541=>"000111101",
  2542=>"000111101",
  2543=>"001000111",
  2544=>"011010001",
  2545=>"101111110",
  2546=>"110111001",
  2547=>"111000000",
  2548=>"010101100",
  2549=>"101000000",
  2550=>"000110101",
  2551=>"001000101",
  2552=>"000010101",
  2553=>"101100001",
  2554=>"101000111",
  2555=>"101111111",
  2556=>"111101101",
  2557=>"100011101",
  2558=>"110011000",
  2559=>"000100111",
  2560=>"111110110",
  2561=>"100101100",
  2562=>"001001101",
  2563=>"011010111",
  2564=>"100001001",
  2565=>"100010111",
  2566=>"100111111",
  2567=>"000000100",
  2568=>"010001001",
  2569=>"100110101",
  2570=>"100001111",
  2571=>"010010111",
  2572=>"100111101",
  2573=>"111000110",
  2574=>"000011101",
  2575=>"011011101",
  2576=>"001011111",
  2577=>"001110001",
  2578=>"011011111",
  2579=>"101111111",
  2580=>"010001010",
  2581=>"111100001",
  2582=>"000001011",
  2583=>"101011111",
  2584=>"101001111",
  2585=>"101001111",
  2586=>"111011000",
  2587=>"100011101",
  2588=>"011001110",
  2589=>"111101011",
  2590=>"100001011",
  2591=>"111100101",
  2592=>"010100110",
  2593=>"101111011",
  2594=>"000011111",
  2595=>"011001010",
  2596=>"010110001",
  2597=>"101001101",
  2598=>"100011010",
  2599=>"100111011",
  2600=>"011010101",
  2601=>"011100011",
  2602=>"011001011",
  2603=>"010110110",
  2604=>"010110110",
  2605=>"111100100",
  2606=>"111011101",
  2607=>"001000000",
  2608=>"111101001",
  2609=>"010001000",
  2610=>"101100000",
  2611=>"111101010",
  2612=>"100100110",
  2613=>"011111010",
  2614=>"010100010",
  2615=>"011000101",
  2616=>"110000110",
  2617=>"101100100",
  2618=>"001011010",
  2619=>"010111011",
  2620=>"010001111",
  2621=>"010010000",
  2622=>"101011110",
  2623=>"010101001",
  2624=>"101110000",
  2625=>"110101110",
  2626=>"111100100",
  2627=>"100001100",
  2628=>"000000100",
  2629=>"110000101",
  2630=>"011000110",
  2631=>"100011000",
  2632=>"000010001",
  2633=>"111011100",
  2634=>"001010110",
  2635=>"001111111",
  2636=>"011101100",
  2637=>"010000010",
  2638=>"111100010",
  2639=>"101011000",
  2640=>"001011101",
  2641=>"111101111",
  2642=>"000011000",
  2643=>"001000011",
  2644=>"101100011",
  2645=>"111111101",
  2646=>"001100011",
  2647=>"101110110",
  2648=>"110101011",
  2649=>"101010010",
  2650=>"100110001",
  2651=>"010001100",
  2652=>"000001010",
  2653=>"000111111",
  2654=>"111001110",
  2655=>"110001000",
  2656=>"111011001",
  2657=>"110010000",
  2658=>"100010110",
  2659=>"101100111",
  2660=>"010001010",
  2661=>"001111001",
  2662=>"000111011",
  2663=>"001101011",
  2664=>"111001001",
  2665=>"101000011",
  2666=>"010011111",
  2667=>"010011100",
  2668=>"100001011",
  2669=>"000000110",
  2670=>"100111111",
  2671=>"010111101",
  2672=>"001010100",
  2673=>"010000000",
  2674=>"010000001",
  2675=>"111100110",
  2676=>"110111110",
  2677=>"000010011",
  2678=>"001100101",
  2679=>"110111101",
  2680=>"111001000",
  2681=>"000011111",
  2682=>"001101000",
  2683=>"001111111",
  2684=>"001110010",
  2685=>"111111111",
  2686=>"000000001",
  2687=>"111100101",
  2688=>"101000010",
  2689=>"100110111",
  2690=>"001111110",
  2691=>"010001011",
  2692=>"111000010",
  2693=>"000000110",
  2694=>"101111010",
  2695=>"110100101",
  2696=>"110000001",
  2697=>"101111110",
  2698=>"010110001",
  2699=>"010111111",
  2700=>"110110010",
  2701=>"011111110",
  2702=>"111000011",
  2703=>"011010000",
  2704=>"101100011",
  2705=>"011100010",
  2706=>"000001100",
  2707=>"010010101",
  2708=>"001000010",
  2709=>"110000100",
  2710=>"001000000",
  2711=>"101001100",
  2712=>"001101101",
  2713=>"110100000",
  2714=>"101110101",
  2715=>"100100100",
  2716=>"011011001",
  2717=>"001100010",
  2718=>"111001010",
  2719=>"000110011",
  2720=>"010101101",
  2721=>"110000110",
  2722=>"100000110",
  2723=>"101101110",
  2724=>"010101010",
  2725=>"011111111",
  2726=>"110000110",
  2727=>"110111100",
  2728=>"100010101",
  2729=>"001010011",
  2730=>"000100111",
  2731=>"110000010",
  2732=>"100001010",
  2733=>"011000100",
  2734=>"110100100",
  2735=>"110100011",
  2736=>"110000001",
  2737=>"001010001",
  2738=>"000111110",
  2739=>"011100111",
  2740=>"010000001",
  2741=>"011011011",
  2742=>"111100011",
  2743=>"110110100",
  2744=>"100111001",
  2745=>"011111000",
  2746=>"110110001",
  2747=>"000001111",
  2748=>"101100100",
  2749=>"111000110",
  2750=>"100101011",
  2751=>"011110011",
  2752=>"111110101",
  2753=>"101101100",
  2754=>"000000101",
  2755=>"111100010",
  2756=>"101001100",
  2757=>"110101100",
  2758=>"010010001",
  2759=>"100000110",
  2760=>"000100000",
  2761=>"111110101",
  2762=>"010101101",
  2763=>"100110011",
  2764=>"111001100",
  2765=>"000001000",
  2766=>"110000100",
  2767=>"111010001",
  2768=>"010100000",
  2769=>"001010111",
  2770=>"011000101",
  2771=>"011001001",
  2772=>"000110010",
  2773=>"000001110",
  2774=>"010000000",
  2775=>"100101100",
  2776=>"000011111",
  2777=>"010001101",
  2778=>"111010001",
  2779=>"001000110",
  2780=>"000111110",
  2781=>"110001000",
  2782=>"100100101",
  2783=>"101011000",
  2784=>"111000111",
  2785=>"000000100",
  2786=>"011010011",
  2787=>"010111010",
  2788=>"001110001",
  2789=>"111110100",
  2790=>"101101000",
  2791=>"000011001",
  2792=>"001110010",
  2793=>"111011101",
  2794=>"101001111",
  2795=>"111011011",
  2796=>"000000000",
  2797=>"101010001",
  2798=>"010000000",
  2799=>"001110111",
  2800=>"011110100",
  2801=>"000101011",
  2802=>"010011011",
  2803=>"101011011",
  2804=>"000101100",
  2805=>"001001011",
  2806=>"001001110",
  2807=>"100000111",
  2808=>"100111110",
  2809=>"101111010",
  2810=>"010100001",
  2811=>"001100011",
  2812=>"110101100",
  2813=>"111000001",
  2814=>"101100000",
  2815=>"000000111",
  2816=>"111001101",
  2817=>"111010000",
  2818=>"011101001",
  2819=>"111001000",
  2820=>"101010000",
  2821=>"001100010",
  2822=>"001001010",
  2823=>"111011101",
  2824=>"001011011",
  2825=>"000100111",
  2826=>"101100001",
  2827=>"010100001",
  2828=>"001111010",
  2829=>"100010100",
  2830=>"100010010",
  2831=>"001100101",
  2832=>"010100110",
  2833=>"000001101",
  2834=>"110011110",
  2835=>"100111000",
  2836=>"101101101",
  2837=>"100100101",
  2838=>"101101110",
  2839=>"111001101",
  2840=>"010010100",
  2841=>"000100101",
  2842=>"000000101",
  2843=>"111101100",
  2844=>"000001100",
  2845=>"110000111",
  2846=>"001100110",
  2847=>"111010000",
  2848=>"001011100",
  2849=>"011110010",
  2850=>"110000000",
  2851=>"111111101",
  2852=>"011000100",
  2853=>"111000111",
  2854=>"110100001",
  2855=>"010111000",
  2856=>"001010001",
  2857=>"111100100",
  2858=>"000010000",
  2859=>"100010100",
  2860=>"010110001",
  2861=>"000001000",
  2862=>"011100011",
  2863=>"000100101",
  2864=>"000100000",
  2865=>"101000101",
  2866=>"100111101",
  2867=>"000111011",
  2868=>"101000101",
  2869=>"001010100",
  2870=>"000001000",
  2871=>"001000111",
  2872=>"101111011",
  2873=>"000111111",
  2874=>"111000000",
  2875=>"001000010",
  2876=>"000111100",
  2877=>"001011110",
  2878=>"011100100",
  2879=>"011011001",
  2880=>"101001000",
  2881=>"111111111",
  2882=>"110110101",
  2883=>"100000001",
  2884=>"100001100",
  2885=>"010101001",
  2886=>"000001011",
  2887=>"110011111",
  2888=>"001000100",
  2889=>"111101001",
  2890=>"101110111",
  2891=>"000001010",
  2892=>"111100010",
  2893=>"110111010",
  2894=>"001010100",
  2895=>"110101001",
  2896=>"111010110",
  2897=>"110001101",
  2898=>"100001000",
  2899=>"000000111",
  2900=>"010111010",
  2901=>"011111011",
  2902=>"001011110",
  2903=>"010100110",
  2904=>"111011110",
  2905=>"111010001",
  2906=>"101100010",
  2907=>"111100110",
  2908=>"101100000",
  2909=>"111101000",
  2910=>"101001100",
  2911=>"011000101",
  2912=>"011110010",
  2913=>"001011010",
  2914=>"110111100",
  2915=>"010000010",
  2916=>"001101000",
  2917=>"000001001",
  2918=>"011000101",
  2919=>"110101111",
  2920=>"010100100",
  2921=>"111001111",
  2922=>"000000100",
  2923=>"000000101",
  2924=>"101011100",
  2925=>"000100101",
  2926=>"000010010",
  2927=>"111011111",
  2928=>"111011000",
  2929=>"101010011",
  2930=>"100010101",
  2931=>"101010110",
  2932=>"001101111",
  2933=>"000010010",
  2934=>"111101000",
  2935=>"100100100",
  2936=>"111000000",
  2937=>"111010111",
  2938=>"010100001",
  2939=>"100111010",
  2940=>"000010100",
  2941=>"011000011",
  2942=>"100001110",
  2943=>"100001111",
  2944=>"011101011",
  2945=>"111111001",
  2946=>"101000100",
  2947=>"010001110",
  2948=>"000000100",
  2949=>"100101001",
  2950=>"100111010",
  2951=>"010010101",
  2952=>"011010110",
  2953=>"111011000",
  2954=>"001010000",
  2955=>"111010110",
  2956=>"011010010",
  2957=>"101000000",
  2958=>"110001001",
  2959=>"100110101",
  2960=>"101101101",
  2961=>"111100001",
  2962=>"000110110",
  2963=>"010010101",
  2964=>"100011110",
  2965=>"010110011",
  2966=>"110100001",
  2967=>"101010100",
  2968=>"100101101",
  2969=>"100010111",
  2970=>"000011111",
  2971=>"001010000",
  2972=>"011000010",
  2973=>"011100000",
  2974=>"111011001",
  2975=>"000101011",
  2976=>"101001001",
  2977=>"101110000",
  2978=>"000011000",
  2979=>"111100100",
  2980=>"010000100",
  2981=>"011101100",
  2982=>"110110101",
  2983=>"100000001",
  2984=>"000011101",
  2985=>"010111010",
  2986=>"001101000",
  2987=>"011100000",
  2988=>"100100000",
  2989=>"101010101",
  2990=>"000010110",
  2991=>"011011110",
  2992=>"011010011",
  2993=>"011110011",
  2994=>"011110000",
  2995=>"101111110",
  2996=>"110000010",
  2997=>"110100010",
  2998=>"101111110",
  2999=>"000000110",
  3000=>"010101100",
  3001=>"101110010",
  3002=>"000001111",
  3003=>"111010011",
  3004=>"010001000",
  3005=>"001000000",
  3006=>"010111011",
  3007=>"100101001",
  3008=>"001111100",
  3009=>"110010011",
  3010=>"000101001",
  3011=>"000000000",
  3012=>"110110011",
  3013=>"001101000",
  3014=>"000010000",
  3015=>"000000100",
  3016=>"001100000",
  3017=>"001100100",
  3018=>"010011101",
  3019=>"111001000",
  3020=>"001100110",
  3021=>"011000000",
  3022=>"100000000",
  3023=>"000111111",
  3024=>"100011110",
  3025=>"001001011",
  3026=>"001110101",
  3027=>"110010110",
  3028=>"110111001",
  3029=>"111101011",
  3030=>"110000011",
  3031=>"011101111",
  3032=>"011110001",
  3033=>"111100101",
  3034=>"110110000",
  3035=>"011011010",
  3036=>"110011101",
  3037=>"110101101",
  3038=>"110011001",
  3039=>"100000110",
  3040=>"001001010",
  3041=>"011010001",
  3042=>"000001001",
  3043=>"110101110",
  3044=>"000001110",
  3045=>"011101100",
  3046=>"010010010",
  3047=>"000010001",
  3048=>"000100010",
  3049=>"011001100",
  3050=>"111001110",
  3051=>"101000101",
  3052=>"110010100",
  3053=>"011010011",
  3054=>"000110100",
  3055=>"110110011",
  3056=>"000010100",
  3057=>"001111101",
  3058=>"001010111",
  3059=>"111100011",
  3060=>"010101111",
  3061=>"011011111",
  3062=>"000000100",
  3063=>"100111111",
  3064=>"011001111",
  3065=>"001000000",
  3066=>"011111100",
  3067=>"010010010",
  3068=>"100011011",
  3069=>"010011100",
  3070=>"110000010",
  3071=>"111111101",
  3072=>"000001011",
  3073=>"010110010",
  3074=>"110100001",
  3075=>"110000001",
  3076=>"111011000",
  3077=>"100001000",
  3078=>"010111110",
  3079=>"100101001",
  3080=>"111001001",
  3081=>"010011000",
  3082=>"000011110",
  3083=>"100011010",
  3084=>"100001011",
  3085=>"011100101",
  3086=>"001111001",
  3087=>"111101010",
  3088=>"100000010",
  3089=>"001011001",
  3090=>"100001100",
  3091=>"100100010",
  3092=>"011100011",
  3093=>"100101111",
  3094=>"011100100",
  3095=>"101000001",
  3096=>"001000010",
  3097=>"111000010",
  3098=>"010101110",
  3099=>"111111001",
  3100=>"101101101",
  3101=>"100011000",
  3102=>"011011111",
  3103=>"001000000",
  3104=>"010100011",
  3105=>"000100000",
  3106=>"000110000",
  3107=>"010111011",
  3108=>"010010100",
  3109=>"110011111",
  3110=>"101011000",
  3111=>"100001000",
  3112=>"011110000",
  3113=>"010010001",
  3114=>"110000011",
  3115=>"110011111",
  3116=>"010110010",
  3117=>"010000010",
  3118=>"100011001",
  3119=>"000010011",
  3120=>"110100011",
  3121=>"010100111",
  3122=>"001010011",
  3123=>"111011111",
  3124=>"010011010",
  3125=>"110101000",
  3126=>"000010000",
  3127=>"000001011",
  3128=>"001110100",
  3129=>"000111101",
  3130=>"000100000",
  3131=>"000010110",
  3132=>"000011111",
  3133=>"000011011",
  3134=>"010011110",
  3135=>"001010101",
  3136=>"110100000",
  3137=>"101110101",
  3138=>"001110000",
  3139=>"000011110",
  3140=>"010010111",
  3141=>"110011110",
  3142=>"010001111",
  3143=>"010000010",
  3144=>"001000000",
  3145=>"001100010",
  3146=>"100011101",
  3147=>"100111110",
  3148=>"100101000",
  3149=>"111001011",
  3150=>"101110010",
  3151=>"100100001",
  3152=>"000001111",
  3153=>"110000000",
  3154=>"101000001",
  3155=>"100101110",
  3156=>"001001001",
  3157=>"101011000",
  3158=>"110001000",
  3159=>"011011110",
  3160=>"111011001",
  3161=>"001010101",
  3162=>"010011100",
  3163=>"100100100",
  3164=>"010101110",
  3165=>"000001101",
  3166=>"000110111",
  3167=>"001000001",
  3168=>"101110111",
  3169=>"101000010",
  3170=>"001000011",
  3171=>"001011011",
  3172=>"000110111",
  3173=>"100010100",
  3174=>"100010000",
  3175=>"000111110",
  3176=>"000101100",
  3177=>"000011101",
  3178=>"100111101",
  3179=>"100100011",
  3180=>"001001111",
  3181=>"101001000",
  3182=>"110000000",
  3183=>"100001110",
  3184=>"100001000",
  3185=>"100000011",
  3186=>"001110111",
  3187=>"111011111",
  3188=>"000011100",
  3189=>"010110111",
  3190=>"101101100",
  3191=>"000111001",
  3192=>"000100110",
  3193=>"110101101",
  3194=>"011101100",
  3195=>"100000111",
  3196=>"101100001",
  3197=>"011001010",
  3198=>"010101011",
  3199=>"100001010",
  3200=>"101010010",
  3201=>"010000010",
  3202=>"001001110",
  3203=>"101111011",
  3204=>"010111010",
  3205=>"101110000",
  3206=>"000010011",
  3207=>"110110111",
  3208=>"001010010",
  3209=>"110001011",
  3210=>"111000001",
  3211=>"011000010",
  3212=>"101111111",
  3213=>"001110010",
  3214=>"001111000",
  3215=>"111001011",
  3216=>"101111010",
  3217=>"010011010",
  3218=>"001010000",
  3219=>"101100001",
  3220=>"101001101",
  3221=>"010110000",
  3222=>"001001010",
  3223=>"010110001",
  3224=>"011110000",
  3225=>"000110010",
  3226=>"001001110",
  3227=>"100100100",
  3228=>"001011000",
  3229=>"010010101",
  3230=>"110010111",
  3231=>"101100011",
  3232=>"000111111",
  3233=>"011001111",
  3234=>"000100111",
  3235=>"101101111",
  3236=>"011011000",
  3237=>"111101101",
  3238=>"111110001",
  3239=>"110110011",
  3240=>"111101100",
  3241=>"110110001",
  3242=>"000000111",
  3243=>"101110011",
  3244=>"101111100",
  3245=>"110101011",
  3246=>"001001010",
  3247=>"000010100",
  3248=>"000101010",
  3249=>"011000100",
  3250=>"011100111",
  3251=>"000000110",
  3252=>"110100110",
  3253=>"101111111",
  3254=>"010110000",
  3255=>"000110001",
  3256=>"000111111",
  3257=>"010111111",
  3258=>"010100001",
  3259=>"100110110",
  3260=>"100001000",
  3261=>"100010111",
  3262=>"011011101",
  3263=>"011010111",
  3264=>"111011100",
  3265=>"010000111",
  3266=>"001111010",
  3267=>"011111110",
  3268=>"111011010",
  3269=>"001100111",
  3270=>"101011101",
  3271=>"111011101",
  3272=>"111101100",
  3273=>"101111010",
  3274=>"111011111",
  3275=>"011101011",
  3276=>"000010001",
  3277=>"010000001",
  3278=>"100001010",
  3279=>"111110101",
  3280=>"000101010",
  3281=>"101000000",
  3282=>"001000101",
  3283=>"101101100",
  3284=>"101100100",
  3285=>"110101100",
  3286=>"110000101",
  3287=>"111100100",
  3288=>"101101000",
  3289=>"100110011",
  3290=>"010000101",
  3291=>"011110101",
  3292=>"001001110",
  3293=>"100001100",
  3294=>"000010001",
  3295=>"001100010",
  3296=>"100000011",
  3297=>"010001101",
  3298=>"010110111",
  3299=>"101111001",
  3300=>"001010001",
  3301=>"110101110",
  3302=>"000110010",
  3303=>"100111010",
  3304=>"110110110",
  3305=>"001100000",
  3306=>"010101111",
  3307=>"101101010",
  3308=>"001010010",
  3309=>"111100010",
  3310=>"110101000",
  3311=>"110011000",
  3312=>"110110100",
  3313=>"100010111",
  3314=>"011110111",
  3315=>"001100101",
  3316=>"110010110",
  3317=>"111100000",
  3318=>"000000001",
  3319=>"000001000",
  3320=>"000001010",
  3321=>"101111110",
  3322=>"001111001",
  3323=>"010001111",
  3324=>"011111110",
  3325=>"001101100",
  3326=>"111011101",
  3327=>"010000101",
  3328=>"110111011",
  3329=>"101000001",
  3330=>"111101101",
  3331=>"111101110",
  3332=>"101001000",
  3333=>"111000000",
  3334=>"100010000",
  3335=>"101011101",
  3336=>"000110010",
  3337=>"010110011",
  3338=>"100000100",
  3339=>"111001000",
  3340=>"100100111",
  3341=>"000101111",
  3342=>"011111100",
  3343=>"000101001",
  3344=>"011110101",
  3345=>"000001011",
  3346=>"111110011",
  3347=>"011011110",
  3348=>"000111111",
  3349=>"011001000",
  3350=>"011010110",
  3351=>"011101110",
  3352=>"011010111",
  3353=>"110001101",
  3354=>"001001111",
  3355=>"111110001",
  3356=>"010010010",
  3357=>"100000001",
  3358=>"011100000",
  3359=>"000010001",
  3360=>"000000111",
  3361=>"001101100",
  3362=>"011111001",
  3363=>"001010100",
  3364=>"111100000",
  3365=>"010001110",
  3366=>"110101000",
  3367=>"101100100",
  3368=>"100100110",
  3369=>"000111001",
  3370=>"010000000",
  3371=>"011111000",
  3372=>"101011011",
  3373=>"100100111",
  3374=>"011001000",
  3375=>"111110110",
  3376=>"011011000",
  3377=>"100001110",
  3378=>"000100100",
  3379=>"000011101",
  3380=>"111000001",
  3381=>"011111000",
  3382=>"011111100",
  3383=>"101111101",
  3384=>"000000110",
  3385=>"011101011",
  3386=>"111011101",
  3387=>"111101000",
  3388=>"100011101",
  3389=>"001100000",
  3390=>"110111101",
  3391=>"110100001",
  3392=>"101101010",
  3393=>"101011001",
  3394=>"100111110",
  3395=>"011010000",
  3396=>"010010111",
  3397=>"101100011",
  3398=>"111010010",
  3399=>"011101101",
  3400=>"110110111",
  3401=>"111011000",
  3402=>"101101011",
  3403=>"101001011",
  3404=>"101111100",
  3405=>"000011010",
  3406=>"111110010",
  3407=>"001010101",
  3408=>"001101010",
  3409=>"011011000",
  3410=>"111101100",
  3411=>"100110001",
  3412=>"011111100",
  3413=>"000010010",
  3414=>"011111101",
  3415=>"010010110",
  3416=>"000010100",
  3417=>"000101101",
  3418=>"001100010",
  3419=>"001000000",
  3420=>"110011000",
  3421=>"001111111",
  3422=>"111011111",
  3423=>"000000101",
  3424=>"010010001",
  3425=>"110110010",
  3426=>"010011001",
  3427=>"010001111",
  3428=>"110110101",
  3429=>"010100000",
  3430=>"110000110",
  3431=>"000100011",
  3432=>"001111011",
  3433=>"010001111",
  3434=>"100001111",
  3435=>"011010010",
  3436=>"111111111",
  3437=>"101011100",
  3438=>"010001100",
  3439=>"101010111",
  3440=>"000010000",
  3441=>"010100100",
  3442=>"010010110",
  3443=>"111100011",
  3444=>"000101000",
  3445=>"010001101",
  3446=>"100110010",
  3447=>"010000011",
  3448=>"001000111",
  3449=>"001010011",
  3450=>"101010110",
  3451=>"100110011",
  3452=>"101010001",
  3453=>"111001110",
  3454=>"110010001",
  3455=>"011000011",
  3456=>"001001111",
  3457=>"000100101",
  3458=>"100101000",
  3459=>"000000011",
  3460=>"100011101",
  3461=>"100111101",
  3462=>"010100111",
  3463=>"000111001",
  3464=>"101110001",
  3465=>"101110111",
  3466=>"101110010",
  3467=>"011111111",
  3468=>"110111001",
  3469=>"001001000",
  3470=>"011111001",
  3471=>"100000110",
  3472=>"010111101",
  3473=>"000011011",
  3474=>"100011101",
  3475=>"010000100",
  3476=>"010000001",
  3477=>"011101010",
  3478=>"111101011",
  3479=>"110111111",
  3480=>"100101000",
  3481=>"001001011",
  3482=>"110101101",
  3483=>"101111011",
  3484=>"100000001",
  3485=>"000000000",
  3486=>"011011111",
  3487=>"011011111",
  3488=>"110010111",
  3489=>"101011110",
  3490=>"000011011",
  3491=>"111101010",
  3492=>"110111110",
  3493=>"010000110",
  3494=>"110110001",
  3495=>"111011010",
  3496=>"100001010",
  3497=>"111101101",
  3498=>"000101001",
  3499=>"100000000",
  3500=>"100010111",
  3501=>"101001100",
  3502=>"010111011",
  3503=>"100011101",
  3504=>"100010111",
  3505=>"101111001",
  3506=>"110100100",
  3507=>"111101111",
  3508=>"001011010",
  3509=>"011110010",
  3510=>"000010010",
  3511=>"111100100",
  3512=>"001001001",
  3513=>"110101111",
  3514=>"011011111",
  3515=>"101010110",
  3516=>"111110101",
  3517=>"110110011",
  3518=>"000001100",
  3519=>"100111100",
  3520=>"101011111",
  3521=>"010001100",
  3522=>"001101001",
  3523=>"110010000",
  3524=>"110001000",
  3525=>"111001110",
  3526=>"000100101",
  3527=>"001101111",
  3528=>"011101111",
  3529=>"111101001",
  3530=>"001100111",
  3531=>"100101110",
  3532=>"001101110",
  3533=>"010100111",
  3534=>"010110100",
  3535=>"010001010",
  3536=>"001001001",
  3537=>"001011000",
  3538=>"101001011",
  3539=>"001001000",
  3540=>"010000000",
  3541=>"111001000",
  3542=>"111000000",
  3543=>"111011001",
  3544=>"000101010",
  3545=>"110010100",
  3546=>"001010010",
  3547=>"000111001",
  3548=>"101101000",
  3549=>"000100011",
  3550=>"111100001",
  3551=>"100010010",
  3552=>"101111100",
  3553=>"111100110",
  3554=>"110011111",
  3555=>"111001010",
  3556=>"111000100",
  3557=>"011111000",
  3558=>"010111100",
  3559=>"000101000",
  3560=>"000000011",
  3561=>"000100101",
  3562=>"000010010",
  3563=>"010101000",
  3564=>"010110101",
  3565=>"111100100",
  3566=>"111111011",
  3567=>"110111000",
  3568=>"010110100",
  3569=>"001111111",
  3570=>"010001000",
  3571=>"001011110",
  3572=>"100001010",
  3573=>"101010011",
  3574=>"101101111",
  3575=>"000100011",
  3576=>"111011011",
  3577=>"011111000",
  3578=>"011111111",
  3579=>"010111110",
  3580=>"101101001",
  3581=>"001110000",
  3582=>"101000000",
  3583=>"100110111",
  3584=>"101010101",
  3585=>"010100111",
  3586=>"100100000",
  3587=>"011000100",
  3588=>"101110111",
  3589=>"001011011",
  3590=>"000100100",
  3591=>"010011100",
  3592=>"011100101",
  3593=>"100010110",
  3594=>"100010111",
  3595=>"000110110",
  3596=>"011011111",
  3597=>"100101100",
  3598=>"100100101",
  3599=>"100010010",
  3600=>"100010100",
  3601=>"010011000",
  3602=>"001010101",
  3603=>"011101000",
  3604=>"101010010",
  3605=>"000010000",
  3606=>"101100010",
  3607=>"011111011",
  3608=>"101100110",
  3609=>"001011110",
  3610=>"100001111",
  3611=>"110001111",
  3612=>"010001010",
  3613=>"111010010",
  3614=>"110100010",
  3615=>"101110111",
  3616=>"010010000",
  3617=>"101100101",
  3618=>"000000100",
  3619=>"101001011",
  3620=>"001010100",
  3621=>"010111011",
  3622=>"110110111",
  3623=>"100001010",
  3624=>"000101100",
  3625=>"001011000",
  3626=>"100011111",
  3627=>"010011110",
  3628=>"100010110",
  3629=>"101111110",
  3630=>"000001001",
  3631=>"010011010",
  3632=>"110101110",
  3633=>"110111111",
  3634=>"101101011",
  3635=>"110010000",
  3636=>"010011111",
  3637=>"110111000",
  3638=>"011110000",
  3639=>"011100010",
  3640=>"111010100",
  3641=>"111100011",
  3642=>"100101100",
  3643=>"101100111",
  3644=>"000001110",
  3645=>"000010011",
  3646=>"000000100",
  3647=>"010001000",
  3648=>"011010011",
  3649=>"100000101",
  3650=>"111001101",
  3651=>"000011111",
  3652=>"001000010",
  3653=>"000100100",
  3654=>"011001010",
  3655=>"000011001",
  3656=>"000011111",
  3657=>"001001110",
  3658=>"010100000",
  3659=>"100101010",
  3660=>"101010001",
  3661=>"011011011",
  3662=>"101100111",
  3663=>"101111100",
  3664=>"101101101",
  3665=>"011110000",
  3666=>"011101010",
  3667=>"000100011",
  3668=>"010111101",
  3669=>"100011100",
  3670=>"001010111",
  3671=>"010110111",
  3672=>"100001010",
  3673=>"000001011",
  3674=>"111110010",
  3675=>"001000111",
  3676=>"011000101",
  3677=>"111101001",
  3678=>"000001001",
  3679=>"110110000",
  3680=>"101000111",
  3681=>"001011001",
  3682=>"011011001",
  3683=>"011010110",
  3684=>"000100101",
  3685=>"110101000",
  3686=>"111010000",
  3687=>"001110110",
  3688=>"000010011",
  3689=>"001010110",
  3690=>"001110001",
  3691=>"001001000",
  3692=>"010000111",
  3693=>"001011000",
  3694=>"100110001",
  3695=>"100110100",
  3696=>"111100000",
  3697=>"000001110",
  3698=>"001111011",
  3699=>"001101111",
  3700=>"101011111",
  3701=>"111011100",
  3702=>"110001100",
  3703=>"010110111",
  3704=>"101101001",
  3705=>"000110011",
  3706=>"011000000",
  3707=>"111010100",
  3708=>"001001100",
  3709=>"110011010",
  3710=>"101111111",
  3711=>"100100010",
  3712=>"101000110",
  3713=>"110100011",
  3714=>"101010001",
  3715=>"001010101",
  3716=>"010010110",
  3717=>"110101001",
  3718=>"110101101",
  3719=>"101101010",
  3720=>"011101000",
  3721=>"111001001",
  3722=>"010100101",
  3723=>"011110000",
  3724=>"100001100",
  3725=>"010011110",
  3726=>"100100011",
  3727=>"000010000",
  3728=>"111010000",
  3729=>"010010101",
  3730=>"110100110",
  3731=>"010110011",
  3732=>"100000011",
  3733=>"000000100",
  3734=>"111001100",
  3735=>"111100110",
  3736=>"110110010",
  3737=>"101101111",
  3738=>"000101110",
  3739=>"110010011",
  3740=>"011101110",
  3741=>"001110011",
  3742=>"111000100",
  3743=>"111011110",
  3744=>"101110110",
  3745=>"011000110",
  3746=>"101110100",
  3747=>"010010010",
  3748=>"111110011",
  3749=>"111111111",
  3750=>"101001011",
  3751=>"110101000",
  3752=>"101100001",
  3753=>"100000001",
  3754=>"001100101",
  3755=>"110110110",
  3756=>"101101011",
  3757=>"100001111",
  3758=>"011101011",
  3759=>"000001111",
  3760=>"001011000",
  3761=>"001000010",
  3762=>"011100100",
  3763=>"010000001",
  3764=>"010000001",
  3765=>"110110100",
  3766=>"100010000",
  3767=>"101000110",
  3768=>"011100001",
  3769=>"010111000",
  3770=>"011000111",
  3771=>"100001100",
  3772=>"010000011",
  3773=>"011111011",
  3774=>"011010011",
  3775=>"011110000",
  3776=>"010111100",
  3777=>"110000101",
  3778=>"111010110",
  3779=>"010111111",
  3780=>"111100000",
  3781=>"111010110",
  3782=>"111110110",
  3783=>"100011110",
  3784=>"011010011",
  3785=>"000000010",
  3786=>"011100010",
  3787=>"011011110",
  3788=>"110100000",
  3789=>"110101010",
  3790=>"011010000",
  3791=>"011110110",
  3792=>"111000010",
  3793=>"110110110",
  3794=>"010001111",
  3795=>"000001011",
  3796=>"001110110",
  3797=>"101100101",
  3798=>"101101111",
  3799=>"011001110",
  3800=>"000000001",
  3801=>"110111100",
  3802=>"111101001",
  3803=>"101010010",
  3804=>"111101100",
  3805=>"100110111",
  3806=>"001111100",
  3807=>"111111101",
  3808=>"001011001",
  3809=>"011110110",
  3810=>"000100110",
  3811=>"011001110",
  3812=>"101010010",
  3813=>"011000111",
  3814=>"011010010",
  3815=>"110110011",
  3816=>"010100011",
  3817=>"100001101",
  3818=>"111000011",
  3819=>"110100110",
  3820=>"001110111",
  3821=>"101000100",
  3822=>"000110000",
  3823=>"000000010",
  3824=>"010001011",
  3825=>"000111100",
  3826=>"001011100",
  3827=>"010011000",
  3828=>"101100001",
  3829=>"001100111",
  3830=>"001010100",
  3831=>"010010001",
  3832=>"011011110",
  3833=>"011000111",
  3834=>"110111000",
  3835=>"011000000",
  3836=>"010000000",
  3837=>"000011001",
  3838=>"000111001",
  3839=>"000011000",
  3840=>"110010100",
  3841=>"000000010",
  3842=>"000011001",
  3843=>"011001101",
  3844=>"011000001",
  3845=>"110001101",
  3846=>"000011100",
  3847=>"111000100",
  3848=>"110010010",
  3849=>"101111100",
  3850=>"101111011",
  3851=>"010001011",
  3852=>"010111001",
  3853=>"000100111",
  3854=>"000111110",
  3855=>"110100110",
  3856=>"110011101",
  3857=>"111011110",
  3858=>"111101011",
  3859=>"010000111",
  3860=>"100001011",
  3861=>"100010001",
  3862=>"111110001",
  3863=>"010000011",
  3864=>"010011010",
  3865=>"000011111",
  3866=>"010110010",
  3867=>"100000001",
  3868=>"011101001",
  3869=>"000111001",
  3870=>"011001100",
  3871=>"100000000",
  3872=>"101000000",
  3873=>"111010101",
  3874=>"101100011",
  3875=>"011011000",
  3876=>"011101110",
  3877=>"001100100",
  3878=>"100011001",
  3879=>"101011011",
  3880=>"000111111",
  3881=>"101000011",
  3882=>"011110110",
  3883=>"111110100",
  3884=>"101100100",
  3885=>"001011101",
  3886=>"000010001",
  3887=>"110101101",
  3888=>"011000011",
  3889=>"100010111",
  3890=>"111111001",
  3891=>"011101100",
  3892=>"111000111",
  3893=>"001101000",
  3894=>"100011000",
  3895=>"101010101",
  3896=>"000001111",
  3897=>"101111110",
  3898=>"111111111",
  3899=>"110010110",
  3900=>"011101011",
  3901=>"010110001",
  3902=>"001001010",
  3903=>"000101001",
  3904=>"111101100",
  3905=>"111111111",
  3906=>"100001000",
  3907=>"011110100",
  3908=>"111111001",
  3909=>"010011110",
  3910=>"001101000",
  3911=>"100110101",
  3912=>"110011101",
  3913=>"011101011",
  3914=>"000111110",
  3915=>"000010001",
  3916=>"001111101",
  3917=>"101110000",
  3918=>"111110010",
  3919=>"000010000",
  3920=>"010011101",
  3921=>"001001101",
  3922=>"001110001",
  3923=>"011011111",
  3924=>"011011010",
  3925=>"010101101",
  3926=>"100011010",
  3927=>"010101010",
  3928=>"000000100",
  3929=>"010011010",
  3930=>"001111101",
  3931=>"000100111",
  3932=>"101001111",
  3933=>"001001010",
  3934=>"100001100",
  3935=>"000111100",
  3936=>"010010000",
  3937=>"000010101",
  3938=>"000100011",
  3939=>"010001101",
  3940=>"110000000",
  3941=>"001011001",
  3942=>"001111101",
  3943=>"110100001",
  3944=>"110001010",
  3945=>"100110111",
  3946=>"111000010",
  3947=>"101000001",
  3948=>"100100111",
  3949=>"111000101",
  3950=>"010111001",
  3951=>"101111110",
  3952=>"001111111",
  3953=>"010111101",
  3954=>"011111010",
  3955=>"011110111",
  3956=>"001101110",
  3957=>"110000111",
  3958=>"101100110",
  3959=>"101000001",
  3960=>"011010111",
  3961=>"000110111",
  3962=>"001000011",
  3963=>"001101010",
  3964=>"000010010",
  3965=>"111110000",
  3966=>"110011111",
  3967=>"111100000",
  3968=>"110001011",
  3969=>"011110110",
  3970=>"010110010",
  3971=>"111000001",
  3972=>"000110100",
  3973=>"110010011",
  3974=>"110010110",
  3975=>"111010111",
  3976=>"001100100",
  3977=>"001101000",
  3978=>"111011100",
  3979=>"110111011",
  3980=>"100101001",
  3981=>"001001001",
  3982=>"110111101",
  3983=>"100100000",
  3984=>"011110100",
  3985=>"100000111",
  3986=>"010000000",
  3987=>"101101100",
  3988=>"110110001",
  3989=>"010001000",
  3990=>"101110111",
  3991=>"011101000",
  3992=>"101000100",
  3993=>"100101100",
  3994=>"000110001",
  3995=>"101001110",
  3996=>"101001100",
  3997=>"011011110",
  3998=>"111010010",
  3999=>"001100100",
  4000=>"010110110",
  4001=>"111110001",
  4002=>"001110111",
  4003=>"101001011",
  4004=>"011000011",
  4005=>"011000010",
  4006=>"001100101",
  4007=>"010101010",
  4008=>"000100110",
  4009=>"110101111",
  4010=>"100110100",
  4011=>"100111110",
  4012=>"011101001",
  4013=>"101111000",
  4014=>"010011100",
  4015=>"001000001",
  4016=>"000010110",
  4017=>"111110101",
  4018=>"000010101",
  4019=>"001011010",
  4020=>"100110011",
  4021=>"100011110",
  4022=>"110011011",
  4023=>"110011000",
  4024=>"100111100",
  4025=>"000101110",
  4026=>"101001000",
  4027=>"101010000",
  4028=>"111001010",
  4029=>"110101111",
  4030=>"000100011",
  4031=>"010001110",
  4032=>"011111111",
  4033=>"000001111",
  4034=>"100101111",
  4035=>"111011011",
  4036=>"000001100",
  4037=>"110010101",
  4038=>"100011111",
  4039=>"000100000",
  4040=>"111100011",
  4041=>"000111010",
  4042=>"001110010",
  4043=>"011110000",
  4044=>"001010011",
  4045=>"001001101",
  4046=>"000011000",
  4047=>"101000010",
  4048=>"000100010",
  4049=>"000111101",
  4050=>"101000001",
  4051=>"100110011",
  4052=>"010001111",
  4053=>"110000100",
  4054=>"000100011",
  4055=>"010000010",
  4056=>"010101010",
  4057=>"011110100",
  4058=>"000010010",
  4059=>"100101100",
  4060=>"111101110",
  4061=>"001000110",
  4062=>"000111110",
  4063=>"000100100",
  4064=>"000101111",
  4065=>"111111100",
  4066=>"000011110",
  4067=>"011101101",
  4068=>"011000001",
  4069=>"010111100",
  4070=>"101101010",
  4071=>"110011111",
  4072=>"001110101",
  4073=>"010000011",
  4074=>"111100100",
  4075=>"100000011",
  4076=>"011011111",
  4077=>"011111100",
  4078=>"000101101",
  4079=>"111111100",
  4080=>"010011011",
  4081=>"110010101",
  4082=>"000000110",
  4083=>"010110100",
  4084=>"101000000",
  4085=>"111001000",
  4086=>"101011110",
  4087=>"011010001",
  4088=>"111101100",
  4089=>"100100101",
  4090=>"011110110",
  4091=>"110011001",
  4092=>"100111011",
  4093=>"101110001",
  4094=>"010100111",
  4095=>"110100100",
  4096=>"111111101",
  4097=>"111110111",
  4098=>"010101110",
  4099=>"010010100",
  4100=>"101100010",
  4101=>"001000001",
  4102=>"001000100",
  4103=>"000100001",
  4104=>"011001111",
  4105=>"011000010",
  4106=>"001000110",
  4107=>"010010000",
  4108=>"010111111",
  4109=>"110011000",
  4110=>"101101111",
  4111=>"001001101",
  4112=>"011010000",
  4113=>"010001110",
  4114=>"111111000",
  4115=>"000100010",
  4116=>"000100001",
  4117=>"100110000",
  4118=>"010010001",
  4119=>"110100010",
  4120=>"101111100",
  4121=>"001001111",
  4122=>"101011110",
  4123=>"001100011",
  4124=>"111011000",
  4125=>"000100100",
  4126=>"100010000",
  4127=>"110011011",
  4128=>"000011100",
  4129=>"101001010",
  4130=>"001110101",
  4131=>"100001110",
  4132=>"000100000",
  4133=>"101010111",
  4134=>"110000001",
  4135=>"111011100",
  4136=>"011011011",
  4137=>"000010101",
  4138=>"111111010",
  4139=>"001000111",
  4140=>"010011001",
  4141=>"011001001",
  4142=>"100011001",
  4143=>"110101011",
  4144=>"100111110",
  4145=>"010110001",
  4146=>"011111110",
  4147=>"010010001",
  4148=>"000010110",
  4149=>"101110011",
  4150=>"010101101",
  4151=>"111110000",
  4152=>"110100000",
  4153=>"000011001",
  4154=>"000100110",
  4155=>"000111110",
  4156=>"011101001",
  4157=>"110110110",
  4158=>"000000000",
  4159=>"001001001",
  4160=>"001010011",
  4161=>"000000010",
  4162=>"100010111",
  4163=>"111011001",
  4164=>"001011110",
  4165=>"000000100",
  4166=>"110111011",
  4167=>"001000010",
  4168=>"000011011",
  4169=>"100011110",
  4170=>"000011000",
  4171=>"001100001",
  4172=>"011101111",
  4173=>"100011110",
  4174=>"110101111",
  4175=>"110100000",
  4176=>"010111000",
  4177=>"010000011",
  4178=>"110110001",
  4179=>"111100001",
  4180=>"011101000",
  4181=>"111100000",
  4182=>"010000100",
  4183=>"010011111",
  4184=>"111100100",
  4185=>"011011100",
  4186=>"000101001",
  4187=>"001111110",
  4188=>"111011001",
  4189=>"010101110",
  4190=>"100101001",
  4191=>"010011001",
  4192=>"011001000",
  4193=>"101010101",
  4194=>"011111010",
  4195=>"100010111",
  4196=>"010010010",
  4197=>"001100000",
  4198=>"101000110",
  4199=>"011101000",
  4200=>"100111110",
  4201=>"110111111",
  4202=>"010011111",
  4203=>"110011101",
  4204=>"011011111",
  4205=>"011110110",
  4206=>"110100101",
  4207=>"111111101",
  4208=>"100111111",
  4209=>"110101010",
  4210=>"011111111",
  4211=>"100101111",
  4212=>"000011110",
  4213=>"110101100",
  4214=>"101101111",
  4215=>"110111000",
  4216=>"010000000",
  4217=>"001111011",
  4218=>"100000000",
  4219=>"100000010",
  4220=>"011111001",
  4221=>"010000111",
  4222=>"111111001",
  4223=>"010111000",
  4224=>"110010110",
  4225=>"101101111",
  4226=>"011110010",
  4227=>"110101001",
  4228=>"011100000",
  4229=>"011001001",
  4230=>"000010100",
  4231=>"101111000",
  4232=>"011101101",
  4233=>"001010001",
  4234=>"000001010",
  4235=>"011001011",
  4236=>"000001011",
  4237=>"010011101",
  4238=>"110010101",
  4239=>"100000101",
  4240=>"010010011",
  4241=>"111011111",
  4242=>"010001111",
  4243=>"001110001",
  4244=>"000110101",
  4245=>"110011101",
  4246=>"011110100",
  4247=>"010110110",
  4248=>"101001011",
  4249=>"000000100",
  4250=>"010011000",
  4251=>"100011111",
  4252=>"100010010",
  4253=>"111111011",
  4254=>"000100001",
  4255=>"101000101",
  4256=>"100100001",
  4257=>"101110110",
  4258=>"111110010",
  4259=>"000100011",
  4260=>"001100111",
  4261=>"100001100",
  4262=>"011010000",
  4263=>"000100001",
  4264=>"001110010",
  4265=>"111100110",
  4266=>"110011100",
  4267=>"111101001",
  4268=>"100100110",
  4269=>"000001101",
  4270=>"011011101",
  4271=>"010100000",
  4272=>"100000000",
  4273=>"001000110",
  4274=>"001011001",
  4275=>"110000001",
  4276=>"110001100",
  4277=>"000010100",
  4278=>"000000110",
  4279=>"111010110",
  4280=>"111010111",
  4281=>"001010111",
  4282=>"000000011",
  4283=>"110010000",
  4284=>"001010010",
  4285=>"011110000",
  4286=>"010101010",
  4287=>"010101001",
  4288=>"100010010",
  4289=>"011110111",
  4290=>"110110000",
  4291=>"010101010",
  4292=>"111111011",
  4293=>"000100000",
  4294=>"011010111",
  4295=>"000111111",
  4296=>"011000001",
  4297=>"010111100",
  4298=>"100010001",
  4299=>"101110011",
  4300=>"101010011",
  4301=>"101111111",
  4302=>"100101110",
  4303=>"111101000",
  4304=>"110000110",
  4305=>"010000000",
  4306=>"111111110",
  4307=>"001010001",
  4308=>"110001000",
  4309=>"000010111",
  4310=>"011101010",
  4311=>"011100000",
  4312=>"100010000",
  4313=>"101000011",
  4314=>"110100010",
  4315=>"111010010",
  4316=>"101111110",
  4317=>"011101101",
  4318=>"110110110",
  4319=>"101000010",
  4320=>"011000010",
  4321=>"000010111",
  4322=>"000101001",
  4323=>"100110110",
  4324=>"100111110",
  4325=>"111100111",
  4326=>"001111010",
  4327=>"000110111",
  4328=>"000110100",
  4329=>"001000000",
  4330=>"001010000",
  4331=>"111000111",
  4332=>"110010101",
  4333=>"010011010",
  4334=>"101111001",
  4335=>"010011111",
  4336=>"011000000",
  4337=>"100001000",
  4338=>"111001000",
  4339=>"100010110",
  4340=>"101000100",
  4341=>"011111101",
  4342=>"010001000",
  4343=>"110010111",
  4344=>"000111111",
  4345=>"001010111",
  4346=>"010101111",
  4347=>"100001000",
  4348=>"001111011",
  4349=>"111101110",
  4350=>"101000001",
  4351=>"001010110",
  4352=>"100001111",
  4353=>"101110110",
  4354=>"101111110",
  4355=>"000110110",
  4356=>"111100101",
  4357=>"010010000",
  4358=>"101000011",
  4359=>"011100000",
  4360=>"001001100",
  4361=>"111101000",
  4362=>"010011100",
  4363=>"110000100",
  4364=>"001011000",
  4365=>"011010110",
  4366=>"011010110",
  4367=>"111100011",
  4368=>"000001101",
  4369=>"011000111",
  4370=>"011011011",
  4371=>"011101000",
  4372=>"101001111",
  4373=>"001010010",
  4374=>"011001001",
  4375=>"000100011",
  4376=>"110101001",
  4377=>"000000000",
  4378=>"010101000",
  4379=>"010000010",
  4380=>"000100110",
  4381=>"100100101",
  4382=>"101010110",
  4383=>"100111100",
  4384=>"111010100",
  4385=>"101111101",
  4386=>"010101101",
  4387=>"110100101",
  4388=>"111001111",
  4389=>"101110111",
  4390=>"111111100",
  4391=>"110010010",
  4392=>"110001011",
  4393=>"110000000",
  4394=>"101101011",
  4395=>"111110000",
  4396=>"101111001",
  4397=>"001010010",
  4398=>"000101000",
  4399=>"010010000",
  4400=>"011101101",
  4401=>"111001000",
  4402=>"001110000",
  4403=>"111110110",
  4404=>"000100000",
  4405=>"000100111",
  4406=>"110000101",
  4407=>"111111110",
  4408=>"000011000",
  4409=>"001001001",
  4410=>"011000101",
  4411=>"111111001",
  4412=>"101000110",
  4413=>"001011101",
  4414=>"001100101",
  4415=>"111000101",
  4416=>"100010010",
  4417=>"011111110",
  4418=>"000110111",
  4419=>"110000100",
  4420=>"011010010",
  4421=>"010010010",
  4422=>"110111100",
  4423=>"111111000",
  4424=>"100000000",
  4425=>"010111101",
  4426=>"100100000",
  4427=>"111101000",
  4428=>"101110000",
  4429=>"000110101",
  4430=>"101000110",
  4431=>"001011010",
  4432=>"111110011",
  4433=>"001000101",
  4434=>"000110000",
  4435=>"011101110",
  4436=>"101000010",
  4437=>"111011101",
  4438=>"110111101",
  4439=>"011001110",
  4440=>"101100111",
  4441=>"110011011",
  4442=>"101111100",
  4443=>"110110111",
  4444=>"001011000",
  4445=>"001100101",
  4446=>"010100001",
  4447=>"000001100",
  4448=>"000011000",
  4449=>"100111110",
  4450=>"111001101",
  4451=>"001000010",
  4452=>"101111101",
  4453=>"100110000",
  4454=>"100000000",
  4455=>"100000110",
  4456=>"110001101",
  4457=>"110001000",
  4458=>"011011011",
  4459=>"111011010",
  4460=>"110010110",
  4461=>"110010001",
  4462=>"011111011",
  4463=>"001001100",
  4464=>"000000110",
  4465=>"100101010",
  4466=>"100110110",
  4467=>"101100111",
  4468=>"001011001",
  4469=>"111010111",
  4470=>"101010001",
  4471=>"000001000",
  4472=>"100001011",
  4473=>"101010001",
  4474=>"100011001",
  4475=>"000101110",
  4476=>"001100110",
  4477=>"100100110",
  4478=>"000011011",
  4479=>"010101000",
  4480=>"110100101",
  4481=>"000111001",
  4482=>"111110000",
  4483=>"111100111",
  4484=>"110100010",
  4485=>"010111000",
  4486=>"000111011",
  4487=>"000100100",
  4488=>"000000011",
  4489=>"101000100",
  4490=>"001000101",
  4491=>"101001010",
  4492=>"111010100",
  4493=>"000011010",
  4494=>"011101100",
  4495=>"101111111",
  4496=>"111010101",
  4497=>"000100000",
  4498=>"100111101",
  4499=>"000110101",
  4500=>"100110011",
  4501=>"000010110",
  4502=>"100010111",
  4503=>"001001101",
  4504=>"001000100",
  4505=>"110000010",
  4506=>"101011101",
  4507=>"100101001",
  4508=>"110011110",
  4509=>"000101100",
  4510=>"001011011",
  4511=>"000101110",
  4512=>"100100000",
  4513=>"000111011",
  4514=>"000000010",
  4515=>"011111011",
  4516=>"100100000",
  4517=>"101010110",
  4518=>"101010110",
  4519=>"111110111",
  4520=>"000010011",
  4521=>"011110111",
  4522=>"010011000",
  4523=>"001011001",
  4524=>"001010001",
  4525=>"101000001",
  4526=>"100011110",
  4527=>"110001100",
  4528=>"011000101",
  4529=>"100000101",
  4530=>"000011101",
  4531=>"001101110",
  4532=>"010011001",
  4533=>"001010111",
  4534=>"010110110",
  4535=>"101111000",
  4536=>"101101100",
  4537=>"111000110",
  4538=>"111111111",
  4539=>"011111000",
  4540=>"011100010",
  4541=>"010001010",
  4542=>"110010011",
  4543=>"110111000",
  4544=>"100111011",
  4545=>"010010000",
  4546=>"101100111",
  4547=>"101000011",
  4548=>"111101000",
  4549=>"010110000",
  4550=>"000000001",
  4551=>"001000000",
  4552=>"100110001",
  4553=>"100111101",
  4554=>"000110000",
  4555=>"011101100",
  4556=>"111101110",
  4557=>"111010110",
  4558=>"000000100",
  4559=>"101100010",
  4560=>"110001111",
  4561=>"100001010",
  4562=>"100110010",
  4563=>"111110110",
  4564=>"101010111",
  4565=>"110101111",
  4566=>"001111010",
  4567=>"010100110",
  4568=>"111001011",
  4569=>"011110110",
  4570=>"010001000",
  4571=>"100100010",
  4572=>"010001001",
  4573=>"011110110",
  4574=>"000110111",
  4575=>"000010000",
  4576=>"000001100",
  4577=>"010100100",
  4578=>"010101000",
  4579=>"010101010",
  4580=>"111111111",
  4581=>"011111011",
  4582=>"110101000",
  4583=>"000001001",
  4584=>"000011000",
  4585=>"110011000",
  4586=>"000100010",
  4587=>"011110010",
  4588=>"010100110",
  4589=>"101111100",
  4590=>"011011000",
  4591=>"010100011",
  4592=>"010101100",
  4593=>"011010001",
  4594=>"000100010",
  4595=>"000001000",
  4596=>"010001011",
  4597=>"000001001",
  4598=>"101001010",
  4599=>"101101111",
  4600=>"110100100",
  4601=>"011111111",
  4602=>"010100000",
  4603=>"100000010",
  4604=>"111010110",
  4605=>"111011010",
  4606=>"011101111",
  4607=>"110001111",
  4608=>"000011111",
  4609=>"010000111",
  4610=>"011011110",
  4611=>"000101101",
  4612=>"110000110",
  4613=>"000111100",
  4614=>"110111011",
  4615=>"000100100",
  4616=>"111000000",
  4617=>"101000100",
  4618=>"001000010",
  4619=>"011111101",
  4620=>"100000001",
  4621=>"011100111",
  4622=>"111110110",
  4623=>"010011001",
  4624=>"001011001",
  4625=>"100011110",
  4626=>"000110111",
  4627=>"110001100",
  4628=>"000010010",
  4629=>"001010001",
  4630=>"001010101",
  4631=>"001010111",
  4632=>"000110010",
  4633=>"101101111",
  4634=>"101000011",
  4635=>"010000011",
  4636=>"001001000",
  4637=>"011100100",
  4638=>"110100010",
  4639=>"010000111",
  4640=>"111011011",
  4641=>"001000110",
  4642=>"001001101",
  4643=>"100100100",
  4644=>"001110001",
  4645=>"101001111",
  4646=>"100110000",
  4647=>"001000111",
  4648=>"001111110",
  4649=>"001101001",
  4650=>"100000000",
  4651=>"010111110",
  4652=>"100101000",
  4653=>"000000001",
  4654=>"100001001",
  4655=>"000110111",
  4656=>"110101001",
  4657=>"111010100",
  4658=>"111010001",
  4659=>"101101011",
  4660=>"100011000",
  4661=>"111101101",
  4662=>"100100010",
  4663=>"100011000",
  4664=>"011100101",
  4665=>"011111111",
  4666=>"011101001",
  4667=>"110001101",
  4668=>"011001111",
  4669=>"000011010",
  4670=>"010110110",
  4671=>"111010001",
  4672=>"010100011",
  4673=>"010010010",
  4674=>"011101011",
  4675=>"101000101",
  4676=>"100100011",
  4677=>"111101011",
  4678=>"001000001",
  4679=>"100101110",
  4680=>"110101101",
  4681=>"111101110",
  4682=>"101001001",
  4683=>"100010010",
  4684=>"110010010",
  4685=>"100110000",
  4686=>"001011101",
  4687=>"010010011",
  4688=>"010010000",
  4689=>"101010111",
  4690=>"111110111",
  4691=>"001111010",
  4692=>"001100110",
  4693=>"001100010",
  4694=>"010010000",
  4695=>"111111011",
  4696=>"110111111",
  4697=>"100011001",
  4698=>"110110100",
  4699=>"001101110",
  4700=>"101010000",
  4701=>"000110011",
  4702=>"010000111",
  4703=>"000100000",
  4704=>"010100100",
  4705=>"100000100",
  4706=>"001111101",
  4707=>"010000110",
  4708=>"011011100",
  4709=>"011000110",
  4710=>"111010111",
  4711=>"100101010",
  4712=>"001000111",
  4713=>"011000110",
  4714=>"001111111",
  4715=>"110001000",
  4716=>"101000100",
  4717=>"001101010",
  4718=>"110110000",
  4719=>"101011101",
  4720=>"000000000",
  4721=>"000101101",
  4722=>"011100101",
  4723=>"000000011",
  4724=>"110010001",
  4725=>"000111100",
  4726=>"000001100",
  4727=>"011001001",
  4728=>"110101000",
  4729=>"010011000",
  4730=>"000000001",
  4731=>"110000110",
  4732=>"000110011",
  4733=>"010101111",
  4734=>"100001110",
  4735=>"111111000",
  4736=>"010110010",
  4737=>"011010001",
  4738=>"111110111",
  4739=>"001110010",
  4740=>"011101110",
  4741=>"100010000",
  4742=>"000010110",
  4743=>"011001100",
  4744=>"011110101",
  4745=>"000011100",
  4746=>"100100111",
  4747=>"011111101",
  4748=>"110101100",
  4749=>"111111011",
  4750=>"010001111",
  4751=>"101101111",
  4752=>"011111011",
  4753=>"101001100",
  4754=>"000101010",
  4755=>"011110001",
  4756=>"100000110",
  4757=>"000001100",
  4758=>"011111011",
  4759=>"001010111",
  4760=>"011001111",
  4761=>"000011101",
  4762=>"000110011",
  4763=>"110010001",
  4764=>"010001101",
  4765=>"111011000",
  4766=>"110011101",
  4767=>"101001110",
  4768=>"110111101",
  4769=>"000110111",
  4770=>"010101000",
  4771=>"111010010",
  4772=>"010001010",
  4773=>"101111101",
  4774=>"100100100",
  4775=>"110101000",
  4776=>"101001100",
  4777=>"011000000",
  4778=>"101001001",
  4779=>"100101101",
  4780=>"110001110",
  4781=>"101011011",
  4782=>"010110010",
  4783=>"011101100",
  4784=>"111110000",
  4785=>"001001001",
  4786=>"101000100",
  4787=>"101111110",
  4788=>"100101110",
  4789=>"101010111",
  4790=>"010100010",
  4791=>"100110111",
  4792=>"100011110",
  4793=>"110011101",
  4794=>"010000010",
  4795=>"111001010",
  4796=>"110111001",
  4797=>"110011100",
  4798=>"110011011",
  4799=>"111100001",
  4800=>"001110000",
  4801=>"111011010",
  4802=>"000111011",
  4803=>"011110011",
  4804=>"110011110",
  4805=>"000001110",
  4806=>"000000000",
  4807=>"110011011",
  4808=>"011101111",
  4809=>"111011000",
  4810=>"101111110",
  4811=>"110011101",
  4812=>"000010101",
  4813=>"110000111",
  4814=>"011100110",
  4815=>"001000001",
  4816=>"100011111",
  4817=>"101110001",
  4818=>"100110110",
  4819=>"111101111",
  4820=>"001110101",
  4821=>"100100001",
  4822=>"011000010",
  4823=>"100101000",
  4824=>"101001011",
  4825=>"110101100",
  4826=>"110111010",
  4827=>"001110000",
  4828=>"110101111",
  4829=>"100000011",
  4830=>"000000110",
  4831=>"010100100",
  4832=>"110110111",
  4833=>"111101001",
  4834=>"111011100",
  4835=>"100110111",
  4836=>"010110100",
  4837=>"111101000",
  4838=>"111011111",
  4839=>"100101111",
  4840=>"001011001",
  4841=>"000000101",
  4842=>"110010101",
  4843=>"100001000",
  4844=>"100101110",
  4845=>"010100011",
  4846=>"101110010",
  4847=>"111010110",
  4848=>"110111000",
  4849=>"111000001",
  4850=>"100001001",
  4851=>"111011010",
  4852=>"000111101",
  4853=>"111101000",
  4854=>"000010000",
  4855=>"001111111",
  4856=>"101011101",
  4857=>"100111000",
  4858=>"010110010",
  4859=>"101011011",
  4860=>"010101001",
  4861=>"100001111",
  4862=>"010010101",
  4863=>"111111011",
  4864=>"101000100",
  4865=>"110010000",
  4866=>"101100110",
  4867=>"011110100",
  4868=>"101000000",
  4869=>"010000100",
  4870=>"001001010",
  4871=>"001101110",
  4872=>"001000101",
  4873=>"101100110",
  4874=>"100011101",
  4875=>"111011101",
  4876=>"111011000",
  4877=>"000110110",
  4878=>"011011110",
  4879=>"000000101",
  4880=>"011001000",
  4881=>"000010111",
  4882=>"011111010",
  4883=>"000000110",
  4884=>"001110011",
  4885=>"111110000",
  4886=>"000010111",
  4887=>"100011111",
  4888=>"001101101",
  4889=>"100101110",
  4890=>"000101101",
  4891=>"011001110",
  4892=>"111101110",
  4893=>"011110110",
  4894=>"000010100",
  4895=>"110100110",
  4896=>"100011111",
  4897=>"011000010",
  4898=>"010111011",
  4899=>"000001001",
  4900=>"000000101",
  4901=>"010001000",
  4902=>"101101011",
  4903=>"000110000",
  4904=>"111101101",
  4905=>"101101011",
  4906=>"001011000",
  4907=>"000010000",
  4908=>"001101011",
  4909=>"111111111",
  4910=>"001110011",
  4911=>"101011111",
  4912=>"011001010",
  4913=>"000100101",
  4914=>"101111000",
  4915=>"111101011",
  4916=>"010000000",
  4917=>"000101001",
  4918=>"101100111",
  4919=>"111011001",
  4920=>"101010001",
  4921=>"011101101",
  4922=>"001000100",
  4923=>"011000100",
  4924=>"000001100",
  4925=>"110101001",
  4926=>"110011110",
  4927=>"111000000",
  4928=>"001111111",
  4929=>"101010000",
  4930=>"000011000",
  4931=>"010101010",
  4932=>"100010111",
  4933=>"000110110",
  4934=>"101100000",
  4935=>"100100111",
  4936=>"111000101",
  4937=>"111111101",
  4938=>"101000010",
  4939=>"100111000",
  4940=>"110010011",
  4941=>"101010001",
  4942=>"000100010",
  4943=>"000000010",
  4944=>"101101001",
  4945=>"110000101",
  4946=>"001110110",
  4947=>"001000010",
  4948=>"111111101",
  4949=>"010001111",
  4950=>"111010010",
  4951=>"011011010",
  4952=>"000010010",
  4953=>"111100100",
  4954=>"011011101",
  4955=>"010000100",
  4956=>"100001100",
  4957=>"011000000",
  4958=>"111011100",
  4959=>"111010010",
  4960=>"111010101",
  4961=>"100011111",
  4962=>"000100000",
  4963=>"111101000",
  4964=>"110011111",
  4965=>"010111001",
  4966=>"101010000",
  4967=>"110100011",
  4968=>"101010100",
  4969=>"110011110",
  4970=>"001011110",
  4971=>"110101010",
  4972=>"111100000",
  4973=>"110111110",
  4974=>"101110001",
  4975=>"111110000",
  4976=>"110010101",
  4977=>"110110000",
  4978=>"001000000",
  4979=>"100101111",
  4980=>"101111111",
  4981=>"100001101",
  4982=>"111010001",
  4983=>"010110100",
  4984=>"100111000",
  4985=>"111111010",
  4986=>"010010010",
  4987=>"111110011",
  4988=>"111001100",
  4989=>"111110000",
  4990=>"000110011",
  4991=>"001011000",
  4992=>"100100000",
  4993=>"010001011",
  4994=>"000010110",
  4995=>"001101101",
  4996=>"111101111",
  4997=>"111111111",
  4998=>"000100001",
  4999=>"100010000",
  5000=>"111010001",
  5001=>"101100010",
  5002=>"101111101",
  5003=>"100001100",
  5004=>"010010100",
  5005=>"010000110",
  5006=>"111101110",
  5007=>"001011010",
  5008=>"110010110",
  5009=>"100011101",
  5010=>"110000100",
  5011=>"110100010",
  5012=>"011111101",
  5013=>"010011001",
  5014=>"010111010",
  5015=>"001110000",
  5016=>"000000011",
  5017=>"011001011",
  5018=>"000100010",
  5019=>"111001110",
  5020=>"011011110",
  5021=>"110011111",
  5022=>"110010010",
  5023=>"001010111",
  5024=>"011000100",
  5025=>"111011010",
  5026=>"000110110",
  5027=>"000100000",
  5028=>"111001101",
  5029=>"111010111",
  5030=>"010010111",
  5031=>"110011010",
  5032=>"000100111",
  5033=>"000101100",
  5034=>"010111001",
  5035=>"000001000",
  5036=>"011101001",
  5037=>"100001101",
  5038=>"001010101",
  5039=>"001101001",
  5040=>"111000000",
  5041=>"001110010",
  5042=>"100010001",
  5043=>"111100100",
  5044=>"111011110",
  5045=>"011010110",
  5046=>"110110001",
  5047=>"100111000",
  5048=>"001000000",
  5049=>"011011100",
  5050=>"110010001",
  5051=>"101011011",
  5052=>"110110100",
  5053=>"111000000",
  5054=>"101100111",
  5055=>"010101000",
  5056=>"101010111",
  5057=>"101110010",
  5058=>"101001000",
  5059=>"110001110",
  5060=>"000110111",
  5061=>"110011110",
  5062=>"110010111",
  5063=>"010110010",
  5064=>"010100011",
  5065=>"101101001",
  5066=>"111000000",
  5067=>"000111110",
  5068=>"000111111",
  5069=>"111101000",
  5070=>"011001000",
  5071=>"100000000",
  5072=>"111110111",
  5073=>"000100011",
  5074=>"100011111",
  5075=>"000001000",
  5076=>"000011010",
  5077=>"001110110",
  5078=>"111110110",
  5079=>"101010111",
  5080=>"100111000",
  5081=>"100100000",
  5082=>"101000001",
  5083=>"011101010",
  5084=>"000100111",
  5085=>"111111011",
  5086=>"000001111",
  5087=>"100101001",
  5088=>"001100010",
  5089=>"010000000",
  5090=>"010000111",
  5091=>"111001011",
  5092=>"000100110",
  5093=>"001101011",
  5094=>"011001101",
  5095=>"101101010",
  5096=>"011000100",
  5097=>"110100000",
  5098=>"101011111",
  5099=>"001001111",
  5100=>"111000010",
  5101=>"001111101",
  5102=>"000111001",
  5103=>"010001100",
  5104=>"011001000",
  5105=>"001001110",
  5106=>"000000011",
  5107=>"001011001",
  5108=>"001110101",
  5109=>"010100001",
  5110=>"000011011",
  5111=>"111011011",
  5112=>"100111110",
  5113=>"001111011",
  5114=>"011100010",
  5115=>"001010000",
  5116=>"101001111",
  5117=>"110011000",
  5118=>"111101111",
  5119=>"010010000",
  5120=>"111001011",
  5121=>"001001011",
  5122=>"110010110",
  5123=>"110010001",
  5124=>"010111101",
  5125=>"100000110",
  5126=>"010010011",
  5127=>"100000000",
  5128=>"010101011",
  5129=>"110110001",
  5130=>"011001001",
  5131=>"101100101",
  5132=>"010100000",
  5133=>"010111011",
  5134=>"001110101",
  5135=>"100000100",
  5136=>"100111010",
  5137=>"100101001",
  5138=>"110110111",
  5139=>"000001111",
  5140=>"010011100",
  5141=>"000110101",
  5142=>"011010000",
  5143=>"010110111",
  5144=>"011101001",
  5145=>"000001010",
  5146=>"001001011",
  5147=>"110000010",
  5148=>"011101111",
  5149=>"111011101",
  5150=>"101010100",
  5151=>"000000010",
  5152=>"110111011",
  5153=>"100111000",
  5154=>"111111001",
  5155=>"001011010",
  5156=>"011001111",
  5157=>"001000100",
  5158=>"111000010",
  5159=>"111100011",
  5160=>"001111100",
  5161=>"000110010",
  5162=>"011011110",
  5163=>"011110111",
  5164=>"111111100",
  5165=>"110000001",
  5166=>"100011011",
  5167=>"011111101",
  5168=>"001101011",
  5169=>"010001010",
  5170=>"011100000",
  5171=>"010101101",
  5172=>"000000001",
  5173=>"010000000",
  5174=>"001110001",
  5175=>"111100010",
  5176=>"010000000",
  5177=>"110101101",
  5178=>"000000111",
  5179=>"000110110",
  5180=>"101110000",
  5181=>"101111111",
  5182=>"111001100",
  5183=>"111001101",
  5184=>"000110011",
  5185=>"000001110",
  5186=>"100101110",
  5187=>"101100110",
  5188=>"001001101",
  5189=>"000111010",
  5190=>"111100000",
  5191=>"000001111",
  5192=>"000011111",
  5193=>"111010101",
  5194=>"001001110",
  5195=>"011000111",
  5196=>"001100001",
  5197=>"001001111",
  5198=>"101110111",
  5199=>"111101001",
  5200=>"011100100",
  5201=>"111110001",
  5202=>"111001101",
  5203=>"001001000",
  5204=>"011000001",
  5205=>"011001011",
  5206=>"101110100",
  5207=>"001011011",
  5208=>"100011000",
  5209=>"101100011",
  5210=>"111010101",
  5211=>"101011101",
  5212=>"111100110",
  5213=>"000001001",
  5214=>"001010100",
  5215=>"010111100",
  5216=>"000100000",
  5217=>"011101101",
  5218=>"111101111",
  5219=>"010010000",
  5220=>"010111000",
  5221=>"111011011",
  5222=>"100000111",
  5223=>"100001001",
  5224=>"010000011",
  5225=>"111111111",
  5226=>"101100111",
  5227=>"111001110",
  5228=>"111101010",
  5229=>"100100010",
  5230=>"001001111",
  5231=>"110101110",
  5232=>"001110110",
  5233=>"000001011",
  5234=>"011100010",
  5235=>"010011100",
  5236=>"110010001",
  5237=>"110111010",
  5238=>"111101001",
  5239=>"000010001",
  5240=>"101011010",
  5241=>"001111001",
  5242=>"010000000",
  5243=>"010110010",
  5244=>"101111101",
  5245=>"101100111",
  5246=>"110011001",
  5247=>"101101101",
  5248=>"110010100",
  5249=>"100111111",
  5250=>"101010110",
  5251=>"010000011",
  5252=>"110000010",
  5253=>"010100101",
  5254=>"010101110",
  5255=>"010111011",
  5256=>"011011011",
  5257=>"000010001",
  5258=>"000001000",
  5259=>"001110100",
  5260=>"011100011",
  5261=>"010011000",
  5262=>"010000010",
  5263=>"100011010",
  5264=>"010100011",
  5265=>"110100110",
  5266=>"000001110",
  5267=>"001111010",
  5268=>"011101001",
  5269=>"011000010",
  5270=>"111001010",
  5271=>"111011110",
  5272=>"110010000",
  5273=>"011100011",
  5274=>"110100111",
  5275=>"000100000",
  5276=>"010101110",
  5277=>"011110111",
  5278=>"100101001",
  5279=>"000010000",
  5280=>"000000101",
  5281=>"001100111",
  5282=>"101001111",
  5283=>"010110010",
  5284=>"011011101",
  5285=>"101011101",
  5286=>"101010011",
  5287=>"111101100",
  5288=>"111011101",
  5289=>"101001001",
  5290=>"010000000",
  5291=>"000100000",
  5292=>"000111111",
  5293=>"100111101",
  5294=>"011001111",
  5295=>"110110010",
  5296=>"000100010",
  5297=>"100100001",
  5298=>"001101001",
  5299=>"100110110",
  5300=>"011010111",
  5301=>"111111010",
  5302=>"110001001",
  5303=>"000100100",
  5304=>"111110001",
  5305=>"000000010",
  5306=>"010011111",
  5307=>"001111010",
  5308=>"000001100",
  5309=>"001101010",
  5310=>"000010001",
  5311=>"111101001",
  5312=>"001011000",
  5313=>"101010000",
  5314=>"101111011",
  5315=>"111110000",
  5316=>"001010001",
  5317=>"110000011",
  5318=>"000010010",
  5319=>"000000110",
  5320=>"011010011",
  5321=>"000011011",
  5322=>"000111011",
  5323=>"010110011",
  5324=>"111001101",
  5325=>"011101000",
  5326=>"100111001",
  5327=>"101001001",
  5328=>"000101000",
  5329=>"000000011",
  5330=>"010101000",
  5331=>"011101010",
  5332=>"100101010",
  5333=>"001001100",
  5334=>"001101101",
  5335=>"101100010",
  5336=>"000011000",
  5337=>"101001101",
  5338=>"101010000",
  5339=>"010000000",
  5340=>"111111010",
  5341=>"110100110",
  5342=>"101000001",
  5343=>"111001100",
  5344=>"101000101",
  5345=>"010010001",
  5346=>"010110110",
  5347=>"000001000",
  5348=>"100000100",
  5349=>"000101010",
  5350=>"010110100",
  5351=>"111000111",
  5352=>"101011010",
  5353=>"100011011",
  5354=>"110111111",
  5355=>"100000000",
  5356=>"010010101",
  5357=>"001000000",
  5358=>"010010111",
  5359=>"010000000",
  5360=>"010101100",
  5361=>"010000110",
  5362=>"101001101",
  5363=>"100011110",
  5364=>"011001111",
  5365=>"110111111",
  5366=>"111110111",
  5367=>"101001110",
  5368=>"111001110",
  5369=>"010101101",
  5370=>"101001001",
  5371=>"010000100",
  5372=>"001000100",
  5373=>"111111011",
  5374=>"011001100",
  5375=>"101011100",
  5376=>"100000110",
  5377=>"011000010",
  5378=>"011000000",
  5379=>"000011111",
  5380=>"110000100",
  5381=>"011111100",
  5382=>"100111010",
  5383=>"011110010",
  5384=>"101100001",
  5385=>"010011110",
  5386=>"100001110",
  5387=>"101111010",
  5388=>"110010001",
  5389=>"000010010",
  5390=>"100100000",
  5391=>"001000110",
  5392=>"101100000",
  5393=>"000001001",
  5394=>"010111011",
  5395=>"111010101",
  5396=>"001010101",
  5397=>"110111101",
  5398=>"000001100",
  5399=>"100001011",
  5400=>"111000100",
  5401=>"111110011",
  5402=>"010001110",
  5403=>"000111001",
  5404=>"000001011",
  5405=>"101001110",
  5406=>"111101101",
  5407=>"111110100",
  5408=>"111110000",
  5409=>"100101101",
  5410=>"101000011",
  5411=>"001000011",
  5412=>"110110101",
  5413=>"110000110",
  5414=>"011100111",
  5415=>"000110011",
  5416=>"011001000",
  5417=>"000111100",
  5418=>"001100100",
  5419=>"101000000",
  5420=>"111000010",
  5421=>"010110001",
  5422=>"101100111",
  5423=>"110010000",
  5424=>"001110000",
  5425=>"111111001",
  5426=>"110110100",
  5427=>"110111100",
  5428=>"001000110",
  5429=>"001011000",
  5430=>"100111110",
  5431=>"011110000",
  5432=>"010000100",
  5433=>"010100000",
  5434=>"111101001",
  5435=>"110110010",
  5436=>"010000100",
  5437=>"000000010",
  5438=>"001110111",
  5439=>"000000111",
  5440=>"111010001",
  5441=>"010011100",
  5442=>"100000000",
  5443=>"100101101",
  5444=>"011111010",
  5445=>"000100011",
  5446=>"100101011",
  5447=>"110011000",
  5448=>"001011101",
  5449=>"001111111",
  5450=>"101010111",
  5451=>"000001100",
  5452=>"101100010",
  5453=>"010100000",
  5454=>"101111110",
  5455=>"111001101",
  5456=>"001000111",
  5457=>"011001010",
  5458=>"101101100",
  5459=>"000101110",
  5460=>"000101010",
  5461=>"001000010",
  5462=>"100001001",
  5463=>"001001100",
  5464=>"000110101",
  5465=>"100001100",
  5466=>"111111000",
  5467=>"110001010",
  5468=>"100011000",
  5469=>"011101011",
  5470=>"111010001",
  5471=>"100000101",
  5472=>"101001110",
  5473=>"101001101",
  5474=>"011110110",
  5475=>"001100101",
  5476=>"000111011",
  5477=>"011000000",
  5478=>"001100001",
  5479=>"011110001",
  5480=>"011101100",
  5481=>"000110101",
  5482=>"000100111",
  5483=>"001001101",
  5484=>"110101101",
  5485=>"001000101",
  5486=>"000100100",
  5487=>"101110001",
  5488=>"100000010",
  5489=>"110111111",
  5490=>"010101111",
  5491=>"010111000",
  5492=>"000001010",
  5493=>"011000000",
  5494=>"010111010",
  5495=>"110101100",
  5496=>"111111101",
  5497=>"000111101",
  5498=>"001101111",
  5499=>"111110100",
  5500=>"100001110",
  5501=>"111110110",
  5502=>"001001000",
  5503=>"100010000",
  5504=>"000010000",
  5505=>"011000000",
  5506=>"111101001",
  5507=>"110010101",
  5508=>"000110110",
  5509=>"000101110",
  5510=>"000000011",
  5511=>"000011101",
  5512=>"110110000",
  5513=>"100111010",
  5514=>"000010111",
  5515=>"111011111",
  5516=>"110010001",
  5517=>"000001110",
  5518=>"110010010",
  5519=>"111100101",
  5520=>"100001011",
  5521=>"000111001",
  5522=>"111110000",
  5523=>"010111000",
  5524=>"100110110",
  5525=>"111100001",
  5526=>"000000000",
  5527=>"100000100",
  5528=>"010110001",
  5529=>"011100011",
  5530=>"010011001",
  5531=>"111111000",
  5532=>"001100101",
  5533=>"110010010",
  5534=>"101110110",
  5535=>"100011100",
  5536=>"010000011",
  5537=>"001101001",
  5538=>"110101001",
  5539=>"000110010",
  5540=>"000001111",
  5541=>"111101000",
  5542=>"101110101",
  5543=>"111011110",
  5544=>"010011000",
  5545=>"100001101",
  5546=>"011010100",
  5547=>"011101100",
  5548=>"101000101",
  5549=>"101001001",
  5550=>"001111111",
  5551=>"000100111",
  5552=>"111100111",
  5553=>"110001011",
  5554=>"000111000",
  5555=>"000101110",
  5556=>"111100111",
  5557=>"100000001",
  5558=>"100010010",
  5559=>"000001000",
  5560=>"101010111",
  5561=>"111110110",
  5562=>"000000110",
  5563=>"010000001",
  5564=>"001110110",
  5565=>"000010011",
  5566=>"000000110",
  5567=>"011000100",
  5568=>"101001010",
  5569=>"010010101",
  5570=>"100000000",
  5571=>"001001101",
  5572=>"101111101",
  5573=>"010000111",
  5574=>"110010111",
  5575=>"010001100",
  5576=>"111010111",
  5577=>"110101101",
  5578=>"111000111",
  5579=>"000111001",
  5580=>"110111110",
  5581=>"100000111",
  5582=>"001000000",
  5583=>"100010000",
  5584=>"111100010",
  5585=>"011011110",
  5586=>"000111010",
  5587=>"000011111",
  5588=>"010100001",
  5589=>"001101010",
  5590=>"000000001",
  5591=>"011000100",
  5592=>"000000011",
  5593=>"111111000",
  5594=>"000000100",
  5595=>"100010100",
  5596=>"000101111",
  5597=>"110110111",
  5598=>"100000000",
  5599=>"100000001",
  5600=>"001010010",
  5601=>"100101110",
  5602=>"001111111",
  5603=>"000000000",
  5604=>"011001111",
  5605=>"010001111",
  5606=>"011011111",
  5607=>"101100000",
  5608=>"001001111",
  5609=>"001110101",
  5610=>"011100101",
  5611=>"110000100",
  5612=>"011011011",
  5613=>"010010111",
  5614=>"001011101",
  5615=>"001010110",
  5616=>"110001111",
  5617=>"100010110",
  5618=>"010100101",
  5619=>"001111110",
  5620=>"110011011",
  5621=>"000011110",
  5622=>"011011110",
  5623=>"110101000",
  5624=>"001010000",
  5625=>"111001100",
  5626=>"010001100",
  5627=>"000101010",
  5628=>"111111111",
  5629=>"111111100",
  5630=>"110100110",
  5631=>"100000111",
  5632=>"101000010",
  5633=>"110010010",
  5634=>"110000111",
  5635=>"101101110",
  5636=>"001000101",
  5637=>"111001111",
  5638=>"101110010",
  5639=>"000100000",
  5640=>"110011011",
  5641=>"100101010",
  5642=>"001001010",
  5643=>"101100100",
  5644=>"001010100",
  5645=>"001111010",
  5646=>"000010101",
  5647=>"001110000",
  5648=>"000001010",
  5649=>"100011001",
  5650=>"100000010",
  5651=>"010000100",
  5652=>"110011110",
  5653=>"000000011",
  5654=>"011011101",
  5655=>"101010110",
  5656=>"010100100",
  5657=>"001111111",
  5658=>"001101011",
  5659=>"101110100",
  5660=>"010000001",
  5661=>"111011010",
  5662=>"101110001",
  5663=>"101101011",
  5664=>"110011111",
  5665=>"100110110",
  5666=>"111101000",
  5667=>"001001011",
  5668=>"011110111",
  5669=>"001001010",
  5670=>"000000011",
  5671=>"111011110",
  5672=>"001011100",
  5673=>"011001110",
  5674=>"111111000",
  5675=>"010011011",
  5676=>"011001111",
  5677=>"010010001",
  5678=>"110001011",
  5679=>"110010011",
  5680=>"100110001",
  5681=>"000000000",
  5682=>"001011000",
  5683=>"100010010",
  5684=>"110000100",
  5685=>"100010010",
  5686=>"101011000",
  5687=>"110001111",
  5688=>"100101011",
  5689=>"110111111",
  5690=>"101010100",
  5691=>"111010100",
  5692=>"111001100",
  5693=>"011100010",
  5694=>"110001000",
  5695=>"001110010",
  5696=>"110111110",
  5697=>"100111001",
  5698=>"100011000",
  5699=>"011111111",
  5700=>"100100100",
  5701=>"101011101",
  5702=>"000001100",
  5703=>"101111010",
  5704=>"010100110",
  5705=>"111111101",
  5706=>"001001011",
  5707=>"010000000",
  5708=>"110111111",
  5709=>"100001100",
  5710=>"101001111",
  5711=>"101001000",
  5712=>"100010101",
  5713=>"011111000",
  5714=>"000001001",
  5715=>"010011010",
  5716=>"010000100",
  5717=>"110000000",
  5718=>"011101010",
  5719=>"110000111",
  5720=>"111001001",
  5721=>"100000001",
  5722=>"100010101",
  5723=>"000001000",
  5724=>"010110000",
  5725=>"100001100",
  5726=>"110110011",
  5727=>"000000001",
  5728=>"100110011",
  5729=>"100000000",
  5730=>"110011101",
  5731=>"111111100",
  5732=>"010001100",
  5733=>"111000110",
  5734=>"000110111",
  5735=>"000101010",
  5736=>"000100111",
  5737=>"111111011",
  5738=>"110011110",
  5739=>"011111000",
  5740=>"011010100",
  5741=>"110011101",
  5742=>"010111011",
  5743=>"010001100",
  5744=>"101110101",
  5745=>"110011010",
  5746=>"001111111",
  5747=>"010100110",
  5748=>"110100101",
  5749=>"001100010",
  5750=>"011100000",
  5751=>"010101001",
  5752=>"101100110",
  5753=>"000010110",
  5754=>"010100101",
  5755=>"110100010",
  5756=>"110011111",
  5757=>"110011010",
  5758=>"110101110",
  5759=>"100011000",
  5760=>"010001001",
  5761=>"010110100",
  5762=>"110101111",
  5763=>"100100010",
  5764=>"001110001",
  5765=>"100011011",
  5766=>"010001101",
  5767=>"101000101",
  5768=>"101100100",
  5769=>"111111001",
  5770=>"101100100",
  5771=>"110011101",
  5772=>"000111111",
  5773=>"001011000",
  5774=>"010001111",
  5775=>"001010010",
  5776=>"011110100",
  5777=>"101100011",
  5778=>"001111001",
  5779=>"101110010",
  5780=>"111101000",
  5781=>"101100010",
  5782=>"010001000",
  5783=>"011100001",
  5784=>"100010011",
  5785=>"011100101",
  5786=>"000110111",
  5787=>"010110010",
  5788=>"011001001",
  5789=>"110000110",
  5790=>"101101100",
  5791=>"001111100",
  5792=>"000010010",
  5793=>"010101111",
  5794=>"100000000",
  5795=>"100011110",
  5796=>"001100110",
  5797=>"000111111",
  5798=>"001101010",
  5799=>"100100110",
  5800=>"010000100",
  5801=>"100000010",
  5802=>"101010010",
  5803=>"111010001",
  5804=>"111000110",
  5805=>"010000010",
  5806=>"011000101",
  5807=>"111010000",
  5808=>"000111010",
  5809=>"010100000",
  5810=>"010000101",
  5811=>"111111100",
  5812=>"101001011",
  5813=>"000001100",
  5814=>"101100110",
  5815=>"001111111",
  5816=>"011001110",
  5817=>"001111101",
  5818=>"110111000",
  5819=>"010000110",
  5820=>"001010011",
  5821=>"100101100",
  5822=>"001111010",
  5823=>"111110111",
  5824=>"000001011",
  5825=>"010101000",
  5826=>"001111100",
  5827=>"111000000",
  5828=>"110101111",
  5829=>"010110000",
  5830=>"110011111",
  5831=>"110000000",
  5832=>"100101110",
  5833=>"000010111",
  5834=>"110101010",
  5835=>"000100001",
  5836=>"101111101",
  5837=>"101010011",
  5838=>"110000000",
  5839=>"001111111",
  5840=>"001011111",
  5841=>"111010111",
  5842=>"101001101",
  5843=>"111000000",
  5844=>"000111011",
  5845=>"000011010",
  5846=>"110100011",
  5847=>"111000000",
  5848=>"010100001",
  5849=>"001100001",
  5850=>"001101101",
  5851=>"101000000",
  5852=>"101110000",
  5853=>"101110000",
  5854=>"100000100",
  5855=>"011000001",
  5856=>"110100110",
  5857=>"101010110",
  5858=>"011100001",
  5859=>"001010011",
  5860=>"000100010",
  5861=>"010010000",
  5862=>"001011011",
  5863=>"101111000",
  5864=>"111011000",
  5865=>"001010011",
  5866=>"001111000",
  5867=>"000000000",
  5868=>"011111000",
  5869=>"010010100",
  5870=>"111010100",
  5871=>"100010001",
  5872=>"111010010",
  5873=>"110111110",
  5874=>"111000000",
  5875=>"101101000",
  5876=>"010101100",
  5877=>"000101000",
  5878=>"000010110",
  5879=>"111000110",
  5880=>"010000110",
  5881=>"110010010",
  5882=>"111011111",
  5883=>"001010010",
  5884=>"110001010",
  5885=>"101110001",
  5886=>"000111010",
  5887=>"000111110",
  5888=>"101111001",
  5889=>"011110011",
  5890=>"010110111",
  5891=>"001001000",
  5892=>"111111111",
  5893=>"100000011",
  5894=>"010001110",
  5895=>"110111001",
  5896=>"111001010",
  5897=>"100011110",
  5898=>"011101001",
  5899=>"011111110",
  5900=>"000100111",
  5901=>"111100111",
  5902=>"100000000",
  5903=>"110000000",
  5904=>"000011110",
  5905=>"001011110",
  5906=>"001010110",
  5907=>"000110010",
  5908=>"010000010",
  5909=>"000110110",
  5910=>"010110011",
  5911=>"001000011",
  5912=>"000101011",
  5913=>"111111100",
  5914=>"000001110",
  5915=>"111011010",
  5916=>"110100111",
  5917=>"000000000",
  5918=>"001001010",
  5919=>"000011110",
  5920=>"100101011",
  5921=>"100101101",
  5922=>"010010010",
  5923=>"011111100",
  5924=>"010000000",
  5925=>"111011011",
  5926=>"111110001",
  5927=>"000101101",
  5928=>"101001010",
  5929=>"001011111",
  5930=>"001101110",
  5931=>"111000000",
  5932=>"000100110",
  5933=>"011111000",
  5934=>"000111010",
  5935=>"000101110",
  5936=>"001001110",
  5937=>"101010001",
  5938=>"001001110",
  5939=>"111110000",
  5940=>"100110100",
  5941=>"111110110",
  5942=>"100110101",
  5943=>"101011001",
  5944=>"110111110",
  5945=>"100001111",
  5946=>"010010011",
  5947=>"001011011",
  5948=>"000001001",
  5949=>"001101101",
  5950=>"010110000",
  5951=>"110010011",
  5952=>"000110101",
  5953=>"001000100",
  5954=>"001110010",
  5955=>"000011000",
  5956=>"011001010",
  5957=>"111110111",
  5958=>"010001010",
  5959=>"111101111",
  5960=>"001000100",
  5961=>"111111010",
  5962=>"001110011",
  5963=>"000111010",
  5964=>"110110100",
  5965=>"010100001",
  5966=>"001101011",
  5967=>"000000101",
  5968=>"100100110",
  5969=>"001011101",
  5970=>"001000100",
  5971=>"101010001",
  5972=>"111111000",
  5973=>"010000011",
  5974=>"000010000",
  5975=>"000110010",
  5976=>"000110100",
  5977=>"000010010",
  5978=>"111011011",
  5979=>"001010001",
  5980=>"101000001",
  5981=>"111111111",
  5982=>"000011001",
  5983=>"010010111",
  5984=>"010001101",
  5985=>"111111111",
  5986=>"001001000",
  5987=>"101011111",
  5988=>"100011110",
  5989=>"110110011",
  5990=>"100010101",
  5991=>"110001000",
  5992=>"010110111",
  5993=>"011111111",
  5994=>"011001111",
  5995=>"000000111",
  5996=>"110100011",
  5997=>"111001000",
  5998=>"111110100",
  5999=>"100000010",
  6000=>"110000000",
  6001=>"101100100",
  6002=>"111011111",
  6003=>"001010110",
  6004=>"101010111",
  6005=>"001101000",
  6006=>"001010111",
  6007=>"011101101",
  6008=>"100111100",
  6009=>"001001010",
  6010=>"110010010",
  6011=>"111111100",
  6012=>"111101010",
  6013=>"001010010",
  6014=>"110110000",
  6015=>"010100010",
  6016=>"111011101",
  6017=>"011001100",
  6018=>"011101111",
  6019=>"011011011",
  6020=>"010111000",
  6021=>"100000100",
  6022=>"111111101",
  6023=>"000100000",
  6024=>"110110001",
  6025=>"000111101",
  6026=>"010010110",
  6027=>"011110111",
  6028=>"101111100",
  6029=>"111100111",
  6030=>"001000101",
  6031=>"110101110",
  6032=>"111100110",
  6033=>"001100010",
  6034=>"101100000",
  6035=>"010100001",
  6036=>"010101100",
  6037=>"111010110",
  6038=>"011011101",
  6039=>"100010001",
  6040=>"010111011",
  6041=>"010100000",
  6042=>"111110001",
  6043=>"010000111",
  6044=>"001101000",
  6045=>"111010010",
  6046=>"010000001",
  6047=>"010010010",
  6048=>"011000100",
  6049=>"001010100",
  6050=>"000111101",
  6051=>"010010001",
  6052=>"100101011",
  6053=>"111110000",
  6054=>"111110000",
  6055=>"010110101",
  6056=>"110001100",
  6057=>"101110111",
  6058=>"110110111",
  6059=>"011101001",
  6060=>"100000100",
  6061=>"011100010",
  6062=>"010101110",
  6063=>"111111110",
  6064=>"010011110",
  6065=>"100101100",
  6066=>"100100011",
  6067=>"000000110",
  6068=>"010001010",
  6069=>"001000001",
  6070=>"010011100",
  6071=>"011110100",
  6072=>"011100100",
  6073=>"111000101",
  6074=>"001000110",
  6075=>"011001001",
  6076=>"110110111",
  6077=>"100110111",
  6078=>"011110001",
  6079=>"101110111",
  6080=>"101100111",
  6081=>"111111001",
  6082=>"001000011",
  6083=>"100001011",
  6084=>"101100111",
  6085=>"011000010",
  6086=>"000001101",
  6087=>"011010100",
  6088=>"100111110",
  6089=>"010101100",
  6090=>"010010101",
  6091=>"110011010",
  6092=>"000001101",
  6093=>"010001001",
  6094=>"101111001",
  6095=>"100111110",
  6096=>"100101111",
  6097=>"001011101",
  6098=>"010101001",
  6099=>"111110100",
  6100=>"001010011",
  6101=>"000011110",
  6102=>"110110111",
  6103=>"111101010",
  6104=>"000000111",
  6105=>"101110010",
  6106=>"001000100",
  6107=>"000100101",
  6108=>"110111011",
  6109=>"111111010",
  6110=>"001110100",
  6111=>"011100100",
  6112=>"000011101",
  6113=>"000010100",
  6114=>"100001001",
  6115=>"111110010",
  6116=>"000111100",
  6117=>"000000101",
  6118=>"011011000",
  6119=>"000100110",
  6120=>"110111110",
  6121=>"111110100",
  6122=>"001011100",
  6123=>"101000100",
  6124=>"100101001",
  6125=>"001100111",
  6126=>"111110111",
  6127=>"010000111",
  6128=>"110110000",
  6129=>"000011000",
  6130=>"000000110",
  6131=>"000000010",
  6132=>"001111101",
  6133=>"011111101",
  6134=>"010110110",
  6135=>"000010101",
  6136=>"010110000",
  6137=>"111010100",
  6138=>"000110111",
  6139=>"110111001",
  6140=>"100010111",
  6141=>"110000011",
  6142=>"111001001",
  6143=>"000011101",
  6144=>"110110111",
  6145=>"100111011",
  6146=>"000010100",
  6147=>"010110000",
  6148=>"101100111",
  6149=>"011000001",
  6150=>"101011110",
  6151=>"011001001",
  6152=>"011001111",
  6153=>"001100110",
  6154=>"001010011",
  6155=>"001110111",
  6156=>"001111011",
  6157=>"100101000",
  6158=>"000100001",
  6159=>"101100001",
  6160=>"010001111",
  6161=>"000100101",
  6162=>"010010111",
  6163=>"011100000",
  6164=>"011101011",
  6165=>"111100110",
  6166=>"111110101",
  6167=>"101011111",
  6168=>"111000000",
  6169=>"001101000",
  6170=>"111010011",
  6171=>"000011000",
  6172=>"100010011",
  6173=>"101111001",
  6174=>"010101001",
  6175=>"101000100",
  6176=>"111001011",
  6177=>"010111111",
  6178=>"111010011",
  6179=>"100111011",
  6180=>"101111100",
  6181=>"000011000",
  6182=>"000011001",
  6183=>"011000101",
  6184=>"011101111",
  6185=>"001100000",
  6186=>"110111100",
  6187=>"110100110",
  6188=>"000000100",
  6189=>"001000100",
  6190=>"110010000",
  6191=>"110101000",
  6192=>"010111000",
  6193=>"010110110",
  6194=>"011101101",
  6195=>"100000001",
  6196=>"010111100",
  6197=>"001001110",
  6198=>"011010010",
  6199=>"101101100",
  6200=>"101001010",
  6201=>"110011011",
  6202=>"000101111",
  6203=>"010100110",
  6204=>"000111000",
  6205=>"000011110",
  6206=>"010001000",
  6207=>"010101101",
  6208=>"001101101",
  6209=>"010001011",
  6210=>"000101000",
  6211=>"101111010",
  6212=>"110000001",
  6213=>"010011010",
  6214=>"011010101",
  6215=>"100000010",
  6216=>"101110110",
  6217=>"100001111",
  6218=>"110101010",
  6219=>"110010110",
  6220=>"010000010",
  6221=>"111001000",
  6222=>"111101100",
  6223=>"010000001",
  6224=>"100101100",
  6225=>"001101101",
  6226=>"010000110",
  6227=>"101001100",
  6228=>"110111010",
  6229=>"010011000",
  6230=>"011101011",
  6231=>"101001011",
  6232=>"000000111",
  6233=>"110101110",
  6234=>"011010010",
  6235=>"001111100",
  6236=>"011101111",
  6237=>"101111110",
  6238=>"010110100",
  6239=>"100101000",
  6240=>"101111011",
  6241=>"010111111",
  6242=>"110001001",
  6243=>"000000000",
  6244=>"000010101",
  6245=>"111010111",
  6246=>"011001001",
  6247=>"100100001",
  6248=>"010001110",
  6249=>"111101001",
  6250=>"110101100",
  6251=>"000010000",
  6252=>"100011100",
  6253=>"100100001",
  6254=>"100000100",
  6255=>"111101000",
  6256=>"000010011",
  6257=>"000010011",
  6258=>"100111110",
  6259=>"010111111",
  6260=>"001010011",
  6261=>"100010010",
  6262=>"011001111",
  6263=>"110111110",
  6264=>"100111110",
  6265=>"000000111",
  6266=>"000111011",
  6267=>"100001110",
  6268=>"010010111",
  6269=>"000001111",
  6270=>"100000101",
  6271=>"001000101",
  6272=>"001100010",
  6273=>"110110111",
  6274=>"011011100",
  6275=>"001001100",
  6276=>"100000010",
  6277=>"110011101",
  6278=>"100000111",
  6279=>"111110010",
  6280=>"010101001",
  6281=>"001001000",
  6282=>"110001010",
  6283=>"111101111",
  6284=>"100001001",
  6285=>"111001000",
  6286=>"000011000",
  6287=>"101010110",
  6288=>"011101110",
  6289=>"101011111",
  6290=>"110100011",
  6291=>"110111110",
  6292=>"011101010",
  6293=>"000110101",
  6294=>"011101111",
  6295=>"100011101",
  6296=>"011011111",
  6297=>"110011111",
  6298=>"101010100",
  6299=>"111100101",
  6300=>"111001010",
  6301=>"111100010",
  6302=>"000001000",
  6303=>"011000101",
  6304=>"010100101",
  6305=>"111101111",
  6306=>"111111011",
  6307=>"011101010",
  6308=>"010111001",
  6309=>"100111111",
  6310=>"011101101",
  6311=>"001000100",
  6312=>"101101001",
  6313=>"111101001",
  6314=>"101111000",
  6315=>"100111011",
  6316=>"011011101",
  6317=>"010100000",
  6318=>"000000110",
  6319=>"001111010",
  6320=>"100101100",
  6321=>"000011000",
  6322=>"111000011",
  6323=>"001111010",
  6324=>"010111011",
  6325=>"001001001",
  6326=>"010000110",
  6327=>"100101110",
  6328=>"110110001",
  6329=>"000100011",
  6330=>"101111010",
  6331=>"110100010",
  6332=>"000000001",
  6333=>"001111111",
  6334=>"010100110",
  6335=>"101100101",
  6336=>"011110010",
  6337=>"001111000",
  6338=>"000111110",
  6339=>"111111110",
  6340=>"110110110",
  6341=>"101111011",
  6342=>"010010100",
  6343=>"011011011",
  6344=>"101111001",
  6345=>"101001110",
  6346=>"000000011",
  6347=>"110001100",
  6348=>"111011101",
  6349=>"111111000",
  6350=>"001001000",
  6351=>"001110111",
  6352=>"001010110",
  6353=>"111100100",
  6354=>"001101000",
  6355=>"011010010",
  6356=>"111101110",
  6357=>"001111000",
  6358=>"110000101",
  6359=>"011010010",
  6360=>"000111011",
  6361=>"010110000",
  6362=>"011000100",
  6363=>"010000110",
  6364=>"001011000",
  6365=>"000110111",
  6366=>"110010000",
  6367=>"110101000",
  6368=>"111000111",
  6369=>"001000101",
  6370=>"100011000",
  6371=>"111011111",
  6372=>"111011100",
  6373=>"100111110",
  6374=>"001101100",
  6375=>"000011001",
  6376=>"100110111",
  6377=>"101111110",
  6378=>"000010100",
  6379=>"001011001",
  6380=>"010001110",
  6381=>"100110001",
  6382=>"110101111",
  6383=>"010101001",
  6384=>"111101101",
  6385=>"001010111",
  6386=>"000100101",
  6387=>"001011010",
  6388=>"111001100",
  6389=>"010001111",
  6390=>"011000000",
  6391=>"111101001",
  6392=>"000111101",
  6393=>"111010000",
  6394=>"011000001",
  6395=>"001010000",
  6396=>"000010111",
  6397=>"001111011",
  6398=>"101000101",
  6399=>"101101110",
  6400=>"000110001",
  6401=>"111000000",
  6402=>"001011100",
  6403=>"001011101",
  6404=>"010110111",
  6405=>"000001010",
  6406=>"111100011",
  6407=>"000101100",
  6408=>"000100100",
  6409=>"011110101",
  6410=>"110111110",
  6411=>"110011101",
  6412=>"010011110",
  6413=>"000101011",
  6414=>"110101001",
  6415=>"111010100",
  6416=>"000101101",
  6417=>"101101111",
  6418=>"100010110",
  6419=>"110110111",
  6420=>"000001111",
  6421=>"010011110",
  6422=>"010111100",
  6423=>"101100101",
  6424=>"000001111",
  6425=>"001010000",
  6426=>"101011001",
  6427=>"000100100",
  6428=>"100010110",
  6429=>"000000110",
  6430=>"011001000",
  6431=>"101000011",
  6432=>"101110010",
  6433=>"110100100",
  6434=>"011101011",
  6435=>"010111100",
  6436=>"100111011",
  6437=>"000110001",
  6438=>"000011010",
  6439=>"000111110",
  6440=>"100101000",
  6441=>"011000100",
  6442=>"011110010",
  6443=>"110110101",
  6444=>"001011001",
  6445=>"001010000",
  6446=>"111100111",
  6447=>"101000010",
  6448=>"100101110",
  6449=>"001010001",
  6450=>"100111011",
  6451=>"101111110",
  6452=>"001000111",
  6453=>"110000111",
  6454=>"001010100",
  6455=>"111001000",
  6456=>"101101110",
  6457=>"101001110",
  6458=>"101011101",
  6459=>"110100001",
  6460=>"011010010",
  6461=>"111000110",
  6462=>"001001010",
  6463=>"110110110",
  6464=>"111110100",
  6465=>"011100001",
  6466=>"010000111",
  6467=>"001000100",
  6468=>"100100001",
  6469=>"010111010",
  6470=>"010011111",
  6471=>"011111101",
  6472=>"010111111",
  6473=>"101100010",
  6474=>"111111101",
  6475=>"000101001",
  6476=>"011111110",
  6477=>"111110101",
  6478=>"010000010",
  6479=>"000100000",
  6480=>"010000101",
  6481=>"111101101",
  6482=>"010010010",
  6483=>"000100101",
  6484=>"100111110",
  6485=>"010010000",
  6486=>"001010110",
  6487=>"011011001",
  6488=>"000011111",
  6489=>"101100110",
  6490=>"111011010",
  6491=>"011101001",
  6492=>"011110100",
  6493=>"100001111",
  6494=>"110100001",
  6495=>"001110111",
  6496=>"100101001",
  6497=>"100010000",
  6498=>"011010000",
  6499=>"011100001",
  6500=>"101100011",
  6501=>"010111001",
  6502=>"100100001",
  6503=>"000100001",
  6504=>"101111111",
  6505=>"001001100",
  6506=>"010101000",
  6507=>"111111111",
  6508=>"110000110",
  6509=>"101110010",
  6510=>"110011111",
  6511=>"010011011",
  6512=>"110010100",
  6513=>"110011110",
  6514=>"000100101",
  6515=>"111011110",
  6516=>"010011001",
  6517=>"001011110",
  6518=>"111100111",
  6519=>"011011010",
  6520=>"001110010",
  6521=>"011101001",
  6522=>"111110101",
  6523=>"011110000",
  6524=>"110111000",
  6525=>"110110000",
  6526=>"001010000",
  6527=>"010101010",
  6528=>"101001110",
  6529=>"100111100",
  6530=>"100010000",
  6531=>"000001001",
  6532=>"101110011",
  6533=>"101010001",
  6534=>"110111001",
  6535=>"111111000",
  6536=>"001000010",
  6537=>"000010010",
  6538=>"111110011",
  6539=>"101000100",
  6540=>"010000100",
  6541=>"001001101",
  6542=>"101001010",
  6543=>"010110110",
  6544=>"010011110",
  6545=>"000001110",
  6546=>"111111010",
  6547=>"000101110",
  6548=>"101100001",
  6549=>"100011001",
  6550=>"110010011",
  6551=>"100111011",
  6552=>"110010101",
  6553=>"000001001",
  6554=>"000011101",
  6555=>"010001011",
  6556=>"101011010",
  6557=>"010100000",
  6558=>"101010011",
  6559=>"011101010",
  6560=>"100100100",
  6561=>"001011111",
  6562=>"000000111",
  6563=>"000010001",
  6564=>"011111101",
  6565=>"001101000",
  6566=>"001111110",
  6567=>"110000010",
  6568=>"100110011",
  6569=>"011001100",
  6570=>"011111011",
  6571=>"001001101",
  6572=>"001011101",
  6573=>"000010111",
  6574=>"011010100",
  6575=>"110111011",
  6576=>"000101111",
  6577=>"011001101",
  6578=>"000010100",
  6579=>"011110111",
  6580=>"010011011",
  6581=>"110111000",
  6582=>"011001001",
  6583=>"110000110",
  6584=>"010011101",
  6585=>"001011000",
  6586=>"010100000",
  6587=>"011101101",
  6588=>"000001000",
  6589=>"110111011",
  6590=>"010101111",
  6591=>"100110111",
  6592=>"110110000",
  6593=>"011101101",
  6594=>"101101110",
  6595=>"011101111",
  6596=>"101010101",
  6597=>"000000011",
  6598=>"111000101",
  6599=>"010011010",
  6600=>"110101101",
  6601=>"000001100",
  6602=>"100010010",
  6603=>"010010101",
  6604=>"001000010",
  6605=>"001010101",
  6606=>"001110000",
  6607=>"010000011",
  6608=>"000100111",
  6609=>"011110001",
  6610=>"000010011",
  6611=>"110100001",
  6612=>"111011100",
  6613=>"110000100",
  6614=>"100001010",
  6615=>"110101011",
  6616=>"001011001",
  6617=>"110110111",
  6618=>"110000011",
  6619=>"000101100",
  6620=>"110110100",
  6621=>"011001001",
  6622=>"111100101",
  6623=>"100110111",
  6624=>"100111110",
  6625=>"001011101",
  6626=>"100010011",
  6627=>"100010010",
  6628=>"011011011",
  6629=>"110011011",
  6630=>"000001101",
  6631=>"010001000",
  6632=>"010101100",
  6633=>"011000110",
  6634=>"001100001",
  6635=>"100000010",
  6636=>"011001011",
  6637=>"111000111",
  6638=>"001111100",
  6639=>"010110111",
  6640=>"001010010",
  6641=>"010110110",
  6642=>"110101111",
  6643=>"111111001",
  6644=>"100110100",
  6645=>"011001111",
  6646=>"111000110",
  6647=>"100011100",
  6648=>"101110000",
  6649=>"010111010",
  6650=>"010000110",
  6651=>"101011111",
  6652=>"001101000",
  6653=>"100111100",
  6654=>"011001111",
  6655=>"101111010",
  6656=>"111111100",
  6657=>"110110100",
  6658=>"011010110",
  6659=>"010110100",
  6660=>"100011111",
  6661=>"001010100",
  6662=>"110010101",
  6663=>"100010110",
  6664=>"011110010",
  6665=>"110110111",
  6666=>"101001111",
  6667=>"110111100",
  6668=>"000010111",
  6669=>"111011000",
  6670=>"111000001",
  6671=>"101001111",
  6672=>"111010011",
  6673=>"000011000",
  6674=>"010101011",
  6675=>"011111000",
  6676=>"100100011",
  6677=>"111111011",
  6678=>"010000101",
  6679=>"110010011",
  6680=>"010001011",
  6681=>"111001101",
  6682=>"101101000",
  6683=>"111011010",
  6684=>"010000110",
  6685=>"001010111",
  6686=>"000011011",
  6687=>"100110111",
  6688=>"111111011",
  6689=>"010111000",
  6690=>"110001101",
  6691=>"001110101",
  6692=>"000100001",
  6693=>"100111000",
  6694=>"001100001",
  6695=>"111010011",
  6696=>"011001101",
  6697=>"100110000",
  6698=>"110101100",
  6699=>"110011100",
  6700=>"100010010",
  6701=>"000001000",
  6702=>"010100100",
  6703=>"100100110",
  6704=>"001001111",
  6705=>"111110011",
  6706=>"111111000",
  6707=>"100001110",
  6708=>"110001101",
  6709=>"011000001",
  6710=>"010100011",
  6711=>"101000000",
  6712=>"100100011",
  6713=>"100101100",
  6714=>"111110010",
  6715=>"111110101",
  6716=>"100100110",
  6717=>"110111101",
  6718=>"100000011",
  6719=>"000011100",
  6720=>"001000010",
  6721=>"000000000",
  6722=>"010110110",
  6723=>"100110111",
  6724=>"100101101",
  6725=>"000100111",
  6726=>"001001110",
  6727=>"101111000",
  6728=>"100101111",
  6729=>"010001101",
  6730=>"011011000",
  6731=>"011001100",
  6732=>"000001100",
  6733=>"010000111",
  6734=>"110101010",
  6735=>"000110011",
  6736=>"100100111",
  6737=>"000111101",
  6738=>"100001011",
  6739=>"100110001",
  6740=>"000101100",
  6741=>"101111010",
  6742=>"000100000",
  6743=>"001010100",
  6744=>"001111011",
  6745=>"010111110",
  6746=>"010001100",
  6747=>"100001101",
  6748=>"110010111",
  6749=>"001000110",
  6750=>"111111010",
  6751=>"110011011",
  6752=>"000011111",
  6753=>"101001111",
  6754=>"110100101",
  6755=>"000011101",
  6756=>"010011110",
  6757=>"111000111",
  6758=>"100011101",
  6759=>"000010010",
  6760=>"011111101",
  6761=>"111000100",
  6762=>"101001110",
  6763=>"000000001",
  6764=>"101011000",
  6765=>"100111010",
  6766=>"011011010",
  6767=>"111011001",
  6768=>"001011000",
  6769=>"011000101",
  6770=>"110100011",
  6771=>"011010010",
  6772=>"001111001",
  6773=>"000111001",
  6774=>"100000010",
  6775=>"101100110",
  6776=>"110110110",
  6777=>"101101010",
  6778=>"001010010",
  6779=>"111001100",
  6780=>"010110101",
  6781=>"110101100",
  6782=>"110101100",
  6783=>"000100111",
  6784=>"110001001",
  6785=>"011110111",
  6786=>"000110001",
  6787=>"110001101",
  6788=>"100101011",
  6789=>"010101101",
  6790=>"011101111",
  6791=>"010001011",
  6792=>"001100001",
  6793=>"000001011",
  6794=>"100101011",
  6795=>"111011110",
  6796=>"000111011",
  6797=>"001010111",
  6798=>"010101101",
  6799=>"010111011",
  6800=>"100100100",
  6801=>"110011010",
  6802=>"000110011",
  6803=>"111101111",
  6804=>"001111110",
  6805=>"100101101",
  6806=>"100101010",
  6807=>"011100111",
  6808=>"001101110",
  6809=>"111010110",
  6810=>"010011011",
  6811=>"000010100",
  6812=>"101011100",
  6813=>"001010010",
  6814=>"000001100",
  6815=>"100101100",
  6816=>"001000011",
  6817=>"111001000",
  6818=>"111111011",
  6819=>"001110000",
  6820=>"000010010",
  6821=>"010010100",
  6822=>"011110100",
  6823=>"010100110",
  6824=>"011001000",
  6825=>"101000100",
  6826=>"000010001",
  6827=>"100000000",
  6828=>"001111000",
  6829=>"110101110",
  6830=>"111101100",
  6831=>"010101010",
  6832=>"101011111",
  6833=>"001100011",
  6834=>"010011001",
  6835=>"011011111",
  6836=>"000010000",
  6837=>"110111101",
  6838=>"101011101",
  6839=>"110000000",
  6840=>"111010000",
  6841=>"110001000",
  6842=>"001100101",
  6843=>"010100011",
  6844=>"000001111",
  6845=>"001001111",
  6846=>"001011010",
  6847=>"110000111",
  6848=>"000010001",
  6849=>"110001011",
  6850=>"110111011",
  6851=>"110011111",
  6852=>"101011101",
  6853=>"001000111",
  6854=>"111100010",
  6855=>"100010000",
  6856=>"101111001",
  6857=>"111111011",
  6858=>"101100011",
  6859=>"000100011",
  6860=>"010010111",
  6861=>"100000001",
  6862=>"001000000",
  6863=>"111011110",
  6864=>"110001111",
  6865=>"001001010",
  6866=>"011001010",
  6867=>"110001110",
  6868=>"000010101",
  6869=>"100010111",
  6870=>"101010000",
  6871=>"010001101",
  6872=>"111011111",
  6873=>"111001101",
  6874=>"111011011",
  6875=>"101001101",
  6876=>"111101010",
  6877=>"000000101",
  6878=>"111000010",
  6879=>"111010101",
  6880=>"000101010",
  6881=>"110001000",
  6882=>"011000111",
  6883=>"101111010",
  6884=>"000011000",
  6885=>"001000001",
  6886=>"110010000",
  6887=>"001001111",
  6888=>"001111101",
  6889=>"000111100",
  6890=>"001100101",
  6891=>"010111110",
  6892=>"000001010",
  6893=>"011100111",
  6894=>"101010110",
  6895=>"001011111",
  6896=>"101000111",
  6897=>"100010001",
  6898=>"110111000",
  6899=>"000110110",
  6900=>"110010000",
  6901=>"101100010",
  6902=>"101000001",
  6903=>"011011100",
  6904=>"010100001",
  6905=>"101101100",
  6906=>"101111101",
  6907=>"011000110",
  6908=>"000010111",
  6909=>"101000111",
  6910=>"111011011",
  6911=>"100111000",
  6912=>"110011011",
  6913=>"011110111",
  6914=>"000111010",
  6915=>"101010100",
  6916=>"000110101",
  6917=>"000000100",
  6918=>"000111100",
  6919=>"011111110",
  6920=>"111001111",
  6921=>"011110010",
  6922=>"100101011",
  6923=>"010000100",
  6924=>"100110100",
  6925=>"111000111",
  6926=>"001100111",
  6927=>"111001100",
  6928=>"111110110",
  6929=>"011101111",
  6930=>"010110000",
  6931=>"011110011",
  6932=>"100100001",
  6933=>"100100001",
  6934=>"011100010",
  6935=>"000011110",
  6936=>"001111100",
  6937=>"000010000",
  6938=>"101010010",
  6939=>"111111000",
  6940=>"001010111",
  6941=>"110000010",
  6942=>"000000001",
  6943=>"010110100",
  6944=>"110010111",
  6945=>"000101011",
  6946=>"001000000",
  6947=>"010101101",
  6948=>"110101111",
  6949=>"011010000",
  6950=>"000111110",
  6951=>"010110101",
  6952=>"110111111",
  6953=>"111101111",
  6954=>"000010111",
  6955=>"011011010",
  6956=>"001000101",
  6957=>"100010101",
  6958=>"101001010",
  6959=>"100000100",
  6960=>"001101110",
  6961=>"000100111",
  6962=>"000000001",
  6963=>"110001111",
  6964=>"010111011",
  6965=>"101101011",
  6966=>"001001101",
  6967=>"001011100",
  6968=>"010110101",
  6969=>"000111101",
  6970=>"110100101",
  6971=>"000000101",
  6972=>"010101010",
  6973=>"011001111",
  6974=>"000100011",
  6975=>"001011111",
  6976=>"000000000",
  6977=>"000000100",
  6978=>"000011000",
  6979=>"110000011",
  6980=>"111101111",
  6981=>"010110100",
  6982=>"111001001",
  6983=>"010000010",
  6984=>"000000010",
  6985=>"010101100",
  6986=>"011011111",
  6987=>"111111110",
  6988=>"011101101",
  6989=>"110110100",
  6990=>"101101010",
  6991=>"110100110",
  6992=>"010010010",
  6993=>"000001111",
  6994=>"001111011",
  6995=>"001011101",
  6996=>"010000001",
  6997=>"001111111",
  6998=>"111100100",
  6999=>"000110010",
  7000=>"101100100",
  7001=>"111111001",
  7002=>"010001100",
  7003=>"101000001",
  7004=>"111011000",
  7005=>"001001011",
  7006=>"011010001",
  7007=>"000010101",
  7008=>"111111010",
  7009=>"100101011",
  7010=>"001000100",
  7011=>"100010010",
  7012=>"011010100",
  7013=>"111011001",
  7014=>"111100011",
  7015=>"100000010",
  7016=>"000100111",
  7017=>"011101110",
  7018=>"110100010",
  7019=>"101110000",
  7020=>"011100100",
  7021=>"001001010",
  7022=>"100010011",
  7023=>"011111010",
  7024=>"110110101",
  7025=>"110100000",
  7026=>"011011001",
  7027=>"011101101",
  7028=>"011011110",
  7029=>"011110100",
  7030=>"010000111",
  7031=>"101101101",
  7032=>"011110000",
  7033=>"010110011",
  7034=>"101000001",
  7035=>"111000010",
  7036=>"001111001",
  7037=>"110101000",
  7038=>"010010010",
  7039=>"110000100",
  7040=>"101100110",
  7041=>"110111001",
  7042=>"000110111",
  7043=>"011010101",
  7044=>"111010001",
  7045=>"010111000",
  7046=>"100100001",
  7047=>"100100001",
  7048=>"001010011",
  7049=>"110010100",
  7050=>"011101000",
  7051=>"010110101",
  7052=>"110110111",
  7053=>"110111101",
  7054=>"001110010",
  7055=>"010110100",
  7056=>"010001100",
  7057=>"111000000",
  7058=>"001111011",
  7059=>"010000100",
  7060=>"001110101",
  7061=>"000100001",
  7062=>"000000101",
  7063=>"011111011",
  7064=>"010000110",
  7065=>"001000010",
  7066=>"110011001",
  7067=>"000110101",
  7068=>"001111110",
  7069=>"110100111",
  7070=>"110111010",
  7071=>"001010110",
  7072=>"001110011",
  7073=>"000000010",
  7074=>"011100100",
  7075=>"101101101",
  7076=>"001001100",
  7077=>"001010011",
  7078=>"001010111",
  7079=>"101110001",
  7080=>"000001111",
  7081=>"010011101",
  7082=>"101010010",
  7083=>"111011011",
  7084=>"110000100",
  7085=>"000110110",
  7086=>"101001110",
  7087=>"010010110",
  7088=>"111110111",
  7089=>"011001010",
  7090=>"101011010",
  7091=>"101000000",
  7092=>"000001110",
  7093=>"111100101",
  7094=>"011111110",
  7095=>"110000101",
  7096=>"100111010",
  7097=>"011011000",
  7098=>"011011100",
  7099=>"111111100",
  7100=>"110001101",
  7101=>"010011001",
  7102=>"010010010",
  7103=>"000000100",
  7104=>"110001001",
  7105=>"010111011",
  7106=>"100111001",
  7107=>"011000011",
  7108=>"100001001",
  7109=>"000101010",
  7110=>"010110000",
  7111=>"010100100",
  7112=>"101000100",
  7113=>"011001000",
  7114=>"111010010",
  7115=>"011101110",
  7116=>"100110100",
  7117=>"011111011",
  7118=>"110000100",
  7119=>"111000101",
  7120=>"111011010",
  7121=>"111111010",
  7122=>"011111010",
  7123=>"110000110",
  7124=>"011111110",
  7125=>"010101011",
  7126=>"000010110",
  7127=>"011101101",
  7128=>"010001001",
  7129=>"011111010",
  7130=>"010101100",
  7131=>"010110100",
  7132=>"001010101",
  7133=>"101100110",
  7134=>"000100001",
  7135=>"110001000",
  7136=>"000011101",
  7137=>"001001100",
  7138=>"000111001",
  7139=>"000101110",
  7140=>"000001010",
  7141=>"011111011",
  7142=>"011011001",
  7143=>"110001000",
  7144=>"110001101",
  7145=>"111011010",
  7146=>"000001100",
  7147=>"000010011",
  7148=>"100100111",
  7149=>"010011001",
  7150=>"011010111",
  7151=>"010011110",
  7152=>"011001100",
  7153=>"001010010",
  7154=>"111011110",
  7155=>"100010100",
  7156=>"100111100",
  7157=>"100001101",
  7158=>"101001001",
  7159=>"011000001",
  7160=>"001000101",
  7161=>"111010110",
  7162=>"110000001",
  7163=>"110000000",
  7164=>"011001110",
  7165=>"001001111",
  7166=>"110100110",
  7167=>"010110011",
  7168=>"111110000",
  7169=>"011101100",
  7170=>"001001001",
  7171=>"110111111",
  7172=>"101110111",
  7173=>"111010010",
  7174=>"101011010",
  7175=>"000001000",
  7176=>"101000001",
  7177=>"010110110",
  7178=>"000010011",
  7179=>"001010000",
  7180=>"011000000",
  7181=>"101001011",
  7182=>"000000111",
  7183=>"110001110",
  7184=>"000100101",
  7185=>"001001000",
  7186=>"100110101",
  7187=>"100000001",
  7188=>"110101001",
  7189=>"001110100",
  7190=>"100000101",
  7191=>"011000000",
  7192=>"000011011",
  7193=>"001000000",
  7194=>"110000101",
  7195=>"101100000",
  7196=>"111111001",
  7197=>"000101100",
  7198=>"011111001",
  7199=>"110011100",
  7200=>"111010010",
  7201=>"011010010",
  7202=>"101111110",
  7203=>"011100000",
  7204=>"110011100",
  7205=>"001000001",
  7206=>"111001101",
  7207=>"010011011",
  7208=>"010111000",
  7209=>"000000001",
  7210=>"001001010",
  7211=>"111001110",
  7212=>"010101011",
  7213=>"001100111",
  7214=>"010101000",
  7215=>"011001101",
  7216=>"011011111",
  7217=>"011110100",
  7218=>"111101000",
  7219=>"100111010",
  7220=>"010000100",
  7221=>"011001001",
  7222=>"100011100",
  7223=>"111000110",
  7224=>"100010011",
  7225=>"111110000",
  7226=>"000111000",
  7227=>"100111010",
  7228=>"001011000",
  7229=>"110100010",
  7230=>"011101101",
  7231=>"111100010",
  7232=>"000011110",
  7233=>"011111000",
  7234=>"000001001",
  7235=>"100011000",
  7236=>"001001111",
  7237=>"100101110",
  7238=>"100011000",
  7239=>"000111101",
  7240=>"111010000",
  7241=>"100010000",
  7242=>"100010010",
  7243=>"100100111",
  7244=>"001100101",
  7245=>"010001011",
  7246=>"110010001",
  7247=>"010001001",
  7248=>"011001101",
  7249=>"100001101",
  7250=>"111101110",
  7251=>"000010000",
  7252=>"110001101",
  7253=>"011110100",
  7254=>"001110111",
  7255=>"111101111",
  7256=>"000101101",
  7257=>"111011000",
  7258=>"010101000",
  7259=>"001110111",
  7260=>"100110011",
  7261=>"010010110",
  7262=>"001000000",
  7263=>"101010000",
  7264=>"000111111",
  7265=>"000001010",
  7266=>"111111111",
  7267=>"011101111",
  7268=>"101010101",
  7269=>"110001001",
  7270=>"000110101",
  7271=>"010001011",
  7272=>"011100000",
  7273=>"011110011",
  7274=>"110011110",
  7275=>"011100011",
  7276=>"101001001",
  7277=>"100101100",
  7278=>"111000101",
  7279=>"010101100",
  7280=>"000001011",
  7281=>"010110010",
  7282=>"100100001",
  7283=>"111000100",
  7284=>"110101101",
  7285=>"111000111",
  7286=>"110111111",
  7287=>"101010001",
  7288=>"001110101",
  7289=>"110110101",
  7290=>"010100001",
  7291=>"110011011",
  7292=>"000100011",
  7293=>"010001100",
  7294=>"110100000",
  7295=>"001110000",
  7296=>"010001000",
  7297=>"000010101",
  7298=>"001101010",
  7299=>"100010000",
  7300=>"011111011",
  7301=>"011111001",
  7302=>"000001100",
  7303=>"111000101",
  7304=>"011110111",
  7305=>"011110101",
  7306=>"101011011",
  7307=>"000010111",
  7308=>"011100100",
  7309=>"010100110",
  7310=>"011001100",
  7311=>"100001100",
  7312=>"110011110",
  7313=>"100011011",
  7314=>"001110100",
  7315=>"011010110",
  7316=>"101100101",
  7317=>"001010010",
  7318=>"010111000",
  7319=>"010101001",
  7320=>"001000000",
  7321=>"001010110",
  7322=>"111000101",
  7323=>"100011011",
  7324=>"100111000",
  7325=>"111111110",
  7326=>"110101011",
  7327=>"001011000",
  7328=>"010100101",
  7329=>"011110011",
  7330=>"001001000",
  7331=>"110000001",
  7332=>"110001011",
  7333=>"000001010",
  7334=>"010100111",
  7335=>"011110100",
  7336=>"100010001",
  7337=>"110010111",
  7338=>"000100000",
  7339=>"010000010",
  7340=>"111011110",
  7341=>"111110101",
  7342=>"001011100",
  7343=>"011101101",
  7344=>"010010101",
  7345=>"000101111",
  7346=>"001000010",
  7347=>"101000110",
  7348=>"110111101",
  7349=>"010010011",
  7350=>"011110001",
  7351=>"100111110",
  7352=>"001101010",
  7353=>"110111111",
  7354=>"101000010",
  7355=>"001111000",
  7356=>"111010010",
  7357=>"011101100",
  7358=>"111100011",
  7359=>"000000100",
  7360=>"011010100",
  7361=>"000100010",
  7362=>"110000110",
  7363=>"010011000",
  7364=>"011100010",
  7365=>"100111101",
  7366=>"110110100",
  7367=>"000011100",
  7368=>"001010111",
  7369=>"000001101",
  7370=>"100010000",
  7371=>"000001011",
  7372=>"010000001",
  7373=>"100101101",
  7374=>"001001001",
  7375=>"010110010",
  7376=>"011010110",
  7377=>"110011110",
  7378=>"001111110",
  7379=>"010000000",
  7380=>"110101010",
  7381=>"000001011",
  7382=>"110011000",
  7383=>"100000011",
  7384=>"100001001",
  7385=>"011000011",
  7386=>"111111001",
  7387=>"001111000",
  7388=>"111100010",
  7389=>"100100101",
  7390=>"011110010",
  7391=>"110111010",
  7392=>"000001000",
  7393=>"010010010",
  7394=>"000111101",
  7395=>"101111110",
  7396=>"110010101",
  7397=>"101000011",
  7398=>"011100011",
  7399=>"010110100",
  7400=>"100101110",
  7401=>"101101101",
  7402=>"101111000",
  7403=>"000101010",
  7404=>"111111100",
  7405=>"010011111",
  7406=>"001010000",
  7407=>"010001110",
  7408=>"101111011",
  7409=>"110111011",
  7410=>"001111110",
  7411=>"000101000",
  7412=>"000001100",
  7413=>"110111001",
  7414=>"010001000",
  7415=>"110010000",
  7416=>"011110111",
  7417=>"010001010",
  7418=>"010010101",
  7419=>"111001000",
  7420=>"011011111",
  7421=>"101111110",
  7422=>"001110100",
  7423=>"010111110",
  7424=>"000001100",
  7425=>"011100010",
  7426=>"100111101",
  7427=>"110001110",
  7428=>"010000000",
  7429=>"010010100",
  7430=>"011100000",
  7431=>"101000011",
  7432=>"000101000",
  7433=>"000010100",
  7434=>"010111011",
  7435=>"011100101",
  7436=>"100101110",
  7437=>"001111101",
  7438=>"010010111",
  7439=>"010000101",
  7440=>"101101110",
  7441=>"110110000",
  7442=>"011001011",
  7443=>"110000110",
  7444=>"000101010",
  7445=>"111101000",
  7446=>"101101110",
  7447=>"001011001",
  7448=>"111100010",
  7449=>"100001101",
  7450=>"000100011",
  7451=>"110011100",
  7452=>"000101100",
  7453=>"111010111",
  7454=>"011100001",
  7455=>"000001000",
  7456=>"000010101",
  7457=>"011010010",
  7458=>"110100101",
  7459=>"101100111",
  7460=>"010100100",
  7461=>"011101111",
  7462=>"000111110",
  7463=>"011101011",
  7464=>"010001010",
  7465=>"010000100",
  7466=>"000001000",
  7467=>"100111111",
  7468=>"101101110",
  7469=>"000101001",
  7470=>"010111000",
  7471=>"010100101",
  7472=>"110100001",
  7473=>"100101110",
  7474=>"000000100",
  7475=>"101010111",
  7476=>"111100101",
  7477=>"111000010",
  7478=>"001101111",
  7479=>"000101010",
  7480=>"110110001",
  7481=>"110001111",
  7482=>"111101111",
  7483=>"111000101",
  7484=>"010110011",
  7485=>"010010100",
  7486=>"000101001",
  7487=>"100000111",
  7488=>"000000011",
  7489=>"000100000",
  7490=>"010001001",
  7491=>"111000111",
  7492=>"010100010",
  7493=>"111111110",
  7494=>"000110100",
  7495=>"110111110",
  7496=>"110101001",
  7497=>"111111011",
  7498=>"011001010",
  7499=>"011001110",
  7500=>"011110000",
  7501=>"001100111",
  7502=>"001010000",
  7503=>"001111011",
  7504=>"101111111",
  7505=>"101101001",
  7506=>"111110001",
  7507=>"011010101",
  7508=>"110110011",
  7509=>"011110000",
  7510=>"111010000",
  7511=>"111101100",
  7512=>"011111101",
  7513=>"011101011",
  7514=>"100101110",
  7515=>"010010001",
  7516=>"100011100",
  7517=>"110111000",
  7518=>"000001000",
  7519=>"010111100",
  7520=>"111011110",
  7521=>"100010001",
  7522=>"001100000",
  7523=>"101110000",
  7524=>"010101110",
  7525=>"110100010",
  7526=>"101111111",
  7527=>"111010000",
  7528=>"000000010",
  7529=>"000010000",
  7530=>"001100000",
  7531=>"101000010",
  7532=>"011101101",
  7533=>"001101011",
  7534=>"000010000",
  7535=>"101011101",
  7536=>"000000100",
  7537=>"111111101",
  7538=>"011010011",
  7539=>"010010011",
  7540=>"110101111",
  7541=>"110111101",
  7542=>"110111111",
  7543=>"001111101",
  7544=>"101110011",
  7545=>"001101010",
  7546=>"010100010",
  7547=>"010100010",
  7548=>"011100100",
  7549=>"011111101",
  7550=>"110101011",
  7551=>"110100110",
  7552=>"111100111",
  7553=>"000100001",
  7554=>"100010000",
  7555=>"000111101",
  7556=>"101110010",
  7557=>"011101000",
  7558=>"001001011",
  7559=>"000001111",
  7560=>"000001000",
  7561=>"010000110",
  7562=>"001000000",
  7563=>"000111110",
  7564=>"101110001",
  7565=>"101111101",
  7566=>"000010100",
  7567=>"000011011",
  7568=>"011011111",
  7569=>"000001110",
  7570=>"010110000",
  7571=>"001110010",
  7572=>"100011111",
  7573=>"101000010",
  7574=>"010111110",
  7575=>"010011111",
  7576=>"111011100",
  7577=>"000000000",
  7578=>"011111101",
  7579=>"111100100",
  7580=>"100101010",
  7581=>"000000010",
  7582=>"110111110",
  7583=>"000000111",
  7584=>"111101010",
  7585=>"000001000",
  7586=>"111101110",
  7587=>"010110000",
  7588=>"000010011",
  7589=>"000111110",
  7590=>"110100000",
  7591=>"001100101",
  7592=>"010111110",
  7593=>"101000011",
  7594=>"101001111",
  7595=>"010011100",
  7596=>"110111111",
  7597=>"001111010",
  7598=>"011111100",
  7599=>"010111010",
  7600=>"111110000",
  7601=>"000000010",
  7602=>"110000000",
  7603=>"100001110",
  7604=>"000100000",
  7605=>"010000010",
  7606=>"010101010",
  7607=>"010100000",
  7608=>"111110001",
  7609=>"011110011",
  7610=>"010001000",
  7611=>"101010000",
  7612=>"100111001",
  7613=>"000101110",
  7614=>"111111110",
  7615=>"100101111",
  7616=>"111111100",
  7617=>"101111111",
  7618=>"110111001",
  7619=>"101011000",
  7620=>"001011000",
  7621=>"001010110",
  7622=>"111010001",
  7623=>"000110000",
  7624=>"101001111",
  7625=>"010100010",
  7626=>"011000011",
  7627=>"101111010",
  7628=>"111100011",
  7629=>"101110101",
  7630=>"000001011",
  7631=>"000010010",
  7632=>"100110011",
  7633=>"100101010",
  7634=>"110011100",
  7635=>"110000000",
  7636=>"101010000",
  7637=>"010111101",
  7638=>"010111001",
  7639=>"000110100",
  7640=>"101111100",
  7641=>"111011101",
  7642=>"001011001",
  7643=>"111110101",
  7644=>"010101100",
  7645=>"011101101",
  7646=>"111111110",
  7647=>"110111110",
  7648=>"101100010",
  7649=>"011000100",
  7650=>"011101110",
  7651=>"000010110",
  7652=>"001101000",
  7653=>"000001111",
  7654=>"011100001",
  7655=>"001000001",
  7656=>"111111111",
  7657=>"111111010",
  7658=>"011000011",
  7659=>"011000000",
  7660=>"101010100",
  7661=>"110110010",
  7662=>"001110111",
  7663=>"010010000",
  7664=>"101110011",
  7665=>"111101010",
  7666=>"111110100",
  7667=>"000000100",
  7668=>"001010100",
  7669=>"110000100",
  7670=>"101001110",
  7671=>"010110010",
  7672=>"111100010",
  7673=>"100101001",
  7674=>"010010001",
  7675=>"111010100",
  7676=>"110000110",
  7677=>"100000111",
  7678=>"000100001",
  7679=>"111111010",
  7680=>"000000111",
  7681=>"110111001",
  7682=>"011101101",
  7683=>"001100110",
  7684=>"001110101",
  7685=>"000011010",
  7686=>"010110101",
  7687=>"111111011",
  7688=>"110100101",
  7689=>"110011010",
  7690=>"100111011",
  7691=>"001110010",
  7692=>"001100001",
  7693=>"111111001",
  7694=>"000101101",
  7695=>"100011010",
  7696=>"010010100",
  7697=>"000000010",
  7698=>"001100011",
  7699=>"100110001",
  7700=>"011110001",
  7701=>"100011001",
  7702=>"110111010",
  7703=>"010000110",
  7704=>"111100011",
  7705=>"001110001",
  7706=>"100011110",
  7707=>"001000100",
  7708=>"100100001",
  7709=>"000000010",
  7710=>"111111101",
  7711=>"111010110",
  7712=>"100100100",
  7713=>"101100100",
  7714=>"100100100",
  7715=>"100010101",
  7716=>"010110110",
  7717=>"110010111",
  7718=>"000100101",
  7719=>"100101101",
  7720=>"010110100",
  7721=>"011100110",
  7722=>"111110101",
  7723=>"100111101",
  7724=>"011011001",
  7725=>"101111100",
  7726=>"100000010",
  7727=>"010010101",
  7728=>"111011111",
  7729=>"001010000",
  7730=>"000001001",
  7731=>"100000010",
  7732=>"111001001",
  7733=>"111111111",
  7734=>"111101110",
  7735=>"111010110",
  7736=>"111001011",
  7737=>"110000010",
  7738=>"101010011",
  7739=>"011000011",
  7740=>"101100001",
  7741=>"000010010",
  7742=>"100011000",
  7743=>"000010100",
  7744=>"011110001",
  7745=>"001011101",
  7746=>"001110011",
  7747=>"010111100",
  7748=>"001011101",
  7749=>"111000001",
  7750=>"001011000",
  7751=>"101101011",
  7752=>"101010001",
  7753=>"001000101",
  7754=>"111010101",
  7755=>"101101101",
  7756=>"111010011",
  7757=>"010100001",
  7758=>"110011111",
  7759=>"110111010",
  7760=>"100001010",
  7761=>"111000110",
  7762=>"000101110",
  7763=>"000010111",
  7764=>"101110100",
  7765=>"010001011",
  7766=>"011101010",
  7767=>"000010111",
  7768=>"000011101",
  7769=>"111101011",
  7770=>"010000000",
  7771=>"101000010",
  7772=>"010000000",
  7773=>"001000010",
  7774=>"000111001",
  7775=>"000010101",
  7776=>"100101001",
  7777=>"001100111",
  7778=>"000111111",
  7779=>"101110100",
  7780=>"011111111",
  7781=>"101101100",
  7782=>"111001000",
  7783=>"011011111",
  7784=>"100001010",
  7785=>"000000001",
  7786=>"101000110",
  7787=>"011100010",
  7788=>"101000110",
  7789=>"001111010",
  7790=>"110111010",
  7791=>"101110101",
  7792=>"010010110",
  7793=>"111011011",
  7794=>"110100100",
  7795=>"110010100",
  7796=>"001101101",
  7797=>"101000111",
  7798=>"010000011",
  7799=>"010111101",
  7800=>"111111100",
  7801=>"011011000",
  7802=>"111101101",
  7803=>"011101101",
  7804=>"101001001",
  7805=>"000011010",
  7806=>"111011011",
  7807=>"111001010",
  7808=>"001011010",
  7809=>"101010010",
  7810=>"110111001",
  7811=>"001010010",
  7812=>"011110011",
  7813=>"001001000",
  7814=>"011110111",
  7815=>"010010111",
  7816=>"011111100",
  7817=>"000111000",
  7818=>"000100000",
  7819=>"000100101",
  7820=>"001010101",
  7821=>"010111111",
  7822=>"010000111",
  7823=>"101010000",
  7824=>"111010110",
  7825=>"011111101",
  7826=>"011100101",
  7827=>"000001001",
  7828=>"000111101",
  7829=>"011101110",
  7830=>"111110100",
  7831=>"011101011",
  7832=>"010111111",
  7833=>"101011100",
  7834=>"111100000",
  7835=>"001000001",
  7836=>"000010110",
  7837=>"000100010",
  7838=>"001001100",
  7839=>"011111011",
  7840=>"000111101",
  7841=>"001101011",
  7842=>"001100001",
  7843=>"100011101",
  7844=>"101100010",
  7845=>"101101010",
  7846=>"110111001",
  7847=>"011101110",
  7848=>"100010101",
  7849=>"100010101",
  7850=>"010010100",
  7851=>"111001010",
  7852=>"011100001",
  7853=>"010001001",
  7854=>"101000100",
  7855=>"001000100",
  7856=>"100110110",
  7857=>"101001010",
  7858=>"010110001",
  7859=>"011010101",
  7860=>"111010000",
  7861=>"100000010",
  7862=>"000000010",
  7863=>"010010001",
  7864=>"000100101",
  7865=>"000111010",
  7866=>"010100111",
  7867=>"011001010",
  7868=>"010010100",
  7869=>"001111001",
  7870=>"000100100",
  7871=>"110111010",
  7872=>"000000010",
  7873=>"111111111",
  7874=>"110011010",
  7875=>"011100110",
  7876=>"111111001",
  7877=>"001010000",
  7878=>"101111101",
  7879=>"110000111",
  7880=>"100000010",
  7881=>"010111000",
  7882=>"101010110",
  7883=>"010110001",
  7884=>"000110001",
  7885=>"111110100",
  7886=>"000001100",
  7887=>"000111010",
  7888=>"001110100",
  7889=>"100101011",
  7890=>"101000101",
  7891=>"001100000",
  7892=>"000000101",
  7893=>"100001110",
  7894=>"110101100",
  7895=>"000011000",
  7896=>"010000001",
  7897=>"111110110",
  7898=>"000001111",
  7899=>"111111000",
  7900=>"101110001",
  7901=>"010000011",
  7902=>"110110100",
  7903=>"010001100",
  7904=>"000100101",
  7905=>"010000001",
  7906=>"110111011",
  7907=>"111010001",
  7908=>"101010111",
  7909=>"101110110",
  7910=>"110010010",
  7911=>"001110111",
  7912=>"000101111",
  7913=>"010010110",
  7914=>"011101001",
  7915=>"011110000",
  7916=>"010101011",
  7917=>"010100010",
  7918=>"010010111",
  7919=>"101111110",
  7920=>"101001011",
  7921=>"000011111",
  7922=>"111101011",
  7923=>"001101000",
  7924=>"000011000",
  7925=>"101010111",
  7926=>"110101111",
  7927=>"001110000",
  7928=>"111101111",
  7929=>"010100110",
  7930=>"100000000",
  7931=>"100000101",
  7932=>"011100010",
  7933=>"001101110",
  7934=>"101111010",
  7935=>"111010100",
  7936=>"010101010",
  7937=>"001001001",
  7938=>"110001110",
  7939=>"110010000",
  7940=>"111110010",
  7941=>"010101010",
  7942=>"011111100",
  7943=>"100001110",
  7944=>"000101110",
  7945=>"111110111",
  7946=>"010111011",
  7947=>"111011011",
  7948=>"000000000",
  7949=>"111001000",
  7950=>"001000111",
  7951=>"000101001",
  7952=>"001111110",
  7953=>"001001000",
  7954=>"001001100",
  7955=>"100101010",
  7956=>"010100011",
  7957=>"010000011",
  7958=>"000111000",
  7959=>"111000001",
  7960=>"110110000",
  7961=>"001000110",
  7962=>"010110101",
  7963=>"111100101",
  7964=>"001000011",
  7965=>"101001100",
  7966=>"010111100",
  7967=>"001000110",
  7968=>"101101001",
  7969=>"010110001",
  7970=>"000110011",
  7971=>"010010100",
  7972=>"101010110",
  7973=>"101111000",
  7974=>"000100010",
  7975=>"000000001",
  7976=>"101100101",
  7977=>"000111110",
  7978=>"111111111",
  7979=>"000010011",
  7980=>"111010111",
  7981=>"001011000",
  7982=>"001001101",
  7983=>"111010001",
  7984=>"010000110",
  7985=>"011001011",
  7986=>"000110111",
  7987=>"011101100",
  7988=>"000111011",
  7989=>"101101001",
  7990=>"000000010",
  7991=>"010010001",
  7992=>"001110110",
  7993=>"111111000",
  7994=>"101111001",
  7995=>"110101100",
  7996=>"101010110",
  7997=>"010001001",
  7998=>"000110101",
  7999=>"101111111",
  8000=>"110000111",
  8001=>"000001110",
  8002=>"010101111",
  8003=>"111001111",
  8004=>"001011011",
  8005=>"111110001",
  8006=>"010100111",
  8007=>"010100010",
  8008=>"011010011",
  8009=>"000100010",
  8010=>"101000000",
  8011=>"111101101",
  8012=>"100110011",
  8013=>"000010110",
  8014=>"101111111",
  8015=>"100001001",
  8016=>"101011010",
  8017=>"000101001",
  8018=>"000010111",
  8019=>"000000011",
  8020=>"011110001",
  8021=>"101011011",
  8022=>"111011111",
  8023=>"000001100",
  8024=>"000011001",
  8025=>"111011111",
  8026=>"111011110",
  8027=>"110110000",
  8028=>"011100000",
  8029=>"000111011",
  8030=>"001100110",
  8031=>"001001110",
  8032=>"101001000",
  8033=>"011100010",
  8034=>"111000010",
  8035=>"100100011",
  8036=>"100110100",
  8037=>"010111100",
  8038=>"000011110",
  8039=>"001000111",
  8040=>"110110010",
  8041=>"110010000",
  8042=>"000010000",
  8043=>"010100001",
  8044=>"000000001",
  8045=>"000001110",
  8046=>"001101001",
  8047=>"001100010",
  8048=>"000011110",
  8049=>"110010001",
  8050=>"110111010",
  8051=>"011000110",
  8052=>"011010100",
  8053=>"011000011",
  8054=>"100100000",
  8055=>"110001111",
  8056=>"011100111",
  8057=>"110000001",
  8058=>"011011011",
  8059=>"010100010",
  8060=>"000010001",
  8061=>"101111101",
  8062=>"001110001",
  8063=>"011000011",
  8064=>"110001010",
  8065=>"001101001",
  8066=>"001001000",
  8067=>"001011011",
  8068=>"101001111",
  8069=>"111000011",
  8070=>"001000001",
  8071=>"110110010",
  8072=>"010010011",
  8073=>"101001111",
  8074=>"101110111",
  8075=>"101101110",
  8076=>"110000101",
  8077=>"000000111",
  8078=>"110100111",
  8079=>"110110100",
  8080=>"000101011",
  8081=>"110101000",
  8082=>"001010111",
  8083=>"111011111",
  8084=>"000111010",
  8085=>"111100110",
  8086=>"100001111",
  8087=>"101000011",
  8088=>"011111010",
  8089=>"010001001",
  8090=>"110010000",
  8091=>"011101100",
  8092=>"110111100",
  8093=>"110000111",
  8094=>"110010011",
  8095=>"000110010",
  8096=>"100100001",
  8097=>"111000101",
  8098=>"110001101",
  8099=>"101110010",
  8100=>"100110010",
  8101=>"100001111",
  8102=>"111001111",
  8103=>"001001010",
  8104=>"000101000",
  8105=>"101001001",
  8106=>"100010000",
  8107=>"000111011",
  8108=>"010111101",
  8109=>"010101011",
  8110=>"111101010",
  8111=>"101101000",
  8112=>"011010001",
  8113=>"110010010",
  8114=>"011010011",
  8115=>"111010101",
  8116=>"010111001",
  8117=>"000011011",
  8118=>"000100011",
  8119=>"001110001",
  8120=>"111010111",
  8121=>"111001011",
  8122=>"010001010",
  8123=>"110010101",
  8124=>"011101011",
  8125=>"110100010",
  8126=>"100100001",
  8127=>"010011100",
  8128=>"001100001",
  8129=>"101001000",
  8130=>"111100101",
  8131=>"000011000",
  8132=>"110001011",
  8133=>"011000111",
  8134=>"100110101",
  8135=>"000010101",
  8136=>"000000000",
  8137=>"100101111",
  8138=>"100110101",
  8139=>"100010000",
  8140=>"111010000",
  8141=>"011010101",
  8142=>"100110101",
  8143=>"100111111",
  8144=>"101111000",
  8145=>"100100100",
  8146=>"011011001",
  8147=>"010000000",
  8148=>"011111010",
  8149=>"110010010",
  8150=>"011110110",
  8151=>"000100010",
  8152=>"111111001",
  8153=>"000100000",
  8154=>"111101011",
  8155=>"001101010",
  8156=>"100110001",
  8157=>"100110110",
  8158=>"010000011",
  8159=>"000111110",
  8160=>"010100010",
  8161=>"001111101",
  8162=>"001110000",
  8163=>"010110110",
  8164=>"011100011",
  8165=>"001010101",
  8166=>"011000110",
  8167=>"110100010",
  8168=>"101101111",
  8169=>"000001111",
  8170=>"001001111",
  8171=>"000001000",
  8172=>"011100101",
  8173=>"001001111",
  8174=>"001010100",
  8175=>"010111101",
  8176=>"010000101",
  8177=>"000111010",
  8178=>"101111100",
  8179=>"110100101",
  8180=>"111000111",
  8181=>"000111111",
  8182=>"110000000",
  8183=>"110000011",
  8184=>"000100000",
  8185=>"110001000",
  8186=>"111110111",
  8187=>"001111110",
  8188=>"110000001",
  8189=>"000110001",
  8190=>"101001000",
  8191=>"101100101",
  8192=>"010000101",
  8193=>"100000111",
  8194=>"111110000",
  8195=>"111000101",
  8196=>"111100100",
  8197=>"001011110",
  8198=>"000100010",
  8199=>"111010100",
  8200=>"111000100",
  8201=>"101010110",
  8202=>"111000100",
  8203=>"001100001",
  8204=>"101110010",
  8205=>"100100001",
  8206=>"100011001",
  8207=>"111001001",
  8208=>"001010000",
  8209=>"101111010",
  8210=>"100001011",
  8211=>"010100000",
  8212=>"110011101",
  8213=>"001010000",
  8214=>"001011000",
  8215=>"110000100",
  8216=>"000011001",
  8217=>"110100100",
  8218=>"110100001",
  8219=>"100101111",
  8220=>"101011011",
  8221=>"011000001",
  8222=>"000000101",
  8223=>"110001001",
  8224=>"111110111",
  8225=>"100110100",
  8226=>"010100000",
  8227=>"101101011",
  8228=>"111111100",
  8229=>"101100001",
  8230=>"001100100",
  8231=>"000110011",
  8232=>"101010010",
  8233=>"111110111",
  8234=>"011110111",
  8235=>"010011001",
  8236=>"000111000",
  8237=>"010001110",
  8238=>"001111111",
  8239=>"110101010",
  8240=>"110000000",
  8241=>"101000000",
  8242=>"110100100",
  8243=>"001101000",
  8244=>"011011010",
  8245=>"101101110",
  8246=>"100000011",
  8247=>"110001111",
  8248=>"110011101",
  8249=>"100100000",
  8250=>"000000111",
  8251=>"001111011",
  8252=>"110111111",
  8253=>"000011100",
  8254=>"101011000",
  8255=>"110011100",
  8256=>"001100000",
  8257=>"110111001",
  8258=>"011011101",
  8259=>"010010010",
  8260=>"110111010",
  8261=>"011100111",
  8262=>"101111011",
  8263=>"111101100",
  8264=>"111011001",
  8265=>"100110000",
  8266=>"010001010",
  8267=>"011000010",
  8268=>"011101010",
  8269=>"101000010",
  8270=>"011001000",
  8271=>"011111010",
  8272=>"111010110",
  8273=>"111001011",
  8274=>"110110101",
  8275=>"001101000",
  8276=>"111111101",
  8277=>"100101111",
  8278=>"110101001",
  8279=>"100000010",
  8280=>"100100000",
  8281=>"000000000",
  8282=>"000000010",
  8283=>"000100101",
  8284=>"000110000",
  8285=>"111111010",
  8286=>"001110101",
  8287=>"000101101",
  8288=>"000101000",
  8289=>"001111000",
  8290=>"101001100",
  8291=>"000010001",
  8292=>"111010000",
  8293=>"111101010",
  8294=>"000011110",
  8295=>"000100100",
  8296=>"101001111",
  8297=>"101101100",
  8298=>"000100000",
  8299=>"110110111",
  8300=>"011011101",
  8301=>"000111111",
  8302=>"010101101",
  8303=>"001100011",
  8304=>"000010100",
  8305=>"100101111",
  8306=>"111011100",
  8307=>"100001010",
  8308=>"101010000",
  8309=>"000111010",
  8310=>"011101100",
  8311=>"001110110",
  8312=>"111001010",
  8313=>"100101100",
  8314=>"010000010",
  8315=>"110010110",
  8316=>"111101110",
  8317=>"101110001",
  8318=>"100101100",
  8319=>"110101100",
  8320=>"101110111",
  8321=>"001010110",
  8322=>"110000001",
  8323=>"101010000",
  8324=>"001001111",
  8325=>"111101000",
  8326=>"001101110",
  8327=>"101101110",
  8328=>"111001101",
  8329=>"000110111",
  8330=>"111101100",
  8331=>"011110101",
  8332=>"010101100",
  8333=>"000010110",
  8334=>"101110001",
  8335=>"111101110",
  8336=>"110000100",
  8337=>"101011100",
  8338=>"010000110",
  8339=>"110101000",
  8340=>"101101001",
  8341=>"111000001",
  8342=>"101010001",
  8343=>"010011001",
  8344=>"011111011",
  8345=>"111111011",
  8346=>"110101111",
  8347=>"110011001",
  8348=>"111110101",
  8349=>"100001010",
  8350=>"010010010",
  8351=>"010110101",
  8352=>"101110110",
  8353=>"100110011",
  8354=>"111110011",
  8355=>"000000101",
  8356=>"111010111",
  8357=>"001111011",
  8358=>"110011110",
  8359=>"100000011",
  8360=>"011011100",
  8361=>"010101010",
  8362=>"101110100",
  8363=>"010101000",
  8364=>"100010010",
  8365=>"001110011",
  8366=>"111010110",
  8367=>"011011111",
  8368=>"101001011",
  8369=>"000000000",
  8370=>"011001001",
  8371=>"101101100",
  8372=>"000110110",
  8373=>"101000111",
  8374=>"110111011",
  8375=>"000001000",
  8376=>"110010110",
  8377=>"010110000",
  8378=>"110010111",
  8379=>"000110111",
  8380=>"111111110",
  8381=>"001010001",
  8382=>"111100101",
  8383=>"001001111",
  8384=>"100101110",
  8385=>"100100111",
  8386=>"111110111",
  8387=>"011010111",
  8388=>"101100000",
  8389=>"110111111",
  8390=>"101101110",
  8391=>"111001010",
  8392=>"000010001",
  8393=>"010100011",
  8394=>"000001111",
  8395=>"111101110",
  8396=>"111100000",
  8397=>"111010010",
  8398=>"100010110",
  8399=>"101011110",
  8400=>"000111010",
  8401=>"001110101",
  8402=>"000110000",
  8403=>"011001001",
  8404=>"100011100",
  8405=>"101100110",
  8406=>"000000000",
  8407=>"010111010",
  8408=>"101000011",
  8409=>"010111101",
  8410=>"000001110",
  8411=>"101010110",
  8412=>"001000110",
  8413=>"010111101",
  8414=>"011111111",
  8415=>"011111000",
  8416=>"111010000",
  8417=>"000010111",
  8418=>"111000011",
  8419=>"101001101",
  8420=>"110111010",
  8421=>"010011001",
  8422=>"011010010",
  8423=>"111100110",
  8424=>"000110101",
  8425=>"100101110",
  8426=>"101000011",
  8427=>"101111000",
  8428=>"000000010",
  8429=>"001000100",
  8430=>"011110011",
  8431=>"010011110",
  8432=>"100100111",
  8433=>"100100000",
  8434=>"110011101",
  8435=>"100111101",
  8436=>"011100001",
  8437=>"000001001",
  8438=>"110010101",
  8439=>"010011010",
  8440=>"011000011",
  8441=>"110110101",
  8442=>"101111110",
  8443=>"110000100",
  8444=>"110111001",
  8445=>"011110101",
  8446=>"000010101",
  8447=>"110111001",
  8448=>"000011010",
  8449=>"001111011",
  8450=>"101011000",
  8451=>"111100111",
  8452=>"111001000",
  8453=>"000100100",
  8454=>"110110111",
  8455=>"011000111",
  8456=>"011111100",
  8457=>"001011110",
  8458=>"000101001",
  8459=>"100000000",
  8460=>"100100010",
  8461=>"001001100",
  8462=>"001001010",
  8463=>"011111111",
  8464=>"100100001",
  8465=>"001100001",
  8466=>"111110101",
  8467=>"111101001",
  8468=>"111001001",
  8469=>"110101001",
  8470=>"011000101",
  8471=>"101011101",
  8472=>"110001000",
  8473=>"000101000",
  8474=>"100010110",
  8475=>"110101101",
  8476=>"000011100",
  8477=>"011000011",
  8478=>"111000001",
  8479=>"000000010",
  8480=>"001111100",
  8481=>"011000100",
  8482=>"001000000",
  8483=>"111011001",
  8484=>"101010110",
  8485=>"011111010",
  8486=>"010111000",
  8487=>"000001101",
  8488=>"000010001",
  8489=>"100110111",
  8490=>"100010111",
  8491=>"011100001",
  8492=>"110101101",
  8493=>"000011010",
  8494=>"111100111",
  8495=>"010011000",
  8496=>"110010101",
  8497=>"001000001",
  8498=>"100000011",
  8499=>"011011011",
  8500=>"001001010",
  8501=>"010001010",
  8502=>"000001100",
  8503=>"000100001",
  8504=>"010010110",
  8505=>"100010100",
  8506=>"001100001",
  8507=>"101000010",
  8508=>"111010111",
  8509=>"000010010",
  8510=>"011100000",
  8511=>"100111100",
  8512=>"110001111",
  8513=>"100101010",
  8514=>"000001111",
  8515=>"111011001",
  8516=>"010111000",
  8517=>"011010110",
  8518=>"100100101",
  8519=>"110011111",
  8520=>"110111110",
  8521=>"111000000",
  8522=>"000011010",
  8523=>"010001010",
  8524=>"100100101",
  8525=>"011011100",
  8526=>"110010000",
  8527=>"100011111",
  8528=>"111000111",
  8529=>"101000100",
  8530=>"110100100",
  8531=>"101111110",
  8532=>"110111011",
  8533=>"100111010",
  8534=>"001111110",
  8535=>"010001110",
  8536=>"010010010",
  8537=>"011000100",
  8538=>"010001001",
  8539=>"010100101",
  8540=>"000001111",
  8541=>"111001011",
  8542=>"110100110",
  8543=>"010110100",
  8544=>"011011010",
  8545=>"011111001",
  8546=>"000000100",
  8547=>"110011001",
  8548=>"110100101",
  8549=>"001110110",
  8550=>"101100101",
  8551=>"100001011",
  8552=>"111010010",
  8553=>"000000111",
  8554=>"111111111",
  8555=>"101111001",
  8556=>"001101011",
  8557=>"001111110",
  8558=>"101110110",
  8559=>"010100000",
  8560=>"000011010",
  8561=>"110011000",
  8562=>"111111010",
  8563=>"001111110",
  8564=>"111101110",
  8565=>"000111101",
  8566=>"110111000",
  8567=>"100111000",
  8568=>"001010000",
  8569=>"001111010",
  8570=>"111010010",
  8571=>"100001010",
  8572=>"011111000",
  8573=>"001101100",
  8574=>"110110011",
  8575=>"110111000",
  8576=>"011000011",
  8577=>"000100100",
  8578=>"000101000",
  8579=>"111011001",
  8580=>"101111100",
  8581=>"100000101",
  8582=>"111101100",
  8583=>"110101010",
  8584=>"000000111",
  8585=>"010101111",
  8586=>"110111101",
  8587=>"000101011",
  8588=>"111110100",
  8589=>"010001010",
  8590=>"100111010",
  8591=>"010110001",
  8592=>"001001011",
  8593=>"011110000",
  8594=>"101111000",
  8595=>"001111110",
  8596=>"001010101",
  8597=>"100100000",
  8598=>"000111010",
  8599=>"100101110",
  8600=>"101100000",
  8601=>"101011101",
  8602=>"100100001",
  8603=>"111010111",
  8604=>"010110001",
  8605=>"010100101",
  8606=>"100100101",
  8607=>"100100011",
  8608=>"101001000",
  8609=>"110111111",
  8610=>"100101111",
  8611=>"001010011",
  8612=>"101101000",
  8613=>"100101011",
  8614=>"001001000",
  8615=>"010110000",
  8616=>"010110000",
  8617=>"101100000",
  8618=>"111000011",
  8619=>"000111000",
  8620=>"000101110",
  8621=>"101010110",
  8622=>"001011111",
  8623=>"011111011",
  8624=>"100001000",
  8625=>"101001100",
  8626=>"111001011",
  8627=>"000100010",
  8628=>"001101110",
  8629=>"001100000",
  8630=>"010101100",
  8631=>"001110110",
  8632=>"101100001",
  8633=>"010111100",
  8634=>"000101010",
  8635=>"110101100",
  8636=>"011010001",
  8637=>"000010010",
  8638=>"111111011",
  8639=>"110101001",
  8640=>"000011100",
  8641=>"101111001",
  8642=>"101100110",
  8643=>"100001100",
  8644=>"011000011",
  8645=>"000001111",
  8646=>"111101011",
  8647=>"110011100",
  8648=>"001110010",
  8649=>"010000011",
  8650=>"011110001",
  8651=>"010101110",
  8652=>"000101111",
  8653=>"010110001",
  8654=>"011001001",
  8655=>"111001010",
  8656=>"110011000",
  8657=>"111010010",
  8658=>"100010000",
  8659=>"000001011",
  8660=>"010101010",
  8661=>"110110001",
  8662=>"000101111",
  8663=>"001000010",
  8664=>"111001010",
  8665=>"010000011",
  8666=>"100100000",
  8667=>"000101100",
  8668=>"111111011",
  8669=>"111010100",
  8670=>"010000101",
  8671=>"000001000",
  8672=>"000000111",
  8673=>"000010101",
  8674=>"000100111",
  8675=>"001100100",
  8676=>"100101010",
  8677=>"110010000",
  8678=>"111101001",
  8679=>"010111010",
  8680=>"100001110",
  8681=>"101101111",
  8682=>"000000100",
  8683=>"101100111",
  8684=>"001111010",
  8685=>"100100111",
  8686=>"101110110",
  8687=>"101001000",
  8688=>"000000010",
  8689=>"010100000",
  8690=>"110100111",
  8691=>"001100110",
  8692=>"100011110",
  8693=>"001010011",
  8694=>"101111101",
  8695=>"111111111",
  8696=>"100100100",
  8697=>"000001011",
  8698=>"100111011",
  8699=>"110100100",
  8700=>"000111110",
  8701=>"010011011",
  8702=>"010011001",
  8703=>"001100001",
  8704=>"010000001",
  8705=>"111000000",
  8706=>"010000001",
  8707=>"001001111",
  8708=>"110110110",
  8709=>"111101001",
  8710=>"001000111",
  8711=>"010010111",
  8712=>"110010100",
  8713=>"010010001",
  8714=>"110011101",
  8715=>"111101100",
  8716=>"100101011",
  8717=>"011000000",
  8718=>"000111111",
  8719=>"110000011",
  8720=>"110000001",
  8721=>"000111010",
  8722=>"110101111",
  8723=>"011110000",
  8724=>"101011010",
  8725=>"011000100",
  8726=>"000010111",
  8727=>"010001000",
  8728=>"110001110",
  8729=>"011100101",
  8730=>"100101100",
  8731=>"101101100",
  8732=>"000101101",
  8733=>"101010010",
  8734=>"000001010",
  8735=>"010100101",
  8736=>"001011111",
  8737=>"001100001",
  8738=>"010000111",
  8739=>"000000000",
  8740=>"001000111",
  8741=>"001100011",
  8742=>"110100000",
  8743=>"010110000",
  8744=>"101001100",
  8745=>"000100010",
  8746=>"011001110",
  8747=>"100101101",
  8748=>"000101001",
  8749=>"001100011",
  8750=>"111010100",
  8751=>"011000000",
  8752=>"111011011",
  8753=>"111010011",
  8754=>"000110011",
  8755=>"110011111",
  8756=>"110000111",
  8757=>"111111111",
  8758=>"100010010",
  8759=>"000110010",
  8760=>"110011011",
  8761=>"000110001",
  8762=>"000111111",
  8763=>"011100111",
  8764=>"001000100",
  8765=>"000101001",
  8766=>"001101011",
  8767=>"101110000",
  8768=>"111111110",
  8769=>"100010011",
  8770=>"100111100",
  8771=>"111100000",
  8772=>"011000101",
  8773=>"111001010",
  8774=>"000111010",
  8775=>"000100000",
  8776=>"010000111",
  8777=>"011001101",
  8778=>"101011101",
  8779=>"010011001",
  8780=>"001011100",
  8781=>"110001001",
  8782=>"100001101",
  8783=>"001111110",
  8784=>"010010001",
  8785=>"001010100",
  8786=>"010001101",
  8787=>"011001100",
  8788=>"000101100",
  8789=>"011000101",
  8790=>"001101010",
  8791=>"010111111",
  8792=>"011000111",
  8793=>"000111110",
  8794=>"001101111",
  8795=>"000111000",
  8796=>"000101001",
  8797=>"010111011",
  8798=>"100111000",
  8799=>"001101010",
  8800=>"100110111",
  8801=>"001100001",
  8802=>"011111111",
  8803=>"011111001",
  8804=>"111001011",
  8805=>"101000110",
  8806=>"000111010",
  8807=>"010100000",
  8808=>"011001101",
  8809=>"001100101",
  8810=>"110111011",
  8811=>"010011111",
  8812=>"000011101",
  8813=>"100101111",
  8814=>"000000000",
  8815=>"010101001",
  8816=>"100111101",
  8817=>"101111101",
  8818=>"010011111",
  8819=>"001011001",
  8820=>"100110001",
  8821=>"100101110",
  8822=>"001010110",
  8823=>"101001011",
  8824=>"111010000",
  8825=>"110011011",
  8826=>"000010001",
  8827=>"110000001",
  8828=>"010011010",
  8829=>"011100110",
  8830=>"000000010",
  8831=>"101111110",
  8832=>"000101110",
  8833=>"001011110",
  8834=>"101101110",
  8835=>"000011111",
  8836=>"000001001",
  8837=>"011000100",
  8838=>"111001010",
  8839=>"011000010",
  8840=>"010000111",
  8841=>"111001110",
  8842=>"111001001",
  8843=>"010000101",
  8844=>"010101111",
  8845=>"111100010",
  8846=>"111010100",
  8847=>"010100111",
  8848=>"101000110",
  8849=>"001111011",
  8850=>"000000011",
  8851=>"010011100",
  8852=>"111001110",
  8853=>"011111000",
  8854=>"101011111",
  8855=>"111101000",
  8856=>"001010000",
  8857=>"001001001",
  8858=>"010001010",
  8859=>"101001011",
  8860=>"101111101",
  8861=>"111011110",
  8862=>"010001111",
  8863=>"101110111",
  8864=>"100001010",
  8865=>"000001110",
  8866=>"010010001",
  8867=>"011001010",
  8868=>"000100111",
  8869=>"000111101",
  8870=>"101100010",
  8871=>"010000111",
  8872=>"111000000",
  8873=>"010110011",
  8874=>"010010001",
  8875=>"011110111",
  8876=>"001001100",
  8877=>"011000100",
  8878=>"001111010",
  8879=>"101111010",
  8880=>"000110011",
  8881=>"100010011",
  8882=>"000001110",
  8883=>"100111101",
  8884=>"110001011",
  8885=>"101000010",
  8886=>"110000111",
  8887=>"000101000",
  8888=>"110100010",
  8889=>"010110000",
  8890=>"111100110",
  8891=>"110110110",
  8892=>"010101001",
  8893=>"011011001",
  8894=>"001011111",
  8895=>"110010111",
  8896=>"011010001",
  8897=>"101100110",
  8898=>"011011011",
  8899=>"100010100",
  8900=>"000001011",
  8901=>"011011010",
  8902=>"001110000",
  8903=>"000001100",
  8904=>"011010000",
  8905=>"100110100",
  8906=>"100110101",
  8907=>"111100100",
  8908=>"000011000",
  8909=>"010111100",
  8910=>"001010000",
  8911=>"111010100",
  8912=>"011100011",
  8913=>"111011000",
  8914=>"101000010",
  8915=>"000010100",
  8916=>"001100001",
  8917=>"011001101",
  8918=>"011111100",
  8919=>"101111011",
  8920=>"100101110",
  8921=>"001010110",
  8922=>"100101111",
  8923=>"000110000",
  8924=>"011010110",
  8925=>"111100000",
  8926=>"110110110",
  8927=>"110010110",
  8928=>"110111111",
  8929=>"001100110",
  8930=>"101100000",
  8931=>"100001001",
  8932=>"001001111",
  8933=>"011011000",
  8934=>"011111110",
  8935=>"010100101",
  8936=>"001001010",
  8937=>"011001100",
  8938=>"111110010",
  8939=>"011011100",
  8940=>"011100010",
  8941=>"000001111",
  8942=>"011100100",
  8943=>"011000001",
  8944=>"110101000",
  8945=>"100110010",
  8946=>"101001110",
  8947=>"110010010",
  8948=>"111010011",
  8949=>"010110010",
  8950=>"011011101",
  8951=>"000000000",
  8952=>"111010111",
  8953=>"101110111",
  8954=>"011110000",
  8955=>"110110011",
  8956=>"001001010",
  8957=>"110000001",
  8958=>"010001111",
  8959=>"001111101",
  8960=>"001010110",
  8961=>"110100000",
  8962=>"010110011",
  8963=>"001000110",
  8964=>"000100010",
  8965=>"000111110",
  8966=>"100100001",
  8967=>"100101100",
  8968=>"110101000",
  8969=>"000100110",
  8970=>"111001100",
  8971=>"101101101",
  8972=>"100000000",
  8973=>"100001110",
  8974=>"010001011",
  8975=>"010001111",
  8976=>"000110001",
  8977=>"001010100",
  8978=>"100010000",
  8979=>"010110010",
  8980=>"010110000",
  8981=>"100111001",
  8982=>"010110110",
  8983=>"011010100",
  8984=>"011001000",
  8985=>"000111101",
  8986=>"000001010",
  8987=>"100100010",
  8988=>"001010101",
  8989=>"100100111",
  8990=>"000001000",
  8991=>"010101000",
  8992=>"110100001",
  8993=>"010001100",
  8994=>"010110100",
  8995=>"010010111",
  8996=>"111001101",
  8997=>"010011101",
  8998=>"001000110",
  8999=>"001100110",
  9000=>"000010110",
  9001=>"011111100",
  9002=>"111110000",
  9003=>"111101010",
  9004=>"100111011",
  9005=>"000011010",
  9006=>"001011111",
  9007=>"000111100",
  9008=>"111111101",
  9009=>"111111101",
  9010=>"100011100",
  9011=>"001110010",
  9012=>"001100010",
  9013=>"001101000",
  9014=>"101110000",
  9015=>"111010110",
  9016=>"000101011",
  9017=>"010111100",
  9018=>"100001101",
  9019=>"010001011",
  9020=>"111010101",
  9021=>"011111111",
  9022=>"011011100",
  9023=>"000100001",
  9024=>"010101011",
  9025=>"001010001",
  9026=>"111111000",
  9027=>"110001010",
  9028=>"001010110",
  9029=>"110110110",
  9030=>"011000000",
  9031=>"000001000",
  9032=>"011100110",
  9033=>"111010100",
  9034=>"001110000",
  9035=>"100010100",
  9036=>"100100001",
  9037=>"101100110",
  9038=>"010011100",
  9039=>"010000110",
  9040=>"101111110",
  9041=>"101101010",
  9042=>"111010000",
  9043=>"110010001",
  9044=>"010011111",
  9045=>"000010001",
  9046=>"011100110",
  9047=>"100101000",
  9048=>"000110111",
  9049=>"110101010",
  9050=>"010010100",
  9051=>"011010010",
  9052=>"001010001",
  9053=>"101000011",
  9054=>"100101100",
  9055=>"010000110",
  9056=>"001011010",
  9057=>"101011010",
  9058=>"001100111",
  9059=>"110001100",
  9060=>"111101111",
  9061=>"011000011",
  9062=>"101000111",
  9063=>"101000100",
  9064=>"110010000",
  9065=>"101011111",
  9066=>"000000000",
  9067=>"000101001",
  9068=>"010001110",
  9069=>"110111101",
  9070=>"010010010",
  9071=>"111000011",
  9072=>"100001011",
  9073=>"110111100",
  9074=>"010100000",
  9075=>"111110011",
  9076=>"000100100",
  9077=>"011111001",
  9078=>"110111101",
  9079=>"011111011",
  9080=>"010100000",
  9081=>"011110111",
  9082=>"111010111",
  9083=>"101101110",
  9084=>"100001100",
  9085=>"110001011",
  9086=>"111000010",
  9087=>"011111110",
  9088=>"110001010",
  9089=>"101000010",
  9090=>"000000011",
  9091=>"110000001",
  9092=>"011101011",
  9093=>"010000011",
  9094=>"001000101",
  9095=>"011000001",
  9096=>"010001000",
  9097=>"100101000",
  9098=>"110010010",
  9099=>"111111111",
  9100=>"100100000",
  9101=>"110100011",
  9102=>"100001111",
  9103=>"110111110",
  9104=>"100011111",
  9105=>"001011001",
  9106=>"010110001",
  9107=>"100100011",
  9108=>"111101001",
  9109=>"011111010",
  9110=>"001001000",
  9111=>"000000100",
  9112=>"011010010",
  9113=>"001010011",
  9114=>"010001101",
  9115=>"011101011",
  9116=>"101001100",
  9117=>"010110100",
  9118=>"011011100",
  9119=>"010010010",
  9120=>"011010111",
  9121=>"011101011",
  9122=>"010110001",
  9123=>"111100010",
  9124=>"101111101",
  9125=>"011001011",
  9126=>"100100000",
  9127=>"011000011",
  9128=>"110000100",
  9129=>"111000010",
  9130=>"101000110",
  9131=>"000001010",
  9132=>"101100111",
  9133=>"001101000",
  9134=>"001100000",
  9135=>"001010100",
  9136=>"100101000",
  9137=>"110100110",
  9138=>"011011010",
  9139=>"100000111",
  9140=>"000111010",
  9141=>"111110000",
  9142=>"100011100",
  9143=>"011100100",
  9144=>"100110110",
  9145=>"010111010",
  9146=>"011111101",
  9147=>"000100100",
  9148=>"011001111",
  9149=>"001100011",
  9150=>"010011000",
  9151=>"100110100",
  9152=>"010001101",
  9153=>"011110010",
  9154=>"010001000",
  9155=>"110000101",
  9156=>"001000100",
  9157=>"110111010",
  9158=>"000000100",
  9159=>"101010011",
  9160=>"001100001",
  9161=>"101000000",
  9162=>"111011101",
  9163=>"110001101",
  9164=>"011101101",
  9165=>"100010110",
  9166=>"111010110",
  9167=>"111010010",
  9168=>"101101101",
  9169=>"100100001",
  9170=>"001110000",
  9171=>"101100111",
  9172=>"110010110",
  9173=>"011000110",
  9174=>"000000111",
  9175=>"011100111",
  9176=>"011100000",
  9177=>"110111111",
  9178=>"011010011",
  9179=>"001001111",
  9180=>"101110010",
  9181=>"100110000",
  9182=>"101010010",
  9183=>"100010010",
  9184=>"111010000",
  9185=>"100011100",
  9186=>"101000111",
  9187=>"010110111",
  9188=>"101001111",
  9189=>"000001111",
  9190=>"100001100",
  9191=>"110000000",
  9192=>"000100111",
  9193=>"000111101",
  9194=>"110011010",
  9195=>"111010010",
  9196=>"010110010",
  9197=>"010001010",
  9198=>"011101000",
  9199=>"000111111",
  9200=>"011010011",
  9201=>"100000110",
  9202=>"001111011",
  9203=>"100110011",
  9204=>"000000001",
  9205=>"111101001",
  9206=>"100000110",
  9207=>"101010010",
  9208=>"100110001",
  9209=>"001100011",
  9210=>"101111101",
  9211=>"110001000",
  9212=>"111110010",
  9213=>"110010100",
  9214=>"100011000",
  9215=>"110001111",
  9216=>"010111010",
  9217=>"111110110",
  9218=>"000101111",
  9219=>"000100111",
  9220=>"111001000",
  9221=>"010000001",
  9222=>"110010000",
  9223=>"110101111",
  9224=>"001001100",
  9225=>"010001011",
  9226=>"101100111",
  9227=>"000010001",
  9228=>"100011000",
  9229=>"001001100",
  9230=>"010000011",
  9231=>"011011001",
  9232=>"111001100",
  9233=>"110100101",
  9234=>"011000000",
  9235=>"100001001",
  9236=>"000011110",
  9237=>"101010111",
  9238=>"001010101",
  9239=>"100100110",
  9240=>"001110111",
  9241=>"111011001",
  9242=>"111000011",
  9243=>"010000010",
  9244=>"001001010",
  9245=>"000110110",
  9246=>"010100010",
  9247=>"000000000",
  9248=>"010010000",
  9249=>"101011000",
  9250=>"000110111",
  9251=>"010011101",
  9252=>"010011100",
  9253=>"110101111",
  9254=>"100010000",
  9255=>"100000100",
  9256=>"001110001",
  9257=>"101101111",
  9258=>"110000011",
  9259=>"001111110",
  9260=>"000110010",
  9261=>"011011110",
  9262=>"111101000",
  9263=>"110100011",
  9264=>"100010101",
  9265=>"010010100",
  9266=>"100000010",
  9267=>"100011101",
  9268=>"010111111",
  9269=>"111011100",
  9270=>"000001101",
  9271=>"101010001",
  9272=>"001010100",
  9273=>"100101011",
  9274=>"000110101",
  9275=>"110100000",
  9276=>"110010010",
  9277=>"100101101",
  9278=>"111111101",
  9279=>"110110011",
  9280=>"111011111",
  9281=>"001000000",
  9282=>"001010011",
  9283=>"011101111",
  9284=>"010011111",
  9285=>"000110010",
  9286=>"001011101",
  9287=>"100100010",
  9288=>"101000111",
  9289=>"001010110",
  9290=>"010000101",
  9291=>"100001011",
  9292=>"001001010",
  9293=>"000010101",
  9294=>"110010111",
  9295=>"000001010",
  9296=>"111000100",
  9297=>"000000000",
  9298=>"010100010",
  9299=>"011011011",
  9300=>"100101010",
  9301=>"000000000",
  9302=>"000001110",
  9303=>"111110110",
  9304=>"111100000",
  9305=>"010101100",
  9306=>"101111101",
  9307=>"001011010",
  9308=>"011000101",
  9309=>"101111101",
  9310=>"100000010",
  9311=>"011001110",
  9312=>"010110111",
  9313=>"111001011",
  9314=>"001001001",
  9315=>"101100001",
  9316=>"001000110",
  9317=>"110100010",
  9318=>"011011110",
  9319=>"001011100",
  9320=>"100010010",
  9321=>"000101001",
  9322=>"001101000",
  9323=>"101011010",
  9324=>"101101101",
  9325=>"111101010",
  9326=>"111111111",
  9327=>"001111110",
  9328=>"001101101",
  9329=>"100110111",
  9330=>"001010110",
  9331=>"101010100",
  9332=>"001110110",
  9333=>"001010101",
  9334=>"010111010",
  9335=>"001001101",
  9336=>"001000000",
  9337=>"000001110",
  9338=>"111101100",
  9339=>"100000000",
  9340=>"010101110",
  9341=>"111000101",
  9342=>"010100111",
  9343=>"000110000",
  9344=>"110111111",
  9345=>"001110001",
  9346=>"000000000",
  9347=>"010110101",
  9348=>"011010011",
  9349=>"110000001",
  9350=>"110100101",
  9351=>"011001111",
  9352=>"010000111",
  9353=>"010110001",
  9354=>"001101101",
  9355=>"111110001",
  9356=>"111111010",
  9357=>"111001001",
  9358=>"100111000",
  9359=>"111110010",
  9360=>"111100010",
  9361=>"111111100",
  9362=>"011001100",
  9363=>"001000001",
  9364=>"111001111",
  9365=>"001101100",
  9366=>"111110110",
  9367=>"001010111",
  9368=>"111000010",
  9369=>"110010001",
  9370=>"001101011",
  9371=>"000101001",
  9372=>"001100010",
  9373=>"011101111",
  9374=>"111101011",
  9375=>"100101111",
  9376=>"011111111",
  9377=>"000010110",
  9378=>"010011001",
  9379=>"101110100",
  9380=>"011100011",
  9381=>"000110101",
  9382=>"010101000",
  9383=>"000100010",
  9384=>"100101010",
  9385=>"001000001",
  9386=>"100110001",
  9387=>"010110101",
  9388=>"111101101",
  9389=>"101100001",
  9390=>"100000000",
  9391=>"111101011",
  9392=>"101101111",
  9393=>"101100010",
  9394=>"010110001",
  9395=>"000100110",
  9396=>"000001000",
  9397=>"001101000",
  9398=>"111111011",
  9399=>"111000011",
  9400=>"010001010",
  9401=>"100000010",
  9402=>"010010111",
  9403=>"100000010",
  9404=>"110110110",
  9405=>"000011010",
  9406=>"001110101",
  9407=>"110000011",
  9408=>"011111110",
  9409=>"101001101",
  9410=>"100000000",
  9411=>"110100111",
  9412=>"011111110",
  9413=>"110010110",
  9414=>"111000100",
  9415=>"110101110",
  9416=>"011000111",
  9417=>"001100011",
  9418=>"110010000",
  9419=>"010001001",
  9420=>"100001011",
  9421=>"000000001",
  9422=>"100101011",
  9423=>"110100110",
  9424=>"110001111",
  9425=>"111011000",
  9426=>"000001110",
  9427=>"111000100",
  9428=>"001101000",
  9429=>"010101101",
  9430=>"111011000",
  9431=>"011000010",
  9432=>"000010000",
  9433=>"010101111",
  9434=>"111101001",
  9435=>"001100011",
  9436=>"101000000",
  9437=>"000111000",
  9438=>"011101010",
  9439=>"111110011",
  9440=>"001110111",
  9441=>"000000110",
  9442=>"100010100",
  9443=>"000101001",
  9444=>"101011111",
  9445=>"110010010",
  9446=>"010110011",
  9447=>"110100110",
  9448=>"100011001",
  9449=>"101110110",
  9450=>"011111100",
  9451=>"011011011",
  9452=>"001000100",
  9453=>"001101100",
  9454=>"000110011",
  9455=>"001100110",
  9456=>"101111110",
  9457=>"101000011",
  9458=>"111100011",
  9459=>"010101101",
  9460=>"010101011",
  9461=>"000110001",
  9462=>"011111010",
  9463=>"000010011",
  9464=>"000111111",
  9465=>"001100100",
  9466=>"101010010",
  9467=>"101001110",
  9468=>"110101011",
  9469=>"011110011",
  9470=>"101110101",
  9471=>"001111001",
  9472=>"111111101",
  9473=>"110010011",
  9474=>"001111011",
  9475=>"111000111",
  9476=>"100010001",
  9477=>"000010000",
  9478=>"000010101",
  9479=>"001010010",
  9480=>"000101010",
  9481=>"001111011",
  9482=>"110010111",
  9483=>"111000000",
  9484=>"100010001",
  9485=>"000001000",
  9486=>"101000001",
  9487=>"111110011",
  9488=>"101001100",
  9489=>"111100111",
  9490=>"011000001",
  9491=>"001110110",
  9492=>"111011011",
  9493=>"000100110",
  9494=>"011111111",
  9495=>"100001011",
  9496=>"110001100",
  9497=>"110010110",
  9498=>"110001110",
  9499=>"110100010",
  9500=>"010110100",
  9501=>"011110001",
  9502=>"011110101",
  9503=>"101111000",
  9504=>"000011000",
  9505=>"100100011",
  9506=>"101000000",
  9507=>"111011100",
  9508=>"010001110",
  9509=>"100011001",
  9510=>"110001110",
  9511=>"101110101",
  9512=>"111101101",
  9513=>"001000111",
  9514=>"000011000",
  9515=>"010001100",
  9516=>"101010101",
  9517=>"110111001",
  9518=>"001111110",
  9519=>"001111001",
  9520=>"011111001",
  9521=>"010011000",
  9522=>"000010100",
  9523=>"111010010",
  9524=>"011001001",
  9525=>"100010010",
  9526=>"011101011",
  9527=>"110100000",
  9528=>"011100011",
  9529=>"101001010",
  9530=>"001001011",
  9531=>"001000001",
  9532=>"111111111",
  9533=>"101110111",
  9534=>"000001000",
  9535=>"111011100",
  9536=>"001001001",
  9537=>"110011000",
  9538=>"100010001",
  9539=>"011000001",
  9540=>"001100000",
  9541=>"100100100",
  9542=>"001101100",
  9543=>"100010111",
  9544=>"000000010",
  9545=>"011000000",
  9546=>"111110111",
  9547=>"110011111",
  9548=>"100000011",
  9549=>"010110001",
  9550=>"001010010",
  9551=>"011110011",
  9552=>"011001010",
  9553=>"011010101",
  9554=>"111011010",
  9555=>"011001110",
  9556=>"011000000",
  9557=>"010010011",
  9558=>"110101101",
  9559=>"101100100",
  9560=>"000010010",
  9561=>"110110000",
  9562=>"001001100",
  9563=>"110010000",
  9564=>"001011000",
  9565=>"001110001",
  9566=>"111001001",
  9567=>"111101001",
  9568=>"010101100",
  9569=>"100000000",
  9570=>"110101110",
  9571=>"000010010",
  9572=>"110001010",
  9573=>"111010011",
  9574=>"010000101",
  9575=>"101000000",
  9576=>"010011101",
  9577=>"100011010",
  9578=>"110001101",
  9579=>"010110100",
  9580=>"010010111",
  9581=>"010011110",
  9582=>"101001101",
  9583=>"111011010",
  9584=>"100001110",
  9585=>"111000101",
  9586=>"001001100",
  9587=>"100011001",
  9588=>"111010110",
  9589=>"111001001",
  9590=>"000010111",
  9591=>"010010111",
  9592=>"110000110",
  9593=>"000100110",
  9594=>"100100110",
  9595=>"100101100",
  9596=>"110000011",
  9597=>"100000011",
  9598=>"010110101",
  9599=>"001001101",
  9600=>"011110010",
  9601=>"000000001",
  9602=>"110000001",
  9603=>"100101000",
  9604=>"100010111",
  9605=>"111101011",
  9606=>"110010001",
  9607=>"001111011",
  9608=>"100000100",
  9609=>"000100001",
  9610=>"110010111",
  9611=>"001000111",
  9612=>"100101101",
  9613=>"100010100",
  9614=>"111110101",
  9615=>"000010100",
  9616=>"101010000",
  9617=>"100100011",
  9618=>"110000000",
  9619=>"001001011",
  9620=>"000010111",
  9621=>"110000110",
  9622=>"110011110",
  9623=>"110101110",
  9624=>"011111101",
  9625=>"111010110",
  9626=>"011111000",
  9627=>"101110100",
  9628=>"000010110",
  9629=>"111101111",
  9630=>"011010001",
  9631=>"001101011",
  9632=>"000010110",
  9633=>"111001110",
  9634=>"110000001",
  9635=>"101001110",
  9636=>"111101101",
  9637=>"000100011",
  9638=>"110101011",
  9639=>"000000000",
  9640=>"110101001",
  9641=>"000010001",
  9642=>"000111010",
  9643=>"000010011",
  9644=>"010001111",
  9645=>"011111010",
  9646=>"000000000",
  9647=>"001111001",
  9648=>"100000000",
  9649=>"000000101",
  9650=>"011001010",
  9651=>"000001111",
  9652=>"011010100",
  9653=>"111110100",
  9654=>"100101001",
  9655=>"000100111",
  9656=>"101011111",
  9657=>"000101010",
  9658=>"101111111",
  9659=>"100100100",
  9660=>"001111011",
  9661=>"011010001",
  9662=>"001000000",
  9663=>"111101101",
  9664=>"000000101",
  9665=>"010111011",
  9666=>"001111001",
  9667=>"011000001",
  9668=>"000001110",
  9669=>"000010111",
  9670=>"110100100",
  9671=>"101100111",
  9672=>"110110011",
  9673=>"010101111",
  9674=>"110000000",
  9675=>"100111100",
  9676=>"111111101",
  9677=>"101100101",
  9678=>"011111100",
  9679=>"010011000",
  9680=>"101101110",
  9681=>"011010000",
  9682=>"001101110",
  9683=>"001100010",
  9684=>"011011111",
  9685=>"011101010",
  9686=>"101011101",
  9687=>"001011010",
  9688=>"111001001",
  9689=>"011001011",
  9690=>"011010001",
  9691=>"001101010",
  9692=>"011010101",
  9693=>"010000011",
  9694=>"010001011",
  9695=>"000101001",
  9696=>"011000111",
  9697=>"110110100",
  9698=>"001111100",
  9699=>"100110010",
  9700=>"001101110",
  9701=>"111010101",
  9702=>"101100111",
  9703=>"111000110",
  9704=>"110011110",
  9705=>"011110100",
  9706=>"100001000",
  9707=>"100011001",
  9708=>"001101100",
  9709=>"111001000",
  9710=>"011001001",
  9711=>"011000110",
  9712=>"000100001",
  9713=>"000010101",
  9714=>"101010010",
  9715=>"010110011",
  9716=>"110011101",
  9717=>"011000111",
  9718=>"010101101",
  9719=>"010000000",
  9720=>"000110111",
  9721=>"110010011",
  9722=>"001111011",
  9723=>"010001110",
  9724=>"100011001",
  9725=>"000010110",
  9726=>"001010000",
  9727=>"010111111",
  9728=>"011100001",
  9729=>"100111011",
  9730=>"101011100",
  9731=>"100000001",
  9732=>"010001010",
  9733=>"000111100",
  9734=>"000001110",
  9735=>"011000110",
  9736=>"110100000",
  9737=>"111110000",
  9738=>"101001110",
  9739=>"111001101",
  9740=>"101010100",
  9741=>"111011110",
  9742=>"101101011",
  9743=>"100100000",
  9744=>"101110011",
  9745=>"110111100",
  9746=>"011010100",
  9747=>"001010110",
  9748=>"010110011",
  9749=>"010000001",
  9750=>"001100010",
  9751=>"101111010",
  9752=>"000001001",
  9753=>"000010000",
  9754=>"001010010",
  9755=>"111001001",
  9756=>"010001000",
  9757=>"000100110",
  9758=>"011011110",
  9759=>"101010110",
  9760=>"011001100",
  9761=>"000000001",
  9762=>"101011100",
  9763=>"111010101",
  9764=>"110000100",
  9765=>"111000010",
  9766=>"000100011",
  9767=>"110001110",
  9768=>"000110001",
  9769=>"110111000",
  9770=>"001011000",
  9771=>"011000000",
  9772=>"010000001",
  9773=>"010010010",
  9774=>"000110011",
  9775=>"100111010",
  9776=>"001010010",
  9777=>"111011100",
  9778=>"000000000",
  9779=>"000001011",
  9780=>"110110011",
  9781=>"100010001",
  9782=>"101000110",
  9783=>"011000010",
  9784=>"011110111",
  9785=>"011110100",
  9786=>"000111010",
  9787=>"100101000",
  9788=>"100000000",
  9789=>"000100010",
  9790=>"010010011",
  9791=>"001110011",
  9792=>"011000100",
  9793=>"001001101",
  9794=>"110011011",
  9795=>"010001110",
  9796=>"100010101",
  9797=>"110011101",
  9798=>"110010111",
  9799=>"001001111",
  9800=>"000101101",
  9801=>"100011000",
  9802=>"111011100",
  9803=>"111100110",
  9804=>"101010010",
  9805=>"000001111",
  9806=>"111001100",
  9807=>"011010000",
  9808=>"110110001",
  9809=>"000101100",
  9810=>"000100110",
  9811=>"000011010",
  9812=>"101001101",
  9813=>"010010110",
  9814=>"000000000",
  9815=>"010110010",
  9816=>"011001000",
  9817=>"111011000",
  9818=>"010110101",
  9819=>"100111000",
  9820=>"010100000",
  9821=>"000010101",
  9822=>"100101101",
  9823=>"101010111",
  9824=>"001110111",
  9825=>"111110101",
  9826=>"001000101",
  9827=>"001101010",
  9828=>"000000111",
  9829=>"010110110",
  9830=>"111010100",
  9831=>"111100001",
  9832=>"000101011",
  9833=>"001000110",
  9834=>"001001001",
  9835=>"101001100",
  9836=>"001010000",
  9837=>"110111001",
  9838=>"101010000",
  9839=>"010001010",
  9840=>"100111101",
  9841=>"101010000",
  9842=>"000101010",
  9843=>"110000001",
  9844=>"001010100",
  9845=>"000010000",
  9846=>"000100110",
  9847=>"001110111",
  9848=>"011000100",
  9849=>"011001110",
  9850=>"110001010",
  9851=>"010000100",
  9852=>"011100111",
  9853=>"100000000",
  9854=>"100110010",
  9855=>"000010101",
  9856=>"000101011",
  9857=>"110111010",
  9858=>"111010000",
  9859=>"001011000",
  9860=>"010000001",
  9861=>"110101011",
  9862=>"111100011",
  9863=>"010010111",
  9864=>"010001101",
  9865=>"110011010",
  9866=>"011110111",
  9867=>"110001010",
  9868=>"011000100",
  9869=>"000100000",
  9870=>"000000010",
  9871=>"000101001",
  9872=>"010000110",
  9873=>"000011011",
  9874=>"000100111",
  9875=>"111011000",
  9876=>"000000110",
  9877=>"000000000",
  9878=>"001011011",
  9879=>"111011000",
  9880=>"110100101",
  9881=>"011001001",
  9882=>"111001100",
  9883=>"111001110",
  9884=>"110010001",
  9885=>"001110111",
  9886=>"011111100",
  9887=>"011111001",
  9888=>"001111101",
  9889=>"010010010",
  9890=>"000010001",
  9891=>"001101000",
  9892=>"010101001",
  9893=>"010001101",
  9894=>"110010111",
  9895=>"100000010",
  9896=>"111000111",
  9897=>"100001101",
  9898=>"001001001",
  9899=>"110010100",
  9900=>"011111101",
  9901=>"110011100",
  9902=>"000110000",
  9903=>"010110111",
  9904=>"101111001",
  9905=>"011100100",
  9906=>"000010001",
  9907=>"010011000",
  9908=>"111110101",
  9909=>"101000010",
  9910=>"100011111",
  9911=>"110111010",
  9912=>"101111000",
  9913=>"101111100",
  9914=>"100111000",
  9915=>"011110100",
  9916=>"010111011",
  9917=>"001101110",
  9918=>"001010000",
  9919=>"010000011",
  9920=>"110101110",
  9921=>"000101101",
  9922=>"000000100",
  9923=>"111001000",
  9924=>"101010101",
  9925=>"101000110",
  9926=>"101100011",
  9927=>"010011000",
  9928=>"110110011",
  9929=>"001100010",
  9930=>"101100110",
  9931=>"010100111",
  9932=>"001110100",
  9933=>"101111100",
  9934=>"001111001",
  9935=>"101000100",
  9936=>"111111110",
  9937=>"101110101",
  9938=>"011010011",
  9939=>"000100000",
  9940=>"101010011",
  9941=>"010111000",
  9942=>"000001100",
  9943=>"011101010",
  9944=>"110001111",
  9945=>"101001100",
  9946=>"010101010",
  9947=>"111000000",
  9948=>"000111011",
  9949=>"111011110",
  9950=>"111111011",
  9951=>"000100000",
  9952=>"100101101",
  9953=>"000100111",
  9954=>"001100100",
  9955=>"101100110",
  9956=>"011010001",
  9957=>"011010011",
  9958=>"111011100",
  9959=>"100111010",
  9960=>"110000111",
  9961=>"111100011",
  9962=>"000000011",
  9963=>"110010110",
  9964=>"010000000",
  9965=>"001000011",
  9966=>"110010110",
  9967=>"100111000",
  9968=>"011111110",
  9969=>"001110011",
  9970=>"111100001",
  9971=>"000101010",
  9972=>"000000001",
  9973=>"111110010",
  9974=>"010010001",
  9975=>"010100101",
  9976=>"110111001",
  9977=>"010001100",
  9978=>"011100010",
  9979=>"010001000",
  9980=>"011101011",
  9981=>"110010100",
  9982=>"100110101",
  9983=>"100011011",
  9984=>"111110110",
  9985=>"011100111",
  9986=>"011100110",
  9987=>"100101010",
  9988=>"110010100",
  9989=>"000101100",
  9990=>"000000011",
  9991=>"000110101",
  9992=>"110001010",
  9993=>"110010000",
  9994=>"110011010",
  9995=>"010000100",
  9996=>"111110110",
  9997=>"111000000",
  9998=>"011000110",
  9999=>"101111101",
  10000=>"100110011",
  10001=>"100001011",
  10002=>"101101010",
  10003=>"101100101",
  10004=>"111101101",
  10005=>"000001011",
  10006=>"101000000",
  10007=>"010111000",
  10008=>"111110110",
  10009=>"011010100",
  10010=>"101000000",
  10011=>"111110100",
  10012=>"110000001",
  10013=>"001110101",
  10014=>"010000000",
  10015=>"100110110",
  10016=>"111101001",
  10017=>"110111100",
  10018=>"001011111",
  10019=>"100000111",
  10020=>"101100110",
  10021=>"110111000",
  10022=>"111000101",
  10023=>"000101101",
  10024=>"011001000",
  10025=>"111010110",
  10026=>"011110110",
  10027=>"111110011",
  10028=>"110011110",
  10029=>"010011011",
  10030=>"001000010",
  10031=>"101111001",
  10032=>"100001011",
  10033=>"001010010",
  10034=>"000100100",
  10035=>"100011101",
  10036=>"000011000",
  10037=>"000110101",
  10038=>"011010110",
  10039=>"000111001",
  10040=>"001001011",
  10041=>"010011010",
  10042=>"010110001",
  10043=>"011010000",
  10044=>"000000011",
  10045=>"011010000",
  10046=>"100100101",
  10047=>"101000110",
  10048=>"111100100",
  10049=>"000001100",
  10050=>"111011000",
  10051=>"010111001",
  10052=>"010100001",
  10053=>"001111001",
  10054=>"100010001",
  10055=>"000011000",
  10056=>"011111111",
  10057=>"011111000",
  10058=>"110011010",
  10059=>"010010001",
  10060=>"000100001",
  10061=>"001100010",
  10062=>"110001010",
  10063=>"000011101",
  10064=>"100111111",
  10065=>"100100101",
  10066=>"100111100",
  10067=>"000100111",
  10068=>"100001011",
  10069=>"101101011",
  10070=>"110101101",
  10071=>"011111011",
  10072=>"100000010",
  10073=>"110010110",
  10074=>"010110011",
  10075=>"110111101",
  10076=>"011110111",
  10077=>"111110010",
  10078=>"000100011",
  10079=>"000010100",
  10080=>"101000000",
  10081=>"100000000",
  10082=>"110111110",
  10083=>"001000000",
  10084=>"111110011",
  10085=>"110001010",
  10086=>"010111001",
  10087=>"000001000",
  10088=>"001100100",
  10089=>"110111000",
  10090=>"110000110",
  10091=>"100110101",
  10092=>"001010010",
  10093=>"111010100",
  10094=>"100010010",
  10095=>"000011110",
  10096=>"001001010",
  10097=>"101001001",
  10098=>"100101001",
  10099=>"101111100",
  10100=>"101000101",
  10101=>"111100010",
  10102=>"010100001",
  10103=>"000111101",
  10104=>"111010100",
  10105=>"010011101",
  10106=>"110100110",
  10107=>"100010011",
  10108=>"010111110",
  10109=>"111011001",
  10110=>"101001101",
  10111=>"101110111",
  10112=>"011111100",
  10113=>"011010111",
  10114=>"111000110",
  10115=>"111101100",
  10116=>"011100000",
  10117=>"110000101",
  10118=>"011010000",
  10119=>"110000110",
  10120=>"001010101",
  10121=>"101001000",
  10122=>"011101001",
  10123=>"111111011",
  10124=>"100001010",
  10125=>"011100011",
  10126=>"100010101",
  10127=>"010001011",
  10128=>"110100010",
  10129=>"111011010",
  10130=>"000011100",
  10131=>"001001101",
  10132=>"110000001",
  10133=>"001010100",
  10134=>"110100100",
  10135=>"111111011",
  10136=>"001010011",
  10137=>"111100011",
  10138=>"001101110",
  10139=>"111000011",
  10140=>"001010000",
  10141=>"010000100",
  10142=>"010000001",
  10143=>"111011000",
  10144=>"101011111",
  10145=>"110001110",
  10146=>"010001100",
  10147=>"111000011",
  10148=>"111111101",
  10149=>"010101100",
  10150=>"101010100",
  10151=>"001111110",
  10152=>"010000010",
  10153=>"110100010",
  10154=>"010111110",
  10155=>"100011011",
  10156=>"001000111",
  10157=>"100100001",
  10158=>"000001000",
  10159=>"010000111",
  10160=>"011111010",
  10161=>"010100001",
  10162=>"100010010",
  10163=>"000000000",
  10164=>"101100001",
  10165=>"001000101",
  10166=>"000111101",
  10167=>"001000111",
  10168=>"001011001",
  10169=>"010111011",
  10170=>"101110111",
  10171=>"101000111",
  10172=>"100110100",
  10173=>"001000011",
  10174=>"000101100",
  10175=>"000110100",
  10176=>"101001111",
  10177=>"110111011",
  10178=>"100010010",
  10179=>"001101111",
  10180=>"000100000",
  10181=>"001001001",
  10182=>"100101000",
  10183=>"111010110",
  10184=>"101101101",
  10185=>"111101011",
  10186=>"100010000",
  10187=>"001101000",
  10188=>"111110100",
  10189=>"000110000",
  10190=>"101101010",
  10191=>"000000111",
  10192=>"101011011",
  10193=>"101111000",
  10194=>"010000010",
  10195=>"000000110",
  10196=>"000110100",
  10197=>"010110100",
  10198=>"011010100",
  10199=>"110100011",
  10200=>"000100110",
  10201=>"010111111",
  10202=>"001111101",
  10203=>"111100010",
  10204=>"000111011",
  10205=>"011010001",
  10206=>"100001101",
  10207=>"011111100",
  10208=>"001111111",
  10209=>"111101010",
  10210=>"110111111",
  10211=>"101000001",
  10212=>"110010000",
  10213=>"000000000",
  10214=>"000010111",
  10215=>"011101010",
  10216=>"001001010",
  10217=>"110101101",
  10218=>"000000001",
  10219=>"100001101",
  10220=>"110100011",
  10221=>"100010101",
  10222=>"000011110",
  10223=>"010001000",
  10224=>"111100000",
  10225=>"100110111",
  10226=>"100110011",
  10227=>"001010100",
  10228=>"111101000",
  10229=>"000111011",
  10230=>"011111111",
  10231=>"000101110",
  10232=>"010110010",
  10233=>"011111110",
  10234=>"100011111",
  10235=>"001011111",
  10236=>"010011011",
  10237=>"100001101",
  10238=>"110101000",
  10239=>"011010100",
  10240=>"011110000",
  10241=>"001111111",
  10242=>"101101110",
  10243=>"101001100",
  10244=>"111111101",
  10245=>"000010111",
  10246=>"000100101",
  10247=>"010111110",
  10248=>"001001001",
  10249=>"100010010",
  10250=>"110100101",
  10251=>"111001100",
  10252=>"101000100",
  10253=>"110011100",
  10254=>"000101101",
  10255=>"010101001",
  10256=>"000100100",
  10257=>"100100110",
  10258=>"100110101",
  10259=>"110111101",
  10260=>"010001101",
  10261=>"101111011",
  10262=>"011100110",
  10263=>"000100101",
  10264=>"001010010",
  10265=>"111110111",
  10266=>"100011001",
  10267=>"010101100",
  10268=>"111011101",
  10269=>"010111011",
  10270=>"000001101",
  10271=>"010011010",
  10272=>"011111010",
  10273=>"110100111",
  10274=>"111110100",
  10275=>"101100001",
  10276=>"111110101",
  10277=>"000111101",
  10278=>"010000111",
  10279=>"101100010",
  10280=>"111011110",
  10281=>"100010110",
  10282=>"011111110",
  10283=>"111111000",
  10284=>"010011100",
  10285=>"110000111",
  10286=>"100100101",
  10287=>"000101011",
  10288=>"111001001",
  10289=>"111011110",
  10290=>"100101100",
  10291=>"110101010",
  10292=>"011110010",
  10293=>"001000101",
  10294=>"000101010",
  10295=>"110110111",
  10296=>"101010001",
  10297=>"011001100",
  10298=>"101101100",
  10299=>"010010111",
  10300=>"001101010",
  10301=>"000011101",
  10302=>"101111110",
  10303=>"110101111",
  10304=>"101101010",
  10305=>"111110111",
  10306=>"001001111",
  10307=>"010001100",
  10308=>"101000010",
  10309=>"010010001",
  10310=>"101110011",
  10311=>"111101100",
  10312=>"010101110",
  10313=>"100111000",
  10314=>"000000101",
  10315=>"000100110",
  10316=>"101100110",
  10317=>"101010111",
  10318=>"010100010",
  10319=>"010001001",
  10320=>"111100101",
  10321=>"101101101",
  10322=>"100010000",
  10323=>"101100100",
  10324=>"111101111",
  10325=>"000101001",
  10326=>"011110001",
  10327=>"001000011",
  10328=>"100111101",
  10329=>"101011010",
  10330=>"111001011",
  10331=>"111010111",
  10332=>"000101100",
  10333=>"000110000",
  10334=>"000101101",
  10335=>"111100110",
  10336=>"011101001",
  10337=>"010011010",
  10338=>"000100110",
  10339=>"000010010",
  10340=>"111110101",
  10341=>"101111010",
  10342=>"011010110",
  10343=>"001001111",
  10344=>"011110110",
  10345=>"111110000",
  10346=>"110100100",
  10347=>"100001000",
  10348=>"110101011",
  10349=>"101111110",
  10350=>"010011110",
  10351=>"011100111",
  10352=>"101011011",
  10353=>"111110001",
  10354=>"011101000",
  10355=>"100010010",
  10356=>"100011011",
  10357=>"100101010",
  10358=>"101111100",
  10359=>"000100110",
  10360=>"111101100",
  10361=>"111000011",
  10362=>"010110101",
  10363=>"010010001",
  10364=>"101111111",
  10365=>"100100111",
  10366=>"010100001",
  10367=>"000100100",
  10368=>"011010111",
  10369=>"101111101",
  10370=>"100010011",
  10371=>"101101110",
  10372=>"001000111",
  10373=>"000001010",
  10374=>"100001110",
  10375=>"011111110",
  10376=>"111000000",
  10377=>"110001110",
  10378=>"110001011",
  10379=>"011001001",
  10380=>"111010001",
  10381=>"110001111",
  10382=>"111100000",
  10383=>"111101000",
  10384=>"111010010",
  10385=>"010000110",
  10386=>"001100111",
  10387=>"100011110",
  10388=>"010101100",
  10389=>"001000000",
  10390=>"100000000",
  10391=>"001001111",
  10392=>"111111001",
  10393=>"001010100",
  10394=>"011011110",
  10395=>"101011000",
  10396=>"000100111",
  10397=>"101000000",
  10398=>"001011100",
  10399=>"010011001",
  10400=>"111101010",
  10401=>"101001101",
  10402=>"111000101",
  10403=>"011000001",
  10404=>"111111111",
  10405=>"011011011",
  10406=>"000001101",
  10407=>"000011100",
  10408=>"100010011",
  10409=>"000100101",
  10410=>"100100101",
  10411=>"101111000",
  10412=>"010110111",
  10413=>"100000011",
  10414=>"100111001",
  10415=>"101111100",
  10416=>"011110010",
  10417=>"111000101",
  10418=>"110001000",
  10419=>"101000000",
  10420=>"001111101",
  10421=>"000011100",
  10422=>"100100101",
  10423=>"001010001",
  10424=>"110010111",
  10425=>"001010110",
  10426=>"011010100",
  10427=>"000110101",
  10428=>"011100111",
  10429=>"001111111",
  10430=>"111011011",
  10431=>"111011011",
  10432=>"010011100",
  10433=>"100001101",
  10434=>"110000010",
  10435=>"111110010",
  10436=>"011110110",
  10437=>"110011000",
  10438=>"010001001",
  10439=>"111011010",
  10440=>"010100111",
  10441=>"110001010",
  10442=>"010111111",
  10443=>"010100111",
  10444=>"011101011",
  10445=>"111110111",
  10446=>"101000001",
  10447=>"111010011",
  10448=>"100001000",
  10449=>"101001100",
  10450=>"000000100",
  10451=>"110010101",
  10452=>"010101011",
  10453=>"011010100",
  10454=>"111111100",
  10455=>"011100011",
  10456=>"100000010",
  10457=>"100000111",
  10458=>"011111000",
  10459=>"110010001",
  10460=>"010000100",
  10461=>"000110111",
  10462=>"000100001",
  10463=>"100101000",
  10464=>"111011111",
  10465=>"000011101",
  10466=>"110100100",
  10467=>"101110001",
  10468=>"000111000",
  10469=>"111110100",
  10470=>"100011011",
  10471=>"101101101",
  10472=>"011000101",
  10473=>"010110101",
  10474=>"000011100",
  10475=>"110100011",
  10476=>"100110100",
  10477=>"100110110",
  10478=>"000100010",
  10479=>"001110001",
  10480=>"111101001",
  10481=>"110101110",
  10482=>"111011111",
  10483=>"010111110",
  10484=>"110001101",
  10485=>"011110000",
  10486=>"101001111",
  10487=>"110100010",
  10488=>"100110000",
  10489=>"010100011",
  10490=>"011100101",
  10491=>"100011110",
  10492=>"011111000",
  10493=>"011010101",
  10494=>"001100010",
  10495=>"011110000",
  10496=>"011000000",
  10497=>"001000100",
  10498=>"111110011",
  10499=>"100011110",
  10500=>"101010111",
  10501=>"100001101",
  10502=>"111111010",
  10503=>"100100101",
  10504=>"100001000",
  10505=>"010110011",
  10506=>"010011110",
  10507=>"101011100",
  10508=>"000000101",
  10509=>"111110101",
  10510=>"010101010",
  10511=>"000111100",
  10512=>"011010111",
  10513=>"001111001",
  10514=>"111000111",
  10515=>"100110010",
  10516=>"011011011",
  10517=>"101111001",
  10518=>"010000001",
  10519=>"111111101",
  10520=>"101001010",
  10521=>"100110000",
  10522=>"000011011",
  10523=>"001101000",
  10524=>"101000011",
  10525=>"110100110",
  10526=>"000101011",
  10527=>"000010010",
  10528=>"000000111",
  10529=>"000011101",
  10530=>"011011000",
  10531=>"100001011",
  10532=>"101000011",
  10533=>"000011111",
  10534=>"001101000",
  10535=>"010110100",
  10536=>"001110000",
  10537=>"110100001",
  10538=>"010110111",
  10539=>"100100000",
  10540=>"100100000",
  10541=>"011010001",
  10542=>"100010000",
  10543=>"101110011",
  10544=>"010110000",
  10545=>"101000101",
  10546=>"000010010",
  10547=>"010000000",
  10548=>"001111101",
  10549=>"111111100",
  10550=>"000110100",
  10551=>"010001101",
  10552=>"111101010",
  10553=>"111001010",
  10554=>"011110011",
  10555=>"011100101",
  10556=>"000100011",
  10557=>"001100100",
  10558=>"010111010",
  10559=>"110100000",
  10560=>"111010011",
  10561=>"001100100",
  10562=>"110101100",
  10563=>"000001011",
  10564=>"010100111",
  10565=>"001100110",
  10566=>"110101011",
  10567=>"101111111",
  10568=>"000101101",
  10569=>"011001001",
  10570=>"011001011",
  10571=>"111111001",
  10572=>"011011101",
  10573=>"111100011",
  10574=>"100111110",
  10575=>"101000001",
  10576=>"001011001",
  10577=>"100001011",
  10578=>"011001010",
  10579=>"010101110",
  10580=>"011101110",
  10581=>"111100101",
  10582=>"000000100",
  10583=>"011100011",
  10584=>"000000110",
  10585=>"000101100",
  10586=>"101010100",
  10587=>"101101111",
  10588=>"111111011",
  10589=>"110010011",
  10590=>"011100111",
  10591=>"010111101",
  10592=>"010010011",
  10593=>"011000111",
  10594=>"000000101",
  10595=>"000001000",
  10596=>"101111011",
  10597=>"110010101",
  10598=>"100111111",
  10599=>"000011001",
  10600=>"011001010",
  10601=>"101100101",
  10602=>"110110101",
  10603=>"000011000",
  10604=>"101000101",
  10605=>"101010101",
  10606=>"100011101",
  10607=>"001110111",
  10608=>"111111001",
  10609=>"111010101",
  10610=>"110000000",
  10611=>"110111011",
  10612=>"010100101",
  10613=>"100111100",
  10614=>"011000010",
  10615=>"001101000",
  10616=>"011111100",
  10617=>"101000100",
  10618=>"000111010",
  10619=>"010010111",
  10620=>"110110010",
  10621=>"000100001",
  10622=>"110110000",
  10623=>"011011000",
  10624=>"011100000",
  10625=>"010001101",
  10626=>"011011010",
  10627=>"001010011",
  10628=>"101101101",
  10629=>"100001010",
  10630=>"100001100",
  10631=>"010111101",
  10632=>"100010100",
  10633=>"011101100",
  10634=>"101001101",
  10635=>"010000110",
  10636=>"000111110",
  10637=>"001011100",
  10638=>"010000011",
  10639=>"110111101",
  10640=>"010110000",
  10641=>"000000110",
  10642=>"101010110",
  10643=>"100011101",
  10644=>"101011100",
  10645=>"110100101",
  10646=>"011011011",
  10647=>"000000110",
  10648=>"100001001",
  10649=>"011011100",
  10650=>"010010111",
  10651=>"110011011",
  10652=>"001101010",
  10653=>"010000010",
  10654=>"100111001",
  10655=>"111111100",
  10656=>"000101001",
  10657=>"011011000",
  10658=>"111010100",
  10659=>"110110110",
  10660=>"001011100",
  10661=>"000001001",
  10662=>"100001001",
  10663=>"111011100",
  10664=>"100011010",
  10665=>"001111100",
  10666=>"110101011",
  10667=>"110000001",
  10668=>"000100011",
  10669=>"001000100",
  10670=>"101101101",
  10671=>"111010001",
  10672=>"110010101",
  10673=>"011100100",
  10674=>"110000010",
  10675=>"001100101",
  10676=>"000011110",
  10677=>"101011111",
  10678=>"101010100",
  10679=>"101100100",
  10680=>"101001001",
  10681=>"010011110",
  10682=>"100001010",
  10683=>"011011101",
  10684=>"101001011",
  10685=>"111110011",
  10686=>"111100010",
  10687=>"010100100",
  10688=>"110001000",
  10689=>"111111011",
  10690=>"000101111",
  10691=>"110001011",
  10692=>"001000010",
  10693=>"111101011",
  10694=>"111100001",
  10695=>"011110001",
  10696=>"100110110",
  10697=>"010011010",
  10698=>"011011000",
  10699=>"011101001",
  10700=>"010100011",
  10701=>"010100001",
  10702=>"110010111",
  10703=>"010100000",
  10704=>"001011101",
  10705=>"100111110",
  10706=>"011011011",
  10707=>"000100110",
  10708=>"000010001",
  10709=>"101000010",
  10710=>"011001000",
  10711=>"001000110",
  10712=>"100111001",
  10713=>"100110111",
  10714=>"111101111",
  10715=>"100100010",
  10716=>"110101000",
  10717=>"111001001",
  10718=>"001110111",
  10719=>"001001100",
  10720=>"110101100",
  10721=>"011011001",
  10722=>"110111011",
  10723=>"001000100",
  10724=>"100011101",
  10725=>"000100001",
  10726=>"110001010",
  10727=>"011001000",
  10728=>"101001000",
  10729=>"000101011",
  10730=>"010011100",
  10731=>"111101000",
  10732=>"000101101",
  10733=>"110000010",
  10734=>"010111100",
  10735=>"010011001",
  10736=>"001010111",
  10737=>"001000001",
  10738=>"011010101",
  10739=>"110010001",
  10740=>"111011101",
  10741=>"111000010",
  10742=>"001010000",
  10743=>"000010000",
  10744=>"111110000",
  10745=>"111000000",
  10746=>"000111001",
  10747=>"101101111",
  10748=>"101011001",
  10749=>"001010100",
  10750=>"011001001",
  10751=>"111011011",
  10752=>"000100110",
  10753=>"101011111",
  10754=>"110110000",
  10755=>"010110001",
  10756=>"110111100",
  10757=>"000000011",
  10758=>"100100101",
  10759=>"100010110",
  10760=>"000001101",
  10761=>"110101000",
  10762=>"000101011",
  10763=>"000110011",
  10764=>"110111000",
  10765=>"001011111",
  10766=>"110001110",
  10767=>"010111100",
  10768=>"011100100",
  10769=>"001001111",
  10770=>"101100010",
  10771=>"111001001",
  10772=>"110110000",
  10773=>"000010110",
  10774=>"000010000",
  10775=>"110111101",
  10776=>"010100100",
  10777=>"010110000",
  10778=>"011000010",
  10779=>"111011111",
  10780=>"101001010",
  10781=>"101100011",
  10782=>"101110100",
  10783=>"011111110",
  10784=>"010100110",
  10785=>"100110111",
  10786=>"000001100",
  10787=>"011110111",
  10788=>"001101010",
  10789=>"111111110",
  10790=>"011000010",
  10791=>"101010000",
  10792=>"100001111",
  10793=>"110101000",
  10794=>"011100111",
  10795=>"111000001",
  10796=>"000110010",
  10797=>"011000101",
  10798=>"000000101",
  10799=>"010100010",
  10800=>"001101011",
  10801=>"110011111",
  10802=>"110100100",
  10803=>"000010101",
  10804=>"011000011",
  10805=>"111001111",
  10806=>"101010010",
  10807=>"111111010",
  10808=>"001001111",
  10809=>"111000011",
  10810=>"010111101",
  10811=>"011000000",
  10812=>"101110101",
  10813=>"100110110",
  10814=>"100110010",
  10815=>"001100011",
  10816=>"110101000",
  10817=>"110011000",
  10818=>"011110000",
  10819=>"010011100",
  10820=>"000010100",
  10821=>"010100010",
  10822=>"101110001",
  10823=>"010111001",
  10824=>"000111011",
  10825=>"001011110",
  10826=>"000110001",
  10827=>"100010101",
  10828=>"000011011",
  10829=>"101000111",
  10830=>"111110100",
  10831=>"111011111",
  10832=>"100010001",
  10833=>"010010011",
  10834=>"001001010",
  10835=>"000100010",
  10836=>"010000000",
  10837=>"001111100",
  10838=>"100001100",
  10839=>"001100011",
  10840=>"111100111",
  10841=>"110110011",
  10842=>"001011100",
  10843=>"001011011",
  10844=>"001010000",
  10845=>"110111111",
  10846=>"001000010",
  10847=>"001110100",
  10848=>"000100111",
  10849=>"101000001",
  10850=>"100111101",
  10851=>"001000101",
  10852=>"010010010",
  10853=>"110111010",
  10854=>"011011110",
  10855=>"101111010",
  10856=>"100010010",
  10857=>"010001000",
  10858=>"001011111",
  10859=>"010010111",
  10860=>"100000010",
  10861=>"110000100",
  10862=>"111011100",
  10863=>"001101100",
  10864=>"001001101",
  10865=>"000010101",
  10866=>"010010010",
  10867=>"101000111",
  10868=>"111110001",
  10869=>"011001001",
  10870=>"111001001",
  10871=>"001100110",
  10872=>"110101100",
  10873=>"011111000",
  10874=>"101100000",
  10875=>"111111101",
  10876=>"110101111",
  10877=>"001101010",
  10878=>"101101010",
  10879=>"011101101",
  10880=>"110000011",
  10881=>"001011100",
  10882=>"011110001",
  10883=>"100011101",
  10884=>"000101111",
  10885=>"011000010",
  10886=>"101000000",
  10887=>"000111101",
  10888=>"010101110",
  10889=>"001000000",
  10890=>"101101100",
  10891=>"111001011",
  10892=>"010011110",
  10893=>"101111000",
  10894=>"000000000",
  10895=>"100111001",
  10896=>"001001010",
  10897=>"001001110",
  10898=>"011011110",
  10899=>"110111101",
  10900=>"101101111",
  10901=>"010010000",
  10902=>"110001011",
  10903=>"101100001",
  10904=>"011110000",
  10905=>"000101101",
  10906=>"000000000",
  10907=>"010001101",
  10908=>"011010110",
  10909=>"001010111",
  10910=>"111110001",
  10911=>"110100000",
  10912=>"111001100",
  10913=>"011110000",
  10914=>"100110100",
  10915=>"111000101",
  10916=>"001101100",
  10917=>"001000111",
  10918=>"000001110",
  10919=>"001010100",
  10920=>"110010100",
  10921=>"000100101",
  10922=>"000010000",
  10923=>"011110010",
  10924=>"101001001",
  10925=>"100111101",
  10926=>"011111010",
  10927=>"111100011",
  10928=>"010110001",
  10929=>"100011101",
  10930=>"111111110",
  10931=>"001001010",
  10932=>"101010001",
  10933=>"000101101",
  10934=>"101101101",
  10935=>"001001001",
  10936=>"011011100",
  10937=>"101001101",
  10938=>"110001011",
  10939=>"110100011",
  10940=>"000011111",
  10941=>"010011010",
  10942=>"101001111",
  10943=>"110100011",
  10944=>"101111100",
  10945=>"100100010",
  10946=>"110010000",
  10947=>"000001101",
  10948=>"111111000",
  10949=>"000100111",
  10950=>"000011100",
  10951=>"100010010",
  10952=>"011010110",
  10953=>"110010000",
  10954=>"010010001",
  10955=>"000101001",
  10956=>"010100110",
  10957=>"100101001",
  10958=>"001011001",
  10959=>"010000111",
  10960=>"110110110",
  10961=>"111111001",
  10962=>"011111001",
  10963=>"010111001",
  10964=>"100001111",
  10965=>"101000000",
  10966=>"100001101",
  10967=>"011100011",
  10968=>"100101000",
  10969=>"110100001",
  10970=>"010101100",
  10971=>"001100010",
  10972=>"001001111",
  10973=>"110001010",
  10974=>"000000000",
  10975=>"010110001",
  10976=>"111100110",
  10977=>"100101110",
  10978=>"010100111",
  10979=>"100101010",
  10980=>"110000010",
  10981=>"111111001",
  10982=>"010011001",
  10983=>"001010111",
  10984=>"100010101",
  10985=>"100110011",
  10986=>"011110101",
  10987=>"011110011",
  10988=>"010011000",
  10989=>"101111000",
  10990=>"101100010",
  10991=>"110111100",
  10992=>"111101010",
  10993=>"101111101",
  10994=>"010000010",
  10995=>"010101110",
  10996=>"111010110",
  10997=>"101100111",
  10998=>"111000000",
  10999=>"010000011",
  11000=>"010100011",
  11001=>"110010110",
  11002=>"111011111",
  11003=>"101010101",
  11004=>"000011000",
  11005=>"111101110",
  11006=>"001011000",
  11007=>"000111011",
  11008=>"001110111",
  11009=>"011000110",
  11010=>"001111010",
  11011=>"100100000",
  11012=>"110101001",
  11013=>"110100010",
  11014=>"110010001",
  11015=>"111101111",
  11016=>"101011001",
  11017=>"010000010",
  11018=>"101111110",
  11019=>"001111101",
  11020=>"101000101",
  11021=>"111011100",
  11022=>"111000100",
  11023=>"101011011",
  11024=>"101000111",
  11025=>"000110111",
  11026=>"111001001",
  11027=>"010101101",
  11028=>"100110001",
  11029=>"110011111",
  11030=>"100110110",
  11031=>"101001101",
  11032=>"111001101",
  11033=>"100101010",
  11034=>"010000111",
  11035=>"101010000",
  11036=>"100111010",
  11037=>"111011100",
  11038=>"100011101",
  11039=>"100000010",
  11040=>"011011010",
  11041=>"000010100",
  11042=>"011011010",
  11043=>"000110111",
  11044=>"001000111",
  11045=>"001101001",
  11046=>"000001100",
  11047=>"110101111",
  11048=>"100110001",
  11049=>"111000100",
  11050=>"010110010",
  11051=>"111000111",
  11052=>"100111000",
  11053=>"010100010",
  11054=>"011100110",
  11055=>"100101011",
  11056=>"111001111",
  11057=>"110100101",
  11058=>"110011000",
  11059=>"011111001",
  11060=>"100000110",
  11061=>"100100101",
  11062=>"010010110",
  11063=>"110111000",
  11064=>"000101011",
  11065=>"000000101",
  11066=>"001001101",
  11067=>"101111111",
  11068=>"010101000",
  11069=>"000000111",
  11070=>"000101011",
  11071=>"010010010",
  11072=>"011000110",
  11073=>"000010001",
  11074=>"101010100",
  11075=>"011001000",
  11076=>"101100111",
  11077=>"101011110",
  11078=>"001001011",
  11079=>"100110011",
  11080=>"110000101",
  11081=>"100101010",
  11082=>"110111111",
  11083=>"000110000",
  11084=>"101010111",
  11085=>"100001011",
  11086=>"101001101",
  11087=>"111001100",
  11088=>"110000100",
  11089=>"001100101",
  11090=>"100001001",
  11091=>"000000111",
  11092=>"101010010",
  11093=>"011010000",
  11094=>"100000011",
  11095=>"000000110",
  11096=>"100011110",
  11097=>"000000011",
  11098=>"001100011",
  11099=>"111001000",
  11100=>"100000000",
  11101=>"100001001",
  11102=>"001100100",
  11103=>"000000101",
  11104=>"000000011",
  11105=>"101100000",
  11106=>"101101011",
  11107=>"110010101",
  11108=>"100000001",
  11109=>"110000111",
  11110=>"010110110",
  11111=>"100111111",
  11112=>"010000001",
  11113=>"111001110",
  11114=>"101100111",
  11115=>"011000000",
  11116=>"110000000",
  11117=>"000010000",
  11118=>"100000000",
  11119=>"001001110",
  11120=>"111011011",
  11121=>"100110001",
  11122=>"001101011",
  11123=>"100001100",
  11124=>"100000001",
  11125=>"011110110",
  11126=>"001110010",
  11127=>"110000000",
  11128=>"011011101",
  11129=>"100000000",
  11130=>"000101101",
  11131=>"000011010",
  11132=>"010111000",
  11133=>"000110101",
  11134=>"110101110",
  11135=>"110100101",
  11136=>"001010001",
  11137=>"101011110",
  11138=>"001010110",
  11139=>"100001011",
  11140=>"001010001",
  11141=>"011001001",
  11142=>"001111001",
  11143=>"001111110",
  11144=>"101101001",
  11145=>"000000111",
  11146=>"001010001",
  11147=>"101011111",
  11148=>"100101110",
  11149=>"010100111",
  11150=>"010000010",
  11151=>"110100011",
  11152=>"110011011",
  11153=>"010010001",
  11154=>"100000011",
  11155=>"101010010",
  11156=>"001011111",
  11157=>"101001001",
  11158=>"111101011",
  11159=>"111101000",
  11160=>"010110000",
  11161=>"001100110",
  11162=>"001011101",
  11163=>"110100111",
  11164=>"001000110",
  11165=>"000010111",
  11166=>"100010110",
  11167=>"110110100",
  11168=>"100001000",
  11169=>"100110100",
  11170=>"000011011",
  11171=>"001101010",
  11172=>"000011011",
  11173=>"110010010",
  11174=>"001110100",
  11175=>"001101001",
  11176=>"100010100",
  11177=>"101110100",
  11178=>"111100000",
  11179=>"001011111",
  11180=>"001000001",
  11181=>"011101000",
  11182=>"110010000",
  11183=>"001100100",
  11184=>"100000101",
  11185=>"110101101",
  11186=>"010000011",
  11187=>"011110001",
  11188=>"111000001",
  11189=>"000000010",
  11190=>"110111101",
  11191=>"101010100",
  11192=>"000010011",
  11193=>"101100111",
  11194=>"101000110",
  11195=>"000101111",
  11196=>"111000000",
  11197=>"000010010",
  11198=>"110111101",
  11199=>"110010111",
  11200=>"011100101",
  11201=>"011100110",
  11202=>"011011111",
  11203=>"110011101",
  11204=>"110000010",
  11205=>"110010111",
  11206=>"101001011",
  11207=>"001111001",
  11208=>"001100111",
  11209=>"011101110",
  11210=>"001101101",
  11211=>"011010111",
  11212=>"101010011",
  11213=>"000000100",
  11214=>"110011101",
  11215=>"110011100",
  11216=>"011110001",
  11217=>"000100000",
  11218=>"010101000",
  11219=>"101010110",
  11220=>"111001101",
  11221=>"100001000",
  11222=>"101001001",
  11223=>"000110000",
  11224=>"010011000",
  11225=>"101000110",
  11226=>"111011111",
  11227=>"111001101",
  11228=>"101001100",
  11229=>"101010110",
  11230=>"101001011",
  11231=>"111110011",
  11232=>"000000010",
  11233=>"111100111",
  11234=>"111011000",
  11235=>"111010101",
  11236=>"101010100",
  11237=>"001000111",
  11238=>"100111010",
  11239=>"101100101",
  11240=>"001011000",
  11241=>"100010101",
  11242=>"001100101",
  11243=>"100111000",
  11244=>"100010001",
  11245=>"101100101",
  11246=>"010111000",
  11247=>"110110010",
  11248=>"101101101",
  11249=>"100100001",
  11250=>"100110111",
  11251=>"100101010",
  11252=>"100101101",
  11253=>"000001111",
  11254=>"000111011",
  11255=>"111011010",
  11256=>"110110010",
  11257=>"101111000",
  11258=>"010010010",
  11259=>"111100101",
  11260=>"000110010",
  11261=>"101101100",
  11262=>"111100101",
  11263=>"111001110",
  11264=>"100100000",
  11265=>"101010011",
  11266=>"001111000",
  11267=>"011100110",
  11268=>"011011011",
  11269=>"010001001",
  11270=>"011010011",
  11271=>"010000110",
  11272=>"011101010",
  11273=>"000100101",
  11274=>"001000001",
  11275=>"101101100",
  11276=>"101101001",
  11277=>"000000101",
  11278=>"110100011",
  11279=>"111100111",
  11280=>"000000101",
  11281=>"100011000",
  11282=>"110001101",
  11283=>"011001010",
  11284=>"101111101",
  11285=>"110000001",
  11286=>"101101101",
  11287=>"000110000",
  11288=>"001000000",
  11289=>"001101100",
  11290=>"011100011",
  11291=>"100011110",
  11292=>"110001100",
  11293=>"110111010",
  11294=>"101100001",
  11295=>"110110001",
  11296=>"111011000",
  11297=>"010011001",
  11298=>"001101001",
  11299=>"001101100",
  11300=>"011011110",
  11301=>"001000000",
  11302=>"001100101",
  11303=>"101011010",
  11304=>"100010001",
  11305=>"001101100",
  11306=>"101011010",
  11307=>"110011111",
  11308=>"011101010",
  11309=>"001000000",
  11310=>"100001101",
  11311=>"110010000",
  11312=>"100001111",
  11313=>"010010100",
  11314=>"001010010",
  11315=>"111011100",
  11316=>"111101101",
  11317=>"001011110",
  11318=>"000100111",
  11319=>"101101111",
  11320=>"000001000",
  11321=>"000000100",
  11322=>"111100100",
  11323=>"010010111",
  11324=>"011111000",
  11325=>"000010000",
  11326=>"101111000",
  11327=>"011001100",
  11328=>"101011000",
  11329=>"000000000",
  11330=>"100111110",
  11331=>"011110111",
  11332=>"101010000",
  11333=>"111110111",
  11334=>"101111111",
  11335=>"110101010",
  11336=>"111010000",
  11337=>"001010010",
  11338=>"100001111",
  11339=>"100110001",
  11340=>"000010000",
  11341=>"100001010",
  11342=>"101001101",
  11343=>"000111001",
  11344=>"111011111",
  11345=>"000110010",
  11346=>"000101101",
  11347=>"110010110",
  11348=>"110110000",
  11349=>"011111111",
  11350=>"011001011",
  11351=>"111100101",
  11352=>"100011101",
  11353=>"110000110",
  11354=>"000011110",
  11355=>"000000000",
  11356=>"100110110",
  11357=>"100000011",
  11358=>"010000001",
  11359=>"110000111",
  11360=>"111110111",
  11361=>"001110011",
  11362=>"101100101",
  11363=>"011010100",
  11364=>"110001000",
  11365=>"101111100",
  11366=>"100110110",
  11367=>"010000111",
  11368=>"011000000",
  11369=>"010011100",
  11370=>"100101010",
  11371=>"011001010",
  11372=>"000100111",
  11373=>"110000010",
  11374=>"010000010",
  11375=>"110100011",
  11376=>"010110110",
  11377=>"000100010",
  11378=>"000101110",
  11379=>"001110111",
  11380=>"001011000",
  11381=>"010001011",
  11382=>"011000110",
  11383=>"010011100",
  11384=>"101011011",
  11385=>"000100101",
  11386=>"100010011",
  11387=>"011000100",
  11388=>"110010101",
  11389=>"011110011",
  11390=>"000010110",
  11391=>"011000101",
  11392=>"001101010",
  11393=>"001000100",
  11394=>"101011000",
  11395=>"001001010",
  11396=>"101100010",
  11397=>"101101110",
  11398=>"111101101",
  11399=>"010000000",
  11400=>"011010001",
  11401=>"100010011",
  11402=>"101110001",
  11403=>"101111101",
  11404=>"101100010",
  11405=>"110010010",
  11406=>"110010110",
  11407=>"000101111",
  11408=>"100010010",
  11409=>"001011101",
  11410=>"010011011",
  11411=>"101101001",
  11412=>"111111100",
  11413=>"101000100",
  11414=>"000000111",
  11415=>"100111110",
  11416=>"001111010",
  11417=>"110011011",
  11418=>"111101000",
  11419=>"000000010",
  11420=>"100100110",
  11421=>"100001010",
  11422=>"011100111",
  11423=>"000011000",
  11424=>"111001011",
  11425=>"011001100",
  11426=>"001101110",
  11427=>"101110000",
  11428=>"010011110",
  11429=>"100010000",
  11430=>"000110110",
  11431=>"010111100",
  11432=>"101110001",
  11433=>"000110000",
  11434=>"001010100",
  11435=>"000111010",
  11436=>"011010010",
  11437=>"111000111",
  11438=>"100010100",
  11439=>"101010100",
  11440=>"000100010",
  11441=>"111001101",
  11442=>"111110011",
  11443=>"110010001",
  11444=>"110101011",
  11445=>"000111011",
  11446=>"100001001",
  11447=>"011101011",
  11448=>"000011000",
  11449=>"011000110",
  11450=>"000100100",
  11451=>"010011010",
  11452=>"011110010",
  11453=>"000001100",
  11454=>"011110011",
  11455=>"001000010",
  11456=>"001001000",
  11457=>"100101001",
  11458=>"100111000",
  11459=>"011100101",
  11460=>"111101101",
  11461=>"010001110",
  11462=>"011100100",
  11463=>"111101010",
  11464=>"010001110",
  11465=>"111000111",
  11466=>"001010100",
  11467=>"100111111",
  11468=>"100100100",
  11469=>"100111110",
  11470=>"011100111",
  11471=>"010011111",
  11472=>"101000110",
  11473=>"011011101",
  11474=>"111000111",
  11475=>"001111100",
  11476=>"110011011",
  11477=>"010010000",
  11478=>"110100011",
  11479=>"011101100",
  11480=>"001001000",
  11481=>"110000010",
  11482=>"000001010",
  11483=>"110100000",
  11484=>"100111000",
  11485=>"011110101",
  11486=>"000110010",
  11487=>"111001111",
  11488=>"010001010",
  11489=>"000111011",
  11490=>"001000010",
  11491=>"000010000",
  11492=>"101010110",
  11493=>"110100111",
  11494=>"110001101",
  11495=>"011110110",
  11496=>"111010000",
  11497=>"010111100",
  11498=>"101010011",
  11499=>"101101000",
  11500=>"111110110",
  11501=>"100101010",
  11502=>"010000101",
  11503=>"101110011",
  11504=>"111011110",
  11505=>"100111111",
  11506=>"100001111",
  11507=>"001000100",
  11508=>"111101101",
  11509=>"100111110",
  11510=>"110011011",
  11511=>"111001110",
  11512=>"110101111",
  11513=>"011100001",
  11514=>"110101111",
  11515=>"101101110",
  11516=>"001001100",
  11517=>"100101011",
  11518=>"010010101",
  11519=>"000000011",
  11520=>"001000010",
  11521=>"010011110",
  11522=>"111001110",
  11523=>"001100100",
  11524=>"110011011",
  11525=>"101010101",
  11526=>"110000010",
  11527=>"000001011",
  11528=>"110000100",
  11529=>"111001001",
  11530=>"111110101",
  11531=>"101001100",
  11532=>"001000000",
  11533=>"111000110",
  11534=>"000001110",
  11535=>"111110100",
  11536=>"101001101",
  11537=>"000010010",
  11538=>"110101111",
  11539=>"101010110",
  11540=>"011000111",
  11541=>"011101001",
  11542=>"110011010",
  11543=>"010100011",
  11544=>"000011000",
  11545=>"100000111",
  11546=>"111001111",
  11547=>"100011101",
  11548=>"001000110",
  11549=>"110110100",
  11550=>"010110000",
  11551=>"010010000",
  11552=>"100001010",
  11553=>"011110100",
  11554=>"110111111",
  11555=>"010110110",
  11556=>"110111110",
  11557=>"101110000",
  11558=>"111111100",
  11559=>"101001001",
  11560=>"110000100",
  11561=>"010111000",
  11562=>"011011000",
  11563=>"000100101",
  11564=>"010001000",
  11565=>"011111000",
  11566=>"010011011",
  11567=>"001001011",
  11568=>"111000110",
  11569=>"001101010",
  11570=>"101100111",
  11571=>"011000110",
  11572=>"000000001",
  11573=>"101011110",
  11574=>"001100011",
  11575=>"111100011",
  11576=>"111110010",
  11577=>"111111000",
  11578=>"110100000",
  11579=>"001001011",
  11580=>"010110001",
  11581=>"111010100",
  11582=>"111100100",
  11583=>"010001010",
  11584=>"111011100",
  11585=>"111000000",
  11586=>"011011011",
  11587=>"000100110",
  11588=>"000001000",
  11589=>"010100101",
  11590=>"010010100",
  11591=>"001000110",
  11592=>"110100010",
  11593=>"101110011",
  11594=>"111100011",
  11595=>"011100001",
  11596=>"000001010",
  11597=>"010011100",
  11598=>"010101010",
  11599=>"110001111",
  11600=>"111001000",
  11601=>"100001001",
  11602=>"011101111",
  11603=>"001110011",
  11604=>"100010001",
  11605=>"001010100",
  11606=>"011000111",
  11607=>"011011010",
  11608=>"001100001",
  11609=>"111001001",
  11610=>"000010111",
  11611=>"011111110",
  11612=>"101111111",
  11613=>"010110001",
  11614=>"010000010",
  11615=>"111001111",
  11616=>"100000100",
  11617=>"010011101",
  11618=>"101100001",
  11619=>"111111000",
  11620=>"011110100",
  11621=>"111111101",
  11622=>"010111110",
  11623=>"010100110",
  11624=>"100101010",
  11625=>"100111000",
  11626=>"111001001",
  11627=>"110100001",
  11628=>"010011000",
  11629=>"010010011",
  11630=>"100010111",
  11631=>"011101100",
  11632=>"110110110",
  11633=>"111010010",
  11634=>"100001011",
  11635=>"010110110",
  11636=>"001010001",
  11637=>"011000011",
  11638=>"011001110",
  11639=>"111111001",
  11640=>"100101110",
  11641=>"101011101",
  11642=>"001010011",
  11643=>"010011100",
  11644=>"011000010",
  11645=>"011011111",
  11646=>"010111110",
  11647=>"100010001",
  11648=>"110000100",
  11649=>"000000111",
  11650=>"011100010",
  11651=>"011101111",
  11652=>"100110010",
  11653=>"100111100",
  11654=>"100101001",
  11655=>"010010010",
  11656=>"001011100",
  11657=>"011110011",
  11658=>"100110111",
  11659=>"111111000",
  11660=>"011100100",
  11661=>"101110101",
  11662=>"000011101",
  11663=>"011110011",
  11664=>"001001010",
  11665=>"111000001",
  11666=>"000111011",
  11667=>"100000101",
  11668=>"110000100",
  11669=>"001100101",
  11670=>"000101011",
  11671=>"000001001",
  11672=>"100000101",
  11673=>"001010101",
  11674=>"000110011",
  11675=>"001000001",
  11676=>"101001000",
  11677=>"111000010",
  11678=>"100000000",
  11679=>"111000010",
  11680=>"001110001",
  11681=>"111101110",
  11682=>"001110000",
  11683=>"000100111",
  11684=>"101110111",
  11685=>"100100000",
  11686=>"010101111",
  11687=>"001100110",
  11688=>"100001110",
  11689=>"010001111",
  11690=>"011001000",
  11691=>"011010110",
  11692=>"111111001",
  11693=>"001100101",
  11694=>"001100010",
  11695=>"010101101",
  11696=>"100000000",
  11697=>"111010001",
  11698=>"101110011",
  11699=>"101010101",
  11700=>"100010100",
  11701=>"101000000",
  11702=>"001100110",
  11703=>"101001000",
  11704=>"011100000",
  11705=>"101111100",
  11706=>"111010010",
  11707=>"000111111",
  11708=>"101000111",
  11709=>"111001100",
  11710=>"100101101",
  11711=>"110111111",
  11712=>"011010011",
  11713=>"100000100",
  11714=>"011010000",
  11715=>"010100001",
  11716=>"001010000",
  11717=>"011000000",
  11718=>"010111110",
  11719=>"100110010",
  11720=>"101000111",
  11721=>"011001100",
  11722=>"110110100",
  11723=>"011001110",
  11724=>"001101110",
  11725=>"010101110",
  11726=>"011001011",
  11727=>"110011000",
  11728=>"111100111",
  11729=>"000010110",
  11730=>"010011110",
  11731=>"110110110",
  11732=>"000111010",
  11733=>"110010011",
  11734=>"111101000",
  11735=>"101000011",
  11736=>"111001000",
  11737=>"110000011",
  11738=>"000100100",
  11739=>"111001011",
  11740=>"000001011",
  11741=>"001101111",
  11742=>"100001111",
  11743=>"010010100",
  11744=>"001110110",
  11745=>"000000000",
  11746=>"000101011",
  11747=>"101100101",
  11748=>"110001010",
  11749=>"111010110",
  11750=>"001001010",
  11751=>"010010000",
  11752=>"001000110",
  11753=>"100000111",
  11754=>"101010110",
  11755=>"000001010",
  11756=>"111010111",
  11757=>"111001100",
  11758=>"100101000",
  11759=>"110101110",
  11760=>"100000001",
  11761=>"001110110",
  11762=>"111000001",
  11763=>"011111101",
  11764=>"000110110",
  11765=>"111011110",
  11766=>"000110000",
  11767=>"100101110",
  11768=>"011011010",
  11769=>"110010111",
  11770=>"110110000",
  11771=>"100100111",
  11772=>"111010111",
  11773=>"100111010",
  11774=>"011111000",
  11775=>"101111000",
  11776=>"000100100",
  11777=>"101011111",
  11778=>"100001010",
  11779=>"101010001",
  11780=>"100101101",
  11781=>"100000101",
  11782=>"000101110",
  11783=>"101100110",
  11784=>"111001111",
  11785=>"100001000",
  11786=>"100001111",
  11787=>"010101010",
  11788=>"001011000",
  11789=>"001001101",
  11790=>"001101011",
  11791=>"110110000",
  11792=>"000111101",
  11793=>"110111011",
  11794=>"010010010",
  11795=>"100111010",
  11796=>"110100010",
  11797=>"111100000",
  11798=>"001110011",
  11799=>"111011110",
  11800=>"100100110",
  11801=>"010001001",
  11802=>"001101110",
  11803=>"101000011",
  11804=>"000010101",
  11805=>"111010000",
  11806=>"101100110",
  11807=>"110101010",
  11808=>"000001010",
  11809=>"001110111",
  11810=>"101000011",
  11811=>"100001110",
  11812=>"000100101",
  11813=>"111111000",
  11814=>"100000101",
  11815=>"111001000",
  11816=>"000000110",
  11817=>"100110011",
  11818=>"001001100",
  11819=>"001010100",
  11820=>"110100000",
  11821=>"101010110",
  11822=>"011000100",
  11823=>"100001010",
  11824=>"101010011",
  11825=>"011101111",
  11826=>"100010010",
  11827=>"000100010",
  11828=>"111010011",
  11829=>"100000110",
  11830=>"110100011",
  11831=>"010001011",
  11832=>"111110110",
  11833=>"000011111",
  11834=>"011100101",
  11835=>"110010101",
  11836=>"001101111",
  11837=>"000000100",
  11838=>"001011000",
  11839=>"101001110",
  11840=>"100010001",
  11841=>"010000000",
  11842=>"010100011",
  11843=>"110111100",
  11844=>"001011101",
  11845=>"110111010",
  11846=>"100011100",
  11847=>"010101000",
  11848=>"110111111",
  11849=>"111010011",
  11850=>"001110010",
  11851=>"000111111",
  11852=>"100110011",
  11853=>"101000010",
  11854=>"101101011",
  11855=>"111000011",
  11856=>"101110001",
  11857=>"000011001",
  11858=>"111110000",
  11859=>"110001000",
  11860=>"001111000",
  11861=>"101101010",
  11862=>"110001010",
  11863=>"001011111",
  11864=>"110010010",
  11865=>"100011011",
  11866=>"000101011",
  11867=>"011010000",
  11868=>"101101111",
  11869=>"011101000",
  11870=>"001111110",
  11871=>"010011000",
  11872=>"001100001",
  11873=>"001010011",
  11874=>"011011100",
  11875=>"011111010",
  11876=>"101110101",
  11877=>"111111101",
  11878=>"010000011",
  11879=>"001000001",
  11880=>"110111100",
  11881=>"100000111",
  11882=>"010011101",
  11883=>"100111110",
  11884=>"001101110",
  11885=>"111111010",
  11886=>"010000001",
  11887=>"101010001",
  11888=>"000000111",
  11889=>"010000101",
  11890=>"101110101",
  11891=>"100000110",
  11892=>"111111001",
  11893=>"001000011",
  11894=>"001100111",
  11895=>"110011001",
  11896=>"010000000",
  11897=>"000001010",
  11898=>"011111010",
  11899=>"100100100",
  11900=>"100000101",
  11901=>"101111100",
  11902=>"010100100",
  11903=>"010011001",
  11904=>"110111110",
  11905=>"001110101",
  11906=>"100000100",
  11907=>"010010101",
  11908=>"100011100",
  11909=>"101111001",
  11910=>"010011001",
  11911=>"000001000",
  11912=>"100000110",
  11913=>"000110100",
  11914=>"110100111",
  11915=>"010010111",
  11916=>"000001111",
  11917=>"011010001",
  11918=>"110110101",
  11919=>"010010110",
  11920=>"010111011",
  11921=>"001101011",
  11922=>"001111101",
  11923=>"010111100",
  11924=>"011010111",
  11925=>"010111000",
  11926=>"100011111",
  11927=>"101111110",
  11928=>"010001111",
  11929=>"000101100",
  11930=>"100001101",
  11931=>"111000010",
  11932=>"000110000",
  11933=>"111101101",
  11934=>"100001100",
  11935=>"101001000",
  11936=>"100100111",
  11937=>"110111110",
  11938=>"110111010",
  11939=>"000011111",
  11940=>"001111000",
  11941=>"010000111",
  11942=>"001001000",
  11943=>"001010001",
  11944=>"010001100",
  11945=>"110110010",
  11946=>"001010001",
  11947=>"010011001",
  11948=>"110011000",
  11949=>"111111101",
  11950=>"100001111",
  11951=>"000000011",
  11952=>"001111000",
  11953=>"010011011",
  11954=>"000010011",
  11955=>"000010000",
  11956=>"111110010",
  11957=>"000000000",
  11958=>"000100010",
  11959=>"101110010",
  11960=>"000011000",
  11961=>"100000000",
  11962=>"100100000",
  11963=>"110111101",
  11964=>"100100111",
  11965=>"011000101",
  11966=>"010001101",
  11967=>"011000000",
  11968=>"011011011",
  11969=>"100101110",
  11970=>"111010011",
  11971=>"101111110",
  11972=>"001010010",
  11973=>"100011001",
  11974=>"111011010",
  11975=>"110000000",
  11976=>"000001110",
  11977=>"111000110",
  11978=>"000001001",
  11979=>"110101010",
  11980=>"011100001",
  11981=>"111101111",
  11982=>"100110110",
  11983=>"001000010",
  11984=>"101111011",
  11985=>"000000110",
  11986=>"111110100",
  11987=>"010001011",
  11988=>"100011001",
  11989=>"111100010",
  11990=>"000100010",
  11991=>"010100011",
  11992=>"100111000",
  11993=>"110101011",
  11994=>"001000011",
  11995=>"100110110",
  11996=>"110000000",
  11997=>"111010001",
  11998=>"110100100",
  11999=>"011001111",
  12000=>"111100110",
  12001=>"010100010",
  12002=>"000110101",
  12003=>"100011010",
  12004=>"010111100",
  12005=>"111101111",
  12006=>"100001001",
  12007=>"000110100",
  12008=>"101100110",
  12009=>"000001000",
  12010=>"111100001",
  12011=>"100011100",
  12012=>"111000010",
  12013=>"010011101",
  12014=>"111111011",
  12015=>"100110110",
  12016=>"101011111",
  12017=>"000010101",
  12018=>"101100001",
  12019=>"101010000",
  12020=>"111100001",
  12021=>"100001010",
  12022=>"000010110",
  12023=>"111010101",
  12024=>"111101111",
  12025=>"110100000",
  12026=>"100001110",
  12027=>"101010100",
  12028=>"101100001",
  12029=>"111100101",
  12030=>"110011100",
  12031=>"101010110",
  12032=>"111100000",
  12033=>"111011111",
  12034=>"000101100",
  12035=>"111011111",
  12036=>"111111100",
  12037=>"010101011",
  12038=>"101001101",
  12039=>"010000001",
  12040=>"111001111",
  12041=>"011100111",
  12042=>"001010001",
  12043=>"000000100",
  12044=>"111110001",
  12045=>"100101011",
  12046=>"111111101",
  12047=>"100010101",
  12048=>"010010111",
  12049=>"010101101",
  12050=>"101001101",
  12051=>"110100011",
  12052=>"100000101",
  12053=>"110100100",
  12054=>"010010001",
  12055=>"010010101",
  12056=>"101100100",
  12057=>"000001110",
  12058=>"100000011",
  12059=>"101100111",
  12060=>"010011000",
  12061=>"011011000",
  12062=>"011100101",
  12063=>"110100001",
  12064=>"010001001",
  12065=>"001110110",
  12066=>"101001111",
  12067=>"100000101",
  12068=>"110001110",
  12069=>"000101011",
  12070=>"101101110",
  12071=>"001100110",
  12072=>"000100001",
  12073=>"100101101",
  12074=>"101000111",
  12075=>"110011010",
  12076=>"110001000",
  12077=>"110101101",
  12078=>"001110000",
  12079=>"101110000",
  12080=>"100100010",
  12081=>"111011101",
  12082=>"011011011",
  12083=>"111100100",
  12084=>"100011000",
  12085=>"101001010",
  12086=>"111100000",
  12087=>"010011101",
  12088=>"000100111",
  12089=>"011110001",
  12090=>"101011100",
  12091=>"101111111",
  12092=>"101110001",
  12093=>"101110010",
  12094=>"011100011",
  12095=>"011111100",
  12096=>"100000000",
  12097=>"010110011",
  12098=>"010001010",
  12099=>"001000110",
  12100=>"011101011",
  12101=>"000100000",
  12102=>"010100001",
  12103=>"000100111",
  12104=>"111101110",
  12105=>"101011001",
  12106=>"110110110",
  12107=>"010010100",
  12108=>"110010110",
  12109=>"100010100",
  12110=>"101000100",
  12111=>"000010001",
  12112=>"110000010",
  12113=>"110111011",
  12114=>"010010000",
  12115=>"111011111",
  12116=>"001010001",
  12117=>"000110000",
  12118=>"100011000",
  12119=>"111100001",
  12120=>"010100000",
  12121=>"101111111",
  12122=>"101100110",
  12123=>"101011001",
  12124=>"011100001",
  12125=>"111111000",
  12126=>"000010101",
  12127=>"010110000",
  12128=>"010000111",
  12129=>"101111111",
  12130=>"111001111",
  12131=>"101110011",
  12132=>"011101110",
  12133=>"111010000",
  12134=>"100010001",
  12135=>"010111011",
  12136=>"101110100",
  12137=>"000101111",
  12138=>"010101111",
  12139=>"000010110",
  12140=>"000101000",
  12141=>"100101100",
  12142=>"011111100",
  12143=>"010001010",
  12144=>"010110101",
  12145=>"010101001",
  12146=>"011001001",
  12147=>"011000111",
  12148=>"010100110",
  12149=>"111111001",
  12150=>"111111000",
  12151=>"100101101",
  12152=>"101010100",
  12153=>"011110110",
  12154=>"010111101",
  12155=>"010010000",
  12156=>"011110010",
  12157=>"001000010",
  12158=>"010010000",
  12159=>"100011111",
  12160=>"010011001",
  12161=>"111111011",
  12162=>"001110111",
  12163=>"100011101",
  12164=>"001000010",
  12165=>"110000011",
  12166=>"011100010",
  12167=>"110101011",
  12168=>"111111101",
  12169=>"001000110",
  12170=>"010010100",
  12171=>"111101000",
  12172=>"100000100",
  12173=>"000100000",
  12174=>"001110101",
  12175=>"001101010",
  12176=>"111011001",
  12177=>"100011111",
  12178=>"001111111",
  12179=>"110111011",
  12180=>"100101011",
  12181=>"100111101",
  12182=>"100010101",
  12183=>"001100011",
  12184=>"100111011",
  12185=>"100100010",
  12186=>"000001000",
  12187=>"000110110",
  12188=>"011000100",
  12189=>"000010101",
  12190=>"000011100",
  12191=>"100101110",
  12192=>"100101110",
  12193=>"101010101",
  12194=>"001011010",
  12195=>"110111010",
  12196=>"101001001",
  12197=>"011001101",
  12198=>"000000000",
  12199=>"100111101",
  12200=>"001101111",
  12201=>"100111011",
  12202=>"000110010",
  12203=>"100110111",
  12204=>"010000010",
  12205=>"000010010",
  12206=>"011011100",
  12207=>"111000011",
  12208=>"111111000",
  12209=>"001010001",
  12210=>"010110111",
  12211=>"101011111",
  12212=>"011000111",
  12213=>"100100001",
  12214=>"010100110",
  12215=>"100010011",
  12216=>"000000100",
  12217=>"100011110",
  12218=>"010001110",
  12219=>"111011101",
  12220=>"000010110",
  12221=>"111011011",
  12222=>"100101101",
  12223=>"010010001",
  12224=>"110111110",
  12225=>"010011010",
  12226=>"110010000",
  12227=>"000010110",
  12228=>"011001001",
  12229=>"000101010",
  12230=>"001111111",
  12231=>"001110111",
  12232=>"001111101",
  12233=>"001101010",
  12234=>"011101010",
  12235=>"000000001",
  12236=>"010100100",
  12237=>"100101100",
  12238=>"110010011",
  12239=>"000011000",
  12240=>"010111110",
  12241=>"100110111",
  12242=>"001011001",
  12243=>"011101110",
  12244=>"111001101",
  12245=>"110101000",
  12246=>"010110100",
  12247=>"110101111",
  12248=>"001101011",
  12249=>"010001110",
  12250=>"110110101",
  12251=>"111110110",
  12252=>"000000100",
  12253=>"010111110",
  12254=>"010011011",
  12255=>"110000010",
  12256=>"011111111",
  12257=>"101101001",
  12258=>"100101000",
  12259=>"111000010",
  12260=>"001000001",
  12261=>"001100011",
  12262=>"011010011",
  12263=>"111101100",
  12264=>"110100100",
  12265=>"100010101",
  12266=>"011011011",
  12267=>"000000111",
  12268=>"111110011",
  12269=>"000010111",
  12270=>"000000000",
  12271=>"110101011",
  12272=>"010001100",
  12273=>"100010001",
  12274=>"100010111",
  12275=>"000000111",
  12276=>"001100010",
  12277=>"100010100",
  12278=>"010010101",
  12279=>"100010010",
  12280=>"011101111",
  12281=>"011100100",
  12282=>"010111101",
  12283=>"110101010",
  12284=>"110011111",
  12285=>"110110110",
  12286=>"100011010",
  12287=>"001110110",
  12288=>"100101001",
  12289=>"001001101",
  12290=>"111111111",
  12291=>"001100101",
  12292=>"100101011",
  12293=>"111001111",
  12294=>"110111000",
  12295=>"100001110",
  12296=>"001010011",
  12297=>"111010001",
  12298=>"110100010",
  12299=>"110100000",
  12300=>"000111000",
  12301=>"001000001",
  12302=>"100010000",
  12303=>"100000010",
  12304=>"100011111",
  12305=>"001110010",
  12306=>"101101100",
  12307=>"001100001",
  12308=>"111111111",
  12309=>"100110000",
  12310=>"010001010",
  12311=>"111010000",
  12312=>"011101000",
  12313=>"001110011",
  12314=>"101111010",
  12315=>"100100000",
  12316=>"001010011",
  12317=>"001011111",
  12318=>"011011100",
  12319=>"100011101",
  12320=>"101110010",
  12321=>"001110100",
  12322=>"110111010",
  12323=>"111111001",
  12324=>"010011000",
  12325=>"101110010",
  12326=>"101001110",
  12327=>"110011000",
  12328=>"100001110",
  12329=>"111110100",
  12330=>"101101001",
  12331=>"111010010",
  12332=>"000001000",
  12333=>"000101111",
  12334=>"010011010",
  12335=>"000101110",
  12336=>"101010100",
  12337=>"011001001",
  12338=>"101010011",
  12339=>"100100010",
  12340=>"111111111",
  12341=>"000011100",
  12342=>"101010011",
  12343=>"101010101",
  12344=>"001000101",
  12345=>"000000010",
  12346=>"111100011",
  12347=>"101111001",
  12348=>"000010001",
  12349=>"100100001",
  12350=>"100010000",
  12351=>"111100010",
  12352=>"110101110",
  12353=>"100001101",
  12354=>"110000101",
  12355=>"001011100",
  12356=>"101100110",
  12357=>"111100111",
  12358=>"110111001",
  12359=>"011001011",
  12360=>"111100010",
  12361=>"100101100",
  12362=>"101100010",
  12363=>"011100001",
  12364=>"011000001",
  12365=>"101000101",
  12366=>"010010011",
  12367=>"101000001",
  12368=>"111000011",
  12369=>"011001100",
  12370=>"010100111",
  12371=>"000011001",
  12372=>"000110111",
  12373=>"011111111",
  12374=>"101011110",
  12375=>"011001010",
  12376=>"010111110",
  12377=>"001100111",
  12378=>"101010111",
  12379=>"111010000",
  12380=>"111010111",
  12381=>"100101010",
  12382=>"000001101",
  12383=>"001001001",
  12384=>"001000001",
  12385=>"101011101",
  12386=>"011110101",
  12387=>"000010011",
  12388=>"101110010",
  12389=>"100110110",
  12390=>"000101100",
  12391=>"010010100",
  12392=>"100000011",
  12393=>"010111101",
  12394=>"101000100",
  12395=>"100101101",
  12396=>"001010100",
  12397=>"000000101",
  12398=>"000001101",
  12399=>"010101111",
  12400=>"000011001",
  12401=>"101111010",
  12402=>"100010011",
  12403=>"000001001",
  12404=>"110010001",
  12405=>"111100011",
  12406=>"001011010",
  12407=>"001100101",
  12408=>"001010101",
  12409=>"000011110",
  12410=>"100010100",
  12411=>"100100001",
  12412=>"000110110",
  12413=>"010110011",
  12414=>"110011001",
  12415=>"010001010",
  12416=>"010100101",
  12417=>"011000101",
  12418=>"001110000",
  12419=>"100110011",
  12420=>"000001101",
  12421=>"000001001",
  12422=>"001111011",
  12423=>"010000001",
  12424=>"000001010",
  12425=>"010100100",
  12426=>"011101001",
  12427=>"010011010",
  12428=>"111111100",
  12429=>"111100101",
  12430=>"100111111",
  12431=>"011110011",
  12432=>"010000010",
  12433=>"011001000",
  12434=>"000111101",
  12435=>"111110110",
  12436=>"100000011",
  12437=>"000101000",
  12438=>"110011100",
  12439=>"100110110",
  12440=>"101010110",
  12441=>"111001110",
  12442=>"001101001",
  12443=>"000111010",
  12444=>"100001100",
  12445=>"001100000",
  12446=>"001111110",
  12447=>"100101100",
  12448=>"101111010",
  12449=>"100000110",
  12450=>"011101010",
  12451=>"101111101",
  12452=>"010000111",
  12453=>"100010110",
  12454=>"111101001",
  12455=>"001101010",
  12456=>"000001101",
  12457=>"001011010",
  12458=>"001111110",
  12459=>"111101111",
  12460=>"100011010",
  12461=>"100101010",
  12462=>"100110101",
  12463=>"000001000",
  12464=>"101001100",
  12465=>"010111010",
  12466=>"111010110",
  12467=>"100011100",
  12468=>"101001000",
  12469=>"101010110",
  12470=>"101000001",
  12471=>"110100101",
  12472=>"001010001",
  12473=>"101101100",
  12474=>"111110010",
  12475=>"101101011",
  12476=>"001111000",
  12477=>"000101001",
  12478=>"000111001",
  12479=>"101011010",
  12480=>"000001100",
  12481=>"001111001",
  12482=>"101110010",
  12483=>"001010101",
  12484=>"110101001",
  12485=>"001110111",
  12486=>"011010001",
  12487=>"000101001",
  12488=>"001100000",
  12489=>"111010000",
  12490=>"000010010",
  12491=>"110111101",
  12492=>"111111010",
  12493=>"010100001",
  12494=>"001101011",
  12495=>"111011010",
  12496=>"110010100",
  12497=>"110101001",
  12498=>"100111001",
  12499=>"000000101",
  12500=>"111110001",
  12501=>"111110101",
  12502=>"110000001",
  12503=>"100010111",
  12504=>"000010101",
  12505=>"100101101",
  12506=>"000000100",
  12507=>"010100000",
  12508=>"001000010",
  12509=>"110111010",
  12510=>"010100000",
  12511=>"011001101",
  12512=>"101101010",
  12513=>"001011000",
  12514=>"101001111",
  12515=>"000000111",
  12516=>"101101100",
  12517=>"011010000",
  12518=>"100110110",
  12519=>"011101001",
  12520=>"010010101",
  12521=>"000101110",
  12522=>"001000101",
  12523=>"000001111",
  12524=>"011110000",
  12525=>"101101100",
  12526=>"000011001",
  12527=>"010110010",
  12528=>"100110110",
  12529=>"100110010",
  12530=>"000100010",
  12531=>"000000111",
  12532=>"011101101",
  12533=>"000110111",
  12534=>"101011001",
  12535=>"011000100",
  12536=>"101010101",
  12537=>"110101101",
  12538=>"111111000",
  12539=>"100000101",
  12540=>"010011010",
  12541=>"000101101",
  12542=>"000100100",
  12543=>"011001001",
  12544=>"110111011",
  12545=>"010001001",
  12546=>"110000000",
  12547=>"010001101",
  12548=>"111011111",
  12549=>"100101110",
  12550=>"100111010",
  12551=>"100111101",
  12552=>"000010000",
  12553=>"011000000",
  12554=>"000000001",
  12555=>"010010101",
  12556=>"101000111",
  12557=>"000101011",
  12558=>"101100110",
  12559=>"100101000",
  12560=>"001101010",
  12561=>"111011001",
  12562=>"110010000",
  12563=>"100000101",
  12564=>"100000100",
  12565=>"110011000",
  12566=>"001101000",
  12567=>"101110010",
  12568=>"011101101",
  12569=>"101000110",
  12570=>"000000010",
  12571=>"000110000",
  12572=>"001000100",
  12573=>"010000111",
  12574=>"001100000",
  12575=>"010000110",
  12576=>"101000111",
  12577=>"001111110",
  12578=>"101101011",
  12579=>"000101001",
  12580=>"001110111",
  12581=>"010100010",
  12582=>"101110100",
  12583=>"011101101",
  12584=>"010101110",
  12585=>"010010000",
  12586=>"111100010",
  12587=>"111010010",
  12588=>"011101110",
  12589=>"000000101",
  12590=>"011000111",
  12591=>"100010100",
  12592=>"101011110",
  12593=>"011001100",
  12594=>"011010111",
  12595=>"110100011",
  12596=>"111001101",
  12597=>"001001011",
  12598=>"101101110",
  12599=>"101001001",
  12600=>"010001010",
  12601=>"100100010",
  12602=>"110100110",
  12603=>"010000101",
  12604=>"101000011",
  12605=>"100011100",
  12606=>"111001101",
  12607=>"010000101",
  12608=>"011101111",
  12609=>"100100110",
  12610=>"001010011",
  12611=>"100111001",
  12612=>"000111111",
  12613=>"100011000",
  12614=>"101000110",
  12615=>"110101110",
  12616=>"010111010",
  12617=>"101110100",
  12618=>"011001101",
  12619=>"001001100",
  12620=>"000100100",
  12621=>"110000001",
  12622=>"101100110",
  12623=>"011000010",
  12624=>"110100000",
  12625=>"111101100",
  12626=>"100001101",
  12627=>"101010011",
  12628=>"100111000",
  12629=>"001111011",
  12630=>"110110010",
  12631=>"100110110",
  12632=>"001100010",
  12633=>"010111000",
  12634=>"110011000",
  12635=>"010101011",
  12636=>"101101100",
  12637=>"110011010",
  12638=>"101010000",
  12639=>"000010011",
  12640=>"111000001",
  12641=>"011001110",
  12642=>"001101111",
  12643=>"011000000",
  12644=>"111101000",
  12645=>"101000111",
  12646=>"110100011",
  12647=>"111000011",
  12648=>"111111110",
  12649=>"011110001",
  12650=>"010101100",
  12651=>"001110110",
  12652=>"110110000",
  12653=>"111111111",
  12654=>"101000110",
  12655=>"100001111",
  12656=>"000000011",
  12657=>"111011010",
  12658=>"001100101",
  12659=>"100000100",
  12660=>"000001101",
  12661=>"110101111",
  12662=>"011101011",
  12663=>"111010010",
  12664=>"001111111",
  12665=>"000101110",
  12666=>"011111111",
  12667=>"110010000",
  12668=>"001111000",
  12669=>"001001100",
  12670=>"011111010",
  12671=>"010000000",
  12672=>"010010011",
  12673=>"011101010",
  12674=>"010011100",
  12675=>"111010000",
  12676=>"110111100",
  12677=>"010111000",
  12678=>"001100000",
  12679=>"111111110",
  12680=>"101100000",
  12681=>"000110000",
  12682=>"111110100",
  12683=>"100011101",
  12684=>"010010001",
  12685=>"010100001",
  12686=>"100110001",
  12687=>"000010010",
  12688=>"010000001",
  12689=>"010000000",
  12690=>"010101110",
  12691=>"001101000",
  12692=>"000011011",
  12693=>"010011110",
  12694=>"000010000",
  12695=>"110101100",
  12696=>"010000100",
  12697=>"010100000",
  12698=>"101110011",
  12699=>"010100000",
  12700=>"000010000",
  12701=>"101111111",
  12702=>"111100010",
  12703=>"001001010",
  12704=>"000001010",
  12705=>"100000000",
  12706=>"000100101",
  12707=>"110011101",
  12708=>"101000101",
  12709=>"101111110",
  12710=>"000100000",
  12711=>"001110101",
  12712=>"000001001",
  12713=>"001000100",
  12714=>"001001001",
  12715=>"101000111",
  12716=>"101001100",
  12717=>"000101011",
  12718=>"011101100",
  12719=>"001111100",
  12720=>"101101110",
  12721=>"011101100",
  12722=>"111101101",
  12723=>"010110000",
  12724=>"110111111",
  12725=>"101111000",
  12726=>"110000010",
  12727=>"101001100",
  12728=>"011101000",
  12729=>"011001110",
  12730=>"110001111",
  12731=>"001001000",
  12732=>"100000010",
  12733=>"001011100",
  12734=>"011101100",
  12735=>"010001110",
  12736=>"110001110",
  12737=>"000110010",
  12738=>"001000111",
  12739=>"100100000",
  12740=>"100011100",
  12741=>"111011100",
  12742=>"000110011",
  12743=>"111101011",
  12744=>"001010000",
  12745=>"001100000",
  12746=>"001001010",
  12747=>"100110100",
  12748=>"010100101",
  12749=>"101110000",
  12750=>"000100111",
  12751=>"000001100",
  12752=>"110111011",
  12753=>"101111101",
  12754=>"001110101",
  12755=>"111111000",
  12756=>"001111010",
  12757=>"101100100",
  12758=>"100000101",
  12759=>"010101000",
  12760=>"000000000",
  12761=>"010111101",
  12762=>"100101100",
  12763=>"010101111",
  12764=>"110110100",
  12765=>"110110111",
  12766=>"100111010",
  12767=>"011011110",
  12768=>"000101111",
  12769=>"110001000",
  12770=>"111110110",
  12771=>"011000110",
  12772=>"100011100",
  12773=>"011110001",
  12774=>"110000110",
  12775=>"000010000",
  12776=>"111110001",
  12777=>"110000101",
  12778=>"100000010",
  12779=>"100111101",
  12780=>"110101100",
  12781=>"101001101",
  12782=>"110110000",
  12783=>"001000010",
  12784=>"111010110",
  12785=>"001111011",
  12786=>"101100010",
  12787=>"001100101",
  12788=>"110110110",
  12789=>"010101111",
  12790=>"100101000",
  12791=>"111011001",
  12792=>"000110111",
  12793=>"001011011",
  12794=>"001101010",
  12795=>"101110101",
  12796=>"001111011",
  12797=>"110110101",
  12798=>"101100111",
  12799=>"111011111",
  12800=>"100001111",
  12801=>"111100100",
  12802=>"110011011",
  12803=>"010100010",
  12804=>"011100001",
  12805=>"000100110",
  12806=>"000000001",
  12807=>"101101011",
  12808=>"100011111",
  12809=>"111011101",
  12810=>"001010000",
  12811=>"110100111",
  12812=>"000011001",
  12813=>"100101110",
  12814=>"100001000",
  12815=>"111110100",
  12816=>"100100111",
  12817=>"111111011",
  12818=>"111001011",
  12819=>"101101101",
  12820=>"001010011",
  12821=>"101110101",
  12822=>"000100011",
  12823=>"110111101",
  12824=>"111111000",
  12825=>"010101010",
  12826=>"101010110",
  12827=>"111010111",
  12828=>"001011111",
  12829=>"001001011",
  12830=>"100100000",
  12831=>"010110110",
  12832=>"011000010",
  12833=>"101110010",
  12834=>"010000000",
  12835=>"001010010",
  12836=>"010110111",
  12837=>"110000111",
  12838=>"101010001",
  12839=>"100110101",
  12840=>"010110000",
  12841=>"111010000",
  12842=>"000011001",
  12843=>"100000101",
  12844=>"111001110",
  12845=>"001101100",
  12846=>"111000100",
  12847=>"111110111",
  12848=>"010100011",
  12849=>"010100001",
  12850=>"001111001",
  12851=>"000110100",
  12852=>"110011101",
  12853=>"100100100",
  12854=>"001011111",
  12855=>"001101111",
  12856=>"101001010",
  12857=>"101111001",
  12858=>"010000010",
  12859=>"011100010",
  12860=>"000110000",
  12861=>"000110000",
  12862=>"000111000",
  12863=>"111111110",
  12864=>"111101000",
  12865=>"000111100",
  12866=>"011000001",
  12867=>"110000001",
  12868=>"001011000",
  12869=>"010100011",
  12870=>"010110001",
  12871=>"101100101",
  12872=>"010111000",
  12873=>"101010000",
  12874=>"011101111",
  12875=>"111100000",
  12876=>"011000111",
  12877=>"100100010",
  12878=>"111011111",
  12879=>"110100011",
  12880=>"111011111",
  12881=>"101101100",
  12882=>"011011010",
  12883=>"101110000",
  12884=>"010000100",
  12885=>"010100100",
  12886=>"001001101",
  12887=>"011110110",
  12888=>"111000100",
  12889=>"011010011",
  12890=>"010110000",
  12891=>"100110000",
  12892=>"111011001",
  12893=>"100110100",
  12894=>"011011011",
  12895=>"011101111",
  12896=>"011101010",
  12897=>"111111101",
  12898=>"000001100",
  12899=>"011110111",
  12900=>"101011110",
  12901=>"000011011",
  12902=>"000011101",
  12903=>"101001100",
  12904=>"111111000",
  12905=>"100111111",
  12906=>"111000100",
  12907=>"100100101",
  12908=>"000101011",
  12909=>"110000000",
  12910=>"100101111",
  12911=>"110100100",
  12912=>"100001010",
  12913=>"000111011",
  12914=>"101100111",
  12915=>"111011000",
  12916=>"001000101",
  12917=>"011000110",
  12918=>"011100111",
  12919=>"101100111",
  12920=>"101110011",
  12921=>"001000010",
  12922=>"010000001",
  12923=>"100010011",
  12924=>"111001110",
  12925=>"110010001",
  12926=>"110100100",
  12927=>"111100010",
  12928=>"000101101",
  12929=>"111110101",
  12930=>"000000001",
  12931=>"110011010",
  12932=>"001101100",
  12933=>"010111000",
  12934=>"011110010",
  12935=>"000001100",
  12936=>"010110110",
  12937=>"111100001",
  12938=>"101111000",
  12939=>"001110000",
  12940=>"011000001",
  12941=>"000011011",
  12942=>"111011110",
  12943=>"110000111",
  12944=>"000010010",
  12945=>"001110100",
  12946=>"011111111",
  12947=>"001111000",
  12948=>"010000010",
  12949=>"000100011",
  12950=>"010011111",
  12951=>"110000010",
  12952=>"111000000",
  12953=>"111000110",
  12954=>"111001101",
  12955=>"100100100",
  12956=>"010100000",
  12957=>"000111001",
  12958=>"100111010",
  12959=>"110110111",
  12960=>"110101111",
  12961=>"001101111",
  12962=>"001010111",
  12963=>"000101111",
  12964=>"111001011",
  12965=>"000111000",
  12966=>"110010010",
  12967=>"011000000",
  12968=>"000100000",
  12969=>"010100100",
  12970=>"101010100",
  12971=>"011011000",
  12972=>"000000010",
  12973=>"100100100",
  12974=>"010111001",
  12975=>"100001111",
  12976=>"001110110",
  12977=>"011000101",
  12978=>"100101001",
  12979=>"101001011",
  12980=>"001110001",
  12981=>"111111000",
  12982=>"101011101",
  12983=>"000111100",
  12984=>"101000001",
  12985=>"001010111",
  12986=>"010111110",
  12987=>"100011100",
  12988=>"010010101",
  12989=>"111100100",
  12990=>"110101111",
  12991=>"101101101",
  12992=>"000001100",
  12993=>"010100111",
  12994=>"011100100",
  12995=>"001001010",
  12996=>"000000110",
  12997=>"000110101",
  12998=>"101111010",
  12999=>"011010001",
  13000=>"001100011",
  13001=>"010100110",
  13002=>"101010001",
  13003=>"010010111",
  13004=>"101100000",
  13005=>"110110110",
  13006=>"010101101",
  13007=>"111010011",
  13008=>"011001011",
  13009=>"000001000",
  13010=>"010110001",
  13011=>"001000011",
  13012=>"111100111",
  13013=>"001000100",
  13014=>"011011110",
  13015=>"011110101",
  13016=>"101011001",
  13017=>"001000100",
  13018=>"100100110",
  13019=>"010100010",
  13020=>"101101100",
  13021=>"100110011",
  13022=>"001000101",
  13023=>"110000101",
  13024=>"010110010",
  13025=>"111110001",
  13026=>"110011110",
  13027=>"100010000",
  13028=>"110001101",
  13029=>"001010000",
  13030=>"111100011",
  13031=>"000100001",
  13032=>"101111111",
  13033=>"111011110",
  13034=>"011000010",
  13035=>"101001111",
  13036=>"100001000",
  13037=>"100111111",
  13038=>"001011000",
  13039=>"011110101",
  13040=>"110001000",
  13041=>"000001110",
  13042=>"100000011",
  13043=>"111010011",
  13044=>"100000000",
  13045=>"100100000",
  13046=>"000111010",
  13047=>"010110101",
  13048=>"000011111",
  13049=>"110111110",
  13050=>"111111011",
  13051=>"000001111",
  13052=>"000011101",
  13053=>"100111110",
  13054=>"111001100",
  13055=>"011010000",
  13056=>"101001000",
  13057=>"010011110",
  13058=>"000100110",
  13059=>"110010001",
  13060=>"011111110",
  13061=>"101100011",
  13062=>"010000011",
  13063=>"000101011",
  13064=>"011110100",
  13065=>"111111101",
  13066=>"011011011",
  13067=>"000100000",
  13068=>"000101101",
  13069=>"000001111",
  13070=>"010010111",
  13071=>"111101101",
  13072=>"110110100",
  13073=>"111101101",
  13074=>"001011100",
  13075=>"010110100",
  13076=>"110101011",
  13077=>"110101000",
  13078=>"010000111",
  13079=>"100111111",
  13080=>"011010001",
  13081=>"001011101",
  13082=>"000010111",
  13083=>"010010000",
  13084=>"111000011",
  13085=>"110110010",
  13086=>"100010110",
  13087=>"011010110",
  13088=>"000001010",
  13089=>"101000011",
  13090=>"010110101",
  13091=>"101001000",
  13092=>"111100000",
  13093=>"101010000",
  13094=>"110111011",
  13095=>"110000001",
  13096=>"010001100",
  13097=>"101001111",
  13098=>"000010101",
  13099=>"111010110",
  13100=>"110111111",
  13101=>"000011010",
  13102=>"000111000",
  13103=>"101110001",
  13104=>"100111010",
  13105=>"100010000",
  13106=>"010111000",
  13107=>"000001110",
  13108=>"110010111",
  13109=>"100000101",
  13110=>"110101011",
  13111=>"111010010",
  13112=>"000000001",
  13113=>"010111000",
  13114=>"011011100",
  13115=>"000011001",
  13116=>"101101100",
  13117=>"110010000",
  13118=>"110000000",
  13119=>"111111000",
  13120=>"100101001",
  13121=>"101001111",
  13122=>"110001111",
  13123=>"100100100",
  13124=>"001000100",
  13125=>"111010111",
  13126=>"000001011",
  13127=>"001110101",
  13128=>"010101011",
  13129=>"100011111",
  13130=>"011000010",
  13131=>"100011010",
  13132=>"000110111",
  13133=>"110100010",
  13134=>"010000000",
  13135=>"000100110",
  13136=>"110101011",
  13137=>"001000100",
  13138=>"010100011",
  13139=>"010110100",
  13140=>"110011100",
  13141=>"101111111",
  13142=>"011101100",
  13143=>"111000011",
  13144=>"111111010",
  13145=>"111110101",
  13146=>"001001010",
  13147=>"011110000",
  13148=>"100001101",
  13149=>"000110111",
  13150=>"010101000",
  13151=>"000101100",
  13152=>"100001100",
  13153=>"101001101",
  13154=>"101010000",
  13155=>"000000111",
  13156=>"000000011",
  13157=>"101000001",
  13158=>"110011011",
  13159=>"010001011",
  13160=>"101110011",
  13161=>"100101111",
  13162=>"010010010",
  13163=>"000000101",
  13164=>"110010100",
  13165=>"000000001",
  13166=>"110010110",
  13167=>"011111110",
  13168=>"111101001",
  13169=>"010011101",
  13170=>"101101100",
  13171=>"010001111",
  13172=>"011001011",
  13173=>"001010110",
  13174=>"000011100",
  13175=>"110000000",
  13176=>"011111111",
  13177=>"110111000",
  13178=>"100100011",
  13179=>"000111001",
  13180=>"111000100",
  13181=>"100101001",
  13182=>"101000001",
  13183=>"011111110",
  13184=>"100101011",
  13185=>"100100101",
  13186=>"110010011",
  13187=>"011001101",
  13188=>"001100010",
  13189=>"011111000",
  13190=>"110101010",
  13191=>"000001011",
  13192=>"000100101",
  13193=>"000110011",
  13194=>"111001000",
  13195=>"110010011",
  13196=>"101110101",
  13197=>"101011011",
  13198=>"010001011",
  13199=>"000100101",
  13200=>"100100001",
  13201=>"110111101",
  13202=>"010110010",
  13203=>"101110111",
  13204=>"001111110",
  13205=>"100000101",
  13206=>"001011001",
  13207=>"010100010",
  13208=>"011000111",
  13209=>"111100011",
  13210=>"000000000",
  13211=>"010010000",
  13212=>"011110110",
  13213=>"101100001",
  13214=>"110111001",
  13215=>"010101111",
  13216=>"010011111",
  13217=>"010101101",
  13218=>"110011001",
  13219=>"001000100",
  13220=>"001000010",
  13221=>"010000011",
  13222=>"000101101",
  13223=>"001100101",
  13224=>"011010111",
  13225=>"101100000",
  13226=>"101011100",
  13227=>"001001110",
  13228=>"100101011",
  13229=>"100111001",
  13230=>"010100101",
  13231=>"010111001",
  13232=>"111100110",
  13233=>"000000110",
  13234=>"110110111",
  13235=>"110111001",
  13236=>"111101101",
  13237=>"111110000",
  13238=>"101110101",
  13239=>"101000111",
  13240=>"101011010",
  13241=>"001111001",
  13242=>"001010100",
  13243=>"011000110",
  13244=>"110100010",
  13245=>"010000101",
  13246=>"000111110",
  13247=>"100001000",
  13248=>"111101101",
  13249=>"000000001",
  13250=>"010111111",
  13251=>"101011101",
  13252=>"100000011",
  13253=>"101001101",
  13254=>"001011000",
  13255=>"111101110",
  13256=>"011101100",
  13257=>"111000010",
  13258=>"101011111",
  13259=>"100110110",
  13260=>"110011110",
  13261=>"001000000",
  13262=>"101100010",
  13263=>"111101110",
  13264=>"100000010",
  13265=>"001000011",
  13266=>"100110111",
  13267=>"011011010",
  13268=>"010100000",
  13269=>"111011011",
  13270=>"001100101",
  13271=>"001110101",
  13272=>"010111011",
  13273=>"000100000",
  13274=>"111101001",
  13275=>"110110011",
  13276=>"111011001",
  13277=>"111111110",
  13278=>"000000011",
  13279=>"010010100",
  13280=>"011100101",
  13281=>"111101001",
  13282=>"011001001",
  13283=>"101101001",
  13284=>"100011010",
  13285=>"010100100",
  13286=>"111011100",
  13287=>"000000010",
  13288=>"010010110",
  13289=>"010000000",
  13290=>"101000000",
  13291=>"111011001",
  13292=>"001100100",
  13293=>"011011010",
  13294=>"011010010",
  13295=>"101011101",
  13296=>"001000011",
  13297=>"111011100",
  13298=>"000010101",
  13299=>"101101011",
  13300=>"011010111",
  13301=>"001110110",
  13302=>"111000101",
  13303=>"111110000",
  13304=>"011000001",
  13305=>"001000101",
  13306=>"000111011",
  13307=>"110110101",
  13308=>"000001101",
  13309=>"010110010",
  13310=>"001001001",
  13311=>"011100010",
  13312=>"101111001",
  13313=>"111111111",
  13314=>"110001010",
  13315=>"000001010",
  13316=>"100111110",
  13317=>"100101111",
  13318=>"111111101",
  13319=>"011111110",
  13320=>"111111011",
  13321=>"110111111",
  13322=>"010001110",
  13323=>"110101101",
  13324=>"101001000",
  13325=>"001011111",
  13326=>"011000000",
  13327=>"101111000",
  13328=>"100110101",
  13329=>"011001100",
  13330=>"010001000",
  13331=>"001001101",
  13332=>"100110110",
  13333=>"010000011",
  13334=>"011111001",
  13335=>"010011100",
  13336=>"010010100",
  13337=>"010111101",
  13338=>"101011011",
  13339=>"101001111",
  13340=>"111100110",
  13341=>"110000001",
  13342=>"011111110",
  13343=>"100011001",
  13344=>"111101011",
  13345=>"000011101",
  13346=>"100110100",
  13347=>"001010000",
  13348=>"101010010",
  13349=>"001111000",
  13350=>"110111100",
  13351=>"100001000",
  13352=>"010100011",
  13353=>"100110010",
  13354=>"001100000",
  13355=>"011110100",
  13356=>"000010011",
  13357=>"010101100",
  13358=>"001110000",
  13359=>"010111101",
  13360=>"100110101",
  13361=>"111100011",
  13362=>"110100000",
  13363=>"010110001",
  13364=>"101001001",
  13365=>"001101100",
  13366=>"100101101",
  13367=>"100111101",
  13368=>"001000111",
  13369=>"101111110",
  13370=>"111001111",
  13371=>"010011010",
  13372=>"010000110",
  13373=>"111000111",
  13374=>"111000101",
  13375=>"001010101",
  13376=>"111000011",
  13377=>"101001111",
  13378=>"000000110",
  13379=>"001100111",
  13380=>"111101010",
  13381=>"001111110",
  13382=>"010111010",
  13383=>"101101010",
  13384=>"001001110",
  13385=>"110110011",
  13386=>"101110100",
  13387=>"001100110",
  13388=>"000111010",
  13389=>"010000100",
  13390=>"000011000",
  13391=>"000111101",
  13392=>"001001000",
  13393=>"010011100",
  13394=>"010001110",
  13395=>"101111001",
  13396=>"110111000",
  13397=>"111110000",
  13398=>"111111000",
  13399=>"010100101",
  13400=>"000101011",
  13401=>"101111110",
  13402=>"011000110",
  13403=>"000111101",
  13404=>"111001111",
  13405=>"110010100",
  13406=>"011000101",
  13407=>"010000010",
  13408=>"000101000",
  13409=>"011110011",
  13410=>"011001001",
  13411=>"000111101",
  13412=>"100001100",
  13413=>"100000010",
  13414=>"000011000",
  13415=>"001110101",
  13416=>"001111010",
  13417=>"000000101",
  13418=>"111110100",
  13419=>"100110010",
  13420=>"011100110",
  13421=>"110000001",
  13422=>"011011110",
  13423=>"101000111",
  13424=>"000010100",
  13425=>"011100100",
  13426=>"000000100",
  13427=>"001000100",
  13428=>"100000101",
  13429=>"111110100",
  13430=>"100010111",
  13431=>"010010101",
  13432=>"111011001",
  13433=>"111111111",
  13434=>"010110111",
  13435=>"001111110",
  13436=>"000100001",
  13437=>"101000000",
  13438=>"111010011",
  13439=>"100000001",
  13440=>"110100001",
  13441=>"110000110",
  13442=>"111011111",
  13443=>"100110111",
  13444=>"011111011",
  13445=>"000100101",
  13446=>"011110010",
  13447=>"010010101",
  13448=>"011100000",
  13449=>"010000010",
  13450=>"011001100",
  13451=>"000101000",
  13452=>"110100000",
  13453=>"111110101",
  13454=>"010101111",
  13455=>"110001111",
  13456=>"100110101",
  13457=>"000011001",
  13458=>"101010100",
  13459=>"010000100",
  13460=>"000011010",
  13461=>"100101110",
  13462=>"100110111",
  13463=>"001010110",
  13464=>"101010111",
  13465=>"000001100",
  13466=>"100010110",
  13467=>"111100100",
  13468=>"011111001",
  13469=>"100111010",
  13470=>"001100101",
  13471=>"001011111",
  13472=>"011000000",
  13473=>"011010111",
  13474=>"000100110",
  13475=>"101010011",
  13476=>"001000010",
  13477=>"101010011",
  13478=>"110100000",
  13479=>"100000111",
  13480=>"000011101",
  13481=>"110011101",
  13482=>"110100001",
  13483=>"100001011",
  13484=>"000101001",
  13485=>"111111010",
  13486=>"011011111",
  13487=>"000001011",
  13488=>"000100011",
  13489=>"010100001",
  13490=>"110101001",
  13491=>"111011111",
  13492=>"101011101",
  13493=>"100100110",
  13494=>"111000110",
  13495=>"101011111",
  13496=>"111010100",
  13497=>"101011101",
  13498=>"010100110",
  13499=>"000111101",
  13500=>"011100011",
  13501=>"101111000",
  13502=>"011100111",
  13503=>"011001110",
  13504=>"011110111",
  13505=>"110100110",
  13506=>"110101001",
  13507=>"000001100",
  13508=>"111111010",
  13509=>"100111111",
  13510=>"010000100",
  13511=>"011110001",
  13512=>"000010010",
  13513=>"101100100",
  13514=>"001100110",
  13515=>"000001101",
  13516=>"100000100",
  13517=>"111100010",
  13518=>"000110010",
  13519=>"010110110",
  13520=>"101010011",
  13521=>"010111100",
  13522=>"110010000",
  13523=>"110010100",
  13524=>"011111010",
  13525=>"101000001",
  13526=>"111001100",
  13527=>"001000000",
  13528=>"001000000",
  13529=>"100110100",
  13530=>"011111111",
  13531=>"100101110",
  13532=>"101011000",
  13533=>"101011101",
  13534=>"010010010",
  13535=>"010000110",
  13536=>"001100001",
  13537=>"011111000",
  13538=>"110111111",
  13539=>"011100100",
  13540=>"100000000",
  13541=>"110000111",
  13542=>"011100110",
  13543=>"001111100",
  13544=>"001100010",
  13545=>"000101001",
  13546=>"100001000",
  13547=>"111011000",
  13548=>"001000000",
  13549=>"011000110",
  13550=>"011000011",
  13551=>"011110000",
  13552=>"111011110",
  13553=>"100001101",
  13554=>"101111100",
  13555=>"100001000",
  13556=>"100101000",
  13557=>"101111011",
  13558=>"111110110",
  13559=>"001111000",
  13560=>"111001100",
  13561=>"001001010",
  13562=>"110000111",
  13563=>"100111110",
  13564=>"110001001",
  13565=>"011101101",
  13566=>"001011111",
  13567=>"111100100",
  13568=>"011010001",
  13569=>"110110010",
  13570=>"110001111",
  13571=>"111001110",
  13572=>"001010000",
  13573=>"100100000",
  13574=>"111010011",
  13575=>"111001111",
  13576=>"010101001",
  13577=>"010000001",
  13578=>"101100001",
  13579=>"000000000",
  13580=>"100001111",
  13581=>"010001001",
  13582=>"110100101",
  13583=>"001110111",
  13584=>"100001110",
  13585=>"111110100",
  13586=>"001101010",
  13587=>"110000000",
  13588=>"011111010",
  13589=>"000000111",
  13590=>"110101000",
  13591=>"011111110",
  13592=>"011010100",
  13593=>"000111110",
  13594=>"100010000",
  13595=>"111000100",
  13596=>"000001101",
  13597=>"101011111",
  13598=>"110100010",
  13599=>"111010101",
  13600=>"101101111",
  13601=>"111011110",
  13602=>"101010110",
  13603=>"011100110",
  13604=>"000000001",
  13605=>"101101101",
  13606=>"001100000",
  13607=>"010001111",
  13608=>"000001101",
  13609=>"010000101",
  13610=>"001101111",
  13611=>"011001001",
  13612=>"011101001",
  13613=>"000000011",
  13614=>"101001011",
  13615=>"100000001",
  13616=>"101010101",
  13617=>"001000110",
  13618=>"111000101",
  13619=>"100001001",
  13620=>"111000100",
  13621=>"001000001",
  13622=>"110111110",
  13623=>"000010100",
  13624=>"010000110",
  13625=>"011000111",
  13626=>"001001110",
  13627=>"110110111",
  13628=>"111101111",
  13629=>"010000001",
  13630=>"100011000",
  13631=>"101000110",
  13632=>"001111011",
  13633=>"101001100",
  13634=>"010111000",
  13635=>"100010010",
  13636=>"110100010",
  13637=>"001101110",
  13638=>"001100000",
  13639=>"100100100",
  13640=>"111110100",
  13641=>"100010101",
  13642=>"001000111",
  13643=>"010101101",
  13644=>"011001100",
  13645=>"101001001",
  13646=>"101111111",
  13647=>"111111000",
  13648=>"111111100",
  13649=>"101001000",
  13650=>"100001011",
  13651=>"111101011",
  13652=>"111111011",
  13653=>"001111100",
  13654=>"111010001",
  13655=>"011111010",
  13656=>"010010111",
  13657=>"100101011",
  13658=>"000101100",
  13659=>"000100010",
  13660=>"110100111",
  13661=>"000101100",
  13662=>"110101101",
  13663=>"111111101",
  13664=>"011111010",
  13665=>"110100100",
  13666=>"101010001",
  13667=>"100101101",
  13668=>"100111101",
  13669=>"101001010",
  13670=>"010111011",
  13671=>"100010001",
  13672=>"010100110",
  13673=>"110111111",
  13674=>"010011111",
  13675=>"101101100",
  13676=>"100001010",
  13677=>"010101110",
  13678=>"100010100",
  13679=>"111011000",
  13680=>"100011000",
  13681=>"011111011",
  13682=>"110010101",
  13683=>"110001011",
  13684=>"011000000",
  13685=>"001110011",
  13686=>"010000011",
  13687=>"100000010",
  13688=>"010011010",
  13689=>"110101111",
  13690=>"010011110",
  13691=>"101001000",
  13692=>"110110000",
  13693=>"011111010",
  13694=>"111101110",
  13695=>"000100000",
  13696=>"101011001",
  13697=>"101010101",
  13698=>"010000000",
  13699=>"110001100",
  13700=>"000100100",
  13701=>"000101111",
  13702=>"110001100",
  13703=>"100111110",
  13704=>"110011011",
  13705=>"101100101",
  13706=>"110110011",
  13707=>"010011101",
  13708=>"010001000",
  13709=>"111010101",
  13710=>"111111101",
  13711=>"111110011",
  13712=>"001000000",
  13713=>"101110001",
  13714=>"110101001",
  13715=>"001111010",
  13716=>"101101010",
  13717=>"001001000",
  13718=>"000111000",
  13719=>"001000110",
  13720=>"100111111",
  13721=>"101000111",
  13722=>"101100100",
  13723=>"000110101",
  13724=>"001101100",
  13725=>"100110010",
  13726=>"010111101",
  13727=>"000001011",
  13728=>"101001001",
  13729=>"000011001",
  13730=>"111010110",
  13731=>"110111000",
  13732=>"100011101",
  13733=>"101000011",
  13734=>"011101101",
  13735=>"101100010",
  13736=>"000010000",
  13737=>"010011010",
  13738=>"101111011",
  13739=>"010111101",
  13740=>"110001110",
  13741=>"010111010",
  13742=>"101011101",
  13743=>"100001000",
  13744=>"101111111",
  13745=>"011111001",
  13746=>"001101000",
  13747=>"111111100",
  13748=>"000010101",
  13749=>"110111010",
  13750=>"111110011",
  13751=>"101110010",
  13752=>"111000010",
  13753=>"000010101",
  13754=>"001110111",
  13755=>"000000010",
  13756=>"000001110",
  13757=>"010001011",
  13758=>"010011100",
  13759=>"010111000",
  13760=>"110000110",
  13761=>"000101011",
  13762=>"111110010",
  13763=>"110111010",
  13764=>"010010011",
  13765=>"110010011",
  13766=>"110100101",
  13767=>"101001011",
  13768=>"110010111",
  13769=>"111110000",
  13770=>"001000101",
  13771=>"010100010",
  13772=>"101011111",
  13773=>"111101111",
  13774=>"100011111",
  13775=>"110000010",
  13776=>"101001111",
  13777=>"011000001",
  13778=>"110110000",
  13779=>"001110010",
  13780=>"100111100",
  13781=>"001001001",
  13782=>"101110100",
  13783=>"111010010",
  13784=>"100111001",
  13785=>"001110111",
  13786=>"100100110",
  13787=>"011010001",
  13788=>"111001010",
  13789=>"000000001",
  13790=>"110100010",
  13791=>"111101111",
  13792=>"100000000",
  13793=>"101100001",
  13794=>"110110100",
  13795=>"010111110",
  13796=>"101001110",
  13797=>"011110100",
  13798=>"001000100",
  13799=>"010001001",
  13800=>"011101111",
  13801=>"010111101",
  13802=>"110001010",
  13803=>"010100000",
  13804=>"110110000",
  13805=>"000000011",
  13806=>"100100000",
  13807=>"111000001",
  13808=>"001110111",
  13809=>"001101101",
  13810=>"101110101",
  13811=>"101100110",
  13812=>"111110000",
  13813=>"011011011",
  13814=>"101000010",
  13815=>"111110101",
  13816=>"100010111",
  13817=>"011010111",
  13818=>"000001010",
  13819=>"110111110",
  13820=>"111111110",
  13821=>"110000111",
  13822=>"101010001",
  13823=>"000001001",
  13824=>"011010001",
  13825=>"110011110",
  13826=>"001000000",
  13827=>"110010111",
  13828=>"111111111",
  13829=>"010101000",
  13830=>"011001110",
  13831=>"010100101",
  13832=>"101001011",
  13833=>"000101010",
  13834=>"011010010",
  13835=>"111001000",
  13836=>"100100101",
  13837=>"100100011",
  13838=>"000110000",
  13839=>"111010101",
  13840=>"101110001",
  13841=>"010011111",
  13842=>"000111100",
  13843=>"001101010",
  13844=>"111000101",
  13845=>"000000100",
  13846=>"000101110",
  13847=>"001011110",
  13848=>"000111001",
  13849=>"011101000",
  13850=>"111111100",
  13851=>"100100000",
  13852=>"100010111",
  13853=>"010001001",
  13854=>"010100101",
  13855=>"001010111",
  13856=>"100000001",
  13857=>"001011000",
  13858=>"110100110",
  13859=>"101011000",
  13860=>"000011111",
  13861=>"101111011",
  13862=>"000101111",
  13863=>"111100001",
  13864=>"001110011",
  13865=>"111101111",
  13866=>"000010011",
  13867=>"001011101",
  13868=>"100100010",
  13869=>"010101011",
  13870=>"011111000",
  13871=>"010111010",
  13872=>"011110111",
  13873=>"000111001",
  13874=>"001101001",
  13875=>"010010101",
  13876=>"101011100",
  13877=>"011011101",
  13878=>"100100000",
  13879=>"001011110",
  13880=>"001000000",
  13881=>"100101111",
  13882=>"010001101",
  13883=>"110011101",
  13884=>"000010111",
  13885=>"001101011",
  13886=>"001101010",
  13887=>"110100100",
  13888=>"011011010",
  13889=>"101000011",
  13890=>"110000000",
  13891=>"100010110",
  13892=>"111110110",
  13893=>"111111100",
  13894=>"011001000",
  13895=>"101011011",
  13896=>"000000010",
  13897=>"000001110",
  13898=>"000001001",
  13899=>"000011010",
  13900=>"001011111",
  13901=>"111100010",
  13902=>"001100011",
  13903=>"001000110",
  13904=>"010011101",
  13905=>"110011111",
  13906=>"000001111",
  13907=>"000111010",
  13908=>"001000110",
  13909=>"000110110",
  13910=>"111010101",
  13911=>"111110011",
  13912=>"100011000",
  13913=>"011111010",
  13914=>"101110101",
  13915=>"111010110",
  13916=>"010000111",
  13917=>"000000010",
  13918=>"001100111",
  13919=>"000000111",
  13920=>"100001111",
  13921=>"111111010",
  13922=>"000100001",
  13923=>"010100001",
  13924=>"110111110",
  13925=>"110110011",
  13926=>"111010111",
  13927=>"010111111",
  13928=>"101110100",
  13929=>"111010110",
  13930=>"000010110",
  13931=>"001000100",
  13932=>"001010001",
  13933=>"111110010",
  13934=>"001001001",
  13935=>"000100110",
  13936=>"010000000",
  13937=>"001100110",
  13938=>"011001101",
  13939=>"010000111",
  13940=>"011000001",
  13941=>"110000100",
  13942=>"001001110",
  13943=>"111111100",
  13944=>"110001100",
  13945=>"111001001",
  13946=>"111110100",
  13947=>"011011100",
  13948=>"110100010",
  13949=>"000000111",
  13950=>"000010101",
  13951=>"111110001",
  13952=>"110110001",
  13953=>"110011100",
  13954=>"111011010",
  13955=>"010000100",
  13956=>"110000111",
  13957=>"000010001",
  13958=>"100110000",
  13959=>"010100111",
  13960=>"100101111",
  13961=>"011001100",
  13962=>"001111000",
  13963=>"000010011",
  13964=>"011110111",
  13965=>"000010101",
  13966=>"000110100",
  13967=>"111011100",
  13968=>"010010001",
  13969=>"110101110",
  13970=>"010001000",
  13971=>"100010011",
  13972=>"111111111",
  13973=>"001111001",
  13974=>"011001111",
  13975=>"100111111",
  13976=>"010111111",
  13977=>"011110101",
  13978=>"010110010",
  13979=>"101110110",
  13980=>"100010100",
  13981=>"110011000",
  13982=>"101100110",
  13983=>"111000111",
  13984=>"001000000",
  13985=>"010001001",
  13986=>"110111110",
  13987=>"011110100",
  13988=>"001001110",
  13989=>"001100010",
  13990=>"110100010",
  13991=>"011101110",
  13992=>"100011110",
  13993=>"010000000",
  13994=>"010100000",
  13995=>"001000101",
  13996=>"000111111",
  13997=>"000000110",
  13998=>"101100111",
  13999=>"111110111",
  14000=>"011011001",
  14001=>"111111101",
  14002=>"111011010",
  14003=>"000110011",
  14004=>"100000001",
  14005=>"100000101",
  14006=>"110010011",
  14007=>"010000101",
  14008=>"101110100",
  14009=>"100111001",
  14010=>"010110001",
  14011=>"101011111",
  14012=>"001001111",
  14013=>"111100101",
  14014=>"000010000",
  14015=>"011110010",
  14016=>"001111011",
  14017=>"011010101",
  14018=>"010011011",
  14019=>"011010110",
  14020=>"001000111",
  14021=>"110111111",
  14022=>"010010000",
  14023=>"001001000",
  14024=>"000001010",
  14025=>"011101011",
  14026=>"011000011",
  14027=>"101010010",
  14028=>"100001010",
  14029=>"011100101",
  14030=>"110010011",
  14031=>"101101001",
  14032=>"101000100",
  14033=>"001000101",
  14034=>"111101001",
  14035=>"010111110",
  14036=>"100000001",
  14037=>"100101110",
  14038=>"001000101",
  14039=>"010011100",
  14040=>"011101000",
  14041=>"101001000",
  14042=>"001000010",
  14043=>"100100011",
  14044=>"111000010",
  14045=>"011001101",
  14046=>"011111000",
  14047=>"000111000",
  14048=>"100101110",
  14049=>"000010110",
  14050=>"010011111",
  14051=>"111011001",
  14052=>"011000100",
  14053=>"111110110",
  14054=>"010111010",
  14055=>"010000101",
  14056=>"101110011",
  14057=>"111101000",
  14058=>"100000100",
  14059=>"001011110",
  14060=>"000010100",
  14061=>"000100011",
  14062=>"110101000",
  14063=>"110000111",
  14064=>"000101100",
  14065=>"101000110",
  14066=>"001100101",
  14067=>"110101101",
  14068=>"101001110",
  14069=>"110000010",
  14070=>"110010001",
  14071=>"101001101",
  14072=>"100100100",
  14073=>"011000100",
  14074=>"001101101",
  14075=>"100011111",
  14076=>"010110000",
  14077=>"100101000",
  14078=>"011011001",
  14079=>"011110010",
  14080=>"000010111",
  14081=>"111111001",
  14082=>"001111111",
  14083=>"110110111",
  14084=>"110000000",
  14085=>"011111111",
  14086=>"101000001",
  14087=>"101101010",
  14088=>"110111010",
  14089=>"010110010",
  14090=>"101111101",
  14091=>"110110110",
  14092=>"111001010",
  14093=>"000101101",
  14094=>"101100000",
  14095=>"011011001",
  14096=>"111000100",
  14097=>"011101010",
  14098=>"110100100",
  14099=>"010010100",
  14100=>"110000010",
  14101=>"100000100",
  14102=>"110001000",
  14103=>"000000100",
  14104=>"100001111",
  14105=>"101001001",
  14106=>"000010101",
  14107=>"100011000",
  14108=>"111110111",
  14109=>"001100011",
  14110=>"010110110",
  14111=>"101100110",
  14112=>"000010011",
  14113=>"111100111",
  14114=>"010000101",
  14115=>"111101010",
  14116=>"100110000",
  14117=>"001101001",
  14118=>"110011111",
  14119=>"110001100",
  14120=>"101111111",
  14121=>"111011111",
  14122=>"000000110",
  14123=>"100111000",
  14124=>"100011011",
  14125=>"000001101",
  14126=>"000100110",
  14127=>"101010000",
  14128=>"010110011",
  14129=>"100101001",
  14130=>"101111111",
  14131=>"110010111",
  14132=>"010111000",
  14133=>"111101010",
  14134=>"011000010",
  14135=>"000000000",
  14136=>"001100010",
  14137=>"110011111",
  14138=>"000010111",
  14139=>"110110110",
  14140=>"010011110",
  14141=>"111111000",
  14142=>"000001001",
  14143=>"010100011",
  14144=>"111100000",
  14145=>"101011100",
  14146=>"001001011",
  14147=>"001000011",
  14148=>"110000110",
  14149=>"100011100",
  14150=>"100010100",
  14151=>"011001010",
  14152=>"101110010",
  14153=>"010011011",
  14154=>"011100001",
  14155=>"000010000",
  14156=>"010010111",
  14157=>"100010000",
  14158=>"111001111",
  14159=>"000101111",
  14160=>"100001100",
  14161=>"100000010",
  14162=>"010111100",
  14163=>"100001011",
  14164=>"101101101",
  14165=>"011110001",
  14166=>"010001101",
  14167=>"010100111",
  14168=>"100101000",
  14169=>"111000111",
  14170=>"001001001",
  14171=>"000101010",
  14172=>"010011010",
  14173=>"011100101",
  14174=>"111100010",
  14175=>"100000111",
  14176=>"011010111",
  14177=>"111000001",
  14178=>"100010010",
  14179=>"000101001",
  14180=>"001001010",
  14181=>"100010110",
  14182=>"010110111",
  14183=>"110000010",
  14184=>"111000101",
  14185=>"000100110",
  14186=>"011001001",
  14187=>"000110110",
  14188=>"101101100",
  14189=>"011000100",
  14190=>"001010111",
  14191=>"101001110",
  14192=>"110010110",
  14193=>"010101100",
  14194=>"001010001",
  14195=>"000010001",
  14196=>"111101101",
  14197=>"000111101",
  14198=>"010011101",
  14199=>"100101010",
  14200=>"010001000",
  14201=>"010101001",
  14202=>"101111001",
  14203=>"111101000",
  14204=>"110111101",
  14205=>"110110100",
  14206=>"001001111",
  14207=>"000011011",
  14208=>"000001001",
  14209=>"100011111",
  14210=>"101001011",
  14211=>"000101100",
  14212=>"111111110",
  14213=>"001001100",
  14214=>"111011011",
  14215=>"001100000",
  14216=>"011000000",
  14217=>"111111101",
  14218=>"010001010",
  14219=>"101100110",
  14220=>"110010010",
  14221=>"100010110",
  14222=>"110000101",
  14223=>"111111110",
  14224=>"011100111",
  14225=>"101001000",
  14226=>"011010101",
  14227=>"001111101",
  14228=>"101110100",
  14229=>"000100010",
  14230=>"010101000",
  14231=>"101100000",
  14232=>"011101111",
  14233=>"010101001",
  14234=>"101001110",
  14235=>"100001111",
  14236=>"110100011",
  14237=>"101010111",
  14238=>"100110111",
  14239=>"111001101",
  14240=>"001111111",
  14241=>"010111110",
  14242=>"000101100",
  14243=>"000001011",
  14244=>"011111010",
  14245=>"111110011",
  14246=>"001001101",
  14247=>"111011011",
  14248=>"110111100",
  14249=>"101011000",
  14250=>"111111110",
  14251=>"110000101",
  14252=>"101100100",
  14253=>"100100101",
  14254=>"000110001",
  14255=>"010000101",
  14256=>"101010010",
  14257=>"011010110",
  14258=>"110100000",
  14259=>"101101101",
  14260=>"000111011",
  14261=>"101000001",
  14262=>"111110110",
  14263=>"010001110",
  14264=>"100001100",
  14265=>"001110110",
  14266=>"101110011",
  14267=>"100011001",
  14268=>"000001000",
  14269=>"001010010",
  14270=>"000011010",
  14271=>"000000011",
  14272=>"101011001",
  14273=>"001111111",
  14274=>"000001010",
  14275=>"110010111",
  14276=>"101010000",
  14277=>"000011110",
  14278=>"001011000",
  14279=>"010011011",
  14280=>"001101000",
  14281=>"110101001",
  14282=>"011111100",
  14283=>"001011010",
  14284=>"111111001",
  14285=>"111000010",
  14286=>"110001010",
  14287=>"011111010",
  14288=>"100100011",
  14289=>"110110010",
  14290=>"000000011",
  14291=>"000001001",
  14292=>"110110000",
  14293=>"010110111",
  14294=>"111101100",
  14295=>"111000010",
  14296=>"111100001",
  14297=>"001001111",
  14298=>"111100111",
  14299=>"100110010",
  14300=>"111001100",
  14301=>"100110111",
  14302=>"001101100",
  14303=>"111001101",
  14304=>"000011001",
  14305=>"000000110",
  14306=>"000000010",
  14307=>"110001100",
  14308=>"011100000",
  14309=>"100101111",
  14310=>"010100010",
  14311=>"100010010",
  14312=>"111101001",
  14313=>"001010110",
  14314=>"111010001",
  14315=>"111000100",
  14316=>"100111000",
  14317=>"110111011",
  14318=>"011000111",
  14319=>"101011001",
  14320=>"001100110",
  14321=>"100111110",
  14322=>"111101101",
  14323=>"110011111",
  14324=>"111101100",
  14325=>"111110110",
  14326=>"000011011",
  14327=>"111100010",
  14328=>"000001000",
  14329=>"011011101",
  14330=>"000001111",
  14331=>"000100010",
  14332=>"110101101",
  14333=>"101000010",
  14334=>"010101111",
  14335=>"001111011",
  14336=>"111110110",
  14337=>"100001100",
  14338=>"000010110",
  14339=>"111011101",
  14340=>"010110100",
  14341=>"100100111",
  14342=>"000010001",
  14343=>"111011001",
  14344=>"010100001",
  14345=>"000010110",
  14346=>"110110111",
  14347=>"011011111",
  14348=>"111000011",
  14349=>"100100001",
  14350=>"010001001",
  14351=>"110010011",
  14352=>"110011100",
  14353=>"100111111",
  14354=>"100110001",
  14355=>"000001000",
  14356=>"100101111",
  14357=>"000000100",
  14358=>"111010110",
  14359=>"001000000",
  14360=>"000011100",
  14361=>"010101000",
  14362=>"110101111",
  14363=>"111010001",
  14364=>"001100001",
  14365=>"101111011",
  14366=>"100000110",
  14367=>"101111010",
  14368=>"100001011",
  14369=>"100001110",
  14370=>"101100000",
  14371=>"010100101",
  14372=>"111010101",
  14373=>"111100000",
  14374=>"111000100",
  14375=>"000000010",
  14376=>"000110111",
  14377=>"111110010",
  14378=>"101011101",
  14379=>"111101001",
  14380=>"011010111",
  14381=>"110001100",
  14382=>"111001101",
  14383=>"101100001",
  14384=>"110011010",
  14385=>"011110001",
  14386=>"101111110",
  14387=>"000111111",
  14388=>"000100111",
  14389=>"001000111",
  14390=>"001011010",
  14391=>"101010111",
  14392=>"110111011",
  14393=>"110111000",
  14394=>"110000000",
  14395=>"010001111",
  14396=>"000001011",
  14397=>"111010010",
  14398=>"110010111",
  14399=>"100011001",
  14400=>"000111110",
  14401=>"010101111",
  14402=>"000111111",
  14403=>"001000001",
  14404=>"000011000",
  14405=>"010010111",
  14406=>"001000101",
  14407=>"000100011",
  14408=>"100011110",
  14409=>"111111110",
  14410=>"111111110",
  14411=>"110111101",
  14412=>"000101010",
  14413=>"000001011",
  14414=>"111000011",
  14415=>"110111001",
  14416=>"001011101",
  14417=>"001100000",
  14418=>"000010110",
  14419=>"010011011",
  14420=>"101111111",
  14421=>"100001101",
  14422=>"100000101",
  14423=>"101101010",
  14424=>"111101011",
  14425=>"010010101",
  14426=>"111000011",
  14427=>"010111000",
  14428=>"100100111",
  14429=>"100001010",
  14430=>"000001011",
  14431=>"011000110",
  14432=>"110110100",
  14433=>"100010000",
  14434=>"000001010",
  14435=>"111000000",
  14436=>"001001110",
  14437=>"110011000",
  14438=>"000001000",
  14439=>"100000111",
  14440=>"000001111",
  14441=>"100101001",
  14442=>"111101010",
  14443=>"001000001",
  14444=>"110110101",
  14445=>"010101101",
  14446=>"000000010",
  14447=>"000010101",
  14448=>"010001000",
  14449=>"110110110",
  14450=>"001010011",
  14451=>"110000001",
  14452=>"011111011",
  14453=>"010000001",
  14454=>"011000000",
  14455=>"111010001",
  14456=>"001000011",
  14457=>"010001100",
  14458=>"111010000",
  14459=>"010000010",
  14460=>"000100110",
  14461=>"001101011",
  14462=>"001000101",
  14463=>"011111011",
  14464=>"001100111",
  14465=>"000100111",
  14466=>"111110000",
  14467=>"001000010",
  14468=>"100110001",
  14469=>"001011101",
  14470=>"010001111",
  14471=>"011110001",
  14472=>"101110010",
  14473=>"111110111",
  14474=>"110011010",
  14475=>"111101010",
  14476=>"010111010",
  14477=>"101001011",
  14478=>"100010100",
  14479=>"001111101",
  14480=>"110111111",
  14481=>"001001101",
  14482=>"101100101",
  14483=>"111000110",
  14484=>"000000110",
  14485=>"001011100",
  14486=>"000110100",
  14487=>"010010101",
  14488=>"110100111",
  14489=>"000011110",
  14490=>"111010010",
  14491=>"010100101",
  14492=>"010101001",
  14493=>"100011110",
  14494=>"111101010",
  14495=>"010100110",
  14496=>"111011011",
  14497=>"100111110",
  14498=>"000001101",
  14499=>"101011110",
  14500=>"010100100",
  14501=>"110100111",
  14502=>"101101100",
  14503=>"010100000",
  14504=>"001111100",
  14505=>"001000110",
  14506=>"110010110",
  14507=>"011001101",
  14508=>"001101100",
  14509=>"011000000",
  14510=>"110000010",
  14511=>"110110011",
  14512=>"010010001",
  14513=>"110110101",
  14514=>"000101010",
  14515=>"000001000",
  14516=>"010100000",
  14517=>"110110011",
  14518=>"110000001",
  14519=>"010100100",
  14520=>"001000000",
  14521=>"101001011",
  14522=>"101001100",
  14523=>"100010001",
  14524=>"110101110",
  14525=>"011110000",
  14526=>"011110101",
  14527=>"111000001",
  14528=>"010010001",
  14529=>"111100010",
  14530=>"111010100",
  14531=>"111011100",
  14532=>"001010100",
  14533=>"010000000",
  14534=>"101110011",
  14535=>"111110110",
  14536=>"100110101",
  14537=>"101010101",
  14538=>"011111101",
  14539=>"110111010",
  14540=>"111011010",
  14541=>"011010111",
  14542=>"000010010",
  14543=>"010110110",
  14544=>"101001010",
  14545=>"110010110",
  14546=>"000101101",
  14547=>"100100000",
  14548=>"001010100",
  14549=>"110010101",
  14550=>"110010010",
  14551=>"111110101",
  14552=>"110010111",
  14553=>"110000101",
  14554=>"110000000",
  14555=>"010000001",
  14556=>"011000111",
  14557=>"101001010",
  14558=>"000001000",
  14559=>"110101110",
  14560=>"000111101",
  14561=>"011001100",
  14562=>"111111100",
  14563=>"000011011",
  14564=>"000011110",
  14565=>"110100100",
  14566=>"011010000",
  14567=>"001110111",
  14568=>"101100011",
  14569=>"111111001",
  14570=>"101110101",
  14571=>"000011111",
  14572=>"001010110",
  14573=>"110000101",
  14574=>"101001111",
  14575=>"111001000",
  14576=>"001111100",
  14577=>"011111111",
  14578=>"000011001",
  14579=>"100010000",
  14580=>"100100101",
  14581=>"000100110",
  14582=>"010001011",
  14583=>"110101100",
  14584=>"000011101",
  14585=>"110000000",
  14586=>"001110001",
  14587=>"111100011",
  14588=>"001001101",
  14589=>"111000011",
  14590=>"100000101",
  14591=>"000101100",
  14592=>"011111111",
  14593=>"011001001",
  14594=>"001101110",
  14595=>"111100001",
  14596=>"010110010",
  14597=>"001000110",
  14598=>"110001101",
  14599=>"101111011",
  14600=>"000001101",
  14601=>"101001100",
  14602=>"010011000",
  14603=>"111100001",
  14604=>"101010000",
  14605=>"111010010",
  14606=>"101110110",
  14607=>"000000010",
  14608=>"111011111",
  14609=>"101011111",
  14610=>"100000010",
  14611=>"100110011",
  14612=>"000101000",
  14613=>"110111110",
  14614=>"001010011",
  14615=>"001000010",
  14616=>"000100110",
  14617=>"000011011",
  14618=>"010000101",
  14619=>"011101011",
  14620=>"100100101",
  14621=>"111000101",
  14622=>"101001101",
  14623=>"000100100",
  14624=>"001010110",
  14625=>"101001010",
  14626=>"110110011",
  14627=>"001010001",
  14628=>"001111010",
  14629=>"000111011",
  14630=>"000000010",
  14631=>"111001100",
  14632=>"110000010",
  14633=>"110000011",
  14634=>"101001110",
  14635=>"100000000",
  14636=>"100011011",
  14637=>"111011111",
  14638=>"010110010",
  14639=>"100000000",
  14640=>"010110001",
  14641=>"001010010",
  14642=>"111110110",
  14643=>"000100100",
  14644=>"010000100",
  14645=>"011111010",
  14646=>"000000011",
  14647=>"011011011",
  14648=>"111101110",
  14649=>"101110000",
  14650=>"000011001",
  14651=>"001000000",
  14652=>"111100100",
  14653=>"111010011",
  14654=>"011110001",
  14655=>"011101001",
  14656=>"010011110",
  14657=>"111111100",
  14658=>"110010000",
  14659=>"111100010",
  14660=>"111010000",
  14661=>"011110000",
  14662=>"001110011",
  14663=>"110111100",
  14664=>"000110011",
  14665=>"101101101",
  14666=>"000000000",
  14667=>"100100010",
  14668=>"000111011",
  14669=>"001111011",
  14670=>"100110101",
  14671=>"010011111",
  14672=>"110011010",
  14673=>"101110001",
  14674=>"100011011",
  14675=>"001010100",
  14676=>"000100011",
  14677=>"100010010",
  14678=>"000000110",
  14679=>"100001010",
  14680=>"000010001",
  14681=>"000100100",
  14682=>"011010111",
  14683=>"101101000",
  14684=>"011110010",
  14685=>"111111100",
  14686=>"100110011",
  14687=>"011100110",
  14688=>"111001111",
  14689=>"011000100",
  14690=>"001111101",
  14691=>"000010001",
  14692=>"010000010",
  14693=>"000101000",
  14694=>"011011100",
  14695=>"100000100",
  14696=>"110001110",
  14697=>"000101011",
  14698=>"101010000",
  14699=>"111000010",
  14700=>"001010101",
  14701=>"110101111",
  14702=>"101000100",
  14703=>"011101110",
  14704=>"100010100",
  14705=>"011010010",
  14706=>"111101010",
  14707=>"001001001",
  14708=>"110000111",
  14709=>"011001101",
  14710=>"011110110",
  14711=>"101101111",
  14712=>"101110111",
  14713=>"110001001",
  14714=>"111011101",
  14715=>"010011110",
  14716=>"001011001",
  14717=>"111111010",
  14718=>"000010001",
  14719=>"111010110",
  14720=>"100011101",
  14721=>"110101101",
  14722=>"000010111",
  14723=>"011001001",
  14724=>"100110110",
  14725=>"100001010",
  14726=>"100100000",
  14727=>"110110000",
  14728=>"001100111",
  14729=>"000000110",
  14730=>"001000010",
  14731=>"011111110",
  14732=>"010001010",
  14733=>"000010111",
  14734=>"000111001",
  14735=>"000010010",
  14736=>"101010011",
  14737=>"111100011",
  14738=>"001100011",
  14739=>"001111000",
  14740=>"000011010",
  14741=>"010110111",
  14742=>"011100001",
  14743=>"110110001",
  14744=>"001010010",
  14745=>"101111111",
  14746=>"101111111",
  14747=>"111110000",
  14748=>"001100010",
  14749=>"011100111",
  14750=>"011100101",
  14751=>"110010101",
  14752=>"010010010",
  14753=>"110100011",
  14754=>"000101100",
  14755=>"101000010",
  14756=>"011001011",
  14757=>"101101101",
  14758=>"001001100",
  14759=>"000000000",
  14760=>"110110100",
  14761=>"101010010",
  14762=>"000000110",
  14763=>"100100111",
  14764=>"011001010",
  14765=>"110110010",
  14766=>"000001001",
  14767=>"001000110",
  14768=>"111111111",
  14769=>"001110001",
  14770=>"111111010",
  14771=>"111110111",
  14772=>"100100100",
  14773=>"011000011",
  14774=>"011001111",
  14775=>"111100100",
  14776=>"101100111",
  14777=>"000000011",
  14778=>"101000001",
  14779=>"001100000",
  14780=>"011000111",
  14781=>"100010000",
  14782=>"010000001",
  14783=>"001100101",
  14784=>"000011101",
  14785=>"101010011",
  14786=>"111100010",
  14787=>"000011111",
  14788=>"011011000",
  14789=>"100100011",
  14790=>"110101001",
  14791=>"011101111",
  14792=>"011000111",
  14793=>"111101011",
  14794=>"100010000",
  14795=>"101011011",
  14796=>"111001010",
  14797=>"110110111",
  14798=>"110111010",
  14799=>"101101010",
  14800=>"001111000",
  14801=>"111100111",
  14802=>"001101010",
  14803=>"000100111",
  14804=>"011011101",
  14805=>"001101001",
  14806=>"011110110",
  14807=>"101101100",
  14808=>"001001111",
  14809=>"001010000",
  14810=>"111011011",
  14811=>"111011010",
  14812=>"100111000",
  14813=>"101010000",
  14814=>"101110001",
  14815=>"100100010",
  14816=>"100000110",
  14817=>"000000000",
  14818=>"011101100",
  14819=>"111111110",
  14820=>"000001110",
  14821=>"010111001",
  14822=>"010101011",
  14823=>"000000011",
  14824=>"010000100",
  14825=>"011100111",
  14826=>"110100101",
  14827=>"111000001",
  14828=>"101111001",
  14829=>"111000101",
  14830=>"010100010",
  14831=>"101101010",
  14832=>"001001111",
  14833=>"110010111",
  14834=>"111011001",
  14835=>"111101000",
  14836=>"011000100",
  14837=>"010010111",
  14838=>"101000011",
  14839=>"000000100",
  14840=>"100111000",
  14841=>"110000110",
  14842=>"000100101",
  14843=>"010011001",
  14844=>"111000011",
  14845=>"111001000",
  14846=>"100001100",
  14847=>"011101110",
  14848=>"110000110",
  14849=>"001101100",
  14850=>"001100100",
  14851=>"000101100",
  14852=>"001001001",
  14853=>"010000010",
  14854=>"011000010",
  14855=>"111011010",
  14856=>"110110010",
  14857=>"000001010",
  14858=>"000101111",
  14859=>"000001001",
  14860=>"000101101",
  14861=>"111001111",
  14862=>"000001000",
  14863=>"000010101",
  14864=>"110101010",
  14865=>"001011001",
  14866=>"111100110",
  14867=>"001000000",
  14868=>"000011010",
  14869=>"101101110",
  14870=>"110111110",
  14871=>"000111100",
  14872=>"000000010",
  14873=>"111010110",
  14874=>"110011100",
  14875=>"001011010",
  14876=>"010011000",
  14877=>"010001000",
  14878=>"001000101",
  14879=>"111101011",
  14880=>"000010000",
  14881=>"110110100",
  14882=>"110100011",
  14883=>"011110110",
  14884=>"110001010",
  14885=>"010100101",
  14886=>"011111110",
  14887=>"001001001",
  14888=>"100110011",
  14889=>"001011010",
  14890=>"101101001",
  14891=>"010101001",
  14892=>"110011000",
  14893=>"100110001",
  14894=>"000000010",
  14895=>"101010100",
  14896=>"100011110",
  14897=>"001010110",
  14898=>"110010101",
  14899=>"000000110",
  14900=>"101100110",
  14901=>"000010011",
  14902=>"010001110",
  14903=>"101100001",
  14904=>"010000000",
  14905=>"010010000",
  14906=>"011100010",
  14907=>"000100000",
  14908=>"100110001",
  14909=>"010111110",
  14910=>"110001101",
  14911=>"000100010",
  14912=>"000010100",
  14913=>"001100011",
  14914=>"110001011",
  14915=>"000111100",
  14916=>"100011110",
  14917=>"000010000",
  14918=>"100011000",
  14919=>"101101001",
  14920=>"111001101",
  14921=>"000111001",
  14922=>"001101011",
  14923=>"110010000",
  14924=>"010110001",
  14925=>"101011111",
  14926=>"101111111",
  14927=>"001001110",
  14928=>"110011111",
  14929=>"111101100",
  14930=>"001100101",
  14931=>"000010100",
  14932=>"100000001",
  14933=>"001101000",
  14934=>"010000000",
  14935=>"001010000",
  14936=>"101111110",
  14937=>"100011001",
  14938=>"000001010",
  14939=>"000000000",
  14940=>"001010101",
  14941=>"001000100",
  14942=>"000100111",
  14943=>"011010001",
  14944=>"001010000",
  14945=>"111101010",
  14946=>"101001010",
  14947=>"011100000",
  14948=>"110100000",
  14949=>"100000011",
  14950=>"110011111",
  14951=>"000000101",
  14952=>"001000111",
  14953=>"100100010",
  14954=>"111011001",
  14955=>"101100110",
  14956=>"000001110",
  14957=>"010001010",
  14958=>"010111100",
  14959=>"100010111",
  14960=>"110110101",
  14961=>"000010111",
  14962=>"100011000",
  14963=>"001110010",
  14964=>"111010101",
  14965=>"000000100",
  14966=>"010110011",
  14967=>"101010000",
  14968=>"011001110",
  14969=>"010111111",
  14970=>"011011111",
  14971=>"100111000",
  14972=>"001000100",
  14973=>"101001001",
  14974=>"000111010",
  14975=>"000010000",
  14976=>"010100101",
  14977=>"000010010",
  14978=>"010011000",
  14979=>"100000011",
  14980=>"000011010",
  14981=>"101110111",
  14982=>"011000100",
  14983=>"101100001",
  14984=>"110010100",
  14985=>"100001110",
  14986=>"011001000",
  14987=>"101111001",
  14988=>"110110111",
  14989=>"101110001",
  14990=>"011110100",
  14991=>"110110001",
  14992=>"110011010",
  14993=>"001010110",
  14994=>"010011100",
  14995=>"110110101",
  14996=>"000101001",
  14997=>"100110001",
  14998=>"111001100",
  14999=>"000000100",
  15000=>"011100001",
  15001=>"000001010",
  15002=>"111011110",
  15003=>"000010110",
  15004=>"100111110",
  15005=>"011010111",
  15006=>"101100011",
  15007=>"000000010",
  15008=>"101111110",
  15009=>"111101110",
  15010=>"101001110",
  15011=>"001100100",
  15012=>"010111101",
  15013=>"111101111",
  15014=>"101111001",
  15015=>"001110000",
  15016=>"101000010",
  15017=>"000100011",
  15018=>"000011101",
  15019=>"000110110",
  15020=>"000101100",
  15021=>"001010000",
  15022=>"011111100",
  15023=>"000111110",
  15024=>"110110100",
  15025=>"000010010",
  15026=>"110111111",
  15027=>"110111111",
  15028=>"011110010",
  15029=>"101110000",
  15030=>"101011111",
  15031=>"000011000",
  15032=>"000010010",
  15033=>"111100100",
  15034=>"001100101",
  15035=>"111110000",
  15036=>"001000100",
  15037=>"010000000",
  15038=>"010001010",
  15039=>"011000110",
  15040=>"010110111",
  15041=>"010100101",
  15042=>"000110111",
  15043=>"110111110",
  15044=>"000010110",
  15045=>"010011010",
  15046=>"100011101",
  15047=>"010111111",
  15048=>"100001000",
  15049=>"111111111",
  15050=>"000000001",
  15051=>"000101100",
  15052=>"101011110",
  15053=>"111100111",
  15054=>"111011111",
  15055=>"000010000",
  15056=>"100101011",
  15057=>"000000111",
  15058=>"111111001",
  15059=>"100010000",
  15060=>"100110001",
  15061=>"010011110",
  15062=>"111011010",
  15063=>"110011011",
  15064=>"001101010",
  15065=>"110110001",
  15066=>"110000111",
  15067=>"101000001",
  15068=>"001101011",
  15069=>"001100101",
  15070=>"000100010",
  15071=>"111110110",
  15072=>"111001110",
  15073=>"110011110",
  15074=>"111011000",
  15075=>"000110010",
  15076=>"011001000",
  15077=>"000100011",
  15078=>"010101010",
  15079=>"001110011",
  15080=>"001110001",
  15081=>"101011111",
  15082=>"011101110",
  15083=>"101110001",
  15084=>"000000010",
  15085=>"110110000",
  15086=>"111111100",
  15087=>"010110010",
  15088=>"111010000",
  15089=>"000000000",
  15090=>"101100011",
  15091=>"001011010",
  15092=>"011000001",
  15093=>"100111011",
  15094=>"000010001",
  15095=>"010100111",
  15096=>"111100000",
  15097=>"100110111",
  15098=>"010001011",
  15099=>"000000000",
  15100=>"111100001",
  15101=>"000000000",
  15102=>"010000101",
  15103=>"011100011",
  15104=>"001111110",
  15105=>"000110101",
  15106=>"111110010",
  15107=>"110000010",
  15108=>"110101010",
  15109=>"001000110",
  15110=>"101001010",
  15111=>"000101000",
  15112=>"101011111",
  15113=>"000101110",
  15114=>"011100001",
  15115=>"001000001",
  15116=>"000000101",
  15117=>"110100100",
  15118=>"010111101",
  15119=>"100010001",
  15120=>"001111110",
  15121=>"010000111",
  15122=>"101001111",
  15123=>"110100110",
  15124=>"110110000",
  15125=>"001100101",
  15126=>"111111111",
  15127=>"000010001",
  15128=>"110110011",
  15129=>"001111000",
  15130=>"000100010",
  15131=>"110001000",
  15132=>"110100010",
  15133=>"011110111",
  15134=>"001001110",
  15135=>"111001011",
  15136=>"101110000",
  15137=>"111110110",
  15138=>"111010101",
  15139=>"101010100",
  15140=>"000011001",
  15141=>"010100111",
  15142=>"011000110",
  15143=>"111111101",
  15144=>"100011100",
  15145=>"101100000",
  15146=>"000101000",
  15147=>"011100111",
  15148=>"010001000",
  15149=>"101000110",
  15150=>"100000011",
  15151=>"001010001",
  15152=>"001100110",
  15153=>"000111011",
  15154=>"000101111",
  15155=>"000011000",
  15156=>"001101011",
  15157=>"101100010",
  15158=>"111000111",
  15159=>"110100100",
  15160=>"001101111",
  15161=>"110010010",
  15162=>"000101111",
  15163=>"000100001",
  15164=>"111100000",
  15165=>"001011011",
  15166=>"000000000",
  15167=>"110010100",
  15168=>"011000001",
  15169=>"010011011",
  15170=>"001110111",
  15171=>"010111011",
  15172=>"011000010",
  15173=>"010110100",
  15174=>"000101110",
  15175=>"111001001",
  15176=>"100010011",
  15177=>"111101100",
  15178=>"101111111",
  15179=>"001010110",
  15180=>"100110010",
  15181=>"010011010",
  15182=>"101110111",
  15183=>"011111001",
  15184=>"010111010",
  15185=>"010111111",
  15186=>"100000000",
  15187=>"000000000",
  15188=>"100010001",
  15189=>"111001011",
  15190=>"001111100",
  15191=>"010000101",
  15192=>"110001101",
  15193=>"011000000",
  15194=>"011110111",
  15195=>"101010000",
  15196=>"111101101",
  15197=>"111111100",
  15198=>"001101000",
  15199=>"010100110",
  15200=>"010111100",
  15201=>"000110101",
  15202=>"111000100",
  15203=>"011111001",
  15204=>"101010100",
  15205=>"001000101",
  15206=>"001000010",
  15207=>"101000010",
  15208=>"001110100",
  15209=>"011111100",
  15210=>"001000001",
  15211=>"100101000",
  15212=>"010111001",
  15213=>"001101011",
  15214=>"110101111",
  15215=>"011001010",
  15216=>"001010100",
  15217=>"111111000",
  15218=>"011011001",
  15219=>"111101100",
  15220=>"101100011",
  15221=>"101000010",
  15222=>"111101001",
  15223=>"010111010",
  15224=>"101011000",
  15225=>"001001110",
  15226=>"001011010",
  15227=>"101011110",
  15228=>"010011010",
  15229=>"010110000",
  15230=>"111111101",
  15231=>"011011100",
  15232=>"111011010",
  15233=>"110011001",
  15234=>"011010000",
  15235=>"001010010",
  15236=>"100010001",
  15237=>"001100010",
  15238=>"110000110",
  15239=>"000000100",
  15240=>"100011101",
  15241=>"000000111",
  15242=>"011010000",
  15243=>"010011010",
  15244=>"011110101",
  15245=>"111110110",
  15246=>"100011100",
  15247=>"111010010",
  15248=>"000000011",
  15249=>"111010010",
  15250=>"000101011",
  15251=>"011101010",
  15252=>"011111010",
  15253=>"010011000",
  15254=>"011001111",
  15255=>"111100110",
  15256=>"011100010",
  15257=>"101110000",
  15258=>"100110110",
  15259=>"110000000",
  15260=>"101101101",
  15261=>"101001100",
  15262=>"111111110",
  15263=>"110010111",
  15264=>"000001100",
  15265=>"101010111",
  15266=>"111111010",
  15267=>"111001101",
  15268=>"000010110",
  15269=>"001010111",
  15270=>"101111001",
  15271=>"000110010",
  15272=>"111110001",
  15273=>"010111111",
  15274=>"001011000",
  15275=>"110110100",
  15276=>"010010111",
  15277=>"001000010",
  15278=>"100010000",
  15279=>"011001001",
  15280=>"000011000",
  15281=>"110100000",
  15282=>"011101000",
  15283=>"011101001",
  15284=>"100011100",
  15285=>"011001111",
  15286=>"000111001",
  15287=>"100101001",
  15288=>"011110100",
  15289=>"110011011",
  15290=>"000010100",
  15291=>"001111001",
  15292=>"001011110",
  15293=>"010010010",
  15294=>"111011110",
  15295=>"000010000",
  15296=>"010010011",
  15297=>"101110011",
  15298=>"011101111",
  15299=>"111010010",
  15300=>"001011100",
  15301=>"101010001",
  15302=>"110011111",
  15303=>"100000100",
  15304=>"000011000",
  15305=>"100010001",
  15306=>"110011101",
  15307=>"010010100",
  15308=>"111111001",
  15309=>"101001110",
  15310=>"110110000",
  15311=>"110101001",
  15312=>"001010110",
  15313=>"000100001",
  15314=>"010001100",
  15315=>"010111110",
  15316=>"010111000",
  15317=>"000001010",
  15318=>"000001000",
  15319=>"010111000",
  15320=>"011011110",
  15321=>"101101000",
  15322=>"110100111",
  15323=>"101000001",
  15324=>"000001001",
  15325=>"000010010",
  15326=>"110110010",
  15327=>"011100010",
  15328=>"011011111",
  15329=>"100111110",
  15330=>"011011011",
  15331=>"000111011",
  15332=>"111011110",
  15333=>"010110000",
  15334=>"000111000",
  15335=>"000100010",
  15336=>"110100111",
  15337=>"000000001",
  15338=>"101000001",
  15339=>"001100010",
  15340=>"010010001",
  15341=>"010011010",
  15342=>"010000101",
  15343=>"101001000",
  15344=>"000010011",
  15345=>"110100100",
  15346=>"000101000",
  15347=>"111010100",
  15348=>"000010110",
  15349=>"101001110",
  15350=>"110010110",
  15351=>"111001101",
  15352=>"010111111",
  15353=>"000000000",
  15354=>"001101111",
  15355=>"000111100",
  15356=>"000101010",
  15357=>"110101100",
  15358=>"110100100",
  15359=>"100010000",
  15360=>"011011111",
  15361=>"001111100",
  15362=>"011101111",
  15363=>"010110011",
  15364=>"100111100",
  15365=>"000110001",
  15366=>"111011110",
  15367=>"000111100",
  15368=>"010101110",
  15369=>"010010001",
  15370=>"111011010",
  15371=>"111101010",
  15372=>"101001000",
  15373=>"000000110",
  15374=>"011000000",
  15375=>"100101100",
  15376=>"000011011",
  15377=>"110101110",
  15378=>"100100101",
  15379=>"001100101",
  15380=>"111011100",
  15381=>"000000000",
  15382=>"111000110",
  15383=>"011001110",
  15384=>"100101000",
  15385=>"010010010",
  15386=>"010010010",
  15387=>"110100000",
  15388=>"011011100",
  15389=>"000101101",
  15390=>"001101101",
  15391=>"101000010",
  15392=>"110010001",
  15393=>"001100110",
  15394=>"001001010",
  15395=>"011110011",
  15396=>"100100100",
  15397=>"111000101",
  15398=>"100111011",
  15399=>"111101101",
  15400=>"100101100",
  15401=>"001111111",
  15402=>"110111000",
  15403=>"101111111",
  15404=>"110101001",
  15405=>"100010001",
  15406=>"100100111",
  15407=>"001000111",
  15408=>"001111001",
  15409=>"010001001",
  15410=>"111100010",
  15411=>"000100100",
  15412=>"100010111",
  15413=>"000000001",
  15414=>"000100101",
  15415=>"000010100",
  15416=>"011000111",
  15417=>"111100111",
  15418=>"111111111",
  15419=>"001010001",
  15420=>"010101101",
  15421=>"110010000",
  15422=>"001101001",
  15423=>"111010010",
  15424=>"000011100",
  15425=>"001001100",
  15426=>"111100010",
  15427=>"101111011",
  15428=>"110111011",
  15429=>"011111001",
  15430=>"011010111",
  15431=>"111110100",
  15432=>"010100111",
  15433=>"010011001",
  15434=>"000000111",
  15435=>"010110010",
  15436=>"011000000",
  15437=>"001111010",
  15438=>"011001100",
  15439=>"100100000",
  15440=>"110011110",
  15441=>"111101101",
  15442=>"101011000",
  15443=>"101110000",
  15444=>"101010110",
  15445=>"011001010",
  15446=>"100000011",
  15447=>"110100000",
  15448=>"110000101",
  15449=>"000100010",
  15450=>"011001000",
  15451=>"011100100",
  15452=>"110101001",
  15453=>"000000001",
  15454=>"011100010",
  15455=>"110100001",
  15456=>"000011111",
  15457=>"110101000",
  15458=>"001100001",
  15459=>"011010110",
  15460=>"111011100",
  15461=>"100110000",
  15462=>"011100110",
  15463=>"110111100",
  15464=>"011110110",
  15465=>"101101001",
  15466=>"101110100",
  15467=>"000110001",
  15468=>"000100011",
  15469=>"111110001",
  15470=>"100100100",
  15471=>"010101011",
  15472=>"110110000",
  15473=>"110000010",
  15474=>"110111001",
  15475=>"110100010",
  15476=>"001000100",
  15477=>"011000111",
  15478=>"100011111",
  15479=>"001010110",
  15480=>"010000010",
  15481=>"100010000",
  15482=>"110100101",
  15483=>"100000010",
  15484=>"101010010",
  15485=>"101000000",
  15486=>"011111111",
  15487=>"000000001",
  15488=>"111101101",
  15489=>"001100010",
  15490=>"011010000",
  15491=>"000011100",
  15492=>"000000111",
  15493=>"101101010",
  15494=>"001111010",
  15495=>"011011010",
  15496=>"110100000",
  15497=>"010100001",
  15498=>"001000000",
  15499=>"010110110",
  15500=>"101001100",
  15501=>"000010001",
  15502=>"100110001",
  15503=>"011011000",
  15504=>"100101000",
  15505=>"111011010",
  15506=>"010000110",
  15507=>"010111011",
  15508=>"110000000",
  15509=>"011100001",
  15510=>"100110110",
  15511=>"111111000",
  15512=>"111100001",
  15513=>"110101101",
  15514=>"000011011",
  15515=>"101101010",
  15516=>"100010101",
  15517=>"001101100",
  15518=>"100000001",
  15519=>"011111011",
  15520=>"010101110",
  15521=>"111000011",
  15522=>"001111100",
  15523=>"000001111",
  15524=>"101110001",
  15525=>"111110111",
  15526=>"101011010",
  15527=>"101110111",
  15528=>"010001110",
  15529=>"101100000",
  15530=>"101101111",
  15531=>"110010011",
  15532=>"011111100",
  15533=>"111011100",
  15534=>"100010101",
  15535=>"111100011",
  15536=>"001000110",
  15537=>"001110001",
  15538=>"101001111",
  15539=>"000101111",
  15540=>"000000000",
  15541=>"101011001",
  15542=>"000100001",
  15543=>"001101000",
  15544=>"111110000",
  15545=>"101001000",
  15546=>"110110011",
  15547=>"010101101",
  15548=>"111010111",
  15549=>"110110101",
  15550=>"011101010",
  15551=>"111111010",
  15552=>"010001011",
  15553=>"000011111",
  15554=>"101110001",
  15555=>"000010100",
  15556=>"101110001",
  15557=>"000010111",
  15558=>"011010010",
  15559=>"110101001",
  15560=>"000000000",
  15561=>"000010010",
  15562=>"001010100",
  15563=>"111001000",
  15564=>"110001000",
  15565=>"100111100",
  15566=>"101010100",
  15567=>"110000100",
  15568=>"000000110",
  15569=>"011101011",
  15570=>"110011000",
  15571=>"011110000",
  15572=>"010001010",
  15573=>"001101010",
  15574=>"110001110",
  15575=>"100010000",
  15576=>"000000001",
  15577=>"100100000",
  15578=>"100010101",
  15579=>"111110100",
  15580=>"000001101",
  15581=>"100000000",
  15582=>"011000000",
  15583=>"110011111",
  15584=>"001001101",
  15585=>"110000111",
  15586=>"100101101",
  15587=>"010000101",
  15588=>"100101100",
  15589=>"000111001",
  15590=>"100011111",
  15591=>"110101100",
  15592=>"101101101",
  15593=>"100000110",
  15594=>"110011000",
  15595=>"001011000",
  15596=>"010101111",
  15597=>"001000110",
  15598=>"100100010",
  15599=>"011010000",
  15600=>"011011100",
  15601=>"110100101",
  15602=>"000010010",
  15603=>"011110100",
  15604=>"110001010",
  15605=>"000010100",
  15606=>"000011010",
  15607=>"100100001",
  15608=>"111100010",
  15609=>"000111100",
  15610=>"001100000",
  15611=>"000001000",
  15612=>"101110101",
  15613=>"010101101",
  15614=>"001101111",
  15615=>"111100111",
  15616=>"111101100",
  15617=>"010101111",
  15618=>"100000010",
  15619=>"100000000",
  15620=>"110000000",
  15621=>"011100011",
  15622=>"010101100",
  15623=>"110000110",
  15624=>"100100111",
  15625=>"100001110",
  15626=>"100011000",
  15627=>"011101101",
  15628=>"011111010",
  15629=>"101100000",
  15630=>"010011110",
  15631=>"010011000",
  15632=>"101000101",
  15633=>"011010010",
  15634=>"011000000",
  15635=>"100001110",
  15636=>"011110010",
  15637=>"010011011",
  15638=>"100101000",
  15639=>"010110011",
  15640=>"110011001",
  15641=>"101111001",
  15642=>"110111111",
  15643=>"110011010",
  15644=>"010110010",
  15645=>"001010010",
  15646=>"000001101",
  15647=>"001000101",
  15648=>"010000000",
  15649=>"010000000",
  15650=>"011100111",
  15651=>"001001110",
  15652=>"001011011",
  15653=>"100000000",
  15654=>"011110101",
  15655=>"101101000",
  15656=>"110110001",
  15657=>"100011101",
  15658=>"010101011",
  15659=>"101100111",
  15660=>"000111111",
  15661=>"110110000",
  15662=>"100101111",
  15663=>"010100100",
  15664=>"011011010",
  15665=>"101000101",
  15666=>"100100110",
  15667=>"000111110",
  15668=>"000010011",
  15669=>"000001111",
  15670=>"010001011",
  15671=>"000101001",
  15672=>"001101000",
  15673=>"010101110",
  15674=>"111000101",
  15675=>"001000100",
  15676=>"101011001",
  15677=>"110000100",
  15678=>"011001110",
  15679=>"001000001",
  15680=>"100000100",
  15681=>"101010111",
  15682=>"111111000",
  15683=>"101101110",
  15684=>"111010111",
  15685=>"010001011",
  15686=>"001100011",
  15687=>"000000011",
  15688=>"001110011",
  15689=>"100001011",
  15690=>"111010101",
  15691=>"100011010",
  15692=>"010110001",
  15693=>"000000101",
  15694=>"111000100",
  15695=>"101111000",
  15696=>"010110110",
  15697=>"100000010",
  15698=>"111001100",
  15699=>"101110001",
  15700=>"000001100",
  15701=>"110111011",
  15702=>"000111110",
  15703=>"100100010",
  15704=>"000000010",
  15705=>"011001010",
  15706=>"110110001",
  15707=>"100110101",
  15708=>"100010010",
  15709=>"011011000",
  15710=>"111010111",
  15711=>"011110000",
  15712=>"101111110",
  15713=>"100011101",
  15714=>"100010111",
  15715=>"110100110",
  15716=>"010101000",
  15717=>"010110101",
  15718=>"110110111",
  15719=>"000010110",
  15720=>"110110011",
  15721=>"001001110",
  15722=>"110110000",
  15723=>"000110110",
  15724=>"101011010",
  15725=>"001100110",
  15726=>"001111101",
  15727=>"111111100",
  15728=>"110111011",
  15729=>"111111011",
  15730=>"001000000",
  15731=>"010111001",
  15732=>"110001001",
  15733=>"000011010",
  15734=>"110110101",
  15735=>"101000111",
  15736=>"111110000",
  15737=>"100110010",
  15738=>"010101111",
  15739=>"100000011",
  15740=>"010100101",
  15741=>"001000001",
  15742=>"000000010",
  15743=>"001011110",
  15744=>"100100101",
  15745=>"010100100",
  15746=>"011000011",
  15747=>"100110000",
  15748=>"000010010",
  15749=>"100110100",
  15750=>"101001001",
  15751=>"111011001",
  15752=>"000110110",
  15753=>"001111001",
  15754=>"011101001",
  15755=>"101000110",
  15756=>"011010001",
  15757=>"100010111",
  15758=>"111110100",
  15759=>"111110100",
  15760=>"100100111",
  15761=>"000100101",
  15762=>"111011101",
  15763=>"111010100",
  15764=>"100001100",
  15765=>"110101100",
  15766=>"000011000",
  15767=>"011101111",
  15768=>"111101111",
  15769=>"100010010",
  15770=>"100011100",
  15771=>"110011010",
  15772=>"111110111",
  15773=>"111111100",
  15774=>"111001011",
  15775=>"010011110",
  15776=>"001001111",
  15777=>"110111011",
  15778=>"001100100",
  15779=>"001100100",
  15780=>"100001111",
  15781=>"010011000",
  15782=>"111001100",
  15783=>"001010011",
  15784=>"000110111",
  15785=>"100110000",
  15786=>"010110000",
  15787=>"000010011",
  15788=>"000000110",
  15789=>"100010000",
  15790=>"111001011",
  15791=>"110101111",
  15792=>"001100101",
  15793=>"010011110",
  15794=>"101010101",
  15795=>"101110001",
  15796=>"101011111",
  15797=>"010011111",
  15798=>"011000111",
  15799=>"100000011",
  15800=>"011000101",
  15801=>"011011101",
  15802=>"011011000",
  15803=>"100101010",
  15804=>"110100000",
  15805=>"100111110",
  15806=>"000111100",
  15807=>"111011000",
  15808=>"011110111",
  15809=>"101011010",
  15810=>"010010011",
  15811=>"000011111",
  15812=>"100010110",
  15813=>"111011011",
  15814=>"010111100",
  15815=>"111101111",
  15816=>"111100100",
  15817=>"011101010",
  15818=>"000010000",
  15819=>"110101011",
  15820=>"000111011",
  15821=>"101101001",
  15822=>"001100001",
  15823=>"100111011",
  15824=>"100110011",
  15825=>"011101000",
  15826=>"100110111",
  15827=>"111111111",
  15828=>"011011011",
  15829=>"100100010",
  15830=>"011000010",
  15831=>"000110000",
  15832=>"011001001",
  15833=>"111110101",
  15834=>"011011101",
  15835=>"101010111",
  15836=>"110101001",
  15837=>"011110111",
  15838=>"011010111",
  15839=>"011100001",
  15840=>"010101101",
  15841=>"110110101",
  15842=>"011110010",
  15843=>"101101111",
  15844=>"101000100",
  15845=>"110110010",
  15846=>"000100110",
  15847=>"010000111",
  15848=>"000100011",
  15849=>"101111111",
  15850=>"101101011",
  15851=>"110111111",
  15852=>"111100011",
  15853=>"001010011",
  15854=>"110011001",
  15855=>"111110101",
  15856=>"110110000",
  15857=>"100011100",
  15858=>"101001100",
  15859=>"001101100",
  15860=>"000111100",
  15861=>"111010101",
  15862=>"000110101",
  15863=>"100001110",
  15864=>"000100000",
  15865=>"010000011",
  15866=>"001111000",
  15867=>"110001111",
  15868=>"001011110",
  15869=>"010000010",
  15870=>"100010111",
  15871=>"011111111",
  15872=>"000100000",
  15873=>"110100010",
  15874=>"010001111",
  15875=>"111001110",
  15876=>"001110101",
  15877=>"000010010",
  15878=>"100000000",
  15879=>"001101011",
  15880=>"111011010",
  15881=>"100101001",
  15882=>"010001010",
  15883=>"001111000",
  15884=>"100000001",
  15885=>"100110010",
  15886=>"100101110",
  15887=>"111100110",
  15888=>"011111100",
  15889=>"010000100",
  15890=>"000111000",
  15891=>"000111010",
  15892=>"010110001",
  15893=>"010010010",
  15894=>"001001101",
  15895=>"110000011",
  15896=>"111100101",
  15897=>"110110001",
  15898=>"010010110",
  15899=>"111011000",
  15900=>"101010100",
  15901=>"011000110",
  15902=>"001011100",
  15903=>"100101111",
  15904=>"010110001",
  15905=>"101111001",
  15906=>"111000101",
  15907=>"111000010",
  15908=>"001111101",
  15909=>"101001010",
  15910=>"000010101",
  15911=>"001111010",
  15912=>"001101100",
  15913=>"111100010",
  15914=>"110000010",
  15915=>"001110100",
  15916=>"101100001",
  15917=>"000000110",
  15918=>"010000001",
  15919=>"010000000",
  15920=>"100011000",
  15921=>"010011000",
  15922=>"100001111",
  15923=>"100010101",
  15924=>"100101111",
  15925=>"110110011",
  15926=>"101101011",
  15927=>"101101111",
  15928=>"111011100",
  15929=>"011101100",
  15930=>"101001111",
  15931=>"101001010",
  15932=>"001100011",
  15933=>"000001101",
  15934=>"101100100",
  15935=>"111110111",
  15936=>"010111001",
  15937=>"111010110",
  15938=>"101111010",
  15939=>"101101100",
  15940=>"100010000",
  15941=>"001100111",
  15942=>"000000011",
  15943=>"111101001",
  15944=>"100110101",
  15945=>"110010100",
  15946=>"100010110",
  15947=>"100001110",
  15948=>"011001111",
  15949=>"101010110",
  15950=>"110100011",
  15951=>"010001001",
  15952=>"000011000",
  15953=>"000011100",
  15954=>"010001110",
  15955=>"101001001",
  15956=>"100010111",
  15957=>"000000010",
  15958=>"010000011",
  15959=>"111111111",
  15960=>"110111001",
  15961=>"111000111",
  15962=>"110110101",
  15963=>"011010110",
  15964=>"011000111",
  15965=>"000101011",
  15966=>"001011010",
  15967=>"101011110",
  15968=>"000110111",
  15969=>"110001110",
  15970=>"111111110",
  15971=>"101100001",
  15972=>"001010101",
  15973=>"000111010",
  15974=>"001010010",
  15975=>"011001101",
  15976=>"001011100",
  15977=>"011010001",
  15978=>"001110001",
  15979=>"000000011",
  15980=>"000011001",
  15981=>"100111011",
  15982=>"101001010",
  15983=>"001000011",
  15984=>"001010010",
  15985=>"001110010",
  15986=>"110000100",
  15987=>"100110110",
  15988=>"010011010",
  15989=>"011111111",
  15990=>"111010000",
  15991=>"000110010",
  15992=>"110000110",
  15993=>"100001101",
  15994=>"000110111",
  15995=>"110110000",
  15996=>"100010011",
  15997=>"011110100",
  15998=>"001100011",
  15999=>"111011011",
  16000=>"110001001",
  16001=>"111110010",
  16002=>"010101010",
  16003=>"001101101",
  16004=>"110101001",
  16005=>"100101100",
  16006=>"010010010",
  16007=>"111001101",
  16008=>"111000101",
  16009=>"011100111",
  16010=>"000101010",
  16011=>"011011001",
  16012=>"010000011",
  16013=>"110001011",
  16014=>"000100001",
  16015=>"101110100",
  16016=>"101010100",
  16017=>"010011111",
  16018=>"110011011",
  16019=>"011001011",
  16020=>"111000100",
  16021=>"111101111",
  16022=>"010101000",
  16023=>"000010001",
  16024=>"111111100",
  16025=>"001011110",
  16026=>"011101001",
  16027=>"110000101",
  16028=>"101111111",
  16029=>"011101111",
  16030=>"000000001",
  16031=>"101110010",
  16032=>"101011101",
  16033=>"001010110",
  16034=>"010100110",
  16035=>"111011011",
  16036=>"100010001",
  16037=>"001000100",
  16038=>"000000101",
  16039=>"100001000",
  16040=>"111111000",
  16041=>"000010101",
  16042=>"101110101",
  16043=>"110001111",
  16044=>"001101000",
  16045=>"101101111",
  16046=>"011100101",
  16047=>"101011110",
  16048=>"110011101",
  16049=>"011110101",
  16050=>"000010110",
  16051=>"111110010",
  16052=>"001010110",
  16053=>"011110011",
  16054=>"111111000",
  16055=>"111010111",
  16056=>"010011011",
  16057=>"011000001",
  16058=>"011010010",
  16059=>"000001010",
  16060=>"000010101",
  16061=>"001000010",
  16062=>"100001000",
  16063=>"010100101",
  16064=>"001100001",
  16065=>"111011011",
  16066=>"010010011",
  16067=>"001001000",
  16068=>"100000111",
  16069=>"001001110",
  16070=>"110001010",
  16071=>"000011100",
  16072=>"000010101",
  16073=>"010010001",
  16074=>"011011101",
  16075=>"111100101",
  16076=>"011111001",
  16077=>"111010000",
  16078=>"010100100",
  16079=>"101101100",
  16080=>"110101111",
  16081=>"000000101",
  16082=>"001101011",
  16083=>"100010011",
  16084=>"000000000",
  16085=>"011110110",
  16086=>"011100111",
  16087=>"010001001",
  16088=>"101111111",
  16089=>"101100011",
  16090=>"110000100",
  16091=>"010011101",
  16092=>"000100110",
  16093=>"001110001",
  16094=>"011111010",
  16095=>"000110011",
  16096=>"001101001",
  16097=>"100011000",
  16098=>"001100001",
  16099=>"100011111",
  16100=>"001010001",
  16101=>"001100111",
  16102=>"110101001",
  16103=>"111011011",
  16104=>"001100101",
  16105=>"111010001",
  16106=>"010100000",
  16107=>"000010101",
  16108=>"001001000",
  16109=>"011111111",
  16110=>"111000101",
  16111=>"100100000",
  16112=>"001100111",
  16113=>"011110110",
  16114=>"011011000",
  16115=>"111101011",
  16116=>"111111010",
  16117=>"010111010",
  16118=>"000110100",
  16119=>"010001001",
  16120=>"101000000",
  16121=>"010000110",
  16122=>"100000011",
  16123=>"011111111",
  16124=>"101000011",
  16125=>"111010110",
  16126=>"101010110",
  16127=>"111011101",
  16128=>"000001111",
  16129=>"001011011",
  16130=>"111011111",
  16131=>"011100001",
  16132=>"000100011",
  16133=>"001101110",
  16134=>"000010101",
  16135=>"010111110",
  16136=>"001000001",
  16137=>"110001100",
  16138=>"001001111",
  16139=>"110110101",
  16140=>"001111001",
  16141=>"000000010",
  16142=>"100000110",
  16143=>"100100101",
  16144=>"010010001",
  16145=>"110001111",
  16146=>"001000010",
  16147=>"000011111",
  16148=>"101000111",
  16149=>"000010110",
  16150=>"111000011",
  16151=>"001010001",
  16152=>"010101011",
  16153=>"010100000",
  16154=>"110100100",
  16155=>"000110010",
  16156=>"010111111",
  16157=>"001110110",
  16158=>"100001000",
  16159=>"001100100",
  16160=>"101101011",
  16161=>"110011001",
  16162=>"010000111",
  16163=>"010000100",
  16164=>"010101001",
  16165=>"111101101",
  16166=>"000000011",
  16167=>"101111011",
  16168=>"010000000",
  16169=>"101001100",
  16170=>"111000111",
  16171=>"000000111",
  16172=>"010010001",
  16173=>"001011000",
  16174=>"101011110",
  16175=>"011011001",
  16176=>"001101111",
  16177=>"010000101",
  16178=>"001000001",
  16179=>"001100010",
  16180=>"010010011",
  16181=>"101110000",
  16182=>"111010010",
  16183=>"000000011",
  16184=>"100011010",
  16185=>"101110110",
  16186=>"001101010",
  16187=>"110000110",
  16188=>"011001000",
  16189=>"000001001",
  16190=>"101010001",
  16191=>"110100110",
  16192=>"101011100",
  16193=>"100101000",
  16194=>"000000001",
  16195=>"001111000",
  16196=>"101111101",
  16197=>"111101001",
  16198=>"101111111",
  16199=>"111000111",
  16200=>"110011011",
  16201=>"001010010",
  16202=>"010101101",
  16203=>"100111111",
  16204=>"101011001",
  16205=>"100001000",
  16206=>"001101001",
  16207=>"001011100",
  16208=>"010001100",
  16209=>"111111110",
  16210=>"100100010",
  16211=>"100011010",
  16212=>"101110010",
  16213=>"000000101",
  16214=>"000001000",
  16215=>"000000100",
  16216=>"100000010",
  16217=>"000001010",
  16218=>"101000010",
  16219=>"100011011",
  16220=>"011101100",
  16221=>"111110010",
  16222=>"010111010",
  16223=>"101001000",
  16224=>"001111100",
  16225=>"001111000",
  16226=>"100000111",
  16227=>"101101110",
  16228=>"001111011",
  16229=>"011010010",
  16230=>"111101001",
  16231=>"111000111",
  16232=>"101000110",
  16233=>"111000111",
  16234=>"011110111",
  16235=>"100000100",
  16236=>"011001001",
  16237=>"111011010",
  16238=>"110101010",
  16239=>"111000110",
  16240=>"011001110",
  16241=>"010111001",
  16242=>"001010100",
  16243=>"101011110",
  16244=>"011101100",
  16245=>"011100110",
  16246=>"100000001",
  16247=>"101111111",
  16248=>"100001100",
  16249=>"011010100",
  16250=>"111000101",
  16251=>"000011010",
  16252=>"001011111",
  16253=>"001000001",
  16254=>"010111101",
  16255=>"110111110",
  16256=>"011101101",
  16257=>"010101000",
  16258=>"111000000",
  16259=>"010101010",
  16260=>"000010010",
  16261=>"011100110",
  16262=>"100110100",
  16263=>"100111011",
  16264=>"000101100",
  16265=>"011100010",
  16266=>"010111100",
  16267=>"111010101",
  16268=>"100001101",
  16269=>"001011010",
  16270=>"011100001",
  16271=>"001100011",
  16272=>"101101101",
  16273=>"000101010",
  16274=>"000001000",
  16275=>"000101000",
  16276=>"011001100",
  16277=>"000100010",
  16278=>"111001010",
  16279=>"100010111",
  16280=>"101010110",
  16281=>"111101111",
  16282=>"101000000",
  16283=>"100101011",
  16284=>"000101010",
  16285=>"000100100",
  16286=>"111110100",
  16287=>"110000111",
  16288=>"000101100",
  16289=>"000010001",
  16290=>"100111001",
  16291=>"011100011",
  16292=>"010010100",
  16293=>"111101101",
  16294=>"100011010",
  16295=>"100011011",
  16296=>"010011100",
  16297=>"101111110",
  16298=>"111111100",
  16299=>"100110011",
  16300=>"010110100",
  16301=>"110110100",
  16302=>"100100110",
  16303=>"000101111",
  16304=>"011101000",
  16305=>"010001001",
  16306=>"100000011",
  16307=>"111111000",
  16308=>"101110101",
  16309=>"011110110",
  16310=>"010111110",
  16311=>"010010111",
  16312=>"000000011",
  16313=>"011001011",
  16314=>"000111011",
  16315=>"010010100",
  16316=>"110110010",
  16317=>"100010101",
  16318=>"011000000",
  16319=>"010101110",
  16320=>"010010000",
  16321=>"101111011",
  16322=>"100011100",
  16323=>"001001000",
  16324=>"111000001",
  16325=>"011111010",
  16326=>"000010001",
  16327=>"110001010",
  16328=>"011010011",
  16329=>"001000111",
  16330=>"001100001",
  16331=>"101010110",
  16332=>"011111111",
  16333=>"100011001",
  16334=>"000001001",
  16335=>"100000000",
  16336=>"010100001",
  16337=>"110101011",
  16338=>"110001100",
  16339=>"011000011",
  16340=>"100101100",
  16341=>"001001000",
  16342=>"000000010",
  16343=>"110010000",
  16344=>"001001001",
  16345=>"110100110",
  16346=>"111011010",
  16347=>"100001001",
  16348=>"101111101",
  16349=>"010111011",
  16350=>"000100011",
  16351=>"100011000",
  16352=>"001101010",
  16353=>"100011100",
  16354=>"000100010",
  16355=>"101001000",
  16356=>"100000111",
  16357=>"000001001",
  16358=>"111101010",
  16359=>"010111111",
  16360=>"010000011",
  16361=>"000101110",
  16362=>"101111100",
  16363=>"000011011",
  16364=>"100000100",
  16365=>"010001010",
  16366=>"111000011",
  16367=>"110110001",
  16368=>"001011000",
  16369=>"001000001",
  16370=>"110010100",
  16371=>"000001000",
  16372=>"010011100",
  16373=>"101111110",
  16374=>"011000110",
  16375=>"010110111",
  16376=>"111101110",
  16377=>"000000011",
  16378=>"000010111",
  16379=>"111101111",
  16380=>"010011100",
  16381=>"101010100",
  16382=>"111111011",
  16383=>"100101011",
  16384=>"110001010",
  16385=>"100110100",
  16386=>"000000001",
  16387=>"000000000",
  16388=>"000010110",
  16389=>"001010110",
  16390=>"110101101",
  16391=>"110011111",
  16392=>"000011000",
  16393=>"011001101",
  16394=>"110111100",
  16395=>"110010101",
  16396=>"011111001",
  16397=>"011010000",
  16398=>"001110001",
  16399=>"101111101",
  16400=>"111001100",
  16401=>"001101001",
  16402=>"110010001",
  16403=>"111100100",
  16404=>"001001110",
  16405=>"100111101",
  16406=>"101100001",
  16407=>"010100001",
  16408=>"000000110",
  16409=>"111000111",
  16410=>"011001000",
  16411=>"001110100",
  16412=>"110101111",
  16413=>"111111000",
  16414=>"110111110",
  16415=>"010100101",
  16416=>"010001101",
  16417=>"001101111",
  16418=>"100011100",
  16419=>"001010010",
  16420=>"010110101",
  16421=>"100011001",
  16422=>"011110001",
  16423=>"001001110",
  16424=>"100010101",
  16425=>"011011001",
  16426=>"111110111",
  16427=>"011111001",
  16428=>"111111111",
  16429=>"111101111",
  16430=>"101001010",
  16431=>"001011000",
  16432=>"111100110",
  16433=>"001101010",
  16434=>"010101100",
  16435=>"000111010",
  16436=>"111110100",
  16437=>"010101110",
  16438=>"110110001",
  16439=>"111111101",
  16440=>"001111101",
  16441=>"001110110",
  16442=>"111100001",
  16443=>"100000011",
  16444=>"000111111",
  16445=>"100111110",
  16446=>"011011000",
  16447=>"011011111",
  16448=>"000100000",
  16449=>"111011010",
  16450=>"101110100",
  16451=>"100011110",
  16452=>"110110000",
  16453=>"110100100",
  16454=>"011100111",
  16455=>"111101110",
  16456=>"010000000",
  16457=>"010100110",
  16458=>"100000010",
  16459=>"011010110",
  16460=>"001110010",
  16461=>"001101011",
  16462=>"111000111",
  16463=>"111111011",
  16464=>"110110111",
  16465=>"010000111",
  16466=>"010001111",
  16467=>"101010110",
  16468=>"000101000",
  16469=>"100100000",
  16470=>"110110100",
  16471=>"011011010",
  16472=>"001101011",
  16473=>"011111100",
  16474=>"110110001",
  16475=>"111011111",
  16476=>"010100001",
  16477=>"011101110",
  16478=>"101110010",
  16479=>"000011001",
  16480=>"101000010",
  16481=>"110110010",
  16482=>"111100101",
  16483=>"111101001",
  16484=>"011000100",
  16485=>"100110111",
  16486=>"011010110",
  16487=>"011001110",
  16488=>"000010010",
  16489=>"000110011",
  16490=>"100000000",
  16491=>"100101110",
  16492=>"000100000",
  16493=>"011100011",
  16494=>"010001110",
  16495=>"000000101",
  16496=>"011010001",
  16497=>"000111011",
  16498=>"110111001",
  16499=>"000001110",
  16500=>"000111010",
  16501=>"100111111",
  16502=>"110010101",
  16503=>"000110111",
  16504=>"010101111",
  16505=>"111010011",
  16506=>"110010110",
  16507=>"001011110",
  16508=>"010000011",
  16509=>"101010011",
  16510=>"100010010",
  16511=>"101000011",
  16512=>"010010011",
  16513=>"101100011",
  16514=>"001001000",
  16515=>"010000001",
  16516=>"101010000",
  16517=>"111100011",
  16518=>"110100100",
  16519=>"011111101",
  16520=>"110110111",
  16521=>"011101001",
  16522=>"100000101",
  16523=>"110100001",
  16524=>"010100101",
  16525=>"001011110",
  16526=>"110111101",
  16527=>"010111010",
  16528=>"000011110",
  16529=>"000101100",
  16530=>"101000100",
  16531=>"001011110",
  16532=>"111001001",
  16533=>"100010000",
  16534=>"100111111",
  16535=>"100010001",
  16536=>"001011001",
  16537=>"110000000",
  16538=>"000101010",
  16539=>"111001001",
  16540=>"101110001",
  16541=>"001000101",
  16542=>"100111011",
  16543=>"111010000",
  16544=>"000101110",
  16545=>"010011011",
  16546=>"010011101",
  16547=>"111010101",
  16548=>"000111011",
  16549=>"000111111",
  16550=>"101010101",
  16551=>"110001010",
  16552=>"100000001",
  16553=>"010100100",
  16554=>"100110000",
  16555=>"101011100",
  16556=>"010111011",
  16557=>"000010010",
  16558=>"000001101",
  16559=>"011000101",
  16560=>"001001001",
  16561=>"000110000",
  16562=>"101000110",
  16563=>"001001100",
  16564=>"101110110",
  16565=>"011001010",
  16566=>"010101100",
  16567=>"111111101",
  16568=>"111111000",
  16569=>"110011111",
  16570=>"010000000",
  16571=>"111000011",
  16572=>"100101101",
  16573=>"101100111",
  16574=>"110001010",
  16575=>"110110100",
  16576=>"111110000",
  16577=>"110111100",
  16578=>"001101100",
  16579=>"010100011",
  16580=>"001111101",
  16581=>"101100101",
  16582=>"001000111",
  16583=>"111000011",
  16584=>"111001000",
  16585=>"111001001",
  16586=>"110001010",
  16587=>"111101110",
  16588=>"010100010",
  16589=>"100010001",
  16590=>"011001001",
  16591=>"111101011",
  16592=>"101011101",
  16593=>"000001101",
  16594=>"001001001",
  16595=>"101110001",
  16596=>"010000001",
  16597=>"100110110",
  16598=>"001010001",
  16599=>"011001001",
  16600=>"100100000",
  16601=>"010100001",
  16602=>"000010010",
  16603=>"101101011",
  16604=>"101110100",
  16605=>"011000011",
  16606=>"111011111",
  16607=>"010101010",
  16608=>"010110111",
  16609=>"101000000",
  16610=>"111101001",
  16611=>"000001110",
  16612=>"010100010",
  16613=>"100100111",
  16614=>"001110000",
  16615=>"110001000",
  16616=>"011100001",
  16617=>"111011101",
  16618=>"011011111",
  16619=>"010101001",
  16620=>"110001001",
  16621=>"100110110",
  16622=>"001011001",
  16623=>"110111100",
  16624=>"100101110",
  16625=>"000000010",
  16626=>"111110111",
  16627=>"000001011",
  16628=>"011010101",
  16629=>"011110110",
  16630=>"100111000",
  16631=>"111111000",
  16632=>"011101001",
  16633=>"010001001",
  16634=>"000011001",
  16635=>"101001100",
  16636=>"000110000",
  16637=>"001111011",
  16638=>"111111110",
  16639=>"100111000",
  16640=>"100001100",
  16641=>"001001100",
  16642=>"111001100",
  16643=>"011111100",
  16644=>"111010010",
  16645=>"111110000",
  16646=>"110111101",
  16647=>"000111011",
  16648=>"011111010",
  16649=>"000101001",
  16650=>"010011011",
  16651=>"010100000",
  16652=>"111100101",
  16653=>"110011100",
  16654=>"000111010",
  16655=>"110101000",
  16656=>"100111000",
  16657=>"101100111",
  16658=>"110111000",
  16659=>"000000000",
  16660=>"001101010",
  16661=>"110000001",
  16662=>"011010011",
  16663=>"110011110",
  16664=>"101111110",
  16665=>"100001010",
  16666=>"110001001",
  16667=>"000000000",
  16668=>"111101010",
  16669=>"111000101",
  16670=>"110010111",
  16671=>"010011000",
  16672=>"010001111",
  16673=>"010000011",
  16674=>"000100011",
  16675=>"000001100",
  16676=>"001011011",
  16677=>"000000001",
  16678=>"101001110",
  16679=>"001010011",
  16680=>"100111001",
  16681=>"101010001",
  16682=>"010100011",
  16683=>"011110000",
  16684=>"111111101",
  16685=>"001111101",
  16686=>"011111110",
  16687=>"111111010",
  16688=>"010101110",
  16689=>"110111000",
  16690=>"101101110",
  16691=>"001100011",
  16692=>"111000111",
  16693=>"010111001",
  16694=>"111001101",
  16695=>"001001111",
  16696=>"001010111",
  16697=>"010010011",
  16698=>"111101100",
  16699=>"000110001",
  16700=>"110100010",
  16701=>"111110000",
  16702=>"111110001",
  16703=>"111001100",
  16704=>"001101100",
  16705=>"111101010",
  16706=>"011111101",
  16707=>"000110001",
  16708=>"000101010",
  16709=>"110111011",
  16710=>"100010100",
  16711=>"010111001",
  16712=>"000000010",
  16713=>"001111110",
  16714=>"010010110",
  16715=>"010111001",
  16716=>"111111111",
  16717=>"000111111",
  16718=>"000011111",
  16719=>"000010111",
  16720=>"100010001",
  16721=>"001000101",
  16722=>"111001110",
  16723=>"000100000",
  16724=>"110000010",
  16725=>"001011111",
  16726=>"011110110",
  16727=>"010011110",
  16728=>"001101001",
  16729=>"000000100",
  16730=>"110010001",
  16731=>"001001111",
  16732=>"100000101",
  16733=>"101110000",
  16734=>"011001100",
  16735=>"000001111",
  16736=>"000100110",
  16737=>"011110110",
  16738=>"001100100",
  16739=>"000001101",
  16740=>"111101111",
  16741=>"100100101",
  16742=>"000101100",
  16743=>"110000100",
  16744=>"001001010",
  16745=>"101111110",
  16746=>"000000111",
  16747=>"101111111",
  16748=>"101010010",
  16749=>"101011001",
  16750=>"111001000",
  16751=>"101110101",
  16752=>"001011001",
  16753=>"001000111",
  16754=>"101101100",
  16755=>"110011101",
  16756=>"100010001",
  16757=>"101111010",
  16758=>"010010101",
  16759=>"010110100",
  16760=>"100100010",
  16761=>"010010110",
  16762=>"100111111",
  16763=>"101111000",
  16764=>"111101010",
  16765=>"100111100",
  16766=>"011011100",
  16767=>"110100100",
  16768=>"001111111",
  16769=>"111111010",
  16770=>"011001001",
  16771=>"010100011",
  16772=>"011000000",
  16773=>"110001000",
  16774=>"100111100",
  16775=>"101110000",
  16776=>"000001011",
  16777=>"011000101",
  16778=>"010011000",
  16779=>"010001010",
  16780=>"001101110",
  16781=>"100110000",
  16782=>"111011100",
  16783=>"101001000",
  16784=>"111010111",
  16785=>"010011001",
  16786=>"001010100",
  16787=>"101000010",
  16788=>"001000000",
  16789=>"010010011",
  16790=>"011001000",
  16791=>"111101000",
  16792=>"101011110",
  16793=>"010000011",
  16794=>"001010000",
  16795=>"001000100",
  16796=>"110110000",
  16797=>"110010111",
  16798=>"001100101",
  16799=>"001010000",
  16800=>"001110111",
  16801=>"101110010",
  16802=>"101001111",
  16803=>"111001010",
  16804=>"011000001",
  16805=>"000001000",
  16806=>"000010011",
  16807=>"111001010",
  16808=>"100101011",
  16809=>"111100101",
  16810=>"000101000",
  16811=>"001001010",
  16812=>"010110110",
  16813=>"100100001",
  16814=>"011000011",
  16815=>"101010000",
  16816=>"001001110",
  16817=>"100111011",
  16818=>"000101001",
  16819=>"000110000",
  16820=>"010111000",
  16821=>"000010110",
  16822=>"001011001",
  16823=>"011100110",
  16824=>"110101000",
  16825=>"010000101",
  16826=>"110010100",
  16827=>"010001010",
  16828=>"101000000",
  16829=>"001001100",
  16830=>"001100110",
  16831=>"110110010",
  16832=>"100010000",
  16833=>"100010101",
  16834=>"000011101",
  16835=>"111001111",
  16836=>"010111010",
  16837=>"111011010",
  16838=>"011000111",
  16839=>"000010110",
  16840=>"011000111",
  16841=>"011001101",
  16842=>"001010000",
  16843=>"001101101",
  16844=>"000000111",
  16845=>"010000000",
  16846=>"111110011",
  16847=>"000100011",
  16848=>"011100011",
  16849=>"011000100",
  16850=>"001100100",
  16851=>"011000010",
  16852=>"011100111",
  16853=>"101100101",
  16854=>"000010100",
  16855=>"001111000",
  16856=>"101110011",
  16857=>"101010110",
  16858=>"110101110",
  16859=>"011111000",
  16860=>"111011000",
  16861=>"011001101",
  16862=>"110100001",
  16863=>"010100101",
  16864=>"101111111",
  16865=>"011011010",
  16866=>"101100110",
  16867=>"111010010",
  16868=>"101100100",
  16869=>"111111001",
  16870=>"000000001",
  16871=>"011011100",
  16872=>"101111100",
  16873=>"110010001",
  16874=>"100101011",
  16875=>"101001100",
  16876=>"011100010",
  16877=>"101010011",
  16878=>"010111100",
  16879=>"010010111",
  16880=>"010110010",
  16881=>"011011011",
  16882=>"011001100",
  16883=>"101011100",
  16884=>"110001101",
  16885=>"111010101",
  16886=>"010111110",
  16887=>"001111101",
  16888=>"111001111",
  16889=>"001111100",
  16890=>"011001111",
  16891=>"111011010",
  16892=>"000000100",
  16893=>"000100011",
  16894=>"010000101",
  16895=>"100001000",
  16896=>"100110011",
  16897=>"100000110",
  16898=>"111001101",
  16899=>"110001010",
  16900=>"100001100",
  16901=>"111010001",
  16902=>"110011101",
  16903=>"010101111",
  16904=>"010110111",
  16905=>"101111111",
  16906=>"101001110",
  16907=>"010011001",
  16908=>"110001000",
  16909=>"101011110",
  16910=>"110000000",
  16911=>"101001000",
  16912=>"010000000",
  16913=>"001010000",
  16914=>"110000011",
  16915=>"110110000",
  16916=>"001111011",
  16917=>"111111101",
  16918=>"100011111",
  16919=>"011100110",
  16920=>"001001111",
  16921=>"010001011",
  16922=>"000110110",
  16923=>"001010001",
  16924=>"000010111",
  16925=>"101011001",
  16926=>"011011010",
  16927=>"001000110",
  16928=>"110110001",
  16929=>"001101010",
  16930=>"010111111",
  16931=>"101000001",
  16932=>"101111100",
  16933=>"111001110",
  16934=>"000000111",
  16935=>"000010111",
  16936=>"110011101",
  16937=>"111100101",
  16938=>"010111110",
  16939=>"110010111",
  16940=>"011001001",
  16941=>"100001100",
  16942=>"000010100",
  16943=>"001110001",
  16944=>"100100001",
  16945=>"000100011",
  16946=>"000011000",
  16947=>"111110100",
  16948=>"011111001",
  16949=>"111011000",
  16950=>"000100011",
  16951=>"000001000",
  16952=>"111100011",
  16953=>"001110000",
  16954=>"101110100",
  16955=>"001101110",
  16956=>"100011010",
  16957=>"000011000",
  16958=>"101100100",
  16959=>"001110111",
  16960=>"110110100",
  16961=>"100100100",
  16962=>"001110110",
  16963=>"100110111",
  16964=>"110101000",
  16965=>"101101100",
  16966=>"110111010",
  16967=>"110001100",
  16968=>"010001101",
  16969=>"010010101",
  16970=>"011100111",
  16971=>"110000000",
  16972=>"011111000",
  16973=>"010011001",
  16974=>"110010110",
  16975=>"100110011",
  16976=>"101111100",
  16977=>"000100110",
  16978=>"000010101",
  16979=>"101100110",
  16980=>"010110000",
  16981=>"110110111",
  16982=>"001100000",
  16983=>"110101010",
  16984=>"001110011",
  16985=>"001011000",
  16986=>"000001100",
  16987=>"000010000",
  16988=>"000011100",
  16989=>"100011000",
  16990=>"111010011",
  16991=>"111100110",
  16992=>"010100011",
  16993=>"010000011",
  16994=>"000100000",
  16995=>"000101110",
  16996=>"011011001",
  16997=>"011101011",
  16998=>"000101111",
  16999=>"111010100",
  17000=>"101111010",
  17001=>"110110111",
  17002=>"110001001",
  17003=>"101110100",
  17004=>"001100100",
  17005=>"000111000",
  17006=>"001110111",
  17007=>"000011010",
  17008=>"010101001",
  17009=>"100000100",
  17010=>"010011001",
  17011=>"100101001",
  17012=>"010010011",
  17013=>"111111011",
  17014=>"101111000",
  17015=>"111110111",
  17016=>"011000100",
  17017=>"101010011",
  17018=>"111010000",
  17019=>"101101000",
  17020=>"111110010",
  17021=>"111011010",
  17022=>"101111100",
  17023=>"110000110",
  17024=>"100010101",
  17025=>"101001101",
  17026=>"000111001",
  17027=>"001110010",
  17028=>"010001111",
  17029=>"101000011",
  17030=>"011001101",
  17031=>"111101000",
  17032=>"101110000",
  17033=>"001011000",
  17034=>"000001100",
  17035=>"000000000",
  17036=>"010000011",
  17037=>"010000100",
  17038=>"111101011",
  17039=>"010010101",
  17040=>"110110101",
  17041=>"010111001",
  17042=>"010000000",
  17043=>"101100011",
  17044=>"011111001",
  17045=>"100101001",
  17046=>"110010100",
  17047=>"000011011",
  17048=>"100101111",
  17049=>"100101101",
  17050=>"000101101",
  17051=>"100100010",
  17052=>"000010000",
  17053=>"001101111",
  17054=>"110111100",
  17055=>"000111111",
  17056=>"000000010",
  17057=>"100101110",
  17058=>"001110010",
  17059=>"110110100",
  17060=>"101000011",
  17061=>"000011110",
  17062=>"000100010",
  17063=>"000001000",
  17064=>"111111001",
  17065=>"101101111",
  17066=>"100101010",
  17067=>"001010000",
  17068=>"110000101",
  17069=>"100010011",
  17070=>"011110111",
  17071=>"000010000",
  17072=>"000010110",
  17073=>"101000001",
  17074=>"011011101",
  17075=>"001100111",
  17076=>"100001000",
  17077=>"010000110",
  17078=>"110011011",
  17079=>"000001101",
  17080=>"101111011",
  17081=>"101110000",
  17082=>"101110110",
  17083=>"111100001",
  17084=>"101100001",
  17085=>"110000111",
  17086=>"001000000",
  17087=>"111010111",
  17088=>"101111101",
  17089=>"001000111",
  17090=>"011100110",
  17091=>"111101101",
  17092=>"001101111",
  17093=>"000110101",
  17094=>"000011110",
  17095=>"000000101",
  17096=>"010011110",
  17097=>"110110110",
  17098=>"010001101",
  17099=>"010111010",
  17100=>"110011000",
  17101=>"010100010",
  17102=>"111111100",
  17103=>"110011010",
  17104=>"000010000",
  17105=>"100001000",
  17106=>"100011000",
  17107=>"000001001",
  17108=>"111111001",
  17109=>"100101001",
  17110=>"001100001",
  17111=>"111000000",
  17112=>"100111111",
  17113=>"001100100",
  17114=>"011100111",
  17115=>"001010111",
  17116=>"000010110",
  17117=>"011000011",
  17118=>"101001010",
  17119=>"100010010",
  17120=>"111110100",
  17121=>"100000001",
  17122=>"110001100",
  17123=>"010001000",
  17124=>"111111000",
  17125=>"101011101",
  17126=>"010001000",
  17127=>"011001110",
  17128=>"100011110",
  17129=>"001101011",
  17130=>"000001111",
  17131=>"111111011",
  17132=>"000100101",
  17133=>"001000010",
  17134=>"110101100",
  17135=>"101101101",
  17136=>"100111011",
  17137=>"000001010",
  17138=>"010010100",
  17139=>"011001111",
  17140=>"010010000",
  17141=>"010101101",
  17142=>"111101101",
  17143=>"010100010",
  17144=>"000010100",
  17145=>"001111011",
  17146=>"110001100",
  17147=>"100111011",
  17148=>"110010101",
  17149=>"111010011",
  17150=>"011000101",
  17151=>"010011010",
  17152=>"011101000",
  17153=>"001010111",
  17154=>"010111000",
  17155=>"101111111",
  17156=>"001010111",
  17157=>"001000000",
  17158=>"110011010",
  17159=>"111011110",
  17160=>"010001100",
  17161=>"011010110",
  17162=>"110000110",
  17163=>"110010010",
  17164=>"111011110",
  17165=>"101101000",
  17166=>"111100010",
  17167=>"010111110",
  17168=>"100100110",
  17169=>"100100101",
  17170=>"000010001",
  17171=>"111001001",
  17172=>"101010010",
  17173=>"100001110",
  17174=>"010000010",
  17175=>"001011011",
  17176=>"000101010",
  17177=>"100001110",
  17178=>"100000010",
  17179=>"010101011",
  17180=>"000111100",
  17181=>"111010011",
  17182=>"111110111",
  17183=>"100010000",
  17184=>"100100100",
  17185=>"111001101",
  17186=>"000010010",
  17187=>"001110010",
  17188=>"111100111",
  17189=>"111011111",
  17190=>"000010010",
  17191=>"110011100",
  17192=>"011100000",
  17193=>"111001100",
  17194=>"001101101",
  17195=>"011011010",
  17196=>"110010110",
  17197=>"000000100",
  17198=>"011101110",
  17199=>"010010101",
  17200=>"010000101",
  17201=>"111111001",
  17202=>"110000000",
  17203=>"000110000",
  17204=>"110000101",
  17205=>"100100100",
  17206=>"100001010",
  17207=>"001101110",
  17208=>"000101010",
  17209=>"010011101",
  17210=>"110010111",
  17211=>"000011111",
  17212=>"110011100",
  17213=>"011000100",
  17214=>"001000111",
  17215=>"000011011",
  17216=>"001001011",
  17217=>"100011101",
  17218=>"010101100",
  17219=>"110011001",
  17220=>"110101001",
  17221=>"100000111",
  17222=>"111111101",
  17223=>"011000101",
  17224=>"000110000",
  17225=>"010100110",
  17226=>"000100100",
  17227=>"101001001",
  17228=>"111011111",
  17229=>"100011110",
  17230=>"001010110",
  17231=>"001011100",
  17232=>"011010111",
  17233=>"100011010",
  17234=>"000100000",
  17235=>"100010010",
  17236=>"110100110",
  17237=>"011110000",
  17238=>"101111000",
  17239=>"000110001",
  17240=>"010001001",
  17241=>"111001100",
  17242=>"101111111",
  17243=>"001000001",
  17244=>"010100010",
  17245=>"111001100",
  17246=>"000011110",
  17247=>"001010000",
  17248=>"010001111",
  17249=>"111100111",
  17250=>"000010001",
  17251=>"010110111",
  17252=>"001001000",
  17253=>"001010111",
  17254=>"101110001",
  17255=>"001100110",
  17256=>"110000010",
  17257=>"010110010",
  17258=>"010101000",
  17259=>"101100111",
  17260=>"000111100",
  17261=>"000011110",
  17262=>"111100000",
  17263=>"101010000",
  17264=>"011101100",
  17265=>"111110101",
  17266=>"100000001",
  17267=>"011111011",
  17268=>"100110001",
  17269=>"101000000",
  17270=>"111100100",
  17271=>"001000011",
  17272=>"001101110",
  17273=>"110001100",
  17274=>"011011011",
  17275=>"101000100",
  17276=>"100011000",
  17277=>"011100010",
  17278=>"000010001",
  17279=>"000010100",
  17280=>"000010000",
  17281=>"011110101",
  17282=>"001110011",
  17283=>"100100000",
  17284=>"001011001",
  17285=>"011011010",
  17286=>"011010011",
  17287=>"111001101",
  17288=>"011100001",
  17289=>"110011001",
  17290=>"000101101",
  17291=>"100010110",
  17292=>"001100000",
  17293=>"100011100",
  17294=>"001011100",
  17295=>"110000100",
  17296=>"001000111",
  17297=>"100010110",
  17298=>"000110110",
  17299=>"000100000",
  17300=>"101011000",
  17301=>"110101110",
  17302=>"111000011",
  17303=>"101011101",
  17304=>"101010001",
  17305=>"011010011",
  17306=>"001111011",
  17307=>"011110110",
  17308=>"001111111",
  17309=>"000101010",
  17310=>"110110011",
  17311=>"101001000",
  17312=>"000110101",
  17313=>"000111111",
  17314=>"011101000",
  17315=>"000011000",
  17316=>"100011010",
  17317=>"100000100",
  17318=>"101100010",
  17319=>"000110000",
  17320=>"001101100",
  17321=>"000101001",
  17322=>"100111001",
  17323=>"101110000",
  17324=>"101001011",
  17325=>"110010111",
  17326=>"110100001",
  17327=>"100000100",
  17328=>"111111100",
  17329=>"001100011",
  17330=>"000000101",
  17331=>"111111110",
  17332=>"011101110",
  17333=>"000110101",
  17334=>"011111101",
  17335=>"011101011",
  17336=>"001101111",
  17337=>"110100101",
  17338=>"000101001",
  17339=>"000010100",
  17340=>"100101101",
  17341=>"000110111",
  17342=>"101110011",
  17343=>"111011111",
  17344=>"011100100",
  17345=>"001110101",
  17346=>"111101100",
  17347=>"011110011",
  17348=>"110110110",
  17349=>"111101101",
  17350=>"010101011",
  17351=>"101100110",
  17352=>"010011101",
  17353=>"110100110",
  17354=>"101000000",
  17355=>"110101100",
  17356=>"001001011",
  17357=>"011111111",
  17358=>"110000000",
  17359=>"011000110",
  17360=>"011000111",
  17361=>"111011000",
  17362=>"110110110",
  17363=>"111101111",
  17364=>"111100111",
  17365=>"010001100",
  17366=>"010010001",
  17367=>"010100111",
  17368=>"001101101",
  17369=>"001001101",
  17370=>"101110011",
  17371=>"000110101",
  17372=>"110011011",
  17373=>"110011000",
  17374=>"111110111",
  17375=>"011111000",
  17376=>"101001110",
  17377=>"011110110",
  17378=>"111010000",
  17379=>"110000111",
  17380=>"001100110",
  17381=>"111101111",
  17382=>"111111011",
  17383=>"011101101",
  17384=>"011101111",
  17385=>"000100101",
  17386=>"000000111",
  17387=>"111111011",
  17388=>"010001001",
  17389=>"001000111",
  17390=>"011101111",
  17391=>"001010011",
  17392=>"001000011",
  17393=>"101010000",
  17394=>"000010111",
  17395=>"001111100",
  17396=>"100110010",
  17397=>"000111010",
  17398=>"111000000",
  17399=>"010110100",
  17400=>"110110010",
  17401=>"010000011",
  17402=>"010011000",
  17403=>"110011101",
  17404=>"010010001",
  17405=>"100111110",
  17406=>"111110111",
  17407=>"010101001",
  17408=>"010010010",
  17409=>"010011101",
  17410=>"111101111",
  17411=>"001000110",
  17412=>"010011000",
  17413=>"111110000",
  17414=>"010000000",
  17415=>"110001101",
  17416=>"111100110",
  17417=>"000010111",
  17418=>"110110110",
  17419=>"111011100",
  17420=>"100100110",
  17421=>"111101010",
  17422=>"010101101",
  17423=>"101101111",
  17424=>"111011101",
  17425=>"101010100",
  17426=>"011101110",
  17427=>"001001111",
  17428=>"100001000",
  17429=>"000000010",
  17430=>"101110111",
  17431=>"011100010",
  17432=>"010110010",
  17433=>"010001000",
  17434=>"110111110",
  17435=>"001101011",
  17436=>"010111101",
  17437=>"000111111",
  17438=>"111101111",
  17439=>"011110100",
  17440=>"101110111",
  17441=>"111001101",
  17442=>"000000100",
  17443=>"001010001",
  17444=>"001011011",
  17445=>"100100001",
  17446=>"001011101",
  17447=>"010110111",
  17448=>"010010100",
  17449=>"101001010",
  17450=>"111010011",
  17451=>"101011111",
  17452=>"101000111",
  17453=>"101011111",
  17454=>"000011011",
  17455=>"110001010",
  17456=>"110110100",
  17457=>"011101000",
  17458=>"100000111",
  17459=>"100101011",
  17460=>"001001000",
  17461=>"000101011",
  17462=>"111111111",
  17463=>"111011000",
  17464=>"001010010",
  17465=>"110111110",
  17466=>"100011011",
  17467=>"000100100",
  17468=>"001100010",
  17469=>"010100110",
  17470=>"000010010",
  17471=>"111101100",
  17472=>"001000011",
  17473=>"000110110",
  17474=>"011010111",
  17475=>"101000010",
  17476=>"100011110",
  17477=>"010010101",
  17478=>"010100111",
  17479=>"100010000",
  17480=>"001101110",
  17481=>"010110011",
  17482=>"001001011",
  17483=>"100100111",
  17484=>"000000100",
  17485=>"000001100",
  17486=>"111100100",
  17487=>"000101101",
  17488=>"111110110",
  17489=>"111100010",
  17490=>"110001000",
  17491=>"100010110",
  17492=>"000011101",
  17493=>"011101101",
  17494=>"001100000",
  17495=>"101100111",
  17496=>"110110011",
  17497=>"010011001",
  17498=>"010101111",
  17499=>"111100110",
  17500=>"001010011",
  17501=>"011100010",
  17502=>"100100100",
  17503=>"100000111",
  17504=>"100010000",
  17505=>"110111011",
  17506=>"011110111",
  17507=>"111100111",
  17508=>"011101110",
  17509=>"111101110",
  17510=>"100101110",
  17511=>"011011001",
  17512=>"111100010",
  17513=>"110000000",
  17514=>"000010011",
  17515=>"111011011",
  17516=>"101010100",
  17517=>"000111011",
  17518=>"011101110",
  17519=>"101011001",
  17520=>"101101101",
  17521=>"101001100",
  17522=>"110110000",
  17523=>"111110101",
  17524=>"000001100",
  17525=>"110111100",
  17526=>"011001001",
  17527=>"101000100",
  17528=>"001010101",
  17529=>"001101000",
  17530=>"110100101",
  17531=>"010001001",
  17532=>"001100110",
  17533=>"001000111",
  17534=>"110010010",
  17535=>"101101110",
  17536=>"000000100",
  17537=>"111011101",
  17538=>"011011001",
  17539=>"101000001",
  17540=>"111111101",
  17541=>"000001000",
  17542=>"110101011",
  17543=>"111001001",
  17544=>"111100100",
  17545=>"001000001",
  17546=>"010100000",
  17547=>"000001010",
  17548=>"011010001",
  17549=>"110011010",
  17550=>"001010001",
  17551=>"100000111",
  17552=>"011111010",
  17553=>"010100010",
  17554=>"010111011",
  17555=>"011001110",
  17556=>"101001111",
  17557=>"011101011",
  17558=>"111100101",
  17559=>"111011001",
  17560=>"110000000",
  17561=>"001100010",
  17562=>"111010110",
  17563=>"010001101",
  17564=>"000010110",
  17565=>"010001110",
  17566=>"001011000",
  17567=>"011010001",
  17568=>"100000010",
  17569=>"010011011",
  17570=>"101001110",
  17571=>"100101011",
  17572=>"011100100",
  17573=>"101101010",
  17574=>"100101011",
  17575=>"110110000",
  17576=>"101111100",
  17577=>"011000100",
  17578=>"010111000",
  17579=>"000000010",
  17580=>"101000011",
  17581=>"000101100",
  17582=>"101110000",
  17583=>"101100101",
  17584=>"001111001",
  17585=>"010000001",
  17586=>"000010010",
  17587=>"000000101",
  17588=>"010011000",
  17589=>"100100110",
  17590=>"010001110",
  17591=>"101110111",
  17592=>"000111001",
  17593=>"100100111",
  17594=>"000110101",
  17595=>"011011011",
  17596=>"001010010",
  17597=>"100011000",
  17598=>"101100001",
  17599=>"110011100",
  17600=>"011110100",
  17601=>"111011100",
  17602=>"000111011",
  17603=>"110101110",
  17604=>"010100011",
  17605=>"101100000",
  17606=>"000011001",
  17607=>"101011100",
  17608=>"101110111",
  17609=>"101100101",
  17610=>"100101100",
  17611=>"101001011",
  17612=>"000110110",
  17613=>"101110110",
  17614=>"111111011",
  17615=>"111001011",
  17616=>"110000100",
  17617=>"111011110",
  17618=>"100100000",
  17619=>"110111110",
  17620=>"011110110",
  17621=>"010110000",
  17622=>"101001000",
  17623=>"100110001",
  17624=>"111101100",
  17625=>"000011101",
  17626=>"000001010",
  17627=>"101111011",
  17628=>"011010110",
  17629=>"010001001",
  17630=>"110011111",
  17631=>"101000000",
  17632=>"010010111",
  17633=>"111011010",
  17634=>"011011100",
  17635=>"001010101",
  17636=>"001110101",
  17637=>"111101010",
  17638=>"000001001",
  17639=>"101011001",
  17640=>"001111011",
  17641=>"111011001",
  17642=>"000011001",
  17643=>"000100001",
  17644=>"010010111",
  17645=>"100111011",
  17646=>"001001100",
  17647=>"111000000",
  17648=>"001011111",
  17649=>"010100111",
  17650=>"001101111",
  17651=>"010010000",
  17652=>"011111111",
  17653=>"001110101",
  17654=>"110001111",
  17655=>"101011100",
  17656=>"100000001",
  17657=>"011111011",
  17658=>"100101100",
  17659=>"010111110",
  17660=>"110001000",
  17661=>"100000110",
  17662=>"100000111",
  17663=>"101111101",
  17664=>"110001011",
  17665=>"111101101",
  17666=>"000111011",
  17667=>"100100101",
  17668=>"000110000",
  17669=>"101101101",
  17670=>"111101101",
  17671=>"001001000",
  17672=>"000101011",
  17673=>"010010110",
  17674=>"000000001",
  17675=>"011100010",
  17676=>"100010001",
  17677=>"011000010",
  17678=>"110010000",
  17679=>"000100110",
  17680=>"101101100",
  17681=>"101011110",
  17682=>"011000100",
  17683=>"100000111",
  17684=>"110100110",
  17685=>"110011110",
  17686=>"001111111",
  17687=>"111110111",
  17688=>"000100100",
  17689=>"101000110",
  17690=>"101001011",
  17691=>"010101001",
  17692=>"000100111",
  17693=>"101101110",
  17694=>"110010110",
  17695=>"001000100",
  17696=>"101000101",
  17697=>"100111101",
  17698=>"110001010",
  17699=>"010100111",
  17700=>"001101101",
  17701=>"111010101",
  17702=>"001111001",
  17703=>"011100111",
  17704=>"011101011",
  17705=>"011110111",
  17706=>"110000010",
  17707=>"101011111",
  17708=>"101000001",
  17709=>"101111101",
  17710=>"101110100",
  17711=>"011110100",
  17712=>"101111101",
  17713=>"011101001",
  17714=>"001001000",
  17715=>"010111110",
  17716=>"011000100",
  17717=>"001011001",
  17718=>"010111110",
  17719=>"100110010",
  17720=>"000011000",
  17721=>"001011001",
  17722=>"110000000",
  17723=>"000111000",
  17724=>"111001110",
  17725=>"110110101",
  17726=>"001010000",
  17727=>"100001010",
  17728=>"000100110",
  17729=>"100001001",
  17730=>"110111111",
  17731=>"011101111",
  17732=>"111001110",
  17733=>"000101000",
  17734=>"100110111",
  17735=>"010010110",
  17736=>"000100110",
  17737=>"100001001",
  17738=>"110100111",
  17739=>"100001000",
  17740=>"101011001",
  17741=>"110110000",
  17742=>"011011111",
  17743=>"010100100",
  17744=>"011000001",
  17745=>"000101110",
  17746=>"001011000",
  17747=>"000100001",
  17748=>"011010000",
  17749=>"111111100",
  17750=>"011011010",
  17751=>"111000000",
  17752=>"011100101",
  17753=>"000110100",
  17754=>"101111000",
  17755=>"111100001",
  17756=>"010000101",
  17757=>"110000100",
  17758=>"110100010",
  17759=>"010000000",
  17760=>"111110111",
  17761=>"010011111",
  17762=>"101111011",
  17763=>"000001111",
  17764=>"000110110",
  17765=>"000000011",
  17766=>"111100110",
  17767=>"111110000",
  17768=>"001010100",
  17769=>"101101100",
  17770=>"001101110",
  17771=>"001001011",
  17772=>"110111110",
  17773=>"111101001",
  17774=>"101110101",
  17775=>"111010011",
  17776=>"000111001",
  17777=>"010000000",
  17778=>"010101000",
  17779=>"000101101",
  17780=>"110011000",
  17781=>"000000001",
  17782=>"001000000",
  17783=>"000100001",
  17784=>"010000100",
  17785=>"111110001",
  17786=>"001100100",
  17787=>"101101111",
  17788=>"100101011",
  17789=>"101010010",
  17790=>"010111000",
  17791=>"011110100",
  17792=>"000010011",
  17793=>"000100001",
  17794=>"011011101",
  17795=>"100010111",
  17796=>"011001101",
  17797=>"011010011",
  17798=>"111010110",
  17799=>"100000010",
  17800=>"010000101",
  17801=>"111101110",
  17802=>"111100011",
  17803=>"010101010",
  17804=>"001000101",
  17805=>"011000001",
  17806=>"111101110",
  17807=>"111000101",
  17808=>"001100011",
  17809=>"010101000",
  17810=>"001011101",
  17811=>"010100011",
  17812=>"010100000",
  17813=>"011001100",
  17814=>"111111101",
  17815=>"101000101",
  17816=>"100001100",
  17817=>"101001010",
  17818=>"110110001",
  17819=>"111010011",
  17820=>"010001010",
  17821=>"001101110",
  17822=>"110100101",
  17823=>"000110010",
  17824=>"010001111",
  17825=>"000000101",
  17826=>"010110111",
  17827=>"111101100",
  17828=>"011100001",
  17829=>"111101001",
  17830=>"110110000",
  17831=>"010010011",
  17832=>"001001001",
  17833=>"101110101",
  17834=>"110001000",
  17835=>"100000010",
  17836=>"011101011",
  17837=>"000000010",
  17838=>"001110000",
  17839=>"010111011",
  17840=>"000010010",
  17841=>"010111011",
  17842=>"001011000",
  17843=>"110111000",
  17844=>"011111010",
  17845=>"111111111",
  17846=>"111001001",
  17847=>"101010101",
  17848=>"010000001",
  17849=>"000000111",
  17850=>"010010111",
  17851=>"110110011",
  17852=>"011001000",
  17853=>"111001001",
  17854=>"001010110",
  17855=>"111001011",
  17856=>"011001010",
  17857=>"010100000",
  17858=>"111110000",
  17859=>"010100111",
  17860=>"010000100",
  17861=>"011101000",
  17862=>"111110000",
  17863=>"000100000",
  17864=>"110001010",
  17865=>"010101001",
  17866=>"010110111",
  17867=>"111101011",
  17868=>"110100010",
  17869=>"000110001",
  17870=>"000101001",
  17871=>"000100100",
  17872=>"000111100",
  17873=>"111110001",
  17874=>"110111101",
  17875=>"000000101",
  17876=>"010101111",
  17877=>"100001010",
  17878=>"010110101",
  17879=>"011001011",
  17880=>"000111101",
  17881=>"111001010",
  17882=>"000000000",
  17883=>"110010000",
  17884=>"011000100",
  17885=>"011010000",
  17886=>"101010000",
  17887=>"100010111",
  17888=>"110110110",
  17889=>"100001111",
  17890=>"011011100",
  17891=>"100110110",
  17892=>"110111011",
  17893=>"111001101",
  17894=>"001101011",
  17895=>"010010011",
  17896=>"110010010",
  17897=>"011111110",
  17898=>"111000110",
  17899=>"001111000",
  17900=>"001000000",
  17901=>"010001100",
  17902=>"011010000",
  17903=>"110011010",
  17904=>"111110111",
  17905=>"111010000",
  17906=>"011011110",
  17907=>"011000000",
  17908=>"100101011",
  17909=>"000100000",
  17910=>"011101000",
  17911=>"101010000",
  17912=>"010001000",
  17913=>"100100101",
  17914=>"111110010",
  17915=>"000110010",
  17916=>"011010111",
  17917=>"101110101",
  17918=>"110111010",
  17919=>"011111110",
  17920=>"110000000",
  17921=>"111010100",
  17922=>"111101111",
  17923=>"111000011",
  17924=>"111001101",
  17925=>"100011011",
  17926=>"111101011",
  17927=>"010110110",
  17928=>"011010011",
  17929=>"110111100",
  17930=>"001011010",
  17931=>"000011011",
  17932=>"001100001",
  17933=>"010011110",
  17934=>"010100000",
  17935=>"010111011",
  17936=>"010010101",
  17937=>"000110101",
  17938=>"111101000",
  17939=>"110011111",
  17940=>"010100100",
  17941=>"100101000",
  17942=>"111110110",
  17943=>"100100111",
  17944=>"101110111",
  17945=>"110111001",
  17946=>"100110000",
  17947=>"110010000",
  17948=>"110001010",
  17949=>"100110000",
  17950=>"111101011",
  17951=>"111000001",
  17952=>"100001110",
  17953=>"011100110",
  17954=>"000000000",
  17955=>"111011101",
  17956=>"011101010",
  17957=>"000010001",
  17958=>"110010111",
  17959=>"100110100",
  17960=>"000111011",
  17961=>"001111000",
  17962=>"000001010",
  17963=>"011001110",
  17964=>"010100100",
  17965=>"001100011",
  17966=>"111000111",
  17967=>"100110100",
  17968=>"000110001",
  17969=>"000101111",
  17970=>"110000100",
  17971=>"111111101",
  17972=>"011101111",
  17973=>"111100111",
  17974=>"101111000",
  17975=>"110000010",
  17976=>"110101011",
  17977=>"110000000",
  17978=>"000000100",
  17979=>"111011110",
  17980=>"110101000",
  17981=>"111110100",
  17982=>"010011010",
  17983=>"101101101",
  17984=>"111000010",
  17985=>"010110010",
  17986=>"100010010",
  17987=>"011111010",
  17988=>"111110010",
  17989=>"110110000",
  17990=>"000011111",
  17991=>"101110010",
  17992=>"100010011",
  17993=>"010001001",
  17994=>"000110000",
  17995=>"101011000",
  17996=>"100000000",
  17997=>"011101111",
  17998=>"100000110",
  17999=>"100011011",
  18000=>"010100111",
  18001=>"110010010",
  18002=>"100000110",
  18003=>"011100001",
  18004=>"111111110",
  18005=>"101000011",
  18006=>"001100001",
  18007=>"101111000",
  18008=>"010011101",
  18009=>"010101100",
  18010=>"001000010",
  18011=>"110000010",
  18012=>"010010111",
  18013=>"111101010",
  18014=>"010101010",
  18015=>"010001101",
  18016=>"100000101",
  18017=>"110000110",
  18018=>"001100111",
  18019=>"000001101",
  18020=>"101100000",
  18021=>"111111100",
  18022=>"001110000",
  18023=>"101101011",
  18024=>"101100110",
  18025=>"011011100",
  18026=>"011001111",
  18027=>"111101101",
  18028=>"011111010",
  18029=>"011110001",
  18030=>"010010110",
  18031=>"110001011",
  18032=>"010010010",
  18033=>"100001100",
  18034=>"100100010",
  18035=>"111101111",
  18036=>"000000010",
  18037=>"101001001",
  18038=>"010111111",
  18039=>"011110110",
  18040=>"011010000",
  18041=>"001110101",
  18042=>"110110011",
  18043=>"011111100",
  18044=>"101010001",
  18045=>"001111010",
  18046=>"000001001",
  18047=>"010110111",
  18048=>"111000011",
  18049=>"010010110",
  18050=>"010100111",
  18051=>"001001001",
  18052=>"010010100",
  18053=>"010001001",
  18054=>"001000111",
  18055=>"100111010",
  18056=>"010100111",
  18057=>"010010101",
  18058=>"111111001",
  18059=>"100011111",
  18060=>"111001101",
  18061=>"101111010",
  18062=>"000010010",
  18063=>"000100011",
  18064=>"111110101",
  18065=>"011111001",
  18066=>"000000000",
  18067=>"100000011",
  18068=>"111000000",
  18069=>"110011110",
  18070=>"110010000",
  18071=>"000000010",
  18072=>"010111101",
  18073=>"110001111",
  18074=>"011100010",
  18075=>"010100100",
  18076=>"010101100",
  18077=>"110000011",
  18078=>"000110001",
  18079=>"010111111",
  18080=>"000000110",
  18081=>"001011100",
  18082=>"111001110",
  18083=>"000001000",
  18084=>"101101110",
  18085=>"001000010",
  18086=>"001101010",
  18087=>"000011100",
  18088=>"101001001",
  18089=>"000101100",
  18090=>"110011110",
  18091=>"011010000",
  18092=>"000010111",
  18093=>"001000100",
  18094=>"100111110",
  18095=>"100101000",
  18096=>"001000011",
  18097=>"010010011",
  18098=>"000000000",
  18099=>"111001101",
  18100=>"010111011",
  18101=>"001100011",
  18102=>"000010000",
  18103=>"011100001",
  18104=>"001001101",
  18105=>"001101101",
  18106=>"111111110",
  18107=>"110110001",
  18108=>"110110110",
  18109=>"110111101",
  18110=>"110100011",
  18111=>"000111111",
  18112=>"010101111",
  18113=>"111001111",
  18114=>"111101111",
  18115=>"011010000",
  18116=>"000000110",
  18117=>"000010011",
  18118=>"111100111",
  18119=>"111001000",
  18120=>"001011111",
  18121=>"111111010",
  18122=>"101001110",
  18123=>"110001010",
  18124=>"111011000",
  18125=>"000010000",
  18126=>"100000100",
  18127=>"101000100",
  18128=>"000101111",
  18129=>"010011110",
  18130=>"111000110",
  18131=>"010001000",
  18132=>"001001111",
  18133=>"000000011",
  18134=>"111111110",
  18135=>"110111101",
  18136=>"010111010",
  18137=>"101011111",
  18138=>"110101010",
  18139=>"001010001",
  18140=>"001000011",
  18141=>"111010010",
  18142=>"001100011",
  18143=>"110111100",
  18144=>"100000101",
  18145=>"011010001",
  18146=>"010011101",
  18147=>"000010100",
  18148=>"111000001",
  18149=>"110101001",
  18150=>"000010000",
  18151=>"100011100",
  18152=>"000000000",
  18153=>"010101110",
  18154=>"010010110",
  18155=>"011011010",
  18156=>"100010001",
  18157=>"100100000",
  18158=>"100101110",
  18159=>"000101010",
  18160=>"111011111",
  18161=>"011101100",
  18162=>"111111010",
  18163=>"001110011",
  18164=>"000011100",
  18165=>"000010001",
  18166=>"101101100",
  18167=>"000100001",
  18168=>"100111000",
  18169=>"010001100",
  18170=>"010000100",
  18171=>"101011111",
  18172=>"011010010",
  18173=>"000010000",
  18174=>"110011000",
  18175=>"000101000",
  18176=>"101100001",
  18177=>"010100111",
  18178=>"110010101",
  18179=>"000000101",
  18180=>"101011111",
  18181=>"110000100",
  18182=>"011000101",
  18183=>"001110101",
  18184=>"100110001",
  18185=>"101010101",
  18186=>"010000110",
  18187=>"100000010",
  18188=>"001000110",
  18189=>"100100100",
  18190=>"001001100",
  18191=>"100001111",
  18192=>"000000010",
  18193=>"001000001",
  18194=>"011011111",
  18195=>"111110010",
  18196=>"101010101",
  18197=>"000110101",
  18198=>"001100110",
  18199=>"011100001",
  18200=>"000001100",
  18201=>"110101001",
  18202=>"000100111",
  18203=>"000101110",
  18204=>"011111110",
  18205=>"000111010",
  18206=>"111011111",
  18207=>"111000111",
  18208=>"010010010",
  18209=>"000010011",
  18210=>"001111011",
  18211=>"111100000",
  18212=>"110000011",
  18213=>"101110000",
  18214=>"011101110",
  18215=>"110000101",
  18216=>"110101111",
  18217=>"001000101",
  18218=>"010010111",
  18219=>"001001110",
  18220=>"100010011",
  18221=>"101111110",
  18222=>"110111001",
  18223=>"011101101",
  18224=>"101011001",
  18225=>"110011100",
  18226=>"110100001",
  18227=>"001111011",
  18228=>"010110110",
  18229=>"000100110",
  18230=>"101101111",
  18231=>"001000101",
  18232=>"011100110",
  18233=>"010010110",
  18234=>"000100001",
  18235=>"111101010",
  18236=>"000101010",
  18237=>"010110111",
  18238=>"110101010",
  18239=>"001010110",
  18240=>"100111111",
  18241=>"011100100",
  18242=>"110100010",
  18243=>"100010011",
  18244=>"000111100",
  18245=>"111000000",
  18246=>"010111011",
  18247=>"110011010",
  18248=>"010000101",
  18249=>"100010001",
  18250=>"111010110",
  18251=>"001000101",
  18252=>"000101000",
  18253=>"101101000",
  18254=>"001111001",
  18255=>"110101011",
  18256=>"101001111",
  18257=>"000000010",
  18258=>"000000010",
  18259=>"001110110",
  18260=>"010111101",
  18261=>"111011001",
  18262=>"011011110",
  18263=>"110010011",
  18264=>"001000100",
  18265=>"100010100",
  18266=>"010111011",
  18267=>"111000001",
  18268=>"100011110",
  18269=>"100000001",
  18270=>"011111101",
  18271=>"000001100",
  18272=>"001100001",
  18273=>"001010100",
  18274=>"001010000",
  18275=>"111001110",
  18276=>"111000001",
  18277=>"110001110",
  18278=>"100100101",
  18279=>"110100001",
  18280=>"000000100",
  18281=>"010000000",
  18282=>"100010110",
  18283=>"000100011",
  18284=>"001101110",
  18285=>"010011111",
  18286=>"000010010",
  18287=>"111011110",
  18288=>"111111000",
  18289=>"000101000",
  18290=>"111011111",
  18291=>"110100000",
  18292=>"000001100",
  18293=>"000000010",
  18294=>"010111000",
  18295=>"110111111",
  18296=>"111111111",
  18297=>"000100110",
  18298=>"101010101",
  18299=>"101111000",
  18300=>"000100111",
  18301=>"111001110",
  18302=>"001010000",
  18303=>"011101100",
  18304=>"010001110",
  18305=>"110010001",
  18306=>"100010110",
  18307=>"001111111",
  18308=>"011100100",
  18309=>"010111010",
  18310=>"111111110",
  18311=>"000011100",
  18312=>"001101001",
  18313=>"100011111",
  18314=>"000100101",
  18315=>"101101111",
  18316=>"011010111",
  18317=>"000111010",
  18318=>"000000001",
  18319=>"011001010",
  18320=>"000010000",
  18321=>"111100011",
  18322=>"001001000",
  18323=>"101010001",
  18324=>"110110000",
  18325=>"100010101",
  18326=>"101100000",
  18327=>"000000111",
  18328=>"101011011",
  18329=>"000000000",
  18330=>"111100010",
  18331=>"000010010",
  18332=>"001010010",
  18333=>"100110111",
  18334=>"100011110",
  18335=>"100100110",
  18336=>"001010011",
  18337=>"111100111",
  18338=>"110010011",
  18339=>"100000000",
  18340=>"001011011",
  18341=>"011110000",
  18342=>"011110010",
  18343=>"010000010",
  18344=>"000010101",
  18345=>"001001001",
  18346=>"001111101",
  18347=>"001000111",
  18348=>"100111101",
  18349=>"101101101",
  18350=>"011011000",
  18351=>"011001110",
  18352=>"000000001",
  18353=>"011111011",
  18354=>"001011001",
  18355=>"111100011",
  18356=>"011010000",
  18357=>"110010000",
  18358=>"010110000",
  18359=>"111000100",
  18360=>"001001110",
  18361=>"011000010",
  18362=>"111100110",
  18363=>"101011001",
  18364=>"111011110",
  18365=>"000001000",
  18366=>"011110000",
  18367=>"110100011",
  18368=>"111110100",
  18369=>"100110101",
  18370=>"100001100",
  18371=>"001100110",
  18372=>"001101001",
  18373=>"011111001",
  18374=>"010010111",
  18375=>"101010101",
  18376=>"011011111",
  18377=>"111110100",
  18378=>"011011110",
  18379=>"011110100",
  18380=>"111101011",
  18381=>"001001111",
  18382=>"000111111",
  18383=>"001000111",
  18384=>"101000100",
  18385=>"001110110",
  18386=>"011101110",
  18387=>"100000001",
  18388=>"111100001",
  18389=>"101001011",
  18390=>"100111011",
  18391=>"011101101",
  18392=>"110110010",
  18393=>"111001011",
  18394=>"110000001",
  18395=>"001011000",
  18396=>"110011101",
  18397=>"110000011",
  18398=>"001110110",
  18399=>"011100001",
  18400=>"111001111",
  18401=>"111011010",
  18402=>"011001111",
  18403=>"010100110",
  18404=>"011110000",
  18405=>"011101111",
  18406=>"100010111",
  18407=>"100111011",
  18408=>"001011011",
  18409=>"100001100",
  18410=>"000011000",
  18411=>"101001010",
  18412=>"101101011",
  18413=>"110110010",
  18414=>"000010111",
  18415=>"011111011",
  18416=>"011010010",
  18417=>"001100100",
  18418=>"101011100",
  18419=>"110110010",
  18420=>"001000010",
  18421=>"010101000",
  18422=>"011111110",
  18423=>"000001111",
  18424=>"000000100",
  18425=>"101000000",
  18426=>"100000001",
  18427=>"000100010",
  18428=>"100100011",
  18429=>"011011000",
  18430=>"010111010",
  18431=>"010000100",
  18432=>"011001111",
  18433=>"111111010",
  18434=>"110100111",
  18435=>"101101100",
  18436=>"100111111",
  18437=>"011110110",
  18438=>"100011011",
  18439=>"010010100",
  18440=>"111011001",
  18441=>"000101101",
  18442=>"111000100",
  18443=>"101011010",
  18444=>"011101001",
  18445=>"000010100",
  18446=>"101111101",
  18447=>"101101111",
  18448=>"000110010",
  18449=>"000010000",
  18450=>"000011111",
  18451=>"001001001",
  18452=>"000001100",
  18453=>"011100000",
  18454=>"101100000",
  18455=>"100010101",
  18456=>"001001000",
  18457=>"000001111",
  18458=>"110011101",
  18459=>"011101100",
  18460=>"100001101",
  18461=>"000000001",
  18462=>"001000001",
  18463=>"001000110",
  18464=>"000011111",
  18465=>"001110101",
  18466=>"010011110",
  18467=>"101011000",
  18468=>"111011011",
  18469=>"011110011",
  18470=>"111111011",
  18471=>"001101111",
  18472=>"011100010",
  18473=>"001111101",
  18474=>"111001101",
  18475=>"100011011",
  18476=>"011101000",
  18477=>"000111000",
  18478=>"100111101",
  18479=>"110110110",
  18480=>"010001011",
  18481=>"011011000",
  18482=>"101010000",
  18483=>"101111111",
  18484=>"001111011",
  18485=>"001111001",
  18486=>"110001100",
  18487=>"111001011",
  18488=>"011001001",
  18489=>"001000101",
  18490=>"001111001",
  18491=>"110110001",
  18492=>"000010100",
  18493=>"011100111",
  18494=>"010111001",
  18495=>"001100111",
  18496=>"001111111",
  18497=>"000010110",
  18498=>"011111010",
  18499=>"001011100",
  18500=>"110101011",
  18501=>"000111011",
  18502=>"010001010",
  18503=>"101100010",
  18504=>"111000011",
  18505=>"000001000",
  18506=>"011101001",
  18507=>"101001011",
  18508=>"011010010",
  18509=>"001011010",
  18510=>"100101110",
  18511=>"011001001",
  18512=>"001000011",
  18513=>"101010111",
  18514=>"111100000",
  18515=>"110111010",
  18516=>"000000000",
  18517=>"001011111",
  18518=>"000001111",
  18519=>"010011001",
  18520=>"000100010",
  18521=>"010011101",
  18522=>"010001001",
  18523=>"001001010",
  18524=>"001000011",
  18525=>"101001100",
  18526=>"100000001",
  18527=>"000000101",
  18528=>"000100101",
  18529=>"000110101",
  18530=>"000001010",
  18531=>"000001111",
  18532=>"000000011",
  18533=>"111010010",
  18534=>"100100000",
  18535=>"000010011",
  18536=>"011011010",
  18537=>"011110111",
  18538=>"000001100",
  18539=>"010001011",
  18540=>"101001000",
  18541=>"100110101",
  18542=>"101111001",
  18543=>"000110001",
  18544=>"110011010",
  18545=>"001101001",
  18546=>"111011101",
  18547=>"001000000",
  18548=>"010001100",
  18549=>"100111010",
  18550=>"110110101",
  18551=>"000011100",
  18552=>"010111110",
  18553=>"010011101",
  18554=>"011111110",
  18555=>"100100001",
  18556=>"111110100",
  18557=>"111001010",
  18558=>"111100001",
  18559=>"101101000",
  18560=>"111011011",
  18561=>"101010011",
  18562=>"001111100",
  18563=>"010100011",
  18564=>"101001010",
  18565=>"100011110",
  18566=>"101110001",
  18567=>"000001001",
  18568=>"111011000",
  18569=>"101111000",
  18570=>"010001011",
  18571=>"000000111",
  18572=>"111110111",
  18573=>"010101101",
  18574=>"110101100",
  18575=>"101110110",
  18576=>"101010001",
  18577=>"001011111",
  18578=>"000000000",
  18579=>"011010001",
  18580=>"111101101",
  18581=>"010001010",
  18582=>"010000010",
  18583=>"000110110",
  18584=>"010001101",
  18585=>"111001110",
  18586=>"000000101",
  18587=>"011001010",
  18588=>"111100001",
  18589=>"000001010",
  18590=>"000010001",
  18591=>"101100111",
  18592=>"110100000",
  18593=>"010001111",
  18594=>"110101001",
  18595=>"000000000",
  18596=>"011010001",
  18597=>"000001011",
  18598=>"110100100",
  18599=>"000111001",
  18600=>"111001110",
  18601=>"011011010",
  18602=>"100101000",
  18603=>"111001010",
  18604=>"001001001",
  18605=>"011000101",
  18606=>"000001110",
  18607=>"001000010",
  18608=>"111001000",
  18609=>"101000101",
  18610=>"111111001",
  18611=>"010110101",
  18612=>"111000111",
  18613=>"000100010",
  18614=>"001111100",
  18615=>"101010010",
  18616=>"010001111",
  18617=>"000110110",
  18618=>"010111011",
  18619=>"000100010",
  18620=>"000110010",
  18621=>"010010110",
  18622=>"010100101",
  18623=>"000001101",
  18624=>"011010110",
  18625=>"001100111",
  18626=>"001010000",
  18627=>"010110001",
  18628=>"001011000",
  18629=>"100101011",
  18630=>"000100000",
  18631=>"001011111",
  18632=>"111101010",
  18633=>"101011010",
  18634=>"010101110",
  18635=>"000101000",
  18636=>"101011000",
  18637=>"100111010",
  18638=>"101110110",
  18639=>"100010100",
  18640=>"101000000",
  18641=>"100111010",
  18642=>"011100101",
  18643=>"101100100",
  18644=>"100001101",
  18645=>"010001010",
  18646=>"101000011",
  18647=>"000100111",
  18648=>"100001011",
  18649=>"001010000",
  18650=>"100011100",
  18651=>"000011001",
  18652=>"001011011",
  18653=>"001110001",
  18654=>"010011101",
  18655=>"011110011",
  18656=>"001110101",
  18657=>"111110000",
  18658=>"110100111",
  18659=>"100100110",
  18660=>"101110010",
  18661=>"100101000",
  18662=>"010000000",
  18663=>"110010110",
  18664=>"101100000",
  18665=>"001011110",
  18666=>"100000001",
  18667=>"011010100",
  18668=>"111010101",
  18669=>"111011110",
  18670=>"010010101",
  18671=>"001000000",
  18672=>"001011110",
  18673=>"101100010",
  18674=>"000001001",
  18675=>"000010101",
  18676=>"011000001",
  18677=>"001110111",
  18678=>"011101000",
  18679=>"000110101",
  18680=>"101111010",
  18681=>"001000001",
  18682=>"110011010",
  18683=>"100001001",
  18684=>"101011010",
  18685=>"001010110",
  18686=>"001110001",
  18687=>"011001110",
  18688=>"010111110",
  18689=>"011010111",
  18690=>"010101000",
  18691=>"111001101",
  18692=>"011010000",
  18693=>"011001011",
  18694=>"011010011",
  18695=>"101011001",
  18696=>"001010000",
  18697=>"110000000",
  18698=>"100101111",
  18699=>"000010100",
  18700=>"000000110",
  18701=>"100000110",
  18702=>"110000101",
  18703=>"111100001",
  18704=>"011011110",
  18705=>"110001111",
  18706=>"101001100",
  18707=>"000110100",
  18708=>"111111101",
  18709=>"111001011",
  18710=>"101100001",
  18711=>"111111011",
  18712=>"101100011",
  18713=>"111010010",
  18714=>"011110000",
  18715=>"011100111",
  18716=>"110010001",
  18717=>"000100000",
  18718=>"111110101",
  18719=>"110110101",
  18720=>"010010111",
  18721=>"101110011",
  18722=>"010000100",
  18723=>"100100000",
  18724=>"001101101",
  18725=>"111001010",
  18726=>"000000100",
  18727=>"100110100",
  18728=>"000011001",
  18729=>"100110101",
  18730=>"011111110",
  18731=>"101000011",
  18732=>"110000000",
  18733=>"000100100",
  18734=>"111110010",
  18735=>"001011000",
  18736=>"111010010",
  18737=>"100110111",
  18738=>"111000000",
  18739=>"010010010",
  18740=>"001110000",
  18741=>"101011001",
  18742=>"000000010",
  18743=>"100100111",
  18744=>"100110000",
  18745=>"001010101",
  18746=>"001111110",
  18747=>"100010010",
  18748=>"100001010",
  18749=>"011000010",
  18750=>"101001001",
  18751=>"100101000",
  18752=>"110111101",
  18753=>"000101110",
  18754=>"110001101",
  18755=>"100110010",
  18756=>"111111001",
  18757=>"010001010",
  18758=>"101111111",
  18759=>"001010111",
  18760=>"000000010",
  18761=>"001000010",
  18762=>"111001000",
  18763=>"011001110",
  18764=>"100101101",
  18765=>"111100110",
  18766=>"010010001",
  18767=>"010100100",
  18768=>"011110111",
  18769=>"000001111",
  18770=>"010110000",
  18771=>"100101100",
  18772=>"100000111",
  18773=>"110101110",
  18774=>"101011110",
  18775=>"100100110",
  18776=>"010100100",
  18777=>"101110111",
  18778=>"000011110",
  18779=>"101011000",
  18780=>"101111100",
  18781=>"101101011",
  18782=>"110101110",
  18783=>"111110111",
  18784=>"000110111",
  18785=>"011101001",
  18786=>"110001001",
  18787=>"010000110",
  18788=>"010101000",
  18789=>"000100111",
  18790=>"000110000",
  18791=>"001101001",
  18792=>"100000011",
  18793=>"011001011",
  18794=>"000001011",
  18795=>"111110111",
  18796=>"011000100",
  18797=>"110110000",
  18798=>"100000111",
  18799=>"110001101",
  18800=>"000001001",
  18801=>"110001111",
  18802=>"101000011",
  18803=>"111111100",
  18804=>"111100100",
  18805=>"010001110",
  18806=>"101001111",
  18807=>"111010110",
  18808=>"101000000",
  18809=>"110111100",
  18810=>"101001001",
  18811=>"110011110",
  18812=>"010110101",
  18813=>"000010000",
  18814=>"011101000",
  18815=>"011010100",
  18816=>"000000001",
  18817=>"101010011",
  18818=>"101100110",
  18819=>"011011110",
  18820=>"000101111",
  18821=>"010111110",
  18822=>"001011011",
  18823=>"100011001",
  18824=>"000001010",
  18825=>"100101110",
  18826=>"110011111",
  18827=>"000000110",
  18828=>"001011101",
  18829=>"101110011",
  18830=>"001011011",
  18831=>"101111001",
  18832=>"111100001",
  18833=>"000011000",
  18834=>"110101110",
  18835=>"101000011",
  18836=>"000010100",
  18837=>"000101001",
  18838=>"111110010",
  18839=>"100000010",
  18840=>"101101000",
  18841=>"001000010",
  18842=>"000010001",
  18843=>"110011110",
  18844=>"111100010",
  18845=>"110010011",
  18846=>"001001000",
  18847=>"011110010",
  18848=>"010111110",
  18849=>"111000010",
  18850=>"000000111",
  18851=>"001001000",
  18852=>"110000011",
  18853=>"000100101",
  18854=>"001111101",
  18855=>"000110000",
  18856=>"111101110",
  18857=>"011011101",
  18858=>"110000100",
  18859=>"100100010",
  18860=>"101001001",
  18861=>"000100000",
  18862=>"001000110",
  18863=>"110110110",
  18864=>"010111011",
  18865=>"010010100",
  18866=>"110001101",
  18867=>"100011111",
  18868=>"010000000",
  18869=>"110011001",
  18870=>"011110011",
  18871=>"100111000",
  18872=>"010000100",
  18873=>"100000101",
  18874=>"011111000",
  18875=>"010011100",
  18876=>"110101010",
  18877=>"011010101",
  18878=>"000001011",
  18879=>"011001000",
  18880=>"011110001",
  18881=>"000011000",
  18882=>"000000001",
  18883=>"111000101",
  18884=>"010011101",
  18885=>"011111110",
  18886=>"100000110",
  18887=>"111111000",
  18888=>"100000100",
  18889=>"101100001",
  18890=>"001000000",
  18891=>"100001000",
  18892=>"100101110",
  18893=>"000010111",
  18894=>"011011010",
  18895=>"000001101",
  18896=>"101000101",
  18897=>"001101000",
  18898=>"010010000",
  18899=>"101100101",
  18900=>"100110110",
  18901=>"101010101",
  18902=>"001100100",
  18903=>"110111111",
  18904=>"100010100",
  18905=>"010101110",
  18906=>"000000101",
  18907=>"010100110",
  18908=>"010001100",
  18909=>"011100101",
  18910=>"101101100",
  18911=>"000001000",
  18912=>"000110010",
  18913=>"101011010",
  18914=>"100101111",
  18915=>"110101110",
  18916=>"101011111",
  18917=>"000110011",
  18918=>"110000101",
  18919=>"101100000",
  18920=>"010000111",
  18921=>"111100111",
  18922=>"011100000",
  18923=>"111100101",
  18924=>"000000111",
  18925=>"101011001",
  18926=>"011101111",
  18927=>"110010110",
  18928=>"011001110",
  18929=>"000000100",
  18930=>"001001001",
  18931=>"111110111",
  18932=>"000011011",
  18933=>"010011010",
  18934=>"101110011",
  18935=>"000011101",
  18936=>"000000001",
  18937=>"101000011",
  18938=>"010001110",
  18939=>"000100000",
  18940=>"000001011",
  18941=>"010000101",
  18942=>"010110111",
  18943=>"010011111",
  18944=>"110011101",
  18945=>"110011111",
  18946=>"001000010",
  18947=>"111001101",
  18948=>"101100111",
  18949=>"101010111",
  18950=>"010110100",
  18951=>"001110110",
  18952=>"001000001",
  18953=>"100100000",
  18954=>"010101100",
  18955=>"010101111",
  18956=>"001011000",
  18957=>"000000111",
  18958=>"011111111",
  18959=>"010101001",
  18960=>"010111001",
  18961=>"110000100",
  18962=>"000000100",
  18963=>"010110111",
  18964=>"110010101",
  18965=>"011011100",
  18966=>"010111011",
  18967=>"010001111",
  18968=>"111010110",
  18969=>"100100110",
  18970=>"101001111",
  18971=>"101011011",
  18972=>"011110000",
  18973=>"000000111",
  18974=>"110111110",
  18975=>"110001000",
  18976=>"001101111",
  18977=>"111010000",
  18978=>"101000011",
  18979=>"011100010",
  18980=>"001010100",
  18981=>"111111110",
  18982=>"001001010",
  18983=>"001100000",
  18984=>"110100101",
  18985=>"001011000",
  18986=>"010100000",
  18987=>"011000101",
  18988=>"110101111",
  18989=>"001100111",
  18990=>"010001110",
  18991=>"010010010",
  18992=>"001101100",
  18993=>"011101100",
  18994=>"000011110",
  18995=>"111110111",
  18996=>"100110100",
  18997=>"111010011",
  18998=>"101011011",
  18999=>"010111110",
  19000=>"100100101",
  19001=>"111110010",
  19002=>"100001100",
  19003=>"011000100",
  19004=>"111111101",
  19005=>"101101110",
  19006=>"001000010",
  19007=>"010110011",
  19008=>"100110111",
  19009=>"011111111",
  19010=>"001000111",
  19011=>"000110101",
  19012=>"000110011",
  19013=>"111111100",
  19014=>"010010111",
  19015=>"111100111",
  19016=>"100111010",
  19017=>"100000000",
  19018=>"001001011",
  19019=>"000101101",
  19020=>"001101111",
  19021=>"110001101",
  19022=>"011100010",
  19023=>"010001010",
  19024=>"001010111",
  19025=>"001110010",
  19026=>"100001111",
  19027=>"010100001",
  19028=>"100001100",
  19029=>"011000100",
  19030=>"001011110",
  19031=>"001111011",
  19032=>"111001010",
  19033=>"001101011",
  19034=>"010011000",
  19035=>"110111100",
  19036=>"000001010",
  19037=>"100000101",
  19038=>"000000111",
  19039=>"101110000",
  19040=>"100110100",
  19041=>"100100111",
  19042=>"000010101",
  19043=>"101000010",
  19044=>"010001111",
  19045=>"110111101",
  19046=>"100101100",
  19047=>"110101001",
  19048=>"101000111",
  19049=>"001011001",
  19050=>"010000000",
  19051=>"111111101",
  19052=>"000000100",
  19053=>"101000110",
  19054=>"110111111",
  19055=>"000110111",
  19056=>"001000111",
  19057=>"000000111",
  19058=>"100001100",
  19059=>"111100100",
  19060=>"101001111",
  19061=>"101100011",
  19062=>"111011101",
  19063=>"010000011",
  19064=>"000000000",
  19065=>"010011010",
  19066=>"110110001",
  19067=>"000001110",
  19068=>"010110001",
  19069=>"101000010",
  19070=>"110000111",
  19071=>"010011111",
  19072=>"111111010",
  19073=>"101001100",
  19074=>"111011100",
  19075=>"010111100",
  19076=>"001110100",
  19077=>"101101100",
  19078=>"001100100",
  19079=>"111111111",
  19080=>"111001111",
  19081=>"000011010",
  19082=>"001101111",
  19083=>"001100000",
  19084=>"100111010",
  19085=>"101110010",
  19086=>"110101111",
  19087=>"100111000",
  19088=>"101100100",
  19089=>"001001011",
  19090=>"100111011",
  19091=>"110001001",
  19092=>"010110101",
  19093=>"000101000",
  19094=>"100001000",
  19095=>"010000010",
  19096=>"100001010",
  19097=>"010110100",
  19098=>"110111001",
  19099=>"011001110",
  19100=>"000101001",
  19101=>"101011011",
  19102=>"111110101",
  19103=>"011001011",
  19104=>"000000011",
  19105=>"000000111",
  19106=>"110011101",
  19107=>"011000101",
  19108=>"111111000",
  19109=>"000001000",
  19110=>"000010100",
  19111=>"000101101",
  19112=>"000110110",
  19113=>"101100111",
  19114=>"100101000",
  19115=>"011101101",
  19116=>"011100000",
  19117=>"111111110",
  19118=>"100101000",
  19119=>"001000100",
  19120=>"111000101",
  19121=>"100001100",
  19122=>"110100001",
  19123=>"100001111",
  19124=>"000100001",
  19125=>"001010100",
  19126=>"011001001",
  19127=>"000001110",
  19128=>"001101110",
  19129=>"011110000",
  19130=>"001010110",
  19131=>"000010111",
  19132=>"000100011",
  19133=>"001000001",
  19134=>"000010110",
  19135=>"011010111",
  19136=>"111111111",
  19137=>"001100010",
  19138=>"001110110",
  19139=>"101000001",
  19140=>"111001010",
  19141=>"101100101",
  19142=>"010111000",
  19143=>"000000010",
  19144=>"100111111",
  19145=>"011111110",
  19146=>"111111011",
  19147=>"000011011",
  19148=>"010010011",
  19149=>"100010011",
  19150=>"011101001",
  19151=>"001001111",
  19152=>"101101101",
  19153=>"010010011",
  19154=>"001111110",
  19155=>"000010000",
  19156=>"000000111",
  19157=>"011111010",
  19158=>"010000100",
  19159=>"111101010",
  19160=>"000001001",
  19161=>"001101011",
  19162=>"100110110",
  19163=>"001110110",
  19164=>"001011000",
  19165=>"110100100",
  19166=>"111111101",
  19167=>"110001110",
  19168=>"010101010",
  19169=>"010001100",
  19170=>"110100011",
  19171=>"000100000",
  19172=>"001011111",
  19173=>"010100001",
  19174=>"000111011",
  19175=>"010000001",
  19176=>"000101110",
  19177=>"001111001",
  19178=>"101101111",
  19179=>"111001110",
  19180=>"010010011",
  19181=>"110110001",
  19182=>"100000001",
  19183=>"000010111",
  19184=>"111110101",
  19185=>"110001111",
  19186=>"010011100",
  19187=>"000001000",
  19188=>"011001101",
  19189=>"011100001",
  19190=>"111101111",
  19191=>"001011010",
  19192=>"100110111",
  19193=>"011011100",
  19194=>"110000011",
  19195=>"100001110",
  19196=>"111011010",
  19197=>"110000000",
  19198=>"010110011",
  19199=>"100011101",
  19200=>"000000100",
  19201=>"011111100",
  19202=>"010000000",
  19203=>"001100001",
  19204=>"010111101",
  19205=>"100011110",
  19206=>"101100001",
  19207=>"111001111",
  19208=>"110001100",
  19209=>"111111110",
  19210=>"101110000",
  19211=>"011101011",
  19212=>"110111110",
  19213=>"110010100",
  19214=>"110110110",
  19215=>"000010010",
  19216=>"110110110",
  19217=>"001000110",
  19218=>"110010100",
  19219=>"101001110",
  19220=>"011010100",
  19221=>"110111101",
  19222=>"001010000",
  19223=>"110011100",
  19224=>"011011010",
  19225=>"101101011",
  19226=>"011111001",
  19227=>"001000111",
  19228=>"100001110",
  19229=>"011101100",
  19230=>"011100101",
  19231=>"001111010",
  19232=>"101001001",
  19233=>"110101100",
  19234=>"110010010",
  19235=>"111110101",
  19236=>"000100100",
  19237=>"110100001",
  19238=>"101111011",
  19239=>"101010111",
  19240=>"000100011",
  19241=>"101011001",
  19242=>"111000001",
  19243=>"010101001",
  19244=>"001011110",
  19245=>"010000011",
  19246=>"001000101",
  19247=>"000011011",
  19248=>"101101110",
  19249=>"110100011",
  19250=>"101100000",
  19251=>"011111101",
  19252=>"011010000",
  19253=>"110000000",
  19254=>"110011011",
  19255=>"000001110",
  19256=>"110110101",
  19257=>"001110110",
  19258=>"001010000",
  19259=>"111011100",
  19260=>"010010010",
  19261=>"100011101",
  19262=>"001000100",
  19263=>"001010000",
  19264=>"110100010",
  19265=>"110011110",
  19266=>"111101001",
  19267=>"110011010",
  19268=>"011110011",
  19269=>"011000110",
  19270=>"001010010",
  19271=>"011000000",
  19272=>"111011001",
  19273=>"001011001",
  19274=>"100110000",
  19275=>"110000110",
  19276=>"100000010",
  19277=>"000011100",
  19278=>"001001101",
  19279=>"111011100",
  19280=>"000010110",
  19281=>"100011011",
  19282=>"011001010",
  19283=>"000011010",
  19284=>"010010000",
  19285=>"101100011",
  19286=>"000001101",
  19287=>"100000000",
  19288=>"000000011",
  19289=>"111110110",
  19290=>"001001100",
  19291=>"000011101",
  19292=>"001100110",
  19293=>"000011010",
  19294=>"100010011",
  19295=>"100100111",
  19296=>"100111011",
  19297=>"001010001",
  19298=>"101100110",
  19299=>"001110111",
  19300=>"010111101",
  19301=>"111001000",
  19302=>"111101001",
  19303=>"010000110",
  19304=>"010001010",
  19305=>"001110101",
  19306=>"111001101",
  19307=>"111100001",
  19308=>"000111010",
  19309=>"000110000",
  19310=>"010010011",
  19311=>"110010100",
  19312=>"100111010",
  19313=>"111101000",
  19314=>"101100100",
  19315=>"000001110",
  19316=>"111101000",
  19317=>"000101101",
  19318=>"100001101",
  19319=>"011100000",
  19320=>"011000111",
  19321=>"101101001",
  19322=>"110100110",
  19323=>"001110001",
  19324=>"000110110",
  19325=>"011010000",
  19326=>"100010100",
  19327=>"110011110",
  19328=>"110001110",
  19329=>"001010100",
  19330=>"010000100",
  19331=>"011110111",
  19332=>"010110100",
  19333=>"000000010",
  19334=>"111111000",
  19335=>"110001101",
  19336=>"110111100",
  19337=>"111011010",
  19338=>"010010001",
  19339=>"000011011",
  19340=>"111110101",
  19341=>"001101011",
  19342=>"100100110",
  19343=>"111001000",
  19344=>"000111101",
  19345=>"011011001",
  19346=>"010001010",
  19347=>"001010100",
  19348=>"101111010",
  19349=>"010100111",
  19350=>"101111101",
  19351=>"000010001",
  19352=>"111110001",
  19353=>"000110110",
  19354=>"000111010",
  19355=>"001010110",
  19356=>"011101011",
  19357=>"100110001",
  19358=>"101011001",
  19359=>"001010101",
  19360=>"100111110",
  19361=>"000100111",
  19362=>"110101000",
  19363=>"011001111",
  19364=>"001100000",
  19365=>"001000111",
  19366=>"011101011",
  19367=>"100010001",
  19368=>"010100111",
  19369=>"000000010",
  19370=>"111011101",
  19371=>"110000010",
  19372=>"101011010",
  19373=>"100110110",
  19374=>"010000111",
  19375=>"010010000",
  19376=>"000100111",
  19377=>"001011111",
  19378=>"000100011",
  19379=>"101010010",
  19380=>"010010111",
  19381=>"010110101",
  19382=>"110101001",
  19383=>"000101101",
  19384=>"101110100",
  19385=>"110011100",
  19386=>"110101111",
  19387=>"100101010",
  19388=>"100110010",
  19389=>"011010110",
  19390=>"000101110",
  19391=>"100111010",
  19392=>"110001111",
  19393=>"100010100",
  19394=>"000010000",
  19395=>"011001011",
  19396=>"100101011",
  19397=>"001101111",
  19398=>"011000011",
  19399=>"101110010",
  19400=>"101001101",
  19401=>"100111010",
  19402=>"011010101",
  19403=>"111011010",
  19404=>"011111100",
  19405=>"100000001",
  19406=>"111010101",
  19407=>"111011100",
  19408=>"011010001",
  19409=>"111001111",
  19410=>"010101100",
  19411=>"100111111",
  19412=>"001011010",
  19413=>"101101101",
  19414=>"000000001",
  19415=>"000111100",
  19416=>"100101110",
  19417=>"011000011",
  19418=>"011100000",
  19419=>"000000001",
  19420=>"001011011",
  19421=>"100010000",
  19422=>"110100010",
  19423=>"101101011",
  19424=>"100010100",
  19425=>"000011010",
  19426=>"100100111",
  19427=>"100001111",
  19428=>"101001001",
  19429=>"011110110",
  19430=>"100111101",
  19431=>"111010010",
  19432=>"010100111",
  19433=>"100010000",
  19434=>"010001100",
  19435=>"101001101",
  19436=>"100010100",
  19437=>"111111010",
  19438=>"110000011",
  19439=>"101111101",
  19440=>"010101101",
  19441=>"001000001",
  19442=>"111001111",
  19443=>"111101110",
  19444=>"000011111",
  19445=>"000011111",
  19446=>"011011101",
  19447=>"101110111",
  19448=>"000000110",
  19449=>"000110111",
  19450=>"010000111",
  19451=>"010101010",
  19452=>"101000001",
  19453=>"011100001",
  19454=>"000000101",
  19455=>"100001001",
  19456=>"000001100",
  19457=>"101111000",
  19458=>"100111101",
  19459=>"001111110",
  19460=>"001101010",
  19461=>"001011000",
  19462=>"001101010",
  19463=>"001010000",
  19464=>"010110000",
  19465=>"000110001",
  19466=>"001100110",
  19467=>"110010001",
  19468=>"111111010",
  19469=>"100110110",
  19470=>"100101011",
  19471=>"000010011",
  19472=>"001010001",
  19473=>"011111110",
  19474=>"101111001",
  19475=>"001101110",
  19476=>"111111000",
  19477=>"100100011",
  19478=>"111010111",
  19479=>"010101000",
  19480=>"001110110",
  19481=>"101011110",
  19482=>"010000111",
  19483=>"101100111",
  19484=>"101100101",
  19485=>"011011001",
  19486=>"000011110",
  19487=>"000001111",
  19488=>"100011000",
  19489=>"111011110",
  19490=>"010010110",
  19491=>"010001110",
  19492=>"101010100",
  19493=>"111001011",
  19494=>"010100100",
  19495=>"111111011",
  19496=>"111101000",
  19497=>"001111011",
  19498=>"001101000",
  19499=>"000001101",
  19500=>"110101110",
  19501=>"001111111",
  19502=>"001100101",
  19503=>"001001010",
  19504=>"111011011",
  19505=>"100010011",
  19506=>"010001001",
  19507=>"011010111",
  19508=>"010101110",
  19509=>"011101100",
  19510=>"011000111",
  19511=>"001110001",
  19512=>"001000010",
  19513=>"110001010",
  19514=>"111101100",
  19515=>"011111001",
  19516=>"010010010",
  19517=>"001010101",
  19518=>"000001001",
  19519=>"001110010",
  19520=>"010110000",
  19521=>"000011001",
  19522=>"011100011",
  19523=>"011001011",
  19524=>"101110111",
  19525=>"001001011",
  19526=>"000000100",
  19527=>"010110001",
  19528=>"001010010",
  19529=>"110001100",
  19530=>"011101000",
  19531=>"001011001",
  19532=>"000000000",
  19533=>"010000011",
  19534=>"100101111",
  19535=>"111100010",
  19536=>"100101011",
  19537=>"011101000",
  19538=>"010000000",
  19539=>"011101100",
  19540=>"100011010",
  19541=>"101011010",
  19542=>"000100000",
  19543=>"100111101",
  19544=>"000001000",
  19545=>"110110001",
  19546=>"010000110",
  19547=>"100001111",
  19548=>"011110000",
  19549=>"101000101",
  19550=>"111001011",
  19551=>"101001100",
  19552=>"001000111",
  19553=>"001001000",
  19554=>"111100101",
  19555=>"011010000",
  19556=>"011111000",
  19557=>"010101000",
  19558=>"010010101",
  19559=>"001010011",
  19560=>"001010001",
  19561=>"010101001",
  19562=>"010111101",
  19563=>"000100100",
  19564=>"110100100",
  19565=>"101010111",
  19566=>"001010010",
  19567=>"101101011",
  19568=>"001111111",
  19569=>"111111100",
  19570=>"110000110",
  19571=>"011010000",
  19572=>"000010001",
  19573=>"000110110",
  19574=>"010011001",
  19575=>"000000110",
  19576=>"001101001",
  19577=>"010110000",
  19578=>"100010001",
  19579=>"100100001",
  19580=>"001101001",
  19581=>"001101110",
  19582=>"010001011",
  19583=>"100100001",
  19584=>"000111101",
  19585=>"001011111",
  19586=>"101101110",
  19587=>"100011000",
  19588=>"101100000",
  19589=>"101011100",
  19590=>"110001010",
  19591=>"101001000",
  19592=>"000111001",
  19593=>"001001000",
  19594=>"100001001",
  19595=>"111010110",
  19596=>"010010100",
  19597=>"101101110",
  19598=>"011011010",
  19599=>"001011110",
  19600=>"011110011",
  19601=>"000011000",
  19602=>"100011111",
  19603=>"010110001",
  19604=>"000110010",
  19605=>"100001000",
  19606=>"100011010",
  19607=>"101010011",
  19608=>"111000010",
  19609=>"111100111",
  19610=>"111011010",
  19611=>"001000001",
  19612=>"000001100",
  19613=>"100100000",
  19614=>"100111101",
  19615=>"111101100",
  19616=>"101010010",
  19617=>"011100000",
  19618=>"000001000",
  19619=>"101110010",
  19620=>"101111101",
  19621=>"100111000",
  19622=>"001011101",
  19623=>"011001010",
  19624=>"001010000",
  19625=>"010111000",
  19626=>"010110010",
  19627=>"000000000",
  19628=>"011010110",
  19629=>"010001111",
  19630=>"000100111",
  19631=>"110101001",
  19632=>"000000010",
  19633=>"000000101",
  19634=>"000000011",
  19635=>"000010101",
  19636=>"100011010",
  19637=>"111011100",
  19638=>"001100010",
  19639=>"011111010",
  19640=>"110111010",
  19641=>"111101100",
  19642=>"000000100",
  19643=>"010001100",
  19644=>"011101000",
  19645=>"000001000",
  19646=>"010001110",
  19647=>"111100111",
  19648=>"000001110",
  19649=>"101011111",
  19650=>"011100000",
  19651=>"100110001",
  19652=>"100111100",
  19653=>"010011111",
  19654=>"000111011",
  19655=>"011010111",
  19656=>"110111101",
  19657=>"110100110",
  19658=>"011110111",
  19659=>"111100111",
  19660=>"111110101",
  19661=>"011011010",
  19662=>"111110001",
  19663=>"100011000",
  19664=>"100100010",
  19665=>"111111011",
  19666=>"111000001",
  19667=>"000111001",
  19668=>"011001000",
  19669=>"111001000",
  19670=>"111011101",
  19671=>"000001110",
  19672=>"100111000",
  19673=>"011110001",
  19674=>"110001000",
  19675=>"001100111",
  19676=>"101110001",
  19677=>"100000110",
  19678=>"001010000",
  19679=>"110100110",
  19680=>"110110111",
  19681=>"100000110",
  19682=>"000111100",
  19683=>"001001000",
  19684=>"111010111",
  19685=>"001010111",
  19686=>"001010001",
  19687=>"010011011",
  19688=>"100101011",
  19689=>"011100110",
  19690=>"100111110",
  19691=>"100111101",
  19692=>"111110010",
  19693=>"000001100",
  19694=>"100110101",
  19695=>"010011001",
  19696=>"011000111",
  19697=>"100101111",
  19698=>"110100101",
  19699=>"110100000",
  19700=>"011010010",
  19701=>"000000100",
  19702=>"101110000",
  19703=>"000010010",
  19704=>"111101000",
  19705=>"010010001",
  19706=>"000100011",
  19707=>"010010110",
  19708=>"111111001",
  19709=>"000000001",
  19710=>"100110011",
  19711=>"010110011",
  19712=>"110100100",
  19713=>"010101010",
  19714=>"100110001",
  19715=>"011001011",
  19716=>"100101001",
  19717=>"101001010",
  19718=>"101011011",
  19719=>"100101101",
  19720=>"000001001",
  19721=>"001110101",
  19722=>"100101111",
  19723=>"000000010",
  19724=>"001000010",
  19725=>"010111100",
  19726=>"100111000",
  19727=>"101000001",
  19728=>"101100010",
  19729=>"111111001",
  19730=>"110110100",
  19731=>"000111010",
  19732=>"110100001",
  19733=>"101101100",
  19734=>"100001111",
  19735=>"010111111",
  19736=>"000111101",
  19737=>"110110011",
  19738=>"000110001",
  19739=>"000001000",
  19740=>"011011000",
  19741=>"101110101",
  19742=>"110110101",
  19743=>"001001100",
  19744=>"010001011",
  19745=>"001010000",
  19746=>"100011000",
  19747=>"100011111",
  19748=>"000100110",
  19749=>"101000011",
  19750=>"001101100",
  19751=>"110000011",
  19752=>"111101000",
  19753=>"011000110",
  19754=>"111001001",
  19755=>"000011100",
  19756=>"101101111",
  19757=>"011100000",
  19758=>"110001000",
  19759=>"100100001",
  19760=>"100101010",
  19761=>"000011111",
  19762=>"000001011",
  19763=>"101001110",
  19764=>"101001111",
  19765=>"000001101",
  19766=>"011001100",
  19767=>"111101110",
  19768=>"000011001",
  19769=>"011000100",
  19770=>"100100100",
  19771=>"110101000",
  19772=>"010010101",
  19773=>"001010110",
  19774=>"011101001",
  19775=>"000111001",
  19776=>"000100110",
  19777=>"111010111",
  19778=>"011100000",
  19779=>"000110111",
  19780=>"000011100",
  19781=>"010111110",
  19782=>"101100111",
  19783=>"010110100",
  19784=>"110100111",
  19785=>"101001111",
  19786=>"111101011",
  19787=>"001111001",
  19788=>"001000001",
  19789=>"110110110",
  19790=>"010001101",
  19791=>"100111011",
  19792=>"010010011",
  19793=>"100110001",
  19794=>"111011101",
  19795=>"001010010",
  19796=>"001000000",
  19797=>"000010011",
  19798=>"001010000",
  19799=>"110011111",
  19800=>"001011010",
  19801=>"010101111",
  19802=>"110101000",
  19803=>"110110011",
  19804=>"100000000",
  19805=>"101111110",
  19806=>"011100000",
  19807=>"111000100",
  19808=>"111001101",
  19809=>"011101010",
  19810=>"100111111",
  19811=>"111001010",
  19812=>"010100010",
  19813=>"000010001",
  19814=>"011110110",
  19815=>"011010110",
  19816=>"100010010",
  19817=>"000000001",
  19818=>"111111101",
  19819=>"111111010",
  19820=>"000011000",
  19821=>"110101001",
  19822=>"011111100",
  19823=>"010110011",
  19824=>"100111010",
  19825=>"000100100",
  19826=>"010010110",
  19827=>"011010100",
  19828=>"111111000",
  19829=>"101001101",
  19830=>"011000010",
  19831=>"000100111",
  19832=>"010110001",
  19833=>"111111100",
  19834=>"100101001",
  19835=>"011000111",
  19836=>"110010010",
  19837=>"110110111",
  19838=>"001010001",
  19839=>"110111001",
  19840=>"000010000",
  19841=>"011000100",
  19842=>"010110111",
  19843=>"111110111",
  19844=>"101011011",
  19845=>"000111101",
  19846=>"000100011",
  19847=>"111011000",
  19848=>"101110001",
  19849=>"100100100",
  19850=>"100101100",
  19851=>"111110110",
  19852=>"111111100",
  19853=>"000101101",
  19854=>"100000110",
  19855=>"011000100",
  19856=>"110101111",
  19857=>"111101111",
  19858=>"111110111",
  19859=>"011011101",
  19860=>"000010001",
  19861=>"110111010",
  19862=>"000010111",
  19863=>"110111000",
  19864=>"101011100",
  19865=>"111001001",
  19866=>"101100011",
  19867=>"111000100",
  19868=>"001110110",
  19869=>"101110111",
  19870=>"010001011",
  19871=>"010000111",
  19872=>"000101101",
  19873=>"110011000",
  19874=>"001110010",
  19875=>"010010001",
  19876=>"011110000",
  19877=>"110110111",
  19878=>"011111100",
  19879=>"011111111",
  19880=>"111010010",
  19881=>"110111001",
  19882=>"011101101",
  19883=>"010110110",
  19884=>"001011000",
  19885=>"000010101",
  19886=>"011101011",
  19887=>"111011010",
  19888=>"000101010",
  19889=>"000110111",
  19890=>"100001100",
  19891=>"000111100",
  19892=>"101110011",
  19893=>"001111000",
  19894=>"010100111",
  19895=>"110100010",
  19896=>"101000000",
  19897=>"010000000",
  19898=>"001010111",
  19899=>"010001010",
  19900=>"010010101",
  19901=>"101011111",
  19902=>"010110010",
  19903=>"110100010",
  19904=>"000000100",
  19905=>"101000101",
  19906=>"111000000",
  19907=>"100010000",
  19908=>"101111100",
  19909=>"001010111",
  19910=>"101100100",
  19911=>"000000010",
  19912=>"100100010",
  19913=>"110000111",
  19914=>"111110010",
  19915=>"010001000",
  19916=>"111100000",
  19917=>"010110001",
  19918=>"010111100",
  19919=>"011100000",
  19920=>"100000001",
  19921=>"010000101",
  19922=>"110101101",
  19923=>"111001000",
  19924=>"111000111",
  19925=>"101101001",
  19926=>"110111101",
  19927=>"010100001",
  19928=>"111110010",
  19929=>"001000011",
  19930=>"100110011",
  19931=>"101001111",
  19932=>"001001000",
  19933=>"011000100",
  19934=>"000110101",
  19935=>"100001010",
  19936=>"111000011",
  19937=>"111010000",
  19938=>"100000111",
  19939=>"000100111",
  19940=>"100110101",
  19941=>"100101010",
  19942=>"101011110",
  19943=>"100001010",
  19944=>"101001100",
  19945=>"111101101",
  19946=>"110101011",
  19947=>"101011000",
  19948=>"110110000",
  19949=>"111000000",
  19950=>"011100011",
  19951=>"011111010",
  19952=>"000010110",
  19953=>"101100101",
  19954=>"101111100",
  19955=>"000101110",
  19956=>"101010110",
  19957=>"000101010",
  19958=>"110001000",
  19959=>"101101111",
  19960=>"110111000",
  19961=>"110011111",
  19962=>"001010111",
  19963=>"110000101",
  19964=>"110101001",
  19965=>"110100000",
  19966=>"100101010",
  19967=>"011100000",
  19968=>"101011101",
  19969=>"000000111",
  19970=>"010001110",
  19971=>"100000010",
  19972=>"101001111",
  19973=>"001111001",
  19974=>"101101011",
  19975=>"110110011",
  19976=>"110111011",
  19977=>"111010110",
  19978=>"111000101",
  19979=>"111000110",
  19980=>"110001011",
  19981=>"111111011",
  19982=>"001000111",
  19983=>"000000001",
  19984=>"111011100",
  19985=>"000011101",
  19986=>"010111001",
  19987=>"011100000",
  19988=>"000101101",
  19989=>"001011011",
  19990=>"011100101",
  19991=>"011000111",
  19992=>"001000000",
  19993=>"111001100",
  19994=>"010000100",
  19995=>"101010001",
  19996=>"101011010",
  19997=>"110000000",
  19998=>"001001011",
  19999=>"101011011",
  20000=>"011010011",
  20001=>"100111110",
  20002=>"001000101",
  20003=>"111001101",
  20004=>"001011110",
  20005=>"110101001",
  20006=>"001001001",
  20007=>"000110100",
  20008=>"011101111",
  20009=>"000111111",
  20010=>"001000001",
  20011=>"011001111",
  20012=>"010111110",
  20013=>"001110110",
  20014=>"110100110",
  20015=>"001110100",
  20016=>"101010110",
  20017=>"111001110",
  20018=>"100100000",
  20019=>"111010011",
  20020=>"001001010",
  20021=>"000100101",
  20022=>"000101000",
  20023=>"000101000",
  20024=>"011000010",
  20025=>"111100101",
  20026=>"110001011",
  20027=>"111011101",
  20028=>"101000101",
  20029=>"100011110",
  20030=>"110100000",
  20031=>"100110000",
  20032=>"111011000",
  20033=>"111101010",
  20034=>"010000110",
  20035=>"100010001",
  20036=>"110001100",
  20037=>"100111000",
  20038=>"000101010",
  20039=>"111111101",
  20040=>"010011000",
  20041=>"111000110",
  20042=>"000110001",
  20043=>"111101001",
  20044=>"001000000",
  20045=>"000100111",
  20046=>"100111101",
  20047=>"111100100",
  20048=>"011111100",
  20049=>"011001011",
  20050=>"000011100",
  20051=>"100100111",
  20052=>"010011000",
  20053=>"000111011",
  20054=>"101101000",
  20055=>"011001000",
  20056=>"011100101",
  20057=>"100101100",
  20058=>"000100110",
  20059=>"001111001",
  20060=>"000100000",
  20061=>"001010010",
  20062=>"001100101",
  20063=>"101001100",
  20064=>"111010111",
  20065=>"100001010",
  20066=>"000111000",
  20067=>"010011000",
  20068=>"011011100",
  20069=>"111010111",
  20070=>"000111101",
  20071=>"001111101",
  20072=>"110011001",
  20073=>"010000011",
  20074=>"011101101",
  20075=>"100001000",
  20076=>"111001101",
  20077=>"101001001",
  20078=>"111010000",
  20079=>"111001101",
  20080=>"001010100",
  20081=>"000100101",
  20082=>"010001010",
  20083=>"110000000",
  20084=>"010101111",
  20085=>"011010001",
  20086=>"001011001",
  20087=>"110011101",
  20088=>"001011111",
  20089=>"101011011",
  20090=>"000111101",
  20091=>"111110101",
  20092=>"011010101",
  20093=>"100100100",
  20094=>"000101111",
  20095=>"011000100",
  20096=>"000111001",
  20097=>"000111001",
  20098=>"101110000",
  20099=>"111011000",
  20100=>"111111010",
  20101=>"011000101",
  20102=>"110011110",
  20103=>"101110110",
  20104=>"111100100",
  20105=>"100010011",
  20106=>"100011010",
  20107=>"110100001",
  20108=>"111111011",
  20109=>"000001101",
  20110=>"011100000",
  20111=>"001000011",
  20112=>"011111111",
  20113=>"101111111",
  20114=>"111010100",
  20115=>"010010100",
  20116=>"000000100",
  20117=>"111100110",
  20118=>"111001000",
  20119=>"110010011",
  20120=>"111110011",
  20121=>"100000000",
  20122=>"110000011",
  20123=>"111001010",
  20124=>"010010110",
  20125=>"111010110",
  20126=>"101110101",
  20127=>"110100110",
  20128=>"001101000",
  20129=>"101111111",
  20130=>"001000000",
  20131=>"110111101",
  20132=>"110010010",
  20133=>"111001100",
  20134=>"010111101",
  20135=>"000100000",
  20136=>"100010000",
  20137=>"000100111",
  20138=>"111001001",
  20139=>"100110100",
  20140=>"000001011",
  20141=>"111101011",
  20142=>"101000101",
  20143=>"000100001",
  20144=>"111110001",
  20145=>"111100110",
  20146=>"101010000",
  20147=>"100000011",
  20148=>"100001010",
  20149=>"001000001",
  20150=>"100001111",
  20151=>"110101111",
  20152=>"000101011",
  20153=>"100110110",
  20154=>"010010010",
  20155=>"100110010",
  20156=>"100110010",
  20157=>"000110011",
  20158=>"000001001",
  20159=>"100000000",
  20160=>"011011101",
  20161=>"100101110",
  20162=>"000100001",
  20163=>"111110101",
  20164=>"000100001",
  20165=>"001110111",
  20166=>"011101101",
  20167=>"100110100",
  20168=>"010000000",
  20169=>"001111100",
  20170=>"011101010",
  20171=>"000010000",
  20172=>"001010001",
  20173=>"110010101",
  20174=>"001010100",
  20175=>"000101100",
  20176=>"000000101",
  20177=>"100000010",
  20178=>"010010000",
  20179=>"011000101",
  20180=>"010010101",
  20181=>"000000111",
  20182=>"110111010",
  20183=>"110000010",
  20184=>"000001100",
  20185=>"100101110",
  20186=>"000111100",
  20187=>"011001110",
  20188=>"101000111",
  20189=>"000101101",
  20190=>"101100101",
  20191=>"001011001",
  20192=>"110001101",
  20193=>"110010010",
  20194=>"101110001",
  20195=>"110000000",
  20196=>"000101010",
  20197=>"011010101",
  20198=>"000001010",
  20199=>"101110100",
  20200=>"100000101",
  20201=>"000011000",
  20202=>"001000101",
  20203=>"101000011",
  20204=>"100000110",
  20205=>"100001000",
  20206=>"010011000",
  20207=>"011010001",
  20208=>"101001001",
  20209=>"101111111",
  20210=>"001001110",
  20211=>"000100001",
  20212=>"010100000",
  20213=>"010100101",
  20214=>"101001101",
  20215=>"011111110",
  20216=>"000100100",
  20217=>"011011110",
  20218=>"000000100",
  20219=>"111001010",
  20220=>"110100001",
  20221=>"010000101",
  20222=>"001001101",
  20223=>"101111011",
  20224=>"110010100",
  20225=>"010001101",
  20226=>"001000000",
  20227=>"101100000",
  20228=>"011001101",
  20229=>"010000110",
  20230=>"001011010",
  20231=>"110010001",
  20232=>"101111110",
  20233=>"001010000",
  20234=>"101001111",
  20235=>"001100011",
  20236=>"000010001",
  20237=>"110111111",
  20238=>"010100101",
  20239=>"111000110",
  20240=>"000011000",
  20241=>"100001000",
  20242=>"110110110",
  20243=>"010010111",
  20244=>"100010010",
  20245=>"000011100",
  20246=>"110101111",
  20247=>"011111110",
  20248=>"100100000",
  20249=>"000001100",
  20250=>"101110111",
  20251=>"010101011",
  20252=>"000011010",
  20253=>"110011100",
  20254=>"000011101",
  20255=>"011001101",
  20256=>"001100111",
  20257=>"101111110",
  20258=>"011000000",
  20259=>"001110001",
  20260=>"011000101",
  20261=>"101011101",
  20262=>"010110011",
  20263=>"011001100",
  20264=>"100101100",
  20265=>"110010001",
  20266=>"100100110",
  20267=>"101110010",
  20268=>"100101011",
  20269=>"110000000",
  20270=>"010101101",
  20271=>"110110110",
  20272=>"111100101",
  20273=>"011001110",
  20274=>"000101110",
  20275=>"010010010",
  20276=>"111100110",
  20277=>"011000010",
  20278=>"110100100",
  20279=>"111010001",
  20280=>"110110100",
  20281=>"100000010",
  20282=>"101000100",
  20283=>"110100000",
  20284=>"010101011",
  20285=>"101000001",
  20286=>"101001110",
  20287=>"010000001",
  20288=>"010101100",
  20289=>"010100110",
  20290=>"111111011",
  20291=>"001100001",
  20292=>"000001010",
  20293=>"101010011",
  20294=>"111100011",
  20295=>"101101001",
  20296=>"111000100",
  20297=>"001101011",
  20298=>"001111110",
  20299=>"100101000",
  20300=>"000011010",
  20301=>"101011111",
  20302=>"100111010",
  20303=>"010001100",
  20304=>"110111010",
  20305=>"011101001",
  20306=>"100100010",
  20307=>"011001010",
  20308=>"000011100",
  20309=>"100101000",
  20310=>"110101110",
  20311=>"010111100",
  20312=>"010010110",
  20313=>"110000011",
  20314=>"000110101",
  20315=>"101101111",
  20316=>"110001101",
  20317=>"111001111",
  20318=>"100110000",
  20319=>"010101000",
  20320=>"001011001",
  20321=>"110110110",
  20322=>"101000111",
  20323=>"001110101",
  20324=>"001101110",
  20325=>"110000111",
  20326=>"101001001",
  20327=>"010011001",
  20328=>"111110101",
  20329=>"010000111",
  20330=>"111011100",
  20331=>"101111011",
  20332=>"000110111",
  20333=>"100000010",
  20334=>"000000011",
  20335=>"110001101",
  20336=>"000100110",
  20337=>"101100010",
  20338=>"010010001",
  20339=>"011111011",
  20340=>"000001001",
  20341=>"000101011",
  20342=>"001100010",
  20343=>"001000000",
  20344=>"000111111",
  20345=>"110000110",
  20346=>"000010001",
  20347=>"111011100",
  20348=>"001010110",
  20349=>"110011001",
  20350=>"110011111",
  20351=>"110111100",
  20352=>"000011101",
  20353=>"111100011",
  20354=>"111000100",
  20355=>"001001111",
  20356=>"111110001",
  20357=>"000010000",
  20358=>"011101101",
  20359=>"001011100",
  20360=>"000111101",
  20361=>"000001011",
  20362=>"110100000",
  20363=>"000001100",
  20364=>"100101100",
  20365=>"111111101",
  20366=>"000000111",
  20367=>"001011101",
  20368=>"000000011",
  20369=>"110010101",
  20370=>"010101100",
  20371=>"101100010",
  20372=>"010000010",
  20373=>"100100100",
  20374=>"101011100",
  20375=>"111001001",
  20376=>"110001111",
  20377=>"010110101",
  20378=>"100000110",
  20379=>"010101010",
  20380=>"100100110",
  20381=>"010000000",
  20382=>"101111100",
  20383=>"011000001",
  20384=>"100110110",
  20385=>"011101111",
  20386=>"001110101",
  20387=>"110001001",
  20388=>"010100001",
  20389=>"010111111",
  20390=>"001101011",
  20391=>"101101010",
  20392=>"000010101",
  20393=>"101100001",
  20394=>"000010011",
  20395=>"010101010",
  20396=>"011011100",
  20397=>"100001111",
  20398=>"100010101",
  20399=>"000110101",
  20400=>"110111001",
  20401=>"111011011",
  20402=>"011100011",
  20403=>"110101101",
  20404=>"000101100",
  20405=>"010110010",
  20406=>"000010010",
  20407=>"001010010",
  20408=>"010100011",
  20409=>"101111001",
  20410=>"010110001",
  20411=>"011011011",
  20412=>"111101001",
  20413=>"001100110",
  20414=>"000001110",
  20415=>"000100000",
  20416=>"011111010",
  20417=>"111100011",
  20418=>"100010111",
  20419=>"100011101",
  20420=>"011111010",
  20421=>"010111101",
  20422=>"110011111",
  20423=>"001011011",
  20424=>"000001101",
  20425=>"101001111",
  20426=>"100011111",
  20427=>"111001000",
  20428=>"001111110",
  20429=>"100000100",
  20430=>"101101011",
  20431=>"110000110",
  20432=>"111100011",
  20433=>"110100011",
  20434=>"000101000",
  20435=>"000001100",
  20436=>"000101110",
  20437=>"000000000",
  20438=>"000010011",
  20439=>"010011111",
  20440=>"001001001",
  20441=>"001000110",
  20442=>"000101011",
  20443=>"000001011",
  20444=>"111100111",
  20445=>"100000100",
  20446=>"110000011",
  20447=>"011010010",
  20448=>"011110000",
  20449=>"111100011",
  20450=>"001011110",
  20451=>"110101010",
  20452=>"000110101",
  20453=>"000111001",
  20454=>"110010000",
  20455=>"110010111",
  20456=>"100110000",
  20457=>"110100001",
  20458=>"001000010",
  20459=>"100001100",
  20460=>"000000110",
  20461=>"110001010",
  20462=>"101000001",
  20463=>"001000010",
  20464=>"101001010",
  20465=>"101000011",
  20466=>"000000101",
  20467=>"110011101",
  20468=>"101101100",
  20469=>"001110010",
  20470=>"011001010",
  20471=>"100101000",
  20472=>"000000001",
  20473=>"101110010",
  20474=>"111010000",
  20475=>"011101110",
  20476=>"100111110",
  20477=>"010010111",
  20478=>"100010000",
  20479=>"100000010",
  20480=>"011010110",
  20481=>"010111001",
  20482=>"001101101",
  20483=>"001000100",
  20484=>"010001101",
  20485=>"101001101",
  20486=>"101100101",
  20487=>"101001010",
  20488=>"110100001",
  20489=>"000100110",
  20490=>"001101100",
  20491=>"101100111",
  20492=>"001000100",
  20493=>"111010110",
  20494=>"111101000",
  20495=>"100000010",
  20496=>"010010110",
  20497=>"101000001",
  20498=>"010111110",
  20499=>"101001101",
  20500=>"000101111",
  20501=>"010110000",
  20502=>"110010100",
  20503=>"110000001",
  20504=>"111111110",
  20505=>"000000000",
  20506=>"010110110",
  20507=>"011111101",
  20508=>"101001101",
  20509=>"011001100",
  20510=>"101011010",
  20511=>"111101001",
  20512=>"010100100",
  20513=>"101010000",
  20514=>"101000110",
  20515=>"001101001",
  20516=>"010100111",
  20517=>"110000101",
  20518=>"110011110",
  20519=>"000000001",
  20520=>"011010011",
  20521=>"000101011",
  20522=>"001011110",
  20523=>"010101001",
  20524=>"100011000",
  20525=>"111001111",
  20526=>"101101001",
  20527=>"011100011",
  20528=>"101111111",
  20529=>"111010000",
  20530=>"110010010",
  20531=>"110111110",
  20532=>"011101000",
  20533=>"011100010",
  20534=>"001101110",
  20535=>"011010001",
  20536=>"000001010",
  20537=>"111110100",
  20538=>"001010110",
  20539=>"110100101",
  20540=>"010000000",
  20541=>"011101100",
  20542=>"110000010",
  20543=>"000110001",
  20544=>"001011011",
  20545=>"000001001",
  20546=>"000011101",
  20547=>"111111001",
  20548=>"000100110",
  20549=>"100001111",
  20550=>"110010001",
  20551=>"100001100",
  20552=>"101001110",
  20553=>"100011111",
  20554=>"101000111",
  20555=>"010011011",
  20556=>"000011100",
  20557=>"101010111",
  20558=>"001000010",
  20559=>"000001011",
  20560=>"100010011",
  20561=>"010100101",
  20562=>"011111111",
  20563=>"100011101",
  20564=>"100000110",
  20565=>"010111000",
  20566=>"000100010",
  20567=>"000011101",
  20568=>"101000000",
  20569=>"111010000",
  20570=>"101101001",
  20571=>"000000000",
  20572=>"111100111",
  20573=>"000100100",
  20574=>"110001000",
  20575=>"111001111",
  20576=>"100010000",
  20577=>"001010111",
  20578=>"000111000",
  20579=>"001010000",
  20580=>"111010001",
  20581=>"111000100",
  20582=>"000010010",
  20583=>"001110100",
  20584=>"101101100",
  20585=>"000001101",
  20586=>"000101110",
  20587=>"100001101",
  20588=>"000110111",
  20589=>"111100110",
  20590=>"001000111",
  20591=>"110000110",
  20592=>"110101110",
  20593=>"100111100",
  20594=>"000011100",
  20595=>"110011101",
  20596=>"101110111",
  20597=>"010100111",
  20598=>"111111110",
  20599=>"101011101",
  20600=>"100000110",
  20601=>"110101111",
  20602=>"010000010",
  20603=>"000100011",
  20604=>"101000001",
  20605=>"010110101",
  20606=>"011011011",
  20607=>"111110111",
  20608=>"101000101",
  20609=>"000101111",
  20610=>"100100011",
  20611=>"001111000",
  20612=>"001001101",
  20613=>"000111101",
  20614=>"100001111",
  20615=>"101001110",
  20616=>"010111010",
  20617=>"101011100",
  20618=>"000000000",
  20619=>"011011011",
  20620=>"000000110",
  20621=>"000111101",
  20622=>"101001110",
  20623=>"101000111",
  20624=>"001011101",
  20625=>"011000100",
  20626=>"001010001",
  20627=>"101100111",
  20628=>"101010011",
  20629=>"101010000",
  20630=>"000011101",
  20631=>"000001011",
  20632=>"111100011",
  20633=>"110100010",
  20634=>"011001101",
  20635=>"001000101",
  20636=>"010110000",
  20637=>"111010100",
  20638=>"010001011",
  20639=>"000000101",
  20640=>"111001101",
  20641=>"001010101",
  20642=>"110000101",
  20643=>"110110110",
  20644=>"011111111",
  20645=>"011110100",
  20646=>"000010101",
  20647=>"101000100",
  20648=>"100001011",
  20649=>"111001101",
  20650=>"000101101",
  20651=>"001101011",
  20652=>"010111011",
  20653=>"000010101",
  20654=>"001010110",
  20655=>"101000110",
  20656=>"111010111",
  20657=>"100010011",
  20658=>"001101010",
  20659=>"100101110",
  20660=>"100101110",
  20661=>"100000000",
  20662=>"000010111",
  20663=>"000100011",
  20664=>"111001110",
  20665=>"010110100",
  20666=>"001110000",
  20667=>"100101110",
  20668=>"001011001",
  20669=>"100111100",
  20670=>"000111000",
  20671=>"000010100",
  20672=>"111000101",
  20673=>"011001101",
  20674=>"111111110",
  20675=>"111110001",
  20676=>"010111010",
  20677=>"001001100",
  20678=>"010100011",
  20679=>"101101100",
  20680=>"110111100",
  20681=>"000110010",
  20682=>"100000010",
  20683=>"101010010",
  20684=>"111111110",
  20685=>"010100010",
  20686=>"011010010",
  20687=>"000011000",
  20688=>"110000000",
  20689=>"100000001",
  20690=>"001111111",
  20691=>"100000110",
  20692=>"100011100",
  20693=>"000010100",
  20694=>"011110000",
  20695=>"011110100",
  20696=>"000101110",
  20697=>"001010010",
  20698=>"000111000",
  20699=>"100111110",
  20700=>"111111101",
  20701=>"100010001",
  20702=>"001011100",
  20703=>"100111001",
  20704=>"111010010",
  20705=>"001000010",
  20706=>"011001111",
  20707=>"011101110",
  20708=>"110000100",
  20709=>"000001011",
  20710=>"100111100",
  20711=>"001001100",
  20712=>"101010110",
  20713=>"000111000",
  20714=>"001000010",
  20715=>"000110001",
  20716=>"000000000",
  20717=>"001011101",
  20718=>"000001100",
  20719=>"101111110",
  20720=>"010111000",
  20721=>"010101000",
  20722=>"100010111",
  20723=>"101110000",
  20724=>"010110010",
  20725=>"110110110",
  20726=>"011100100",
  20727=>"100110011",
  20728=>"010010101",
  20729=>"011110011",
  20730=>"101101000",
  20731=>"000100001",
  20732=>"010001011",
  20733=>"101011111",
  20734=>"111101100",
  20735=>"110100111",
  20736=>"110010110",
  20737=>"001111101",
  20738=>"011110100",
  20739=>"011011010",
  20740=>"111110111",
  20741=>"001001100",
  20742=>"000000111",
  20743=>"001100100",
  20744=>"000000111",
  20745=>"011110010",
  20746=>"010001001",
  20747=>"111100101",
  20748=>"000101101",
  20749=>"111010001",
  20750=>"101110101",
  20751=>"101001000",
  20752=>"001110010",
  20753=>"000010111",
  20754=>"100110111",
  20755=>"010110010",
  20756=>"011100110",
  20757=>"101111010",
  20758=>"101110100",
  20759=>"110101110",
  20760=>"100101001",
  20761=>"100001101",
  20762=>"000100010",
  20763=>"010001101",
  20764=>"110011110",
  20765=>"111110010",
  20766=>"000101100",
  20767=>"000000000",
  20768=>"001110010",
  20769=>"110100011",
  20770=>"111001110",
  20771=>"000000110",
  20772=>"000111111",
  20773=>"111010011",
  20774=>"110011111",
  20775=>"110001111",
  20776=>"000000010",
  20777=>"011100000",
  20778=>"100010000",
  20779=>"110001010",
  20780=>"111101110",
  20781=>"101111111",
  20782=>"110011010",
  20783=>"111100101",
  20784=>"111111100",
  20785=>"101010100",
  20786=>"111100111",
  20787=>"111101111",
  20788=>"010100110",
  20789=>"010000101",
  20790=>"001100100",
  20791=>"011110111",
  20792=>"000000101",
  20793=>"000101100",
  20794=>"110000110",
  20795=>"111011001",
  20796=>"010010111",
  20797=>"101001111",
  20798=>"001100000",
  20799=>"110111101",
  20800=>"010101101",
  20801=>"110110001",
  20802=>"110001001",
  20803=>"000001100",
  20804=>"111001010",
  20805=>"101011001",
  20806=>"000000000",
  20807=>"111001101",
  20808=>"001101001",
  20809=>"011100110",
  20810=>"001000000",
  20811=>"101101101",
  20812=>"000100101",
  20813=>"101001110",
  20814=>"110010101",
  20815=>"101101101",
  20816=>"011111011",
  20817=>"001000110",
  20818=>"011001010",
  20819=>"010010110",
  20820=>"000000111",
  20821=>"011110010",
  20822=>"010011111",
  20823=>"010000011",
  20824=>"100011001",
  20825=>"010010001",
  20826=>"011101111",
  20827=>"000111101",
  20828=>"111110000",
  20829=>"111011001",
  20830=>"000000110",
  20831=>"011010100",
  20832=>"011111001",
  20833=>"000010101",
  20834=>"111100101",
  20835=>"100011111",
  20836=>"110000000",
  20837=>"110000100",
  20838=>"100101011",
  20839=>"100111111",
  20840=>"111110011",
  20841=>"001000011",
  20842=>"010011000",
  20843=>"001101100",
  20844=>"001110100",
  20845=>"001110111",
  20846=>"011000110",
  20847=>"011110111",
  20848=>"100010111",
  20849=>"101100100",
  20850=>"000110001",
  20851=>"011000101",
  20852=>"011001101",
  20853=>"000100011",
  20854=>"001000011",
  20855=>"101000100",
  20856=>"110101111",
  20857=>"100001010",
  20858=>"111100000",
  20859=>"111101011",
  20860=>"101011100",
  20861=>"110100101",
  20862=>"000111111",
  20863=>"011011110",
  20864=>"110001111",
  20865=>"101110110",
  20866=>"001011100",
  20867=>"010110101",
  20868=>"010001011",
  20869=>"010101111",
  20870=>"001111001",
  20871=>"011100110",
  20872=>"110001011",
  20873=>"000110110",
  20874=>"000111000",
  20875=>"101110001",
  20876=>"110111111",
  20877=>"000011010",
  20878=>"101110110",
  20879=>"110111101",
  20880=>"100001011",
  20881=>"100000000",
  20882=>"010010001",
  20883=>"010110011",
  20884=>"000110001",
  20885=>"000011101",
  20886=>"111100100",
  20887=>"101001011",
  20888=>"010010010",
  20889=>"000000110",
  20890=>"011001000",
  20891=>"100110101",
  20892=>"011111001",
  20893=>"111000000",
  20894=>"110011001",
  20895=>"100011101",
  20896=>"110100010",
  20897=>"011010101",
  20898=>"100110101",
  20899=>"001000000",
  20900=>"101011001",
  20901=>"101101110",
  20902=>"110010110",
  20903=>"001000000",
  20904=>"011011110",
  20905=>"011011100",
  20906=>"010110001",
  20907=>"111110100",
  20908=>"110101100",
  20909=>"101100010",
  20910=>"011110110",
  20911=>"000010000",
  20912=>"010100001",
  20913=>"000000101",
  20914=>"000000010",
  20915=>"111110001",
  20916=>"100000111",
  20917=>"011000001",
  20918=>"111000001",
  20919=>"110101111",
  20920=>"011011011",
  20921=>"100000101",
  20922=>"111100101",
  20923=>"000001001",
  20924=>"111101100",
  20925=>"100100011",
  20926=>"010000001",
  20927=>"011010101",
  20928=>"101100011",
  20929=>"011110111",
  20930=>"001110011",
  20931=>"101110010",
  20932=>"111011100",
  20933=>"000100001",
  20934=>"100001001",
  20935=>"000000101",
  20936=>"110010011",
  20937=>"000000100",
  20938=>"010000101",
  20939=>"010101010",
  20940=>"100000100",
  20941=>"011001010",
  20942=>"110011100",
  20943=>"110001011",
  20944=>"100010101",
  20945=>"101101100",
  20946=>"110011110",
  20947=>"001011010",
  20948=>"110111000",
  20949=>"000000101",
  20950=>"011010010",
  20951=>"100111000",
  20952=>"111001011",
  20953=>"000001011",
  20954=>"001111111",
  20955=>"111100000",
  20956=>"011101010",
  20957=>"100010000",
  20958=>"101010110",
  20959=>"101001101",
  20960=>"100011000",
  20961=>"100001011",
  20962=>"110000000",
  20963=>"001101001",
  20964=>"100111110",
  20965=>"101000101",
  20966=>"110010010",
  20967=>"111100101",
  20968=>"101111101",
  20969=>"111011000",
  20970=>"100001110",
  20971=>"111110001",
  20972=>"010100111",
  20973=>"000110101",
  20974=>"101011011",
  20975=>"000111010",
  20976=>"000010000",
  20977=>"111101111",
  20978=>"110111010",
  20979=>"111001000",
  20980=>"000100011",
  20981=>"111010101",
  20982=>"001000000",
  20983=>"000111110",
  20984=>"011010111",
  20985=>"101110000",
  20986=>"000000000",
  20987=>"001001010",
  20988=>"001000111",
  20989=>"100111010",
  20990=>"001011000",
  20991=>"100110111",
  20992=>"111101101",
  20993=>"110101010",
  20994=>"100011011",
  20995=>"101100011",
  20996=>"010000100",
  20997=>"000000100",
  20998=>"111110010",
  20999=>"010010000",
  21000=>"011101000",
  21001=>"001101011",
  21002=>"110001111",
  21003=>"111001001",
  21004=>"000011010",
  21005=>"011100111",
  21006=>"000010001",
  21007=>"100101011",
  21008=>"100100110",
  21009=>"010011011",
  21010=>"111100111",
  21011=>"111110111",
  21012=>"000110011",
  21013=>"010101111",
  21014=>"111000110",
  21015=>"001110011",
  21016=>"010110010",
  21017=>"111101011",
  21018=>"101101101",
  21019=>"000001101",
  21020=>"010001011",
  21021=>"000100001",
  21022=>"101001110",
  21023=>"111010110",
  21024=>"010001011",
  21025=>"111100011",
  21026=>"001010110",
  21027=>"011111101",
  21028=>"000100011",
  21029=>"111101000",
  21030=>"100101111",
  21031=>"110010110",
  21032=>"010010100",
  21033=>"011110011",
  21034=>"001001001",
  21035=>"100000011",
  21036=>"100010111",
  21037=>"010101010",
  21038=>"011101010",
  21039=>"001110111",
  21040=>"110110011",
  21041=>"110100011",
  21042=>"100110010",
  21043=>"000001110",
  21044=>"110000110",
  21045=>"100110100",
  21046=>"010001000",
  21047=>"010010100",
  21048=>"101100011",
  21049=>"001001011",
  21050=>"100100110",
  21051=>"011111000",
  21052=>"000010000",
  21053=>"000000101",
  21054=>"110001110",
  21055=>"101100000",
  21056=>"000001011",
  21057=>"100001000",
  21058=>"011011000",
  21059=>"001110110",
  21060=>"010011011",
  21061=>"010001111",
  21062=>"010100111",
  21063=>"110100100",
  21064=>"011001001",
  21065=>"100010011",
  21066=>"100000010",
  21067=>"111111111",
  21068=>"110010100",
  21069=>"111000110",
  21070=>"101010110",
  21071=>"101011010",
  21072=>"000100000",
  21073=>"110010011",
  21074=>"110101000",
  21075=>"111100010",
  21076=>"101101100",
  21077=>"000010000",
  21078=>"100100100",
  21079=>"011100010",
  21080=>"010111010",
  21081=>"100010010",
  21082=>"000001111",
  21083=>"111100101",
  21084=>"000111001",
  21085=>"000011110",
  21086=>"000111010",
  21087=>"000000101",
  21088=>"001111001",
  21089=>"110000010",
  21090=>"010010111",
  21091=>"101011011",
  21092=>"111010110",
  21093=>"011111101",
  21094=>"110011101",
  21095=>"111001110",
  21096=>"101000010",
  21097=>"000110100",
  21098=>"100011001",
  21099=>"100111000",
  21100=>"001011111",
  21101=>"000000000",
  21102=>"100111011",
  21103=>"101101111",
  21104=>"101000000",
  21105=>"110100010",
  21106=>"111001100",
  21107=>"101011100",
  21108=>"010001010",
  21109=>"111011110",
  21110=>"011100001",
  21111=>"001001111",
  21112=>"100100100",
  21113=>"011111101",
  21114=>"100110011",
  21115=>"110000100",
  21116=>"011001000",
  21117=>"100111110",
  21118=>"001101011",
  21119=>"101011111",
  21120=>"101110100",
  21121=>"001001011",
  21122=>"110111111",
  21123=>"000111101",
  21124=>"101101011",
  21125=>"111100100",
  21126=>"111000010",
  21127=>"011001010",
  21128=>"111000110",
  21129=>"011110110",
  21130=>"101000011",
  21131=>"001111110",
  21132=>"010110011",
  21133=>"100101000",
  21134=>"100000110",
  21135=>"011111101",
  21136=>"100111001",
  21137=>"110100000",
  21138=>"010001001",
  21139=>"001101111",
  21140=>"010011111",
  21141=>"110001010",
  21142=>"101001101",
  21143=>"100100110",
  21144=>"001001000",
  21145=>"111100001",
  21146=>"101011110",
  21147=>"101110100",
  21148=>"111100001",
  21149=>"110100010",
  21150=>"001011011",
  21151=>"001010101",
  21152=>"111101100",
  21153=>"111001001",
  21154=>"101010010",
  21155=>"111011101",
  21156=>"111011101",
  21157=>"100101110",
  21158=>"100111001",
  21159=>"101011011",
  21160=>"010000000",
  21161=>"100010000",
  21162=>"011001011",
  21163=>"101110111",
  21164=>"011000010",
  21165=>"001011110",
  21166=>"011110000",
  21167=>"100001000",
  21168=>"110011100",
  21169=>"000001001",
  21170=>"010011000",
  21171=>"010110111",
  21172=>"010100101",
  21173=>"110000101",
  21174=>"100110000",
  21175=>"000011101",
  21176=>"000000011",
  21177=>"011000111",
  21178=>"101011011",
  21179=>"100101001",
  21180=>"100011001",
  21181=>"011001010",
  21182=>"010111001",
  21183=>"110011110",
  21184=>"101110010",
  21185=>"001101101",
  21186=>"001011000",
  21187=>"101011000",
  21188=>"010010011",
  21189=>"100001011",
  21190=>"111010101",
  21191=>"100110101",
  21192=>"011101000",
  21193=>"001001010",
  21194=>"000011110",
  21195=>"010011001",
  21196=>"000111111",
  21197=>"001101011",
  21198=>"101110100",
  21199=>"001010011",
  21200=>"101111010",
  21201=>"011011100",
  21202=>"000011001",
  21203=>"000000100",
  21204=>"101101000",
  21205=>"110111000",
  21206=>"101010011",
  21207=>"111001111",
  21208=>"010001000",
  21209=>"000100011",
  21210=>"101010100",
  21211=>"010011001",
  21212=>"011000011",
  21213=>"000011010",
  21214=>"000010100",
  21215=>"111011001",
  21216=>"101011001",
  21217=>"100001101",
  21218=>"010011101",
  21219=>"001001111",
  21220=>"111001010",
  21221=>"010010000",
  21222=>"010101100",
  21223=>"101011110",
  21224=>"000111011",
  21225=>"101001110",
  21226=>"000110011",
  21227=>"101011111",
  21228=>"011110110",
  21229=>"001010101",
  21230=>"000001101",
  21231=>"110101100",
  21232=>"111111111",
  21233=>"111100000",
  21234=>"011101001",
  21235=>"001101100",
  21236=>"111101001",
  21237=>"101101100",
  21238=>"000110101",
  21239=>"101111001",
  21240=>"010100101",
  21241=>"101100000",
  21242=>"001101010",
  21243=>"101001100",
  21244=>"000110111",
  21245=>"110010000",
  21246=>"011101000",
  21247=>"011011110",
  21248=>"001100000",
  21249=>"001101010",
  21250=>"111110010",
  21251=>"011110011",
  21252=>"110110101",
  21253=>"010101010",
  21254=>"010011001",
  21255=>"111000100",
  21256=>"001111111",
  21257=>"110000110",
  21258=>"000011100",
  21259=>"000000000",
  21260=>"001001001",
  21261=>"111111010",
  21262=>"000000111",
  21263=>"110111100",
  21264=>"010110001",
  21265=>"000010110",
  21266=>"001001001",
  21267=>"101000001",
  21268=>"101000110",
  21269=>"011010011",
  21270=>"010110111",
  21271=>"100001000",
  21272=>"100101001",
  21273=>"010010110",
  21274=>"000110001",
  21275=>"010110010",
  21276=>"101001100",
  21277=>"010100101",
  21278=>"010100011",
  21279=>"010111000",
  21280=>"001111100",
  21281=>"111110110",
  21282=>"111111001",
  21283=>"111010001",
  21284=>"100000011",
  21285=>"000111100",
  21286=>"001100110",
  21287=>"010110000",
  21288=>"111000111",
  21289=>"111010111",
  21290=>"010110110",
  21291=>"110001010",
  21292=>"011000000",
  21293=>"111001100",
  21294=>"000011100",
  21295=>"101111001",
  21296=>"000100100",
  21297=>"100101111",
  21298=>"101110100",
  21299=>"010001001",
  21300=>"010000101",
  21301=>"011000101",
  21302=>"011000111",
  21303=>"111110001",
  21304=>"001110111",
  21305=>"000000010",
  21306=>"011110110",
  21307=>"111111000",
  21308=>"001110001",
  21309=>"001011000",
  21310=>"011110000",
  21311=>"111010110",
  21312=>"000101110",
  21313=>"001111011",
  21314=>"111111111",
  21315=>"111011010",
  21316=>"001010001",
  21317=>"110000010",
  21318=>"101101100",
  21319=>"001010111",
  21320=>"101111010",
  21321=>"111110100",
  21322=>"011110111",
  21323=>"111011000",
  21324=>"010111011",
  21325=>"001111000",
  21326=>"000001011",
  21327=>"100000101",
  21328=>"100001000",
  21329=>"000010000",
  21330=>"011111010",
  21331=>"000110001",
  21332=>"100111111",
  21333=>"111111110",
  21334=>"111110010",
  21335=>"000001110",
  21336=>"001000010",
  21337=>"011001101",
  21338=>"100111000",
  21339=>"110110010",
  21340=>"000000001",
  21341=>"000100100",
  21342=>"111100111",
  21343=>"010100011",
  21344=>"100000000",
  21345=>"111001001",
  21346=>"001110011",
  21347=>"101000000",
  21348=>"110010100",
  21349=>"111100111",
  21350=>"110001011",
  21351=>"000101011",
  21352=>"000100000",
  21353=>"010001011",
  21354=>"110001001",
  21355=>"110111101",
  21356=>"110011110",
  21357=>"001111000",
  21358=>"110100111",
  21359=>"101110100",
  21360=>"010000000",
  21361=>"011110111",
  21362=>"101011111",
  21363=>"010010010",
  21364=>"111110111",
  21365=>"000100111",
  21366=>"111000100",
  21367=>"111001111",
  21368=>"010110011",
  21369=>"001111101",
  21370=>"010000010",
  21371=>"000010110",
  21372=>"111000011",
  21373=>"111110101",
  21374=>"011111101",
  21375=>"011000010",
  21376=>"000011011",
  21377=>"011010100",
  21378=>"110111100",
  21379=>"110100000",
  21380=>"101000000",
  21381=>"000101101",
  21382=>"100111011",
  21383=>"000010000",
  21384=>"001010000",
  21385=>"011000101",
  21386=>"111011011",
  21387=>"110010010",
  21388=>"100110111",
  21389=>"000011011",
  21390=>"011111111",
  21391=>"011001110",
  21392=>"100111001",
  21393=>"011110011",
  21394=>"000010000",
  21395=>"010110010",
  21396=>"010111001",
  21397=>"100101000",
  21398=>"111011000",
  21399=>"110011111",
  21400=>"001110010",
  21401=>"101011100",
  21402=>"111101110",
  21403=>"010000101",
  21404=>"001011101",
  21405=>"001100111",
  21406=>"000001000",
  21407=>"101101001",
  21408=>"001110010",
  21409=>"010101010",
  21410=>"000000110",
  21411=>"000100010",
  21412=>"000100001",
  21413=>"110111011",
  21414=>"000111011",
  21415=>"011001000",
  21416=>"000001100",
  21417=>"001010110",
  21418=>"101101011",
  21419=>"110100011",
  21420=>"001100100",
  21421=>"100010000",
  21422=>"011001001",
  21423=>"111010010",
  21424=>"101101100",
  21425=>"011011001",
  21426=>"101101011",
  21427=>"111111001",
  21428=>"000101111",
  21429=>"011010000",
  21430=>"111000001",
  21431=>"001110011",
  21432=>"110001000",
  21433=>"011010011",
  21434=>"011110111",
  21435=>"000011100",
  21436=>"011101110",
  21437=>"000110010",
  21438=>"111010100",
  21439=>"000010000",
  21440=>"101000100",
  21441=>"110001011",
  21442=>"110110001",
  21443=>"010011000",
  21444=>"110010010",
  21445=>"011110001",
  21446=>"101010100",
  21447=>"110110011",
  21448=>"110100011",
  21449=>"111100001",
  21450=>"101111110",
  21451=>"111011101",
  21452=>"011011101",
  21453=>"011110100",
  21454=>"100110101",
  21455=>"000011010",
  21456=>"111110011",
  21457=>"000100110",
  21458=>"011110100",
  21459=>"101000011",
  21460=>"001010010",
  21461=>"111010010",
  21462=>"110001011",
  21463=>"011001100",
  21464=>"010010001",
  21465=>"001110000",
  21466=>"100101110",
  21467=>"111100100",
  21468=>"100111010",
  21469=>"110110011",
  21470=>"000000111",
  21471=>"011110010",
  21472=>"101011001",
  21473=>"111110001",
  21474=>"110000010",
  21475=>"011100111",
  21476=>"111100010",
  21477=>"100010001",
  21478=>"000010001",
  21479=>"001000011",
  21480=>"001111011",
  21481=>"101010100",
  21482=>"011100100",
  21483=>"100010110",
  21484=>"100000101",
  21485=>"100100101",
  21486=>"100011001",
  21487=>"100111001",
  21488=>"010011001",
  21489=>"010010110",
  21490=>"000000100",
  21491=>"000101100",
  21492=>"111001100",
  21493=>"000000011",
  21494=>"001011000",
  21495=>"010110000",
  21496=>"101000110",
  21497=>"000001011",
  21498=>"000001111",
  21499=>"000100011",
  21500=>"111001111",
  21501=>"011111000",
  21502=>"011000010",
  21503=>"101011111",
  21504=>"000001001",
  21505=>"011110001",
  21506=>"101101111",
  21507=>"001101110",
  21508=>"101111101",
  21509=>"000111011",
  21510=>"111111110",
  21511=>"101101000",
  21512=>"110011101",
  21513=>"111110100",
  21514=>"101110011",
  21515=>"000001101",
  21516=>"101110010",
  21517=>"010110001",
  21518=>"101011011",
  21519=>"010010101",
  21520=>"101111010",
  21521=>"010011100",
  21522=>"110011000",
  21523=>"111110010",
  21524=>"100111000",
  21525=>"100111010",
  21526=>"101100011",
  21527=>"011000101",
  21528=>"100110011",
  21529=>"101101000",
  21530=>"101111110",
  21531=>"110110010",
  21532=>"011110100",
  21533=>"100111001",
  21534=>"101000011",
  21535=>"110001000",
  21536=>"111001111",
  21537=>"010010100",
  21538=>"001010001",
  21539=>"001100011",
  21540=>"001111010",
  21541=>"111111011",
  21542=>"100011001",
  21543=>"101000100",
  21544=>"001110110",
  21545=>"000000011",
  21546=>"011000111",
  21547=>"001010010",
  21548=>"000111110",
  21549=>"101100111",
  21550=>"100101111",
  21551=>"110011100",
  21552=>"111010000",
  21553=>"101010101",
  21554=>"010101010",
  21555=>"000110111",
  21556=>"110000010",
  21557=>"000110101",
  21558=>"110110101",
  21559=>"001111000",
  21560=>"000100011",
  21561=>"010000010",
  21562=>"111111101",
  21563=>"001001010",
  21564=>"000100110",
  21565=>"010111101",
  21566=>"100001011",
  21567=>"011011010",
  21568=>"101010110",
  21569=>"111011101",
  21570=>"000010100",
  21571=>"001000110",
  21572=>"011001010",
  21573=>"000101100",
  21574=>"010011100",
  21575=>"010001010",
  21576=>"111001011",
  21577=>"110011001",
  21578=>"011001000",
  21579=>"011001111",
  21580=>"011001011",
  21581=>"111011001",
  21582=>"000011110",
  21583=>"101111000",
  21584=>"011011101",
  21585=>"100101100",
  21586=>"101000010",
  21587=>"100101101",
  21588=>"000100011",
  21589=>"010111010",
  21590=>"000100001",
  21591=>"010010000",
  21592=>"110111000",
  21593=>"011001101",
  21594=>"000001001",
  21595=>"110001001",
  21596=>"000100101",
  21597=>"011000010",
  21598=>"111111100",
  21599=>"100110101",
  21600=>"001001000",
  21601=>"010110100",
  21602=>"000001111",
  21603=>"100000011",
  21604=>"010011111",
  21605=>"000000010",
  21606=>"001100001",
  21607=>"010110000",
  21608=>"011111100",
  21609=>"101001000",
  21610=>"000100000",
  21611=>"100110101",
  21612=>"100101101",
  21613=>"100100001",
  21614=>"110000000",
  21615=>"110110100",
  21616=>"000001000",
  21617=>"000000000",
  21618=>"101110001",
  21619=>"100011111",
  21620=>"000101011",
  21621=>"010011101",
  21622=>"111111001",
  21623=>"110100111",
  21624=>"011010101",
  21625=>"010111001",
  21626=>"001100000",
  21627=>"000001111",
  21628=>"011010101",
  21629=>"010101001",
  21630=>"100010011",
  21631=>"011000111",
  21632=>"001001000",
  21633=>"000011000",
  21634=>"011001101",
  21635=>"010101100",
  21636=>"000001111",
  21637=>"011011011",
  21638=>"010010100",
  21639=>"000001010",
  21640=>"111000010",
  21641=>"110101001",
  21642=>"011001110",
  21643=>"110100110",
  21644=>"001001101",
  21645=>"101011101",
  21646=>"110001001",
  21647=>"110111101",
  21648=>"001110100",
  21649=>"000010000",
  21650=>"111100100",
  21651=>"111011001",
  21652=>"101100000",
  21653=>"011111011",
  21654=>"110001100",
  21655=>"011101100",
  21656=>"101001101",
  21657=>"000001101",
  21658=>"000000110",
  21659=>"101111110",
  21660=>"010100110",
  21661=>"001001010",
  21662=>"111010101",
  21663=>"011110011",
  21664=>"001101010",
  21665=>"001101100",
  21666=>"110000000",
  21667=>"001001100",
  21668=>"110001111",
  21669=>"000001100",
  21670=>"110101000",
  21671=>"000110000",
  21672=>"101110100",
  21673=>"101010111",
  21674=>"001010110",
  21675=>"111111101",
  21676=>"001001001",
  21677=>"101010011",
  21678=>"111100011",
  21679=>"010111101",
  21680=>"001000110",
  21681=>"011000100",
  21682=>"111110000",
  21683=>"010001111",
  21684=>"000010010",
  21685=>"000001000",
  21686=>"101111111",
  21687=>"110001111",
  21688=>"010101100",
  21689=>"010010110",
  21690=>"100111110",
  21691=>"101010101",
  21692=>"010000001",
  21693=>"101010000",
  21694=>"001010101",
  21695=>"010111110",
  21696=>"001110101",
  21697=>"100011110",
  21698=>"111111110",
  21699=>"110010100",
  21700=>"110111011",
  21701=>"000000001",
  21702=>"111000001",
  21703=>"100000101",
  21704=>"101001100",
  21705=>"000100001",
  21706=>"011100001",
  21707=>"011100110",
  21708=>"000111100",
  21709=>"100000001",
  21710=>"000101000",
  21711=>"101010101",
  21712=>"010000110",
  21713=>"011000001",
  21714=>"010011000",
  21715=>"111000111",
  21716=>"011011111",
  21717=>"101101011",
  21718=>"101000011",
  21719=>"101101111",
  21720=>"000100101",
  21721=>"001010110",
  21722=>"001000101",
  21723=>"110011100",
  21724=>"000011111",
  21725=>"010111110",
  21726=>"100010101",
  21727=>"010001100",
  21728=>"000111000",
  21729=>"011001001",
  21730=>"101111111",
  21731=>"000110101",
  21732=>"110001111",
  21733=>"000011100",
  21734=>"000001000",
  21735=>"110100110",
  21736=>"011001100",
  21737=>"001111110",
  21738=>"010100000",
  21739=>"011101110",
  21740=>"010001000",
  21741=>"001011110",
  21742=>"000100100",
  21743=>"001111101",
  21744=>"010011000",
  21745=>"111001000",
  21746=>"010100011",
  21747=>"101111100",
  21748=>"110111100",
  21749=>"110110100",
  21750=>"111111101",
  21751=>"000000100",
  21752=>"101011000",
  21753=>"111110011",
  21754=>"001111000",
  21755=>"100000000",
  21756=>"111001111",
  21757=>"110101000",
  21758=>"101000011",
  21759=>"110111010",
  21760=>"111111100",
  21761=>"110001000",
  21762=>"011011010",
  21763=>"001000111",
  21764=>"111101101",
  21765=>"100100111",
  21766=>"001000010",
  21767=>"011010000",
  21768=>"100000011",
  21769=>"010111110",
  21770=>"110101000",
  21771=>"001001110",
  21772=>"000001000",
  21773=>"010111000",
  21774=>"010111001",
  21775=>"000000000",
  21776=>"110000000",
  21777=>"001000100",
  21778=>"000000010",
  21779=>"111110010",
  21780=>"100101000",
  21781=>"110101101",
  21782=>"011101000",
  21783=>"100001111",
  21784=>"000110000",
  21785=>"100001000",
  21786=>"100001100",
  21787=>"001110000",
  21788=>"011001111",
  21789=>"111100000",
  21790=>"010000011",
  21791=>"000001111",
  21792=>"100110110",
  21793=>"111010000",
  21794=>"000000001",
  21795=>"000000101",
  21796=>"110110111",
  21797=>"110000100",
  21798=>"011101011",
  21799=>"000011111",
  21800=>"100101111",
  21801=>"100010011",
  21802=>"011100100",
  21803=>"100101010",
  21804=>"111100010",
  21805=>"011111101",
  21806=>"000010111",
  21807=>"011010001",
  21808=>"111111111",
  21809=>"000001010",
  21810=>"001100010",
  21811=>"000010110",
  21812=>"111011000",
  21813=>"111110111",
  21814=>"010111000",
  21815=>"000011101",
  21816=>"101000110",
  21817=>"111010100",
  21818=>"000101110",
  21819=>"010011011",
  21820=>"101000100",
  21821=>"110000011",
  21822=>"011100111",
  21823=>"101100000",
  21824=>"100000000",
  21825=>"111111011",
  21826=>"001000111",
  21827=>"011100101",
  21828=>"111001101",
  21829=>"000010011",
  21830=>"011101110",
  21831=>"011000000",
  21832=>"100110101",
  21833=>"001111001",
  21834=>"001111011",
  21835=>"001001111",
  21836=>"010011100",
  21837=>"011010001",
  21838=>"100111001",
  21839=>"111110011",
  21840=>"100111100",
  21841=>"100011100",
  21842=>"101000001",
  21843=>"000001011",
  21844=>"111010000",
  21845=>"100011000",
  21846=>"011010010",
  21847=>"000011101",
  21848=>"001000100",
  21849=>"000111111",
  21850=>"100110100",
  21851=>"100101101",
  21852=>"110101100",
  21853=>"110011001",
  21854=>"101011001",
  21855=>"010010101",
  21856=>"001011111",
  21857=>"001101101",
  21858=>"010010010",
  21859=>"001001111",
  21860=>"101010110",
  21861=>"000001011",
  21862=>"111101101",
  21863=>"101011011",
  21864=>"011000101",
  21865=>"010000100",
  21866=>"100011101",
  21867=>"001100111",
  21868=>"101101010",
  21869=>"011101100",
  21870=>"110001101",
  21871=>"000100111",
  21872=>"010100010",
  21873=>"011100011",
  21874=>"110110000",
  21875=>"010001100",
  21876=>"110011100",
  21877=>"001001010",
  21878=>"011101111",
  21879=>"000100111",
  21880=>"000111111",
  21881=>"000010101",
  21882=>"110101010",
  21883=>"111100010",
  21884=>"101000110",
  21885=>"010101011",
  21886=>"101000110",
  21887=>"110000011",
  21888=>"100101101",
  21889=>"000000001",
  21890=>"001101101",
  21891=>"011100010",
  21892=>"011000100",
  21893=>"001100010",
  21894=>"010011110",
  21895=>"111011010",
  21896=>"010111110",
  21897=>"101101001",
  21898=>"000010000",
  21899=>"100100000",
  21900=>"000001010",
  21901=>"100000110",
  21902=>"110110001",
  21903=>"110011111",
  21904=>"011111100",
  21905=>"000001000",
  21906=>"110101010",
  21907=>"100110011",
  21908=>"001011000",
  21909=>"001110000",
  21910=>"111100011",
  21911=>"000000111",
  21912=>"000001010",
  21913=>"000000001",
  21914=>"001001101",
  21915=>"100110101",
  21916=>"000111000",
  21917=>"110001011",
  21918=>"100101011",
  21919=>"000010010",
  21920=>"001010001",
  21921=>"100110010",
  21922=>"010111100",
  21923=>"000000100",
  21924=>"010100100",
  21925=>"000001000",
  21926=>"000001111",
  21927=>"111011010",
  21928=>"100001010",
  21929=>"000000010",
  21930=>"100110010",
  21931=>"001011101",
  21932=>"010011100",
  21933=>"100001110",
  21934=>"110100001",
  21935=>"100111010",
  21936=>"101101110",
  21937=>"100001010",
  21938=>"001011000",
  21939=>"110000101",
  21940=>"101111111",
  21941=>"111100001",
  21942=>"010001010",
  21943=>"100000001",
  21944=>"101101101",
  21945=>"000011110",
  21946=>"001000001",
  21947=>"111101100",
  21948=>"010101100",
  21949=>"011101001",
  21950=>"100001010",
  21951=>"011010000",
  21952=>"100011100",
  21953=>"110110100",
  21954=>"001110001",
  21955=>"100001000",
  21956=>"001000110",
  21957=>"011100001",
  21958=>"001010101",
  21959=>"000100001",
  21960=>"011100011",
  21961=>"001110100",
  21962=>"010001000",
  21963=>"011001111",
  21964=>"011010111",
  21965=>"101011010",
  21966=>"000100001",
  21967=>"100111011",
  21968=>"010011011",
  21969=>"000001010",
  21970=>"001101011",
  21971=>"101111010",
  21972=>"100100110",
  21973=>"110100000",
  21974=>"100100111",
  21975=>"111011100",
  21976=>"101011001",
  21977=>"111011001",
  21978=>"111110010",
  21979=>"001011001",
  21980=>"100011000",
  21981=>"101110001",
  21982=>"011011111",
  21983=>"101010110",
  21984=>"100110010",
  21985=>"101110010",
  21986=>"010110101",
  21987=>"101111111",
  21988=>"001111000",
  21989=>"101101100",
  21990=>"110110010",
  21991=>"101101010",
  21992=>"001010011",
  21993=>"101101011",
  21994=>"110111000",
  21995=>"011011100",
  21996=>"001100100",
  21997=>"001001001",
  21998=>"010001001",
  21999=>"101000010",
  22000=>"000011010",
  22001=>"100011100",
  22002=>"001001001",
  22003=>"001000111",
  22004=>"111110111",
  22005=>"100010101",
  22006=>"001010111",
  22007=>"110100101",
  22008=>"101110101",
  22009=>"010100101",
  22010=>"000100000",
  22011=>"010111000",
  22012=>"000010010",
  22013=>"111001100",
  22014=>"000001010",
  22015=>"001001110",
  22016=>"100011111",
  22017=>"111110110",
  22018=>"010110011",
  22019=>"011101110",
  22020=>"000011000",
  22021=>"010100111",
  22022=>"001000101",
  22023=>"100001110",
  22024=>"101011101",
  22025=>"110010101",
  22026=>"011011101",
  22027=>"100010010",
  22028=>"000001001",
  22029=>"101001111",
  22030=>"110010100",
  22031=>"100111011",
  22032=>"001110111",
  22033=>"111111100",
  22034=>"001011111",
  22035=>"011111110",
  22036=>"001000110",
  22037=>"010111100",
  22038=>"010111011",
  22039=>"110111110",
  22040=>"010001100",
  22041=>"011100100",
  22042=>"100000100",
  22043=>"110001010",
  22044=>"100000101",
  22045=>"001000110",
  22046=>"111101111",
  22047=>"111111000",
  22048=>"111001101",
  22049=>"101010101",
  22050=>"001110110",
  22051=>"110010110",
  22052=>"011001111",
  22053=>"000110010",
  22054=>"101001000",
  22055=>"010001100",
  22056=>"101000000",
  22057=>"111110010",
  22058=>"001010111",
  22059=>"110101000",
  22060=>"111111110",
  22061=>"101000001",
  22062=>"001000000",
  22063=>"111001101",
  22064=>"010010111",
  22065=>"101110001",
  22066=>"001100111",
  22067=>"000000011",
  22068=>"101111101",
  22069=>"101010010",
  22070=>"101001110",
  22071=>"100010110",
  22072=>"100001010",
  22073=>"011011110",
  22074=>"010100101",
  22075=>"000101110",
  22076=>"000111100",
  22077=>"000111101",
  22078=>"001110001",
  22079=>"110111100",
  22080=>"101111110",
  22081=>"101100000",
  22082=>"010100011",
  22083=>"100110101",
  22084=>"000110001",
  22085=>"110101011",
  22086=>"010100101",
  22087=>"010100111",
  22088=>"000000000",
  22089=>"110110011",
  22090=>"111010000",
  22091=>"100011100",
  22092=>"010011001",
  22093=>"100011000",
  22094=>"111001010",
  22095=>"001011110",
  22096=>"101010000",
  22097=>"111010110",
  22098=>"101110110",
  22099=>"001100101",
  22100=>"010011110",
  22101=>"000101110",
  22102=>"000011010",
  22103=>"000010011",
  22104=>"111000110",
  22105=>"000100010",
  22106=>"110011100",
  22107=>"100100100",
  22108=>"100001101",
  22109=>"000101101",
  22110=>"111011010",
  22111=>"111111011",
  22112=>"101001000",
  22113=>"000110111",
  22114=>"101110010",
  22115=>"110110101",
  22116=>"111110111",
  22117=>"101101010",
  22118=>"000101111",
  22119=>"001010011",
  22120=>"000101111",
  22121=>"001011000",
  22122=>"001110110",
  22123=>"111110011",
  22124=>"100110010",
  22125=>"001101000",
  22126=>"101011011",
  22127=>"111111011",
  22128=>"101000010",
  22129=>"000101111",
  22130=>"011110010",
  22131=>"001001111",
  22132=>"110001101",
  22133=>"010011001",
  22134=>"111011011",
  22135=>"110011100",
  22136=>"000001111",
  22137=>"100101001",
  22138=>"101101110",
  22139=>"101101010",
  22140=>"001101111",
  22141=>"010000101",
  22142=>"110100101",
  22143=>"011010000",
  22144=>"011110110",
  22145=>"110110111",
  22146=>"110011111",
  22147=>"011001110",
  22148=>"001010110",
  22149=>"100010000",
  22150=>"001101100",
  22151=>"000001001",
  22152=>"010111010",
  22153=>"000011011",
  22154=>"010011110",
  22155=>"110001010",
  22156=>"000000000",
  22157=>"100001111",
  22158=>"010001001",
  22159=>"011011001",
  22160=>"100010001",
  22161=>"010111000",
  22162=>"111111110",
  22163=>"101111111",
  22164=>"000100100",
  22165=>"000001100",
  22166=>"111110111",
  22167=>"001100011",
  22168=>"011000101",
  22169=>"001010011",
  22170=>"010000000",
  22171=>"100010011",
  22172=>"101011110",
  22173=>"001011001",
  22174=>"001000101",
  22175=>"011001010",
  22176=>"101011011",
  22177=>"111110101",
  22178=>"100101010",
  22179=>"011000010",
  22180=>"111110010",
  22181=>"111010000",
  22182=>"001100110",
  22183=>"111111001",
  22184=>"011010001",
  22185=>"010100001",
  22186=>"011011010",
  22187=>"100100011",
  22188=>"001001010",
  22189=>"000101110",
  22190=>"011011100",
  22191=>"111101100",
  22192=>"010111110",
  22193=>"001000011",
  22194=>"010011000",
  22195=>"101010000",
  22196=>"011010011",
  22197=>"111110101",
  22198=>"100000111",
  22199=>"111100110",
  22200=>"101101011",
  22201=>"011100010",
  22202=>"001111111",
  22203=>"000001101",
  22204=>"101110111",
  22205=>"101110100",
  22206=>"001000001",
  22207=>"011010011",
  22208=>"011110101",
  22209=>"100100011",
  22210=>"100001011",
  22211=>"010010011",
  22212=>"000010101",
  22213=>"010100101",
  22214=>"111100000",
  22215=>"001010001",
  22216=>"110001010",
  22217=>"111010000",
  22218=>"011111111",
  22219=>"100000010",
  22220=>"000111001",
  22221=>"100110000",
  22222=>"011001110",
  22223=>"000110100",
  22224=>"100011010",
  22225=>"111010001",
  22226=>"101011101",
  22227=>"100000011",
  22228=>"000100100",
  22229=>"000001110",
  22230=>"101000000",
  22231=>"011110010",
  22232=>"010000100",
  22233=>"100011111",
  22234=>"101000001",
  22235=>"011011001",
  22236=>"110000110",
  22237=>"000100000",
  22238=>"101100110",
  22239=>"100110111",
  22240=>"000001010",
  22241=>"000101100",
  22242=>"110010110",
  22243=>"111111011",
  22244=>"111101111",
  22245=>"110100010",
  22246=>"000100011",
  22247=>"001110011",
  22248=>"001010011",
  22249=>"111111101",
  22250=>"011010110",
  22251=>"000011111",
  22252=>"100100101",
  22253=>"010101011",
  22254=>"100011110",
  22255=>"001101000",
  22256=>"111100100",
  22257=>"011000011",
  22258=>"011000101",
  22259=>"110000101",
  22260=>"111000101",
  22261=>"110111110",
  22262=>"010000010",
  22263=>"000111010",
  22264=>"111010010",
  22265=>"010010011",
  22266=>"010001000",
  22267=>"000000000",
  22268=>"101110011",
  22269=>"000010011",
  22270=>"111000110",
  22271=>"111100001",
  22272=>"101010111",
  22273=>"000000101",
  22274=>"100011110",
  22275=>"100101111",
  22276=>"101011110",
  22277=>"110011111",
  22278=>"010111101",
  22279=>"110001101",
  22280=>"110110001",
  22281=>"111000111",
  22282=>"100001100",
  22283=>"010000000",
  22284=>"100000110",
  22285=>"011100010",
  22286=>"011011100",
  22287=>"110101001",
  22288=>"011010111",
  22289=>"101000101",
  22290=>"010011101",
  22291=>"011011101",
  22292=>"011011111",
  22293=>"001111110",
  22294=>"011110111",
  22295=>"000110111",
  22296=>"000111100",
  22297=>"000101100",
  22298=>"011110111",
  22299=>"100001101",
  22300=>"110111011",
  22301=>"111001110",
  22302=>"010010100",
  22303=>"111000100",
  22304=>"000100101",
  22305=>"000110111",
  22306=>"111000101",
  22307=>"000000101",
  22308=>"110000110",
  22309=>"101000010",
  22310=>"111101111",
  22311=>"010010000",
  22312=>"110011100",
  22313=>"110000111",
  22314=>"010001101",
  22315=>"111111011",
  22316=>"101101111",
  22317=>"101011011",
  22318=>"000110010",
  22319=>"010111000",
  22320=>"010011010",
  22321=>"100101101",
  22322=>"010010010",
  22323=>"001011111",
  22324=>"110110001",
  22325=>"110101011",
  22326=>"111011110",
  22327=>"110101100",
  22328=>"011101101",
  22329=>"100100001",
  22330=>"101011011",
  22331=>"010010010",
  22332=>"110010111",
  22333=>"001101101",
  22334=>"000000000",
  22335=>"111101110",
  22336=>"010110111",
  22337=>"001000010",
  22338=>"010101011",
  22339=>"010000111",
  22340=>"001111110",
  22341=>"001000101",
  22342=>"001010100",
  22343=>"110101000",
  22344=>"000110001",
  22345=>"110000000",
  22346=>"010111110",
  22347=>"000101001",
  22348=>"111100100",
  22349=>"001001000",
  22350=>"001010000",
  22351=>"011110101",
  22352=>"001101010",
  22353=>"010000010",
  22354=>"011100100",
  22355=>"100100101",
  22356=>"000100010",
  22357=>"101111110",
  22358=>"100000000",
  22359=>"111100001",
  22360=>"001100101",
  22361=>"110111111",
  22362=>"001111111",
  22363=>"110110001",
  22364=>"000011001",
  22365=>"100100100",
  22366=>"011001011",
  22367=>"000110111",
  22368=>"101001000",
  22369=>"110001001",
  22370=>"000010001",
  22371=>"101010110",
  22372=>"000010110",
  22373=>"011001110",
  22374=>"010111110",
  22375=>"110010001",
  22376=>"111001000",
  22377=>"111011110",
  22378=>"000000000",
  22379=>"011010011",
  22380=>"101010110",
  22381=>"010101100",
  22382=>"001011001",
  22383=>"011111100",
  22384=>"000111100",
  22385=>"110011100",
  22386=>"001110011",
  22387=>"100001000",
  22388=>"010010110",
  22389=>"001010010",
  22390=>"000000100",
  22391=>"000101011",
  22392=>"100001101",
  22393=>"011010010",
  22394=>"101110110",
  22395=>"110000101",
  22396=>"000011011",
  22397=>"001010010",
  22398=>"011100010",
  22399=>"111000101",
  22400=>"000010100",
  22401=>"110101100",
  22402=>"000011100",
  22403=>"101010101",
  22404=>"011010111",
  22405=>"001001000",
  22406=>"001100010",
  22407=>"110011000",
  22408=>"110011000",
  22409=>"011110111",
  22410=>"101111000",
  22411=>"011000110",
  22412=>"011010110",
  22413=>"001011001",
  22414=>"110001001",
  22415=>"111110000",
  22416=>"101001101",
  22417=>"111101101",
  22418=>"011000000",
  22419=>"100100100",
  22420=>"101000111",
  22421=>"010101100",
  22422=>"010001100",
  22423=>"010100001",
  22424=>"111000000",
  22425=>"010010100",
  22426=>"100110000",
  22427=>"010000111",
  22428=>"000010100",
  22429=>"101000110",
  22430=>"100010111",
  22431=>"011010111",
  22432=>"010000001",
  22433=>"101011100",
  22434=>"000101010",
  22435=>"100001011",
  22436=>"110000000",
  22437=>"101101000",
  22438=>"101000011",
  22439=>"000110011",
  22440=>"101101000",
  22441=>"000010010",
  22442=>"101101001",
  22443=>"010101001",
  22444=>"001010101",
  22445=>"101101110",
  22446=>"110101111",
  22447=>"111100111",
  22448=>"001000100",
  22449=>"111110100",
  22450=>"110000000",
  22451=>"011000000",
  22452=>"100000111",
  22453=>"011001110",
  22454=>"110101111",
  22455=>"110000010",
  22456=>"101110111",
  22457=>"000110011",
  22458=>"100101000",
  22459=>"110001110",
  22460=>"001110000",
  22461=>"000101101",
  22462=>"110001010",
  22463=>"110110110",
  22464=>"011010110",
  22465=>"011100011",
  22466=>"111010000",
  22467=>"111100010",
  22468=>"101010101",
  22469=>"010001100",
  22470=>"011101001",
  22471=>"110100001",
  22472=>"010000001",
  22473=>"100111001",
  22474=>"111101111",
  22475=>"111001011",
  22476=>"010011010",
  22477=>"010001110",
  22478=>"000111001",
  22479=>"011100000",
  22480=>"111011010",
  22481=>"010111111",
  22482=>"001000000",
  22483=>"011100000",
  22484=>"111001111",
  22485=>"000111000",
  22486=>"110011000",
  22487=>"111110110",
  22488=>"000101001",
  22489=>"100001110",
  22490=>"011110001",
  22491=>"100000111",
  22492=>"001100100",
  22493=>"111101110",
  22494=>"111011011",
  22495=>"001000001",
  22496=>"001111011",
  22497=>"101110101",
  22498=>"101111100",
  22499=>"101001111",
  22500=>"000011010",
  22501=>"111100110",
  22502=>"000101010",
  22503=>"000000000",
  22504=>"000101100",
  22505=>"101011111",
  22506=>"010101100",
  22507=>"010111010",
  22508=>"000000001",
  22509=>"100110000",
  22510=>"001000010",
  22511=>"011110001",
  22512=>"011010101",
  22513=>"101100011",
  22514=>"001110010",
  22515=>"010111110",
  22516=>"100011010",
  22517=>"100010101",
  22518=>"010001111",
  22519=>"110111010",
  22520=>"101000111",
  22521=>"100000110",
  22522=>"010001110",
  22523=>"101100100",
  22524=>"111101100",
  22525=>"111001010",
  22526=>"110100110",
  22527=>"011111001",
  22528=>"000100100",
  22529=>"100101101",
  22530=>"001101100",
  22531=>"010000110",
  22532=>"001010111",
  22533=>"011010001",
  22534=>"101110010",
  22535=>"110011000",
  22536=>"111100101",
  22537=>"100010000",
  22538=>"011100010",
  22539=>"110100100",
  22540=>"000010000",
  22541=>"101010111",
  22542=>"010000100",
  22543=>"001101100",
  22544=>"011010011",
  22545=>"111110000",
  22546=>"011101010",
  22547=>"010110000",
  22548=>"011011101",
  22549=>"000110001",
  22550=>"111110010",
  22551=>"101111110",
  22552=>"010000011",
  22553=>"111001101",
  22554=>"011111000",
  22555=>"011010001",
  22556=>"000010100",
  22557=>"111100011",
  22558=>"100110001",
  22559=>"010100000",
  22560=>"010110000",
  22561=>"110101100",
  22562=>"111111110",
  22563=>"111101111",
  22564=>"000111000",
  22565=>"100001011",
  22566=>"110101011",
  22567=>"011001111",
  22568=>"110110010",
  22569=>"010000000",
  22570=>"100110111",
  22571=>"101110111",
  22572=>"101000110",
  22573=>"110011110",
  22574=>"010101011",
  22575=>"000000011",
  22576=>"101101011",
  22577=>"000010110",
  22578=>"000111100",
  22579=>"001101011",
  22580=>"111110110",
  22581=>"001110101",
  22582=>"101110101",
  22583=>"000000100",
  22584=>"000101110",
  22585=>"110100101",
  22586=>"101000110",
  22587=>"000100100",
  22588=>"110111100",
  22589=>"001000101",
  22590=>"001011100",
  22591=>"110000010",
  22592=>"011111001",
  22593=>"100001000",
  22594=>"111000011",
  22595=>"110101011",
  22596=>"101111000",
  22597=>"111100010",
  22598=>"101111011",
  22599=>"111110111",
  22600=>"010111010",
  22601=>"010111111",
  22602=>"011010000",
  22603=>"111001110",
  22604=>"111101010",
  22605=>"110001010",
  22606=>"111000110",
  22607=>"110011010",
  22608=>"110011111",
  22609=>"010110011",
  22610=>"000001101",
  22611=>"000101110",
  22612=>"000100001",
  22613=>"000001011",
  22614=>"001010000",
  22615=>"010100001",
  22616=>"000110111",
  22617=>"000011011",
  22618=>"011101101",
  22619=>"001000011",
  22620=>"011001100",
  22621=>"000010110",
  22622=>"110001000",
  22623=>"010101110",
  22624=>"111010010",
  22625=>"011011001",
  22626=>"101101001",
  22627=>"110010000",
  22628=>"110111101",
  22629=>"001000000",
  22630=>"101001100",
  22631=>"101011010",
  22632=>"001100111",
  22633=>"001000000",
  22634=>"110110100",
  22635=>"010110110",
  22636=>"111010000",
  22637=>"001011011",
  22638=>"111111111",
  22639=>"100000110",
  22640=>"010010000",
  22641=>"000101111",
  22642=>"010010011",
  22643=>"100101011",
  22644=>"100101000",
  22645=>"110101111",
  22646=>"011110011",
  22647=>"111110010",
  22648=>"010000100",
  22649=>"101111111",
  22650=>"010010110",
  22651=>"001000111",
  22652=>"011100101",
  22653=>"100001010",
  22654=>"011010111",
  22655=>"111110011",
  22656=>"000000001",
  22657=>"100011111",
  22658=>"011110000",
  22659=>"001000001",
  22660=>"101100000",
  22661=>"100110101",
  22662=>"011000010",
  22663=>"101001010",
  22664=>"011111100",
  22665=>"000101101",
  22666=>"011101011",
  22667=>"011011110",
  22668=>"100100111",
  22669=>"110100001",
  22670=>"010111000",
  22671=>"010010101",
  22672=>"001111100",
  22673=>"000001001",
  22674=>"001101110",
  22675=>"101111111",
  22676=>"111010101",
  22677=>"100000001",
  22678=>"000100111",
  22679=>"100011101",
  22680=>"110111100",
  22681=>"011011110",
  22682=>"110101100",
  22683=>"110010100",
  22684=>"010000001",
  22685=>"101010001",
  22686=>"000001110",
  22687=>"000000010",
  22688=>"111001111",
  22689=>"000000011",
  22690=>"110010101",
  22691=>"110010111",
  22692=>"110100101",
  22693=>"010100111",
  22694=>"101011100",
  22695=>"000011000",
  22696=>"000001000",
  22697=>"111111001",
  22698=>"011000000",
  22699=>"011011110",
  22700=>"100110001",
  22701=>"101101011",
  22702=>"101101001",
  22703=>"001110100",
  22704=>"010111100",
  22705=>"111001010",
  22706=>"001001000",
  22707=>"001000001",
  22708=>"011100001",
  22709=>"001110001",
  22710=>"001011011",
  22711=>"111011101",
  22712=>"010010100",
  22713=>"010011011",
  22714=>"111100001",
  22715=>"001010010",
  22716=>"001101111",
  22717=>"010010110",
  22718=>"001000100",
  22719=>"110111100",
  22720=>"110100101",
  22721=>"001001001",
  22722=>"000111110",
  22723=>"111110110",
  22724=>"110101111",
  22725=>"011100000",
  22726=>"010001100",
  22727=>"111010110",
  22728=>"001001000",
  22729=>"100100111",
  22730=>"101101001",
  22731=>"010011011",
  22732=>"010000111",
  22733=>"010001101",
  22734=>"110010101",
  22735=>"110100100",
  22736=>"000010010",
  22737=>"010001001",
  22738=>"010010100",
  22739=>"100000101",
  22740=>"101110111",
  22741=>"101011111",
  22742=>"101110111",
  22743=>"010000101",
  22744=>"001011101",
  22745=>"101000010",
  22746=>"000111001",
  22747=>"001001100",
  22748=>"101100010",
  22749=>"010100100",
  22750=>"000000011",
  22751=>"111110100",
  22752=>"011011001",
  22753=>"000111000",
  22754=>"000101110",
  22755=>"100010111",
  22756=>"011000001",
  22757=>"100110111",
  22758=>"110011110",
  22759=>"001111110",
  22760=>"110111110",
  22761=>"011001001",
  22762=>"100000100",
  22763=>"101111011",
  22764=>"100011010",
  22765=>"101110111",
  22766=>"110110010",
  22767=>"011110001",
  22768=>"101001111",
  22769=>"011111100",
  22770=>"011111011",
  22771=>"001010011",
  22772=>"101101001",
  22773=>"001000010",
  22774=>"111100101",
  22775=>"000100010",
  22776=>"001011110",
  22777=>"010011110",
  22778=>"100001100",
  22779=>"010110111",
  22780=>"110110000",
  22781=>"001000110",
  22782=>"100100101",
  22783=>"011000100",
  22784=>"011011010",
  22785=>"011100111",
  22786=>"111101101",
  22787=>"110101001",
  22788=>"010011001",
  22789=>"001100100",
  22790=>"001110011",
  22791=>"000101011",
  22792=>"011000101",
  22793=>"000011011",
  22794=>"101111110",
  22795=>"110001000",
  22796=>"010010001",
  22797=>"011011100",
  22798=>"101001001",
  22799=>"110010110",
  22800=>"101110011",
  22801=>"010100110",
  22802=>"111001110",
  22803=>"101110011",
  22804=>"000000001",
  22805=>"110001110",
  22806=>"111010000",
  22807=>"001111010",
  22808=>"010000011",
  22809=>"000100000",
  22810=>"100111110",
  22811=>"010100110",
  22812=>"000101011",
  22813=>"100111000",
  22814=>"010101111",
  22815=>"010000010",
  22816=>"000000101",
  22817=>"010100110",
  22818=>"100010110",
  22819=>"110100011",
  22820=>"000010010",
  22821=>"011100010",
  22822=>"001110111",
  22823=>"010101000",
  22824=>"110111110",
  22825=>"110100011",
  22826=>"011010000",
  22827=>"011100101",
  22828=>"110010000",
  22829=>"111100001",
  22830=>"000001111",
  22831=>"110110011",
  22832=>"010001011",
  22833=>"100111011",
  22834=>"111100110",
  22835=>"110001100",
  22836=>"000000010",
  22837=>"011000101",
  22838=>"010110100",
  22839=>"000110110",
  22840=>"101010111",
  22841=>"011100010",
  22842=>"011100101",
  22843=>"010110010",
  22844=>"010100100",
  22845=>"111011010",
  22846=>"000110000",
  22847=>"111111111",
  22848=>"101000001",
  22849=>"101001000",
  22850=>"101110110",
  22851=>"100001001",
  22852=>"000000110",
  22853=>"100101111",
  22854=>"110000111",
  22855=>"010000101",
  22856=>"001001011",
  22857=>"011100111",
  22858=>"000000010",
  22859=>"101000000",
  22860=>"100101001",
  22861=>"111011110",
  22862=>"100010001",
  22863=>"000101101",
  22864=>"111111011",
  22865=>"111011001",
  22866=>"101000101",
  22867=>"011010011",
  22868=>"110010010",
  22869=>"001111000",
  22870=>"100000011",
  22871=>"010010100",
  22872=>"000010000",
  22873=>"101111000",
  22874=>"010111010",
  22875=>"111111100",
  22876=>"101100111",
  22877=>"000101101",
  22878=>"101000001",
  22879=>"000110001",
  22880=>"110100001",
  22881=>"000101000",
  22882=>"110111110",
  22883=>"000000001",
  22884=>"000100000",
  22885=>"111100010",
  22886=>"111100001",
  22887=>"110010111",
  22888=>"011010011",
  22889=>"000010001",
  22890=>"101100100",
  22891=>"010110110",
  22892=>"011101111",
  22893=>"111011000",
  22894=>"101011001",
  22895=>"100010000",
  22896=>"111011000",
  22897=>"101101111",
  22898=>"001001100",
  22899=>"101000110",
  22900=>"000000011",
  22901=>"101111001",
  22902=>"010111011",
  22903=>"111111111",
  22904=>"000000010",
  22905=>"100100110",
  22906=>"011001101",
  22907=>"110000000",
  22908=>"100001110",
  22909=>"101111110",
  22910=>"110010110",
  22911=>"100001100",
  22912=>"011111011",
  22913=>"000100101",
  22914=>"111010100",
  22915=>"110001100",
  22916=>"101011111",
  22917=>"001000111",
  22918=>"011011000",
  22919=>"000111100",
  22920=>"001110000",
  22921=>"001001010",
  22922=>"111101011",
  22923=>"000110100",
  22924=>"111000111",
  22925=>"000000101",
  22926=>"110011001",
  22927=>"100001001",
  22928=>"000000011",
  22929=>"010000000",
  22930=>"010011011",
  22931=>"110100001",
  22932=>"111110111",
  22933=>"000001100",
  22934=>"010000000",
  22935=>"001011101",
  22936=>"110110110",
  22937=>"001000001",
  22938=>"001010011",
  22939=>"010101000",
  22940=>"100110111",
  22941=>"111100010",
  22942=>"101001001",
  22943=>"000100001",
  22944=>"011010001",
  22945=>"111100111",
  22946=>"001100001",
  22947=>"111010100",
  22948=>"100010000",
  22949=>"011111000",
  22950=>"110001100",
  22951=>"011001111",
  22952=>"111101101",
  22953=>"000100001",
  22954=>"000100010",
  22955=>"000101100",
  22956=>"010001100",
  22957=>"111110001",
  22958=>"000001100",
  22959=>"101111101",
  22960=>"110110100",
  22961=>"110010100",
  22962=>"010001011",
  22963=>"111000000",
  22964=>"001010010",
  22965=>"100111001",
  22966=>"001111100",
  22967=>"110011011",
  22968=>"110110110",
  22969=>"010000001",
  22970=>"000111110",
  22971=>"000111001",
  22972=>"110100010",
  22973=>"100111110",
  22974=>"000110111",
  22975=>"111111100",
  22976=>"111001111",
  22977=>"001011001",
  22978=>"100011000",
  22979=>"011010011",
  22980=>"111110110",
  22981=>"001110000",
  22982=>"011000010",
  22983=>"110010000",
  22984=>"110100000",
  22985=>"101010101",
  22986=>"000000010",
  22987=>"001011011",
  22988=>"000100000",
  22989=>"000000100",
  22990=>"010110011",
  22991=>"110100110",
  22992=>"001011101",
  22993=>"101100111",
  22994=>"000000110",
  22995=>"110001010",
  22996=>"000100011",
  22997=>"001101011",
  22998=>"001111101",
  22999=>"000100010",
  23000=>"101000100",
  23001=>"101101001",
  23002=>"011100011",
  23003=>"110000011",
  23004=>"011100011",
  23005=>"001101101",
  23006=>"000100000",
  23007=>"110101001",
  23008=>"101010000",
  23009=>"100001100",
  23010=>"110001010",
  23011=>"010011001",
  23012=>"010100011",
  23013=>"011010001",
  23014=>"001010010",
  23015=>"010001010",
  23016=>"111110110",
  23017=>"000011111",
  23018=>"100010010",
  23019=>"001000000",
  23020=>"110100001",
  23021=>"101000001",
  23022=>"111110101",
  23023=>"001001001",
  23024=>"100100001",
  23025=>"011000001",
  23026=>"010111000",
  23027=>"000100011",
  23028=>"101011101",
  23029=>"100101001",
  23030=>"101111011",
  23031=>"000001001",
  23032=>"101101110",
  23033=>"010111000",
  23034=>"001000101",
  23035=>"000100010",
  23036=>"010010011",
  23037=>"000000010",
  23038=>"110101101",
  23039=>"000011011",
  23040=>"101100001",
  23041=>"011011100",
  23042=>"000001010",
  23043=>"100000110",
  23044=>"101000011",
  23045=>"000010010",
  23046=>"000010101",
  23047=>"010001110",
  23048=>"001100001",
  23049=>"101001011",
  23050=>"100000101",
  23051=>"111100011",
  23052=>"110111111",
  23053=>"000111101",
  23054=>"010000110",
  23055=>"100001111",
  23056=>"000100010",
  23057=>"110100100",
  23058=>"100101011",
  23059=>"001101010",
  23060=>"011111101",
  23061=>"101100100",
  23062=>"100111001",
  23063=>"001011001",
  23064=>"001101110",
  23065=>"100101000",
  23066=>"000011010",
  23067=>"110110001",
  23068=>"110010010",
  23069=>"000111010",
  23070=>"010100111",
  23071=>"011111011",
  23072=>"100111110",
  23073=>"011010010",
  23074=>"110010011",
  23075=>"011100111",
  23076=>"100010110",
  23077=>"101010000",
  23078=>"001001011",
  23079=>"010101000",
  23080=>"101101000",
  23081=>"110111101",
  23082=>"001110011",
  23083=>"000111110",
  23084=>"110000100",
  23085=>"001001001",
  23086=>"001010001",
  23087=>"010011100",
  23088=>"111001001",
  23089=>"001000011",
  23090=>"010000001",
  23091=>"101111011",
  23092=>"000111100",
  23093=>"001011011",
  23094=>"000000010",
  23095=>"110111110",
  23096=>"110101100",
  23097=>"010000100",
  23098=>"100001011",
  23099=>"111111001",
  23100=>"000011101",
  23101=>"110110110",
  23102=>"010001000",
  23103=>"111110111",
  23104=>"110111011",
  23105=>"100000111",
  23106=>"011110101",
  23107=>"001000111",
  23108=>"001100000",
  23109=>"100001100",
  23110=>"000101001",
  23111=>"110100001",
  23112=>"000110011",
  23113=>"110010110",
  23114=>"101111101",
  23115=>"111000000",
  23116=>"100000000",
  23117=>"100011101",
  23118=>"100111100",
  23119=>"001010000",
  23120=>"111101000",
  23121=>"001100110",
  23122=>"100000110",
  23123=>"001001110",
  23124=>"101010000",
  23125=>"010000011",
  23126=>"100001011",
  23127=>"011110011",
  23128=>"110101110",
  23129=>"011010011",
  23130=>"001011000",
  23131=>"000001010",
  23132=>"111100000",
  23133=>"011000011",
  23134=>"011011111",
  23135=>"001011001",
  23136=>"111101111",
  23137=>"101000000",
  23138=>"100111101",
  23139=>"000101110",
  23140=>"010001111",
  23141=>"010000100",
  23142=>"010011001",
  23143=>"001001011",
  23144=>"100011101",
  23145=>"010001001",
  23146=>"011111111",
  23147=>"000110000",
  23148=>"111000111",
  23149=>"011010111",
  23150=>"101101101",
  23151=>"011001111",
  23152=>"000001111",
  23153=>"010110000",
  23154=>"000100001",
  23155=>"001111110",
  23156=>"110011111",
  23157=>"000101101",
  23158=>"011110011",
  23159=>"011110111",
  23160=>"000010001",
  23161=>"101100000",
  23162=>"111011110",
  23163=>"001110010",
  23164=>"000011011",
  23165=>"101110100",
  23166=>"001000000",
  23167=>"101110001",
  23168=>"100101010",
  23169=>"011011010",
  23170=>"110100110",
  23171=>"001100000",
  23172=>"111010100",
  23173=>"101110111",
  23174=>"001011011",
  23175=>"111010000",
  23176=>"100011011",
  23177=>"110010000",
  23178=>"110011110",
  23179=>"001011101",
  23180=>"000010000",
  23181=>"001000001",
  23182=>"001000110",
  23183=>"000100110",
  23184=>"111110101",
  23185=>"110100100",
  23186=>"101110001",
  23187=>"001110111",
  23188=>"100000100",
  23189=>"001010011",
  23190=>"010111110",
  23191=>"101100111",
  23192=>"000000010",
  23193=>"101011111",
  23194=>"110001011",
  23195=>"110011000",
  23196=>"111100100",
  23197=>"100000000",
  23198=>"111100111",
  23199=>"000111010",
  23200=>"111011010",
  23201=>"100001100",
  23202=>"111111111",
  23203=>"101100101",
  23204=>"011000100",
  23205=>"001100000",
  23206=>"010010110",
  23207=>"001000010",
  23208=>"111011011",
  23209=>"011111110",
  23210=>"101001000",
  23211=>"010000010",
  23212=>"011000110",
  23213=>"100011010",
  23214=>"011100111",
  23215=>"010011001",
  23216=>"100010001",
  23217=>"011011101",
  23218=>"100001011",
  23219=>"001011111",
  23220=>"000100010",
  23221=>"111011110",
  23222=>"000010010",
  23223=>"010000011",
  23224=>"101110011",
  23225=>"001011010",
  23226=>"101000000",
  23227=>"000001110",
  23228=>"000100000",
  23229=>"010110011",
  23230=>"110001101",
  23231=>"101011001",
  23232=>"100100101",
  23233=>"001101001",
  23234=>"100100011",
  23235=>"010100001",
  23236=>"001100100",
  23237=>"000100001",
  23238=>"010010111",
  23239=>"010110111",
  23240=>"101100001",
  23241=>"011001111",
  23242=>"100100100",
  23243=>"010111100",
  23244=>"011101101",
  23245=>"111011001",
  23246=>"100111000",
  23247=>"101000111",
  23248=>"111001100",
  23249=>"000001100",
  23250=>"001101101",
  23251=>"001010110",
  23252=>"111100111",
  23253=>"001110111",
  23254=>"001010011",
  23255=>"111000101",
  23256=>"110101010",
  23257=>"111100111",
  23258=>"111000001",
  23259=>"011011001",
  23260=>"000010011",
  23261=>"110111011",
  23262=>"110100101",
  23263=>"011010100",
  23264=>"111101011",
  23265=>"101101110",
  23266=>"100100110",
  23267=>"100110110",
  23268=>"111001001",
  23269=>"000011110",
  23270=>"101011011",
  23271=>"111010101",
  23272=>"010010011",
  23273=>"001001101",
  23274=>"000000001",
  23275=>"110010000",
  23276=>"011010100",
  23277=>"000001110",
  23278=>"010000000",
  23279=>"110111111",
  23280=>"110111011",
  23281=>"010010010",
  23282=>"100111011",
  23283=>"101110111",
  23284=>"011111001",
  23285=>"011011101",
  23286=>"100100011",
  23287=>"110010010",
  23288=>"000101100",
  23289=>"101011010",
  23290=>"101110000",
  23291=>"000011101",
  23292=>"110010101",
  23293=>"100111100",
  23294=>"001110101",
  23295=>"010111010",
  23296=>"000011111",
  23297=>"001110110",
  23298=>"100100101",
  23299=>"101111111",
  23300=>"011100100",
  23301=>"011010001",
  23302=>"110010101",
  23303=>"101011101",
  23304=>"000000001",
  23305=>"100001101",
  23306=>"100010001",
  23307=>"000000010",
  23308=>"111110110",
  23309=>"100011101",
  23310=>"100100111",
  23311=>"110000001",
  23312=>"100110000",
  23313=>"000010000",
  23314=>"111110001",
  23315=>"010110110",
  23316=>"001101011",
  23317=>"001001111",
  23318=>"000101100",
  23319=>"000000001",
  23320=>"000011010",
  23321=>"101110101",
  23322=>"001101111",
  23323=>"000101001",
  23324=>"011001001",
  23325=>"011101110",
  23326=>"011111010",
  23327=>"100100010",
  23328=>"010000010",
  23329=>"000010110",
  23330=>"111110001",
  23331=>"100100110",
  23332=>"101001111",
  23333=>"111110110",
  23334=>"000110011",
  23335=>"100101000",
  23336=>"010011110",
  23337=>"000011110",
  23338=>"011100010",
  23339=>"001001010",
  23340=>"001110101",
  23341=>"100101100",
  23342=>"111010111",
  23343=>"010001111",
  23344=>"100100010",
  23345=>"001000000",
  23346=>"000001001",
  23347=>"001110010",
  23348=>"010110101",
  23349=>"000011010",
  23350=>"111101001",
  23351=>"100100100",
  23352=>"000001011",
  23353=>"100000111",
  23354=>"101001101",
  23355=>"001011110",
  23356=>"001000100",
  23357=>"000100000",
  23358=>"011100110",
  23359=>"100110101",
  23360=>"101011001",
  23361=>"101011011",
  23362=>"100100000",
  23363=>"011011000",
  23364=>"101010001",
  23365=>"100111001",
  23366=>"111111000",
  23367=>"100000010",
  23368=>"000100010",
  23369=>"111111111",
  23370=>"010010100",
  23371=>"101001101",
  23372=>"101100011",
  23373=>"001011010",
  23374=>"000100000",
  23375=>"011000110",
  23376=>"000111000",
  23377=>"101010000",
  23378=>"111101000",
  23379=>"001110010",
  23380=>"001010101",
  23381=>"110001110",
  23382=>"000100110",
  23383=>"101101111",
  23384=>"101000101",
  23385=>"001111101",
  23386=>"011011010",
  23387=>"001100000",
  23388=>"011100111",
  23389=>"010000111",
  23390=>"110000100",
  23391=>"110001000",
  23392=>"000010100",
  23393=>"111111111",
  23394=>"011001110",
  23395=>"010101001",
  23396=>"001111010",
  23397=>"101010000",
  23398=>"010110111",
  23399=>"001011001",
  23400=>"111110101",
  23401=>"110100111",
  23402=>"110011101",
  23403=>"100011101",
  23404=>"101101010",
  23405=>"111011001",
  23406=>"000011101",
  23407=>"010110101",
  23408=>"010011000",
  23409=>"111010111",
  23410=>"110010000",
  23411=>"000100010",
  23412=>"000010001",
  23413=>"101110101",
  23414=>"110100101",
  23415=>"011111001",
  23416=>"100110111",
  23417=>"100100110",
  23418=>"100111001",
  23419=>"010010011",
  23420=>"000101011",
  23421=>"101111110",
  23422=>"011010011",
  23423=>"001001100",
  23424=>"001011101",
  23425=>"010101101",
  23426=>"001011110",
  23427=>"000011110",
  23428=>"001000001",
  23429=>"010011011",
  23430=>"100001000",
  23431=>"010100001",
  23432=>"110101101",
  23433=>"101000101",
  23434=>"111001011",
  23435=>"101111101",
  23436=>"100111100",
  23437=>"111101111",
  23438=>"000111111",
  23439=>"001000010",
  23440=>"000000000",
  23441=>"111111010",
  23442=>"100011011",
  23443=>"001110110",
  23444=>"111110101",
  23445=>"010000111",
  23446=>"011101110",
  23447=>"111011110",
  23448=>"010110001",
  23449=>"100110111",
  23450=>"011001001",
  23451=>"101001000",
  23452=>"100101001",
  23453=>"000010100",
  23454=>"111001000",
  23455=>"110111010",
  23456=>"010111111",
  23457=>"100000110",
  23458=>"111110100",
  23459=>"010110001",
  23460=>"000101100",
  23461=>"101111010",
  23462=>"011000000",
  23463=>"001001001",
  23464=>"110110010",
  23465=>"111110011",
  23466=>"111000101",
  23467=>"100010001",
  23468=>"101101100",
  23469=>"001001001",
  23470=>"011100010",
  23471=>"011000101",
  23472=>"010101000",
  23473=>"001010010",
  23474=>"101100000",
  23475=>"000110000",
  23476=>"111110011",
  23477=>"101111110",
  23478=>"101111011",
  23479=>"000101011",
  23480=>"010010100",
  23481=>"111100001",
  23482=>"000110101",
  23483=>"111101000",
  23484=>"000100101",
  23485=>"110111010",
  23486=>"110101000",
  23487=>"101010010",
  23488=>"111000001",
  23489=>"100001000",
  23490=>"111111111",
  23491=>"010100111",
  23492=>"001000111",
  23493=>"100111101",
  23494=>"000101000",
  23495=>"010110100",
  23496=>"011011001",
  23497=>"011010111",
  23498=>"001100101",
  23499=>"000100101",
  23500=>"000011001",
  23501=>"011101010",
  23502=>"010001011",
  23503=>"100011111",
  23504=>"010001111",
  23505=>"111101001",
  23506=>"010001010",
  23507=>"010100100",
  23508=>"111001101",
  23509=>"110011011",
  23510=>"001000011",
  23511=>"110101110",
  23512=>"110011001",
  23513=>"000001111",
  23514=>"001100010",
  23515=>"010001011",
  23516=>"001010111",
  23517=>"011110100",
  23518=>"010111010",
  23519=>"100111010",
  23520=>"101110111",
  23521=>"100100101",
  23522=>"100001010",
  23523=>"000110000",
  23524=>"010100000",
  23525=>"011110110",
  23526=>"010101010",
  23527=>"101100101",
  23528=>"000000000",
  23529=>"000001001",
  23530=>"001011000",
  23531=>"111011001",
  23532=>"100100011",
  23533=>"011100100",
  23534=>"110111001",
  23535=>"011101110",
  23536=>"000100100",
  23537=>"111100000",
  23538=>"011110000",
  23539=>"001000001",
  23540=>"111111110",
  23541=>"000000001",
  23542=>"011001000",
  23543=>"000001011",
  23544=>"010011101",
  23545=>"110111001",
  23546=>"100101101",
  23547=>"111110000",
  23548=>"110110110",
  23549=>"000001010",
  23550=>"111011101",
  23551=>"000010100",
  23552=>"001010111",
  23553=>"101110001",
  23554=>"100010110",
  23555=>"011011010",
  23556=>"101011100",
  23557=>"001010001",
  23558=>"000011000",
  23559=>"100010111",
  23560=>"011110011",
  23561=>"000111000",
  23562=>"100000010",
  23563=>"111001010",
  23564=>"000000000",
  23565=>"110001110",
  23566=>"010101111",
  23567=>"001101100",
  23568=>"011010011",
  23569=>"010010111",
  23570=>"101011001",
  23571=>"000001100",
  23572=>"011110101",
  23573=>"100011000",
  23574=>"110111011",
  23575=>"111001111",
  23576=>"100100000",
  23577=>"101100111",
  23578=>"011111111",
  23579=>"010101000",
  23580=>"000111011",
  23581=>"101000101",
  23582=>"011000101",
  23583=>"001110000",
  23584=>"101000100",
  23585=>"011111101",
  23586=>"011100101",
  23587=>"110100111",
  23588=>"110011011",
  23589=>"101011000",
  23590=>"011010001",
  23591=>"111111101",
  23592=>"100011010",
  23593=>"000110111",
  23594=>"001111100",
  23595=>"110101110",
  23596=>"110100001",
  23597=>"011011101",
  23598=>"101001010",
  23599=>"111011101",
  23600=>"010101100",
  23601=>"101001000",
  23602=>"011001010",
  23603=>"001000000",
  23604=>"001111101",
  23605=>"000001010",
  23606=>"111100001",
  23607=>"110000110",
  23608=>"101001110",
  23609=>"110110110",
  23610=>"001110100",
  23611=>"010010101",
  23612=>"101011110",
  23613=>"100000100",
  23614=>"100010001",
  23615=>"001101100",
  23616=>"000110111",
  23617=>"110101000",
  23618=>"000111111",
  23619=>"000100111",
  23620=>"001000111",
  23621=>"010101010",
  23622=>"100010001",
  23623=>"000011000",
  23624=>"011011110",
  23625=>"011100110",
  23626=>"001000111",
  23627=>"011101110",
  23628=>"100101100",
  23629=>"101001100",
  23630=>"101110001",
  23631=>"110010001",
  23632=>"110010110",
  23633=>"101000111",
  23634=>"000010011",
  23635=>"101001100",
  23636=>"100001101",
  23637=>"101111111",
  23638=>"001111101",
  23639=>"000000111",
  23640=>"001000011",
  23641=>"111010101",
  23642=>"110101110",
  23643=>"001000010",
  23644=>"010011000",
  23645=>"001011000",
  23646=>"100010110",
  23647=>"111011001",
  23648=>"100011111",
  23649=>"011111010",
  23650=>"000001011",
  23651=>"001010101",
  23652=>"100000100",
  23653=>"111010001",
  23654=>"010100100",
  23655=>"001111110",
  23656=>"110111011",
  23657=>"100101001",
  23658=>"110010111",
  23659=>"001111010",
  23660=>"000110101",
  23661=>"101111100",
  23662=>"010000110",
  23663=>"011101011",
  23664=>"010001000",
  23665=>"101010111",
  23666=>"011001010",
  23667=>"010100000",
  23668=>"110111010",
  23669=>"111010100",
  23670=>"000111000",
  23671=>"011111100",
  23672=>"000001101",
  23673=>"101000001",
  23674=>"000001010",
  23675=>"111110000",
  23676=>"110011100",
  23677=>"100100111",
  23678=>"110010111",
  23679=>"010011101",
  23680=>"001010101",
  23681=>"101011110",
  23682=>"111110001",
  23683=>"001110100",
  23684=>"110000010",
  23685=>"111011111",
  23686=>"011110110",
  23687=>"000101000",
  23688=>"111010110",
  23689=>"010010100",
  23690=>"010000111",
  23691=>"111101100",
  23692=>"010001100",
  23693=>"101101111",
  23694=>"111001000",
  23695=>"010101011",
  23696=>"000000001",
  23697=>"011010100",
  23698=>"111111011",
  23699=>"011011000",
  23700=>"010010011",
  23701=>"110001101",
  23702=>"000001100",
  23703=>"111001100",
  23704=>"110110110",
  23705=>"111001110",
  23706=>"011000110",
  23707=>"101000000",
  23708=>"001111100",
  23709=>"010000000",
  23710=>"100010111",
  23711=>"010011010",
  23712=>"101110101",
  23713=>"111000001",
  23714=>"111110100",
  23715=>"001100001",
  23716=>"111010011",
  23717=>"001001111",
  23718=>"111010011",
  23719=>"010101100",
  23720=>"001011011",
  23721=>"101110100",
  23722=>"100101100",
  23723=>"101001110",
  23724=>"110111000",
  23725=>"101101010",
  23726=>"101011011",
  23727=>"010100110",
  23728=>"001011101",
  23729=>"000001101",
  23730=>"110000111",
  23731=>"011001000",
  23732=>"101100000",
  23733=>"001101001",
  23734=>"001000111",
  23735=>"110110100",
  23736=>"111010110",
  23737=>"011011110",
  23738=>"011100101",
  23739=>"010111111",
  23740=>"100111011",
  23741=>"011000000",
  23742=>"011000101",
  23743=>"110010110",
  23744=>"001001111",
  23745=>"011101010",
  23746=>"000010001",
  23747=>"110101001",
  23748=>"101001001",
  23749=>"000011111",
  23750=>"101111011",
  23751=>"100110000",
  23752=>"101111011",
  23753=>"101011000",
  23754=>"110001101",
  23755=>"001101011",
  23756=>"011011111",
  23757=>"010101010",
  23758=>"000010001",
  23759=>"110100101",
  23760=>"010000001",
  23761=>"000110101",
  23762=>"110011100",
  23763=>"000100010",
  23764=>"010100110",
  23765=>"011100001",
  23766=>"000001010",
  23767=>"011011101",
  23768=>"000001001",
  23769=>"110110111",
  23770=>"110101011",
  23771=>"100010101",
  23772=>"100110100",
  23773=>"000110110",
  23774=>"010101111",
  23775=>"000011110",
  23776=>"011011001",
  23777=>"110001000",
  23778=>"001010010",
  23779=>"000100000",
  23780=>"010010110",
  23781=>"101111111",
  23782=>"010100101",
  23783=>"111111001",
  23784=>"010101010",
  23785=>"101001010",
  23786=>"100000000",
  23787=>"001010100",
  23788=>"000101101",
  23789=>"001000101",
  23790=>"011010001",
  23791=>"100011101",
  23792=>"011000010",
  23793=>"101000010",
  23794=>"010000001",
  23795=>"111001010",
  23796=>"011101001",
  23797=>"110110001",
  23798=>"111101111",
  23799=>"000011101",
  23800=>"110111011",
  23801=>"011100111",
  23802=>"000011010",
  23803=>"011011000",
  23804=>"001101100",
  23805=>"001100011",
  23806=>"101101100",
  23807=>"111100001",
  23808=>"000001000",
  23809=>"101110010",
  23810=>"011101111",
  23811=>"000010101",
  23812=>"001000010",
  23813=>"000101100",
  23814=>"111100111",
  23815=>"100010000",
  23816=>"000110011",
  23817=>"011001110",
  23818=>"011010000",
  23819=>"000001001",
  23820=>"001100111",
  23821=>"001000010",
  23822=>"110101110",
  23823=>"010001111",
  23824=>"010110111",
  23825=>"011000111",
  23826=>"000111001",
  23827=>"010101101",
  23828=>"010010001",
  23829=>"111001001",
  23830=>"101111101",
  23831=>"111001100",
  23832=>"011110011",
  23833=>"001001110",
  23834=>"111101111",
  23835=>"000100111",
  23836=>"000101001",
  23837=>"011100011",
  23838=>"010000000",
  23839=>"000011110",
  23840=>"011000110",
  23841=>"100010010",
  23842=>"100011110",
  23843=>"111101001",
  23844=>"111011000",
  23845=>"010010000",
  23846=>"010001001",
  23847=>"110001111",
  23848=>"111001110",
  23849=>"100010001",
  23850=>"010100011",
  23851=>"110001010",
  23852=>"101000101",
  23853=>"100111110",
  23854=>"011000100",
  23855=>"111101111",
  23856=>"000011011",
  23857=>"011010001",
  23858=>"100111111",
  23859=>"101011111",
  23860=>"100000101",
  23861=>"100100100",
  23862=>"011000101",
  23863=>"011001011",
  23864=>"111010000",
  23865=>"111101100",
  23866=>"110100001",
  23867=>"010111110",
  23868=>"000100111",
  23869=>"101101110",
  23870=>"101101100",
  23871=>"100001110",
  23872=>"100010000",
  23873=>"100001110",
  23874=>"011111111",
  23875=>"011010110",
  23876=>"001101101",
  23877=>"111101110",
  23878=>"001011100",
  23879=>"001000110",
  23880=>"010000101",
  23881=>"011000000",
  23882=>"101101101",
  23883=>"111000101",
  23884=>"010010000",
  23885=>"101111010",
  23886=>"111000010",
  23887=>"101010110",
  23888=>"110001101",
  23889=>"110111110",
  23890=>"111101011",
  23891=>"000111010",
  23892=>"011001010",
  23893=>"001000101",
  23894=>"000111100",
  23895=>"110000100",
  23896=>"011110001",
  23897=>"111100011",
  23898=>"110000110",
  23899=>"001010010",
  23900=>"010111100",
  23901=>"100101000",
  23902=>"000101011",
  23903=>"110111111",
  23904=>"111110100",
  23905=>"111001011",
  23906=>"101000000",
  23907=>"010111111",
  23908=>"101001101",
  23909=>"101011100",
  23910=>"100110100",
  23911=>"100001001",
  23912=>"110110110",
  23913=>"010000110",
  23914=>"011001111",
  23915=>"011111100",
  23916=>"110101010",
  23917=>"001110010",
  23918=>"101110100",
  23919=>"101110111",
  23920=>"110101100",
  23921=>"111110101",
  23922=>"110110010",
  23923=>"110001101",
  23924=>"001100010",
  23925=>"100100110",
  23926=>"101010001",
  23927=>"011100010",
  23928=>"001110010",
  23929=>"011000111",
  23930=>"010111101",
  23931=>"100110100",
  23932=>"110111110",
  23933=>"111101100",
  23934=>"011000000",
  23935=>"111101000",
  23936=>"100100111",
  23937=>"011100111",
  23938=>"001001101",
  23939=>"100010101",
  23940=>"100001001",
  23941=>"010111000",
  23942=>"110110010",
  23943=>"111011100",
  23944=>"100100000",
  23945=>"000000001",
  23946=>"101100110",
  23947=>"100100101",
  23948=>"101100110",
  23949=>"101011001",
  23950=>"100111110",
  23951=>"000111010",
  23952=>"111000111",
  23953=>"000011110",
  23954=>"000101111",
  23955=>"100111100",
  23956=>"111100101",
  23957=>"110011001",
  23958=>"011111001",
  23959=>"100101111",
  23960=>"011100000",
  23961=>"110010011",
  23962=>"010010010",
  23963=>"100111101",
  23964=>"010000110",
  23965=>"011101000",
  23966=>"001110111",
  23967=>"001001111",
  23968=>"111011011",
  23969=>"010000110",
  23970=>"001110100",
  23971=>"000010001",
  23972=>"001011000",
  23973=>"001101100",
  23974=>"111001010",
  23975=>"001001011",
  23976=>"011001000",
  23977=>"110010110",
  23978=>"000001110",
  23979=>"101000011",
  23980=>"111101010",
  23981=>"001111011",
  23982=>"111001110",
  23983=>"011111100",
  23984=>"001000001",
  23985=>"111000101",
  23986=>"100101100",
  23987=>"011111110",
  23988=>"111011000",
  23989=>"001111011",
  23990=>"111100100",
  23991=>"010100010",
  23992=>"010001010",
  23993=>"100010011",
  23994=>"101111001",
  23995=>"010000010",
  23996=>"010100000",
  23997=>"001000101",
  23998=>"000010110",
  23999=>"111011010",
  24000=>"010111011",
  24001=>"110001100",
  24002=>"110011011",
  24003=>"100010001",
  24004=>"000001001",
  24005=>"100000101",
  24006=>"001000011",
  24007=>"101001000",
  24008=>"011110110",
  24009=>"100111111",
  24010=>"000010000",
  24011=>"111011000",
  24012=>"000001110",
  24013=>"100111101",
  24014=>"001110000",
  24015=>"101001001",
  24016=>"111000011",
  24017=>"110000010",
  24018=>"100110010",
  24019=>"100110110",
  24020=>"100110100",
  24021=>"011001001",
  24022=>"111101000",
  24023=>"110110100",
  24024=>"000001110",
  24025=>"100010010",
  24026=>"101010010",
  24027=>"001010111",
  24028=>"111101011",
  24029=>"011110011",
  24030=>"110101010",
  24031=>"000001110",
  24032=>"000000111",
  24033=>"100110011",
  24034=>"100011111",
  24035=>"000010011",
  24036=>"011011101",
  24037=>"011101010",
  24038=>"100000110",
  24039=>"110101000",
  24040=>"001000101",
  24041=>"001111001",
  24042=>"111110100",
  24043=>"100010111",
  24044=>"001101001",
  24045=>"111101010",
  24046=>"100001000",
  24047=>"101001101",
  24048=>"111101101",
  24049=>"010001110",
  24050=>"011101001",
  24051=>"000100111",
  24052=>"010111001",
  24053=>"101000000",
  24054=>"001110110",
  24055=>"000011001",
  24056=>"110110111",
  24057=>"101000111",
  24058=>"010001100",
  24059=>"111010001",
  24060=>"111011011",
  24061=>"011111000",
  24062=>"101010010",
  24063=>"000000010",
  24064=>"111101000",
  24065=>"001000111",
  24066=>"010001110",
  24067=>"000010010",
  24068=>"110101100",
  24069=>"100000111",
  24070=>"000000000",
  24071=>"111110000",
  24072=>"001011110",
  24073=>"111011000",
  24074=>"111001101",
  24075=>"110010101",
  24076=>"101110010",
  24077=>"000001010",
  24078=>"111100111",
  24079=>"000110100",
  24080=>"011011101",
  24081=>"001101011",
  24082=>"011011011",
  24083=>"100110110",
  24084=>"000010100",
  24085=>"000111110",
  24086=>"101110111",
  24087=>"001010011",
  24088=>"111100001",
  24089=>"111011001",
  24090=>"000010011",
  24091=>"011111101",
  24092=>"011101111",
  24093=>"011100101",
  24094=>"011011101",
  24095=>"010011010",
  24096=>"011110101",
  24097=>"000111010",
  24098=>"110100000",
  24099=>"010011011",
  24100=>"000001000",
  24101=>"011000101",
  24102=>"010011011",
  24103=>"101101010",
  24104=>"100001111",
  24105=>"111010000",
  24106=>"000100001",
  24107=>"101111010",
  24108=>"011000000",
  24109=>"111111010",
  24110=>"000010110",
  24111=>"010011000",
  24112=>"001000100",
  24113=>"101111011",
  24114=>"000100110",
  24115=>"111100011",
  24116=>"001110111",
  24117=>"100111000",
  24118=>"101111110",
  24119=>"111001011",
  24120=>"001111100",
  24121=>"001011011",
  24122=>"000001110",
  24123=>"111000010",
  24124=>"010001011",
  24125=>"001100011",
  24126=>"100110101",
  24127=>"100000110",
  24128=>"100010001",
  24129=>"001100001",
  24130=>"101110001",
  24131=>"111101000",
  24132=>"001111100",
  24133=>"100101010",
  24134=>"101110010",
  24135=>"011001101",
  24136=>"011010000",
  24137=>"110000100",
  24138=>"100101000",
  24139=>"000110111",
  24140=>"111001100",
  24141=>"000110111",
  24142=>"100100101",
  24143=>"110110101",
  24144=>"011100110",
  24145=>"011100100",
  24146=>"001001110",
  24147=>"100011101",
  24148=>"011000001",
  24149=>"001101111",
  24150=>"001011010",
  24151=>"011011010",
  24152=>"000000111",
  24153=>"110100011",
  24154=>"001110111",
  24155=>"101101100",
  24156=>"100000011",
  24157=>"100001100",
  24158=>"100110001",
  24159=>"000001011",
  24160=>"111111110",
  24161=>"000101110",
  24162=>"001001111",
  24163=>"010010110",
  24164=>"000101011",
  24165=>"111100000",
  24166=>"010100110",
  24167=>"101111101",
  24168=>"001110011",
  24169=>"101001110",
  24170=>"110010100",
  24171=>"000000000",
  24172=>"101000010",
  24173=>"000000100",
  24174=>"011000111",
  24175=>"011110111",
  24176=>"010110100",
  24177=>"010000010",
  24178=>"111110101",
  24179=>"111100110",
  24180=>"110010110",
  24181=>"001110001",
  24182=>"010010100",
  24183=>"000001100",
  24184=>"100100100",
  24185=>"100110110",
  24186=>"011111010",
  24187=>"001001100",
  24188=>"110100000",
  24189=>"111101111",
  24190=>"000000010",
  24191=>"100000001",
  24192=>"101101111",
  24193=>"111110100",
  24194=>"001000000",
  24195=>"000001001",
  24196=>"101101100",
  24197=>"100101001",
  24198=>"111111010",
  24199=>"111011111",
  24200=>"100010110",
  24201=>"111001011",
  24202=>"100010101",
  24203=>"100101101",
  24204=>"000001001",
  24205=>"011111111",
  24206=>"011000110",
  24207=>"011110010",
  24208=>"011100110",
  24209=>"000011110",
  24210=>"001001000",
  24211=>"011111011",
  24212=>"100011010",
  24213=>"011011000",
  24214=>"001000010",
  24215=>"101011100",
  24216=>"010011000",
  24217=>"010010101",
  24218=>"001010101",
  24219=>"101000010",
  24220=>"110111000",
  24221=>"100000010",
  24222=>"011101110",
  24223=>"111101001",
  24224=>"101000010",
  24225=>"000001000",
  24226=>"011110001",
  24227=>"001100100",
  24228=>"110010101",
  24229=>"011111000",
  24230=>"110011001",
  24231=>"100010001",
  24232=>"110101111",
  24233=>"000001111",
  24234=>"000000110",
  24235=>"101100111",
  24236=>"100110100",
  24237=>"000001001",
  24238=>"010111111",
  24239=>"011100010",
  24240=>"000000000",
  24241=>"110100111",
  24242=>"001100100",
  24243=>"010000100",
  24244=>"111111101",
  24245=>"100101000",
  24246=>"100101111",
  24247=>"100111011",
  24248=>"010101000",
  24249=>"001011011",
  24250=>"100110101",
  24251=>"011000011",
  24252=>"101000100",
  24253=>"001100011",
  24254=>"000000010",
  24255=>"010011011",
  24256=>"000010011",
  24257=>"110000110",
  24258=>"001111111",
  24259=>"001010001",
  24260=>"111000111",
  24261=>"111011010",
  24262=>"110100001",
  24263=>"001001101",
  24264=>"110110101",
  24265=>"001001011",
  24266=>"100011010",
  24267=>"101000110",
  24268=>"010101100",
  24269=>"011001110",
  24270=>"010010111",
  24271=>"001000101",
  24272=>"100101010",
  24273=>"101111100",
  24274=>"000001111",
  24275=>"010100001",
  24276=>"011001001",
  24277=>"111101010",
  24278=>"101101101",
  24279=>"001011111",
  24280=>"110010001",
  24281=>"010000001",
  24282=>"110100111",
  24283=>"101000001",
  24284=>"110110110",
  24285=>"010000001",
  24286=>"110111001",
  24287=>"010001011",
  24288=>"010101001",
  24289=>"101001000",
  24290=>"001110011",
  24291=>"101111011",
  24292=>"100011001",
  24293=>"101010110",
  24294=>"010111011",
  24295=>"011111110",
  24296=>"000111111",
  24297=>"110110111",
  24298=>"110001110",
  24299=>"011101100",
  24300=>"110000110",
  24301=>"111101011",
  24302=>"001111001",
  24303=>"101011001",
  24304=>"001001010",
  24305=>"001000001",
  24306=>"000000011",
  24307=>"100000011",
  24308=>"100101011",
  24309=>"111100111",
  24310=>"110110011",
  24311=>"000110011",
  24312=>"101000010",
  24313=>"110111000",
  24314=>"110110100",
  24315=>"010000001",
  24316=>"011100001",
  24317=>"000001111",
  24318=>"111000101",
  24319=>"101110011",
  24320=>"011010100",
  24321=>"110011111",
  24322=>"000101110",
  24323=>"101110110",
  24324=>"110001010",
  24325=>"100101101",
  24326=>"011000011",
  24327=>"101100100",
  24328=>"000101100",
  24329=>"010010001",
  24330=>"011001101",
  24331=>"110001001",
  24332=>"011001110",
  24333=>"100001000",
  24334=>"000000011",
  24335=>"111111110",
  24336=>"010000001",
  24337=>"000001110",
  24338=>"010111100",
  24339=>"000111111",
  24340=>"101101110",
  24341=>"011111100",
  24342=>"101101011",
  24343=>"011111001",
  24344=>"011000010",
  24345=>"011101000",
  24346=>"000111100",
  24347=>"000011100",
  24348=>"011011100",
  24349=>"100010111",
  24350=>"000001100",
  24351=>"100101100",
  24352=>"000101001",
  24353=>"010011001",
  24354=>"100110010",
  24355=>"000111010",
  24356=>"010001101",
  24357=>"000000000",
  24358=>"000110110",
  24359=>"100001110",
  24360=>"100111010",
  24361=>"111001011",
  24362=>"101011000",
  24363=>"001010111",
  24364=>"010101011",
  24365=>"011011111",
  24366=>"000010000",
  24367=>"010111111",
  24368=>"011011111",
  24369=>"111000110",
  24370=>"010100111",
  24371=>"110000001",
  24372=>"111111000",
  24373=>"111001111",
  24374=>"111100010",
  24375=>"010010001",
  24376=>"110001011",
  24377=>"101000001",
  24378=>"000010111",
  24379=>"000010011",
  24380=>"111110001",
  24381=>"101000110",
  24382=>"010111010",
  24383=>"110010111",
  24384=>"000100001",
  24385=>"001000000",
  24386=>"011101001",
  24387=>"000001101",
  24388=>"110100101",
  24389=>"111100110",
  24390=>"111000011",
  24391=>"100101101",
  24392=>"011101101",
  24393=>"110010001",
  24394=>"011000000",
  24395=>"111101000",
  24396=>"010110001",
  24397=>"100111110",
  24398=>"010110000",
  24399=>"011010110",
  24400=>"100101011",
  24401=>"100010011",
  24402=>"100011101",
  24403=>"010000100",
  24404=>"100001101",
  24405=>"011110011",
  24406=>"111011100",
  24407=>"011110101",
  24408=>"100001001",
  24409=>"001100110",
  24410=>"000100011",
  24411=>"010100101",
  24412=>"101010010",
  24413=>"100110001",
  24414=>"001011000",
  24415=>"100011101",
  24416=>"110011000",
  24417=>"111100010",
  24418=>"000111011",
  24419=>"011101010",
  24420=>"111001011",
  24421=>"101011101",
  24422=>"100011000",
  24423=>"111110101",
  24424=>"111000100",
  24425=>"101110100",
  24426=>"101010111",
  24427=>"010001110",
  24428=>"101100010",
  24429=>"111111011",
  24430=>"101110110",
  24431=>"111110110",
  24432=>"100001110",
  24433=>"000101010",
  24434=>"011100010",
  24435=>"010111010",
  24436=>"000100100",
  24437=>"010001001",
  24438=>"001110001",
  24439=>"110011011",
  24440=>"001100010",
  24441=>"010001110",
  24442=>"011010100",
  24443=>"001110111",
  24444=>"011111011",
  24445=>"111101001",
  24446=>"111001000",
  24447=>"011001000",
  24448=>"000000110",
  24449=>"100001011",
  24450=>"111001111",
  24451=>"011100000",
  24452=>"000011010",
  24453=>"011110101",
  24454=>"000000000",
  24455=>"001111010",
  24456=>"100100000",
  24457=>"010100011",
  24458=>"011001110",
  24459=>"011111111",
  24460=>"000001010",
  24461=>"011100110",
  24462=>"000010001",
  24463=>"000000001",
  24464=>"000000001",
  24465=>"101001110",
  24466=>"011001111",
  24467=>"110111111",
  24468=>"010000110",
  24469=>"000110010",
  24470=>"001000011",
  24471=>"110010001",
  24472=>"101010001",
  24473=>"101101000",
  24474=>"011110000",
  24475=>"001001100",
  24476=>"000000100",
  24477=>"111111000",
  24478=>"100001111",
  24479=>"001110011",
  24480=>"001000111",
  24481=>"101100111",
  24482=>"110101100",
  24483=>"100110010",
  24484=>"000011011",
  24485=>"000101000",
  24486=>"000011100",
  24487=>"101010001",
  24488=>"000011111",
  24489=>"111010101",
  24490=>"111110000",
  24491=>"100101110",
  24492=>"101111000",
  24493=>"101110111",
  24494=>"111000010",
  24495=>"110000100",
  24496=>"111111101",
  24497=>"110001000",
  24498=>"010111111",
  24499=>"010101101",
  24500=>"111010001",
  24501=>"101011000",
  24502=>"001111101",
  24503=>"010000100",
  24504=>"001110111",
  24505=>"110001110",
  24506=>"111000001",
  24507=>"100001010",
  24508=>"010100000",
  24509=>"101111101",
  24510=>"110110101",
  24511=>"101111100",
  24512=>"111011001",
  24513=>"110110111",
  24514=>"000111111",
  24515=>"111110010",
  24516=>"001001000",
  24517=>"010010110",
  24518=>"000011000",
  24519=>"110000000",
  24520=>"010100110",
  24521=>"001000000",
  24522=>"010101110",
  24523=>"110010110",
  24524=>"000010001",
  24525=>"010000111",
  24526=>"110110000",
  24527=>"010100000",
  24528=>"101000100",
  24529=>"100101001",
  24530=>"100100111",
  24531=>"100101100",
  24532=>"101001010",
  24533=>"000110011",
  24534=>"110101101",
  24535=>"000001000",
  24536=>"110010001",
  24537=>"111100011",
  24538=>"111110000",
  24539=>"001000001",
  24540=>"111100001",
  24541=>"101100010",
  24542=>"110111111",
  24543=>"100010001",
  24544=>"011011111",
  24545=>"101110011",
  24546=>"101011111",
  24547=>"100001111",
  24548=>"100011111",
  24549=>"111001011",
  24550=>"111111101",
  24551=>"010101011",
  24552=>"000001110",
  24553=>"111011100",
  24554=>"000000101",
  24555=>"010101111",
  24556=>"110100101",
  24557=>"001101010",
  24558=>"001010000",
  24559=>"001110011",
  24560=>"001100100",
  24561=>"100100011",
  24562=>"100000101",
  24563=>"100010111",
  24564=>"001011010",
  24565=>"100100111",
  24566=>"111100101",
  24567=>"000001001",
  24568=>"001100110",
  24569=>"011101010",
  24570=>"110100011",
  24571=>"011100111",
  24572=>"100000000",
  24573=>"110100111",
  24574=>"000000100",
  24575=>"001110001",
  24576=>"001100010",
  24577=>"100011001",
  24578=>"110100110",
  24579=>"000111111",
  24580=>"000111011",
  24581=>"001111011",
  24582=>"011000101",
  24583=>"011101010",
  24584=>"001100101",
  24585=>"101001010",
  24586=>"000000101",
  24587=>"110110111",
  24588=>"111101010",
  24589=>"000110101",
  24590=>"101110101",
  24591=>"000111011",
  24592=>"101001001",
  24593=>"111001111",
  24594=>"011111011",
  24595=>"000001100",
  24596=>"100010010",
  24597=>"110011011",
  24598=>"110101011",
  24599=>"101101010",
  24600=>"010111001",
  24601=>"100000010",
  24602=>"100011010",
  24603=>"001111001",
  24604=>"001100101",
  24605=>"111011000",
  24606=>"101000011",
  24607=>"100100110",
  24608=>"101000101",
  24609=>"011010110",
  24610=>"110110100",
  24611=>"001010100",
  24612=>"001110101",
  24613=>"111000100",
  24614=>"111011001",
  24615=>"011100001",
  24616=>"110111001",
  24617=>"010111001",
  24618=>"111001011",
  24619=>"001011001",
  24620=>"110100111",
  24621=>"000011101",
  24622=>"000011011",
  24623=>"000111011",
  24624=>"001011011",
  24625=>"101000111",
  24626=>"011011010",
  24627=>"011110111",
  24628=>"001010000",
  24629=>"001111010",
  24630=>"100000000",
  24631=>"010110110",
  24632=>"110011010",
  24633=>"101010100",
  24634=>"100100001",
  24635=>"000000101",
  24636=>"011011011",
  24637=>"001101010",
  24638=>"110101011",
  24639=>"000000100",
  24640=>"000000110",
  24641=>"000100110",
  24642=>"011000101",
  24643=>"101010010",
  24644=>"010101111",
  24645=>"001011011",
  24646=>"010001001",
  24647=>"101010011",
  24648=>"100101010",
  24649=>"110101010",
  24650=>"111110011",
  24651=>"010111000",
  24652=>"110010001",
  24653=>"010100011",
  24654=>"010101001",
  24655=>"000011000",
  24656=>"101010000",
  24657=>"000101000",
  24658=>"110100110",
  24659=>"100001100",
  24660=>"011101100",
  24661=>"101011101",
  24662=>"100011011",
  24663=>"011011000",
  24664=>"000110010",
  24665=>"101110101",
  24666=>"111111101",
  24667=>"100101010",
  24668=>"001111011",
  24669=>"001000011",
  24670=>"111100000",
  24671=>"101100110",
  24672=>"000100110",
  24673=>"010011000",
  24674=>"010001010",
  24675=>"100010011",
  24676=>"000010111",
  24677=>"000101111",
  24678=>"000111111",
  24679=>"110101110",
  24680=>"101111100",
  24681=>"001110000",
  24682=>"001101111",
  24683=>"110011001",
  24684=>"101101100",
  24685=>"011110100",
  24686=>"000001010",
  24687=>"011001000",
  24688=>"001100001",
  24689=>"100011011",
  24690=>"001100011",
  24691=>"000110010",
  24692=>"000000100",
  24693=>"011011100",
  24694=>"000010000",
  24695=>"001000100",
  24696=>"011001110",
  24697=>"100111011",
  24698=>"010011101",
  24699=>"010110010",
  24700=>"010000101",
  24701=>"101010011",
  24702=>"010010000",
  24703=>"101001001",
  24704=>"100100000",
  24705=>"001000000",
  24706=>"010100111",
  24707=>"000000001",
  24708=>"001001011",
  24709=>"110000111",
  24710=>"000100011",
  24711=>"110101010",
  24712=>"110111011",
  24713=>"000100001",
  24714=>"000000111",
  24715=>"010010111",
  24716=>"111110101",
  24717=>"001110001",
  24718=>"110010001",
  24719=>"010011100",
  24720=>"011100101",
  24721=>"010101001",
  24722=>"000111011",
  24723=>"111011111",
  24724=>"001110000",
  24725=>"001101101",
  24726=>"001001100",
  24727=>"100101100",
  24728=>"101100001",
  24729=>"011000010",
  24730=>"111001111",
  24731=>"001011010",
  24732=>"000100101",
  24733=>"011000000",
  24734=>"100000010",
  24735=>"011011010",
  24736=>"111010100",
  24737=>"001010100",
  24738=>"110011101",
  24739=>"100111110",
  24740=>"111001011",
  24741=>"000101000",
  24742=>"001011111",
  24743=>"100000110",
  24744=>"011110100",
  24745=>"111001110",
  24746=>"100011011",
  24747=>"010111111",
  24748=>"110110010",
  24749=>"111001101",
  24750=>"001010000",
  24751=>"010000000",
  24752=>"000001001",
  24753=>"001000101",
  24754=>"011111010",
  24755=>"000101111",
  24756=>"100010001",
  24757=>"001111111",
  24758=>"000100111",
  24759=>"000000111",
  24760=>"011001010",
  24761=>"001001100",
  24762=>"001110001",
  24763=>"110110000",
  24764=>"010110001",
  24765=>"000101001",
  24766=>"111011100",
  24767=>"111001001",
  24768=>"110000110",
  24769=>"101010101",
  24770=>"111111111",
  24771=>"010001010",
  24772=>"111110001",
  24773=>"101000000",
  24774=>"111101101",
  24775=>"101111000",
  24776=>"011001010",
  24777=>"111010001",
  24778=>"101101010",
  24779=>"101011111",
  24780=>"100100101",
  24781=>"101100001",
  24782=>"110010011",
  24783=>"111001101",
  24784=>"110011000",
  24785=>"100000000",
  24786=>"111100011",
  24787=>"001111000",
  24788=>"101101110",
  24789=>"011000010",
  24790=>"101000101",
  24791=>"100111110",
  24792=>"101110010",
  24793=>"100110100",
  24794=>"100111011",
  24795=>"001011101",
  24796=>"110101101",
  24797=>"001101001",
  24798=>"100000000",
  24799=>"111111000",
  24800=>"101001000",
  24801=>"001100111",
  24802=>"011011000",
  24803=>"101010100",
  24804=>"111111000",
  24805=>"001000011",
  24806=>"110010010",
  24807=>"001110011",
  24808=>"000010011",
  24809=>"001010101",
  24810=>"101101001",
  24811=>"011011100",
  24812=>"000010101",
  24813=>"110100000",
  24814=>"001010101",
  24815=>"011001001",
  24816=>"110111100",
  24817=>"011110101",
  24818=>"001010000",
  24819=>"011100111",
  24820=>"110011111",
  24821=>"001010101",
  24822=>"001100000",
  24823=>"000010001",
  24824=>"010001011",
  24825=>"000110111",
  24826=>"111100001",
  24827=>"001011101",
  24828=>"111110111",
  24829=>"111010001",
  24830=>"001001000",
  24831=>"101100010",
  24832=>"011001100",
  24833=>"000100101",
  24834=>"010101001",
  24835=>"000010000",
  24836=>"101001001",
  24837=>"110000001",
  24838=>"101011100",
  24839=>"111011111",
  24840=>"110111110",
  24841=>"000001000",
  24842=>"100000100",
  24843=>"000000011",
  24844=>"011010100",
  24845=>"001011110",
  24846=>"101001101",
  24847=>"010000110",
  24848=>"000000111",
  24849=>"101000100",
  24850=>"101000001",
  24851=>"000001111",
  24852=>"000001011",
  24853=>"000100011",
  24854=>"111100111",
  24855=>"010011001",
  24856=>"000110100",
  24857=>"110010100",
  24858=>"111001000",
  24859=>"110110000",
  24860=>"001100110",
  24861=>"110000110",
  24862=>"101110011",
  24863=>"010100010",
  24864=>"011011011",
  24865=>"010100000",
  24866=>"101101000",
  24867=>"010111111",
  24868=>"101010001",
  24869=>"111111101",
  24870=>"001111100",
  24871=>"100010011",
  24872=>"101011010",
  24873=>"110001010",
  24874=>"101011001",
  24875=>"010000010",
  24876=>"101110000",
  24877=>"100011111",
  24878=>"101010101",
  24879=>"001001001",
  24880=>"011000000",
  24881=>"000100001",
  24882=>"100111001",
  24883=>"100111101",
  24884=>"100101100",
  24885=>"001000011",
  24886=>"001010000",
  24887=>"000111111",
  24888=>"001000111",
  24889=>"001001001",
  24890=>"000100100",
  24891=>"011110111",
  24892=>"010010100",
  24893=>"100010010",
  24894=>"100011101",
  24895=>"000010111",
  24896=>"110001001",
  24897=>"000101000",
  24898=>"101010001",
  24899=>"011010011",
  24900=>"001010101",
  24901=>"001100010",
  24902=>"010000111",
  24903=>"011100001",
  24904=>"011100111",
  24905=>"000001101",
  24906=>"001010101",
  24907=>"100110001",
  24908=>"101011000",
  24909=>"101100001",
  24910=>"001101110",
  24911=>"001110010",
  24912=>"101001110",
  24913=>"000101000",
  24914=>"001100110",
  24915=>"000011111",
  24916=>"110111001",
  24917=>"111101110",
  24918=>"000100100",
  24919=>"100111000",
  24920=>"001001001",
  24921=>"111000010",
  24922=>"001011001",
  24923=>"011110101",
  24924=>"101000000",
  24925=>"111000100",
  24926=>"100000000",
  24927=>"010111101",
  24928=>"100000000",
  24929=>"101111010",
  24930=>"110000101",
  24931=>"011010100",
  24932=>"101111010",
  24933=>"011001011",
  24934=>"001111010",
  24935=>"100101111",
  24936=>"000000000",
  24937=>"101110101",
  24938=>"011101001",
  24939=>"110001111",
  24940=>"111011010",
  24941=>"001010110",
  24942=>"110110000",
  24943=>"100110000",
  24944=>"011001000",
  24945=>"100111001",
  24946=>"111001011",
  24947=>"110111101",
  24948=>"000100110",
  24949=>"101010011",
  24950=>"001110000",
  24951=>"101100010",
  24952=>"010101010",
  24953=>"111000111",
  24954=>"000101010",
  24955=>"100011110",
  24956=>"011011011",
  24957=>"111101111",
  24958=>"001110111",
  24959=>"000010101",
  24960=>"101011101",
  24961=>"111101111",
  24962=>"000001111",
  24963=>"101111101",
  24964=>"001011101",
  24965=>"000101001",
  24966=>"110011101",
  24967=>"111001000",
  24968=>"011000111",
  24969=>"011010000",
  24970=>"011111001",
  24971=>"000100111",
  24972=>"000110011",
  24973=>"000101011",
  24974=>"101010101",
  24975=>"100001110",
  24976=>"100100110",
  24977=>"111010001",
  24978=>"000111000",
  24979=>"100011011",
  24980=>"111011101",
  24981=>"101001001",
  24982=>"110110010",
  24983=>"111101110",
  24984=>"000111100",
  24985=>"111001100",
  24986=>"100010011",
  24987=>"100000100",
  24988=>"001010000",
  24989=>"000111001",
  24990=>"100010101",
  24991=>"010010000",
  24992=>"010100100",
  24993=>"000011101",
  24994=>"111110101",
  24995=>"100000110",
  24996=>"110010110",
  24997=>"111000010",
  24998=>"010010110",
  24999=>"100100111",
  25000=>"001000111",
  25001=>"111010001",
  25002=>"111101011",
  25003=>"010111111",
  25004=>"000000100",
  25005=>"110100000",
  25006=>"100001101",
  25007=>"010000100",
  25008=>"101000011",
  25009=>"100111101",
  25010=>"100111101",
  25011=>"010110110",
  25012=>"100100101",
  25013=>"001101110",
  25014=>"110010011",
  25015=>"111101100",
  25016=>"001101111",
  25017=>"111100000",
  25018=>"011000011",
  25019=>"111011110",
  25020=>"110101001",
  25021=>"010111000",
  25022=>"101001010",
  25023=>"100011010",
  25024=>"010101001",
  25025=>"010000011",
  25026=>"101001101",
  25027=>"110111111",
  25028=>"101000000",
  25029=>"111011001",
  25030=>"010100001",
  25031=>"001011000",
  25032=>"111011100",
  25033=>"100110011",
  25034=>"011011111",
  25035=>"001011000",
  25036=>"101001111",
  25037=>"111111011",
  25038=>"011101101",
  25039=>"100000100",
  25040=>"110110101",
  25041=>"011001100",
  25042=>"110110111",
  25043=>"001110011",
  25044=>"010001111",
  25045=>"111111101",
  25046=>"000101001",
  25047=>"111010011",
  25048=>"111001000",
  25049=>"111001100",
  25050=>"011101010",
  25051=>"001010000",
  25052=>"001010101",
  25053=>"011010100",
  25054=>"110001111",
  25055=>"101001111",
  25056=>"101010000",
  25057=>"100001110",
  25058=>"010000111",
  25059=>"100000000",
  25060=>"111010010",
  25061=>"100010001",
  25062=>"010100000",
  25063=>"111101111",
  25064=>"110011011",
  25065=>"011101101",
  25066=>"100110110",
  25067=>"001101000",
  25068=>"001101111",
  25069=>"001111010",
  25070=>"100010111",
  25071=>"011110010",
  25072=>"101101001",
  25073=>"010100000",
  25074=>"101011001",
  25075=>"000101111",
  25076=>"100001000",
  25077=>"111001011",
  25078=>"111000101",
  25079=>"001010101",
  25080=>"110111010",
  25081=>"111001010",
  25082=>"011001011",
  25083=>"011010011",
  25084=>"111010101",
  25085=>"101111101",
  25086=>"001110110",
  25087=>"011010100",
  25088=>"010111001",
  25089=>"010001100",
  25090=>"000000100",
  25091=>"000000101",
  25092=>"110110110",
  25093=>"011111111",
  25094=>"100110101",
  25095=>"111111100",
  25096=>"110011001",
  25097=>"100111000",
  25098=>"100000011",
  25099=>"001010100",
  25100=>"101000111",
  25101=>"010111000",
  25102=>"000001000",
  25103=>"111001111",
  25104=>"101111010",
  25105=>"010001001",
  25106=>"000010001",
  25107=>"111110111",
  25108=>"011000000",
  25109=>"010111001",
  25110=>"101001111",
  25111=>"100100010",
  25112=>"000010101",
  25113=>"100111101",
  25114=>"001001011",
  25115=>"110001010",
  25116=>"111111000",
  25117=>"011001111",
  25118=>"111011111",
  25119=>"001100011",
  25120=>"111001110",
  25121=>"111011110",
  25122=>"001100010",
  25123=>"110010010",
  25124=>"010000101",
  25125=>"010110111",
  25126=>"100010001",
  25127=>"111110010",
  25128=>"011111001",
  25129=>"110011001",
  25130=>"111110111",
  25131=>"101011010",
  25132=>"010000010",
  25133=>"000010000",
  25134=>"010010101",
  25135=>"000010101",
  25136=>"100111000",
  25137=>"101011111",
  25138=>"111101011",
  25139=>"101000101",
  25140=>"001010010",
  25141=>"000001000",
  25142=>"001000000",
  25143=>"000000010",
  25144=>"100100111",
  25145=>"110001111",
  25146=>"100110001",
  25147=>"100111111",
  25148=>"010010011",
  25149=>"101100100",
  25150=>"010010010",
  25151=>"010111000",
  25152=>"000001011",
  25153=>"011000000",
  25154=>"101010000",
  25155=>"011100100",
  25156=>"100010010",
  25157=>"000101000",
  25158=>"011010000",
  25159=>"011001100",
  25160=>"110111011",
  25161=>"100001111",
  25162=>"111010100",
  25163=>"101000100",
  25164=>"101111111",
  25165=>"101110011",
  25166=>"111011011",
  25167=>"001101111",
  25168=>"111111000",
  25169=>"010000001",
  25170=>"111101011",
  25171=>"000011010",
  25172=>"000101110",
  25173=>"101000110",
  25174=>"000111010",
  25175=>"111000111",
  25176=>"011011111",
  25177=>"010011010",
  25178=>"111011001",
  25179=>"111101101",
  25180=>"001000111",
  25181=>"010000011",
  25182=>"100101101",
  25183=>"010000111",
  25184=>"001110110",
  25185=>"010110111",
  25186=>"001001000",
  25187=>"101100010",
  25188=>"110100100",
  25189=>"101111110",
  25190=>"001101110",
  25191=>"100011100",
  25192=>"000110011",
  25193=>"101111001",
  25194=>"011111100",
  25195=>"011011100",
  25196=>"010001110",
  25197=>"111011000",
  25198=>"010000010",
  25199=>"110011010",
  25200=>"010001010",
  25201=>"100000111",
  25202=>"110000011",
  25203=>"001000110",
  25204=>"010011101",
  25205=>"111000111",
  25206=>"101101010",
  25207=>"110111001",
  25208=>"111111111",
  25209=>"101111010",
  25210=>"010001001",
  25211=>"110110011",
  25212=>"110110011",
  25213=>"111000011",
  25214=>"011001010",
  25215=>"010100010",
  25216=>"011011100",
  25217=>"101010010",
  25218=>"111100001",
  25219=>"100100000",
  25220=>"110111001",
  25221=>"111101100",
  25222=>"000110111",
  25223=>"011011011",
  25224=>"010111000",
  25225=>"000101010",
  25226=>"110011011",
  25227=>"000001010",
  25228=>"011001111",
  25229=>"011100111",
  25230=>"101100111",
  25231=>"010100101",
  25232=>"010000110",
  25233=>"000001101",
  25234=>"101110000",
  25235=>"111001111",
  25236=>"101001001",
  25237=>"000000111",
  25238=>"001110010",
  25239=>"001010001",
  25240=>"010001101",
  25241=>"111111000",
  25242=>"010101001",
  25243=>"111011101",
  25244=>"001011101",
  25245=>"101011101",
  25246=>"111000100",
  25247=>"110011110",
  25248=>"011110111",
  25249=>"110011111",
  25250=>"010001001",
  25251=>"011001000",
  25252=>"000111010",
  25253=>"111011001",
  25254=>"001011110",
  25255=>"010001100",
  25256=>"001110000",
  25257=>"110011110",
  25258=>"011011101",
  25259=>"010000111",
  25260=>"010001000",
  25261=>"100001011",
  25262=>"111101100",
  25263=>"001101101",
  25264=>"010010011",
  25265=>"010010010",
  25266=>"011011110",
  25267=>"010100101",
  25268=>"011000100",
  25269=>"101001110",
  25270=>"111100011",
  25271=>"001011101",
  25272=>"010110011",
  25273=>"010001010",
  25274=>"111000100",
  25275=>"100110101",
  25276=>"111100000",
  25277=>"001010110",
  25278=>"001000011",
  25279=>"100000000",
  25280=>"000111011",
  25281=>"010100101",
  25282=>"100111100",
  25283=>"000011111",
  25284=>"111001101",
  25285=>"111000100",
  25286=>"100100110",
  25287=>"001010001",
  25288=>"110000111",
  25289=>"010100110",
  25290=>"011110000",
  25291=>"000001110",
  25292=>"000111100",
  25293=>"000001100",
  25294=>"111111001",
  25295=>"001010111",
  25296=>"001001001",
  25297=>"111100010",
  25298=>"010001110",
  25299=>"001110111",
  25300=>"110011001",
  25301=>"011100100",
  25302=>"101000101",
  25303=>"010010010",
  25304=>"001110100",
  25305=>"001011001",
  25306=>"001001100",
  25307=>"010010011",
  25308=>"111010000",
  25309=>"110100100",
  25310=>"101101011",
  25311=>"111000110",
  25312=>"000001100",
  25313=>"011101101",
  25314=>"010100111",
  25315=>"101101110",
  25316=>"100000101",
  25317=>"010001100",
  25318=>"111101111",
  25319=>"011010011",
  25320=>"001011010",
  25321=>"010001000",
  25322=>"110011101",
  25323=>"010101101",
  25324=>"011000101",
  25325=>"001100100",
  25326=>"100000101",
  25327=>"100110000",
  25328=>"101110110",
  25329=>"001000100",
  25330=>"101100110",
  25331=>"100100010",
  25332=>"101100110",
  25333=>"101000110",
  25334=>"100100010",
  25335=>"100100111",
  25336=>"010101001",
  25337=>"010111101",
  25338=>"101010010",
  25339=>"000011100",
  25340=>"000110001",
  25341=>"111110001",
  25342=>"001000101",
  25343=>"110110110",
  25344=>"010010111",
  25345=>"001110100",
  25346=>"101111101",
  25347=>"000001110",
  25348=>"100000000",
  25349=>"100000011",
  25350=>"110000011",
  25351=>"100010001",
  25352=>"110110000",
  25353=>"000010000",
  25354=>"101001001",
  25355=>"000000111",
  25356=>"000001011",
  25357=>"111100100",
  25358=>"111000011",
  25359=>"011000111",
  25360=>"000110011",
  25361=>"000111000",
  25362=>"111011100",
  25363=>"011010111",
  25364=>"011100011",
  25365=>"100111100",
  25366=>"011000010",
  25367=>"001011111",
  25368=>"101101001",
  25369=>"111001111",
  25370=>"001111001",
  25371=>"000001101",
  25372=>"001011100",
  25373=>"111000110",
  25374=>"101001010",
  25375=>"100010000",
  25376=>"001110101",
  25377=>"111001010",
  25378=>"011000000",
  25379=>"101011010",
  25380=>"000100000",
  25381=>"000110111",
  25382=>"001111110",
  25383=>"101100000",
  25384=>"011001010",
  25385=>"010010100",
  25386=>"001110111",
  25387=>"100011111",
  25388=>"111000000",
  25389=>"101101101",
  25390=>"011101000",
  25391=>"100100001",
  25392=>"100001100",
  25393=>"110101000",
  25394=>"101110010",
  25395=>"110011101",
  25396=>"101001111",
  25397=>"011110001",
  25398=>"001101010",
  25399=>"111111100",
  25400=>"101011000",
  25401=>"011001110",
  25402=>"011111111",
  25403=>"010001010",
  25404=>"101011111",
  25405=>"111101110",
  25406=>"101011101",
  25407=>"111011011",
  25408=>"101000010",
  25409=>"100001111",
  25410=>"001001110",
  25411=>"001000011",
  25412=>"000111111",
  25413=>"100011011",
  25414=>"100111101",
  25415=>"101001101",
  25416=>"000011001",
  25417=>"010101101",
  25418=>"010111001",
  25419=>"110100101",
  25420=>"100010011",
  25421=>"011101011",
  25422=>"111110100",
  25423=>"100110101",
  25424=>"110001011",
  25425=>"101101110",
  25426=>"001000000",
  25427=>"000110010",
  25428=>"000001111",
  25429=>"000101000",
  25430=>"000001100",
  25431=>"100000000",
  25432=>"001100011",
  25433=>"101111000",
  25434=>"110001100",
  25435=>"101001000",
  25436=>"100011010",
  25437=>"010011100",
  25438=>"001000011",
  25439=>"100011000",
  25440=>"111010010",
  25441=>"111111010",
  25442=>"000111110",
  25443=>"011011011",
  25444=>"100101011",
  25445=>"101000001",
  25446=>"000101011",
  25447=>"010101110",
  25448=>"000000011",
  25449=>"010010000",
  25450=>"010001111",
  25451=>"011101101",
  25452=>"100011101",
  25453=>"010000000",
  25454=>"100111001",
  25455=>"110001011",
  25456=>"000111110",
  25457=>"001101110",
  25458=>"010011010",
  25459=>"010001011",
  25460=>"011111000",
  25461=>"111011010",
  25462=>"010111111",
  25463=>"001110101",
  25464=>"100011101",
  25465=>"001100101",
  25466=>"101111000",
  25467=>"011001011",
  25468=>"011101011",
  25469=>"011110101",
  25470=>"000010111",
  25471=>"000101111",
  25472=>"001000100",
  25473=>"110101100",
  25474=>"100111110",
  25475=>"011100100",
  25476=>"100100010",
  25477=>"111011000",
  25478=>"011010010",
  25479=>"000001101",
  25480=>"101010001",
  25481=>"011011101",
  25482=>"100010101",
  25483=>"010011101",
  25484=>"101000010",
  25485=>"100101001",
  25486=>"101001000",
  25487=>"001100100",
  25488=>"110011111",
  25489=>"100010101",
  25490=>"000011101",
  25491=>"100101100",
  25492=>"000110110",
  25493=>"011100000",
  25494=>"101101110",
  25495=>"001101100",
  25496=>"001001001",
  25497=>"001101000",
  25498=>"111101010",
  25499=>"100110101",
  25500=>"000011110",
  25501=>"100010100",
  25502=>"100101000",
  25503=>"010101001",
  25504=>"100101000",
  25505=>"001110110",
  25506=>"100100101",
  25507=>"101010010",
  25508=>"111001110",
  25509=>"010000101",
  25510=>"101001101",
  25511=>"000010000",
  25512=>"100001100",
  25513=>"010101001",
  25514=>"011001111",
  25515=>"011111101",
  25516=>"111101011",
  25517=>"100101010",
  25518=>"101001011",
  25519=>"100000010",
  25520=>"101110011",
  25521=>"101000011",
  25522=>"010101111",
  25523=>"111001001",
  25524=>"011011110",
  25525=>"110010110",
  25526=>"011011010",
  25527=>"011001100",
  25528=>"110101011",
  25529=>"000010011",
  25530=>"101111111",
  25531=>"001001000",
  25532=>"001001000",
  25533=>"110100011",
  25534=>"100101111",
  25535=>"001010111",
  25536=>"100010011",
  25537=>"010110110",
  25538=>"110100101",
  25539=>"000000000",
  25540=>"101111111",
  25541=>"010111110",
  25542=>"110111011",
  25543=>"111001100",
  25544=>"011000010",
  25545=>"001000000",
  25546=>"010100111",
  25547=>"001111001",
  25548=>"000101011",
  25549=>"100001101",
  25550=>"110001111",
  25551=>"011101000",
  25552=>"111101010",
  25553=>"100010100",
  25554=>"011101100",
  25555=>"101100101",
  25556=>"100111001",
  25557=>"001011000",
  25558=>"100011100",
  25559=>"000101101",
  25560=>"001010011",
  25561=>"110110001",
  25562=>"100101101",
  25563=>"110001001",
  25564=>"001001011",
  25565=>"111001100",
  25566=>"000011011",
  25567=>"101000010",
  25568=>"010110111",
  25569=>"001010110",
  25570=>"000010111",
  25571=>"011011110",
  25572=>"010011010",
  25573=>"000011010",
  25574=>"001110100",
  25575=>"111001000",
  25576=>"101010001",
  25577=>"110001111",
  25578=>"011000101",
  25579=>"000101111",
  25580=>"011010010",
  25581=>"000100111",
  25582=>"010100011",
  25583=>"110111001",
  25584=>"000111111",
  25585=>"000100000",
  25586=>"010001011",
  25587=>"001100101",
  25588=>"000001101",
  25589=>"100011110",
  25590=>"010010001",
  25591=>"000010101",
  25592=>"010011000",
  25593=>"010011111",
  25594=>"110101100",
  25595=>"110010111",
  25596=>"100000001",
  25597=>"100010110",
  25598=>"101000010",
  25599=>"011000100",
  25600=>"101011001",
  25601=>"110110110",
  25602=>"111000010",
  25603=>"000011010",
  25604=>"010100101",
  25605=>"111010110",
  25606=>"011000110",
  25607=>"001000001",
  25608=>"111110010",
  25609=>"110110100",
  25610=>"010000110",
  25611=>"000110110",
  25612=>"010101101",
  25613=>"100000000",
  25614=>"000000110",
  25615=>"001001001",
  25616=>"110000010",
  25617=>"011101010",
  25618=>"010110100",
  25619=>"000001011",
  25620=>"000101110",
  25621=>"001000100",
  25622=>"001111100",
  25623=>"100011011",
  25624=>"011001010",
  25625=>"111100011",
  25626=>"110010000",
  25627=>"000111011",
  25628=>"011100010",
  25629=>"111010100",
  25630=>"010011001",
  25631=>"111111001",
  25632=>"011100110",
  25633=>"100001010",
  25634=>"101111111",
  25635=>"100011110",
  25636=>"001011011",
  25637=>"000110000",
  25638=>"001100110",
  25639=>"101101101",
  25640=>"001101001",
  25641=>"110011011",
  25642=>"010101100",
  25643=>"011000111",
  25644=>"100100000",
  25645=>"001011101",
  25646=>"111101101",
  25647=>"101000110",
  25648=>"010011000",
  25649=>"111101000",
  25650=>"010011000",
  25651=>"000001111",
  25652=>"011111111",
  25653=>"001001111",
  25654=>"111011000",
  25655=>"001010011",
  25656=>"100001000",
  25657=>"001101100",
  25658=>"101110101",
  25659=>"101101001",
  25660=>"011110110",
  25661=>"010100100",
  25662=>"100110001",
  25663=>"011110000",
  25664=>"100111011",
  25665=>"001000011",
  25666=>"011010010",
  25667=>"111101001",
  25668=>"101011001",
  25669=>"111001011",
  25670=>"110110111",
  25671=>"011101111",
  25672=>"101100010",
  25673=>"001111001",
  25674=>"011101101",
  25675=>"010001101",
  25676=>"011011010",
  25677=>"111010011",
  25678=>"101010100",
  25679=>"000001001",
  25680=>"110110011",
  25681=>"111000010",
  25682=>"110100010",
  25683=>"011101000",
  25684=>"011000111",
  25685=>"011000100",
  25686=>"000101101",
  25687=>"011010011",
  25688=>"111101011",
  25689=>"100011000",
  25690=>"101100110",
  25691=>"011101101",
  25692=>"100101001",
  25693=>"001000011",
  25694=>"100100001",
  25695=>"011111011",
  25696=>"111010000",
  25697=>"101010100",
  25698=>"100000101",
  25699=>"010100000",
  25700=>"000011011",
  25701=>"000111010",
  25702=>"001000011",
  25703=>"100010111",
  25704=>"000000000",
  25705=>"101001111",
  25706=>"101101101",
  25707=>"001011100",
  25708=>"101011111",
  25709=>"111001001",
  25710=>"011000000",
  25711=>"011011101",
  25712=>"010010101",
  25713=>"111010001",
  25714=>"100101011",
  25715=>"111001111",
  25716=>"111001001",
  25717=>"111100100",
  25718=>"100001011",
  25719=>"001100010",
  25720=>"001101110",
  25721=>"110001010",
  25722=>"001000010",
  25723=>"110100111",
  25724=>"111101110",
  25725=>"000101011",
  25726=>"101010010",
  25727=>"010100011",
  25728=>"110000011",
  25729=>"100110010",
  25730=>"101101101",
  25731=>"000100100",
  25732=>"010110001",
  25733=>"111010100",
  25734=>"011011001",
  25735=>"110001001",
  25736=>"000000000",
  25737=>"001100101",
  25738=>"001001001",
  25739=>"011110000",
  25740=>"010011101",
  25741=>"111100001",
  25742=>"000001101",
  25743=>"010011100",
  25744=>"011111101",
  25745=>"001110011",
  25746=>"110001101",
  25747=>"011000000",
  25748=>"111101001",
  25749=>"101101111",
  25750=>"100001100",
  25751=>"100000100",
  25752=>"111001000",
  25753=>"101111101",
  25754=>"101110010",
  25755=>"001001100",
  25756=>"111111000",
  25757=>"100110111",
  25758=>"100000000",
  25759=>"101011111",
  25760=>"011011101",
  25761=>"110111000",
  25762=>"100100100",
  25763=>"101000010",
  25764=>"001101111",
  25765=>"001000100",
  25766=>"011011111",
  25767=>"011111001",
  25768=>"001111000",
  25769=>"111101000",
  25770=>"001011100",
  25771=>"110011010",
  25772=>"000010010",
  25773=>"100101011",
  25774=>"110001111",
  25775=>"101101011",
  25776=>"010101010",
  25777=>"001101101",
  25778=>"101111011",
  25779=>"000111010",
  25780=>"100100101",
  25781=>"000000010",
  25782=>"000100000",
  25783=>"001001000",
  25784=>"110001001",
  25785=>"101101001",
  25786=>"001000010",
  25787=>"010000100",
  25788=>"011111000",
  25789=>"010001010",
  25790=>"011110001",
  25791=>"010111010",
  25792=>"011010111",
  25793=>"001011101",
  25794=>"011111101",
  25795=>"111010101",
  25796=>"011110011",
  25797=>"011010101",
  25798=>"101111111",
  25799=>"111010001",
  25800=>"011101101",
  25801=>"100110111",
  25802=>"001110000",
  25803=>"100110111",
  25804=>"011110101",
  25805=>"100100000",
  25806=>"110101011",
  25807=>"101010001",
  25808=>"000001111",
  25809=>"101100001",
  25810=>"101010001",
  25811=>"010000000",
  25812=>"110110001",
  25813=>"011110100",
  25814=>"111100101",
  25815=>"000010011",
  25816=>"000000101",
  25817=>"010001110",
  25818=>"011111101",
  25819=>"110110001",
  25820=>"001000100",
  25821=>"100101011",
  25822=>"101010001",
  25823=>"100111101",
  25824=>"011100100",
  25825=>"100000110",
  25826=>"000101010",
  25827=>"001000101",
  25828=>"111010110",
  25829=>"011000010",
  25830=>"110001110",
  25831=>"000100111",
  25832=>"000110110",
  25833=>"000101110",
  25834=>"001010111",
  25835=>"100010110",
  25836=>"010010001",
  25837=>"100110100",
  25838=>"111100111",
  25839=>"001000111",
  25840=>"101000010",
  25841=>"100001011",
  25842=>"011011100",
  25843=>"100001001",
  25844=>"110110010",
  25845=>"111100001",
  25846=>"101010000",
  25847=>"111001110",
  25848=>"110010100",
  25849=>"111111111",
  25850=>"110011011",
  25851=>"111011000",
  25852=>"111111011",
  25853=>"111110011",
  25854=>"001110110",
  25855=>"010100110",
  25856=>"011111000",
  25857=>"010000101",
  25858=>"011101110",
  25859=>"011001111",
  25860=>"001101111",
  25861=>"101101111",
  25862=>"001011011",
  25863=>"010100100",
  25864=>"111000000",
  25865=>"000111100",
  25866=>"011111011",
  25867=>"100110000",
  25868=>"010011010",
  25869=>"101110100",
  25870=>"001000010",
  25871=>"100100001",
  25872=>"100001110",
  25873=>"110001001",
  25874=>"001001101",
  25875=>"100101101",
  25876=>"001000100",
  25877=>"000000011",
  25878=>"111110100",
  25879=>"011001111",
  25880=>"111100010",
  25881=>"111010001",
  25882=>"101101001",
  25883=>"011100101",
  25884=>"111111100",
  25885=>"011110110",
  25886=>"001000001",
  25887=>"000010000",
  25888=>"100001101",
  25889=>"010000101",
  25890=>"100110100",
  25891=>"001000100",
  25892=>"001111011",
  25893=>"100101110",
  25894=>"111110000",
  25895=>"111011000",
  25896=>"110100101",
  25897=>"010111011",
  25898=>"001111000",
  25899=>"001110111",
  25900=>"101011100",
  25901=>"111100010",
  25902=>"101100110",
  25903=>"101100011",
  25904=>"100001010",
  25905=>"001010101",
  25906=>"110011101",
  25907=>"110011011",
  25908=>"010000010",
  25909=>"000000011",
  25910=>"010111100",
  25911=>"010111000",
  25912=>"000001111",
  25913=>"000000010",
  25914=>"100001000",
  25915=>"011110101",
  25916=>"100000000",
  25917=>"001100111",
  25918=>"110010100",
  25919=>"100110111",
  25920=>"011100101",
  25921=>"110100101",
  25922=>"000000011",
  25923=>"100010100",
  25924=>"000100000",
  25925=>"011001000",
  25926=>"011001011",
  25927=>"100111100",
  25928=>"010010010",
  25929=>"100110111",
  25930=>"100011100",
  25931=>"111100111",
  25932=>"111010111",
  25933=>"100000000",
  25934=>"110001101",
  25935=>"111110111",
  25936=>"000101100",
  25937=>"010111110",
  25938=>"000000001",
  25939=>"101101101",
  25940=>"000001101",
  25941=>"100011010",
  25942=>"001011101",
  25943=>"101111100",
  25944=>"111000100",
  25945=>"111000110",
  25946=>"011111001",
  25947=>"001111001",
  25948=>"100100111",
  25949=>"101011110",
  25950=>"101001111",
  25951=>"000010101",
  25952=>"100101100",
  25953=>"000111011",
  25954=>"110100100",
  25955=>"111110010",
  25956=>"101111100",
  25957=>"000000110",
  25958=>"000000010",
  25959=>"110110111",
  25960=>"000000111",
  25961=>"000001100",
  25962=>"000100111",
  25963=>"010011001",
  25964=>"101101010",
  25965=>"111101111",
  25966=>"111010100",
  25967=>"000001100",
  25968=>"110001011",
  25969=>"011000010",
  25970=>"010101000",
  25971=>"100000000",
  25972=>"110111001",
  25973=>"101010000",
  25974=>"001010100",
  25975=>"100001011",
  25976=>"000100001",
  25977=>"101011111",
  25978=>"111010000",
  25979=>"010011011",
  25980=>"010001000",
  25981=>"000101100",
  25982=>"011011110",
  25983=>"011000001",
  25984=>"101101001",
  25985=>"100001010",
  25986=>"100010110",
  25987=>"011010111",
  25988=>"010011010",
  25989=>"010011110",
  25990=>"110000111",
  25991=>"001110100",
  25992=>"011011011",
  25993=>"101001000",
  25994=>"111110110",
  25995=>"000001010",
  25996=>"010111101",
  25997=>"001101101",
  25998=>"111011110",
  25999=>"001101101",
  26000=>"001010100",
  26001=>"111010111",
  26002=>"111110110",
  26003=>"101011001",
  26004=>"101011110",
  26005=>"011111101",
  26006=>"100011101",
  26007=>"111101101",
  26008=>"001100101",
  26009=>"010000100",
  26010=>"111011001",
  26011=>"010110000",
  26012=>"110010111",
  26013=>"010101000",
  26014=>"111110100",
  26015=>"110010111",
  26016=>"111110110",
  26017=>"110011100",
  26018=>"010111110",
  26019=>"110000010",
  26020=>"011101001",
  26021=>"101011111",
  26022=>"101001110",
  26023=>"000101100",
  26024=>"000001101",
  26025=>"101100000",
  26026=>"001011100",
  26027=>"110111011",
  26028=>"000101111",
  26029=>"111011101",
  26030=>"101011010",
  26031=>"011100111",
  26032=>"110110111",
  26033=>"100001001",
  26034=>"010110110",
  26035=>"110001110",
  26036=>"111110000",
  26037=>"001110000",
  26038=>"110110001",
  26039=>"101011010",
  26040=>"001101011",
  26041=>"100010111",
  26042=>"010000100",
  26043=>"001011110",
  26044=>"001000011",
  26045=>"000001010",
  26046=>"001000000",
  26047=>"000010010",
  26048=>"001100101",
  26049=>"111111000",
  26050=>"111011010",
  26051=>"000100100",
  26052=>"000110001",
  26053=>"000011010",
  26054=>"100000000",
  26055=>"001101011",
  26056=>"000000010",
  26057=>"011110111",
  26058=>"111000000",
  26059=>"100010001",
  26060=>"111111100",
  26061=>"101001011",
  26062=>"011010000",
  26063=>"110100001",
  26064=>"011000001",
  26065=>"111111101",
  26066=>"011011101",
  26067=>"110111000",
  26068=>"111011111",
  26069=>"111110100",
  26070=>"010011001",
  26071=>"010110001",
  26072=>"101010111",
  26073=>"001001010",
  26074=>"111000110",
  26075=>"101011100",
  26076=>"111100111",
  26077=>"010110110",
  26078=>"011001111",
  26079=>"010111101",
  26080=>"010100001",
  26081=>"101100101",
  26082=>"000011010",
  26083=>"101101000",
  26084=>"011011101",
  26085=>"011110100",
  26086=>"110101100",
  26087=>"001000000",
  26088=>"000111010",
  26089=>"110101000",
  26090=>"010100000",
  26091=>"110111111",
  26092=>"101000001",
  26093=>"110111000",
  26094=>"111100000",
  26095=>"110101000",
  26096=>"110111101",
  26097=>"110000101",
  26098=>"001011100",
  26099=>"011110100",
  26100=>"101100101",
  26101=>"000101110",
  26102=>"001000111",
  26103=>"010000010",
  26104=>"111111011",
  26105=>"001110010",
  26106=>"011011001",
  26107=>"101010110",
  26108=>"000011110",
  26109=>"101110110",
  26110=>"000001101",
  26111=>"011110111",
  26112=>"001011010",
  26113=>"100010110",
  26114=>"100000001",
  26115=>"010000110",
  26116=>"011110111",
  26117=>"010111100",
  26118=>"010111110",
  26119=>"011001011",
  26120=>"011111011",
  26121=>"110111111",
  26122=>"100011110",
  26123=>"100000100",
  26124=>"100001010",
  26125=>"110011010",
  26126=>"110110010",
  26127=>"011100100",
  26128=>"100000001",
  26129=>"111001000",
  26130=>"100111100",
  26131=>"000011100",
  26132=>"101101100",
  26133=>"010110011",
  26134=>"001010000",
  26135=>"000011111",
  26136=>"100111101",
  26137=>"011111111",
  26138=>"101110010",
  26139=>"111100000",
  26140=>"011011110",
  26141=>"110111110",
  26142=>"000101101",
  26143=>"101100010",
  26144=>"101000011",
  26145=>"110111111",
  26146=>"100010001",
  26147=>"111111110",
  26148=>"100011111",
  26149=>"010100110",
  26150=>"011011000",
  26151=>"010110101",
  26152=>"010011010",
  26153=>"111110010",
  26154=>"101011000",
  26155=>"000010011",
  26156=>"000101101",
  26157=>"000001010",
  26158=>"111011111",
  26159=>"100110010",
  26160=>"000111000",
  26161=>"001010100",
  26162=>"110001101",
  26163=>"011101100",
  26164=>"011011011",
  26165=>"111101010",
  26166=>"011111001",
  26167=>"011010000",
  26168=>"100010010",
  26169=>"100101000",
  26170=>"011111011",
  26171=>"011100010",
  26172=>"010000011",
  26173=>"010111001",
  26174=>"000111100",
  26175=>"101010000",
  26176=>"011001001",
  26177=>"001100101",
  26178=>"110110011",
  26179=>"111001110",
  26180=>"110011101",
  26181=>"001011111",
  26182=>"100010011",
  26183=>"000011011",
  26184=>"010010000",
  26185=>"111000101",
  26186=>"011011011",
  26187=>"001111001",
  26188=>"001100110",
  26189=>"111111001",
  26190=>"001111000",
  26191=>"010101111",
  26192=>"110000110",
  26193=>"010011110",
  26194=>"101000100",
  26195=>"010011111",
  26196=>"101110010",
  26197=>"111101010",
  26198=>"101011000",
  26199=>"001100001",
  26200=>"101110001",
  26201=>"010101010",
  26202=>"101001100",
  26203=>"010000100",
  26204=>"111111010",
  26205=>"111011000",
  26206=>"110001000",
  26207=>"100101001",
  26208=>"100100111",
  26209=>"111111010",
  26210=>"111001010",
  26211=>"001110010",
  26212=>"001000011",
  26213=>"011001110",
  26214=>"001100000",
  26215=>"001110000",
  26216=>"100100111",
  26217=>"000000001",
  26218=>"111100100",
  26219=>"000010001",
  26220=>"001001111",
  26221=>"001101110",
  26222=>"010010000",
  26223=>"111110010",
  26224=>"011100100",
  26225=>"110011001",
  26226=>"111001110",
  26227=>"101010101",
  26228=>"001010000",
  26229=>"010111110",
  26230=>"101100101",
  26231=>"101100001",
  26232=>"111111100",
  26233=>"011000001",
  26234=>"011111000",
  26235=>"101011101",
  26236=>"011110001",
  26237=>"101001110",
  26238=>"110101000",
  26239=>"001110000",
  26240=>"110100001",
  26241=>"001010111",
  26242=>"011111010",
  26243=>"010110110",
  26244=>"001001111",
  26245=>"100011001",
  26246=>"100100110",
  26247=>"110000001",
  26248=>"010111110",
  26249=>"101110010",
  26250=>"001111001",
  26251=>"101011100",
  26252=>"100110010",
  26253=>"001111111",
  26254=>"000101110",
  26255=>"001111101",
  26256=>"000000110",
  26257=>"101001011",
  26258=>"100011101",
  26259=>"101000001",
  26260=>"110000100",
  26261=>"110011110",
  26262=>"011101110",
  26263=>"110010011",
  26264=>"010100101",
  26265=>"011100000",
  26266=>"011100000",
  26267=>"000001010",
  26268=>"111000001",
  26269=>"111101100",
  26270=>"000001001",
  26271=>"011000011",
  26272=>"011001010",
  26273=>"100000011",
  26274=>"001010100",
  26275=>"001010001",
  26276=>"100001000",
  26277=>"100010000",
  26278=>"101111111",
  26279=>"101011100",
  26280=>"100101111",
  26281=>"010010111",
  26282=>"101001011",
  26283=>"100111010",
  26284=>"011011000",
  26285=>"000001101",
  26286=>"110011111",
  26287=>"111100100",
  26288=>"011100000",
  26289=>"101110000",
  26290=>"111110000",
  26291=>"011000000",
  26292=>"001000010",
  26293=>"100101011",
  26294=>"110001110",
  26295=>"010111101",
  26296=>"101111111",
  26297=>"100010010",
  26298=>"011000110",
  26299=>"000000110",
  26300=>"111011111",
  26301=>"101111101",
  26302=>"001010000",
  26303=>"100100111",
  26304=>"101010011",
  26305=>"111111110",
  26306=>"101011000",
  26307=>"100010101",
  26308=>"101100011",
  26309=>"100111110",
  26310=>"101011000",
  26311=>"001000110",
  26312=>"100000010",
  26313=>"110100010",
  26314=>"011101000",
  26315=>"100101111",
  26316=>"000010011",
  26317=>"111010011",
  26318=>"010011010",
  26319=>"100010111",
  26320=>"100100011",
  26321=>"111010110",
  26322=>"001011001",
  26323=>"111011001",
  26324=>"100101001",
  26325=>"010001011",
  26326=>"011111010",
  26327=>"111100110",
  26328=>"100100001",
  26329=>"100000011",
  26330=>"101010111",
  26331=>"001001010",
  26332=>"000011001",
  26333=>"101111001",
  26334=>"010001100",
  26335=>"110100101",
  26336=>"111110110",
  26337=>"110000100",
  26338=>"001011011",
  26339=>"000001100",
  26340=>"011011011",
  26341=>"000110100",
  26342=>"000011011",
  26343=>"011011110",
  26344=>"100011101",
  26345=>"001000111",
  26346=>"010010101",
  26347=>"001101010",
  26348=>"011110011",
  26349=>"110011111",
  26350=>"111101000",
  26351=>"000011010",
  26352=>"000011001",
  26353=>"010010001",
  26354=>"100111101",
  26355=>"110100100",
  26356=>"111100000",
  26357=>"000001000",
  26358=>"101010111",
  26359=>"000111011",
  26360=>"110110110",
  26361=>"110011100",
  26362=>"010101110",
  26363=>"111101110",
  26364=>"000000100",
  26365=>"010110110",
  26366=>"011011001",
  26367=>"111100100",
  26368=>"000000000",
  26369=>"010001000",
  26370=>"111111111",
  26371=>"010100011",
  26372=>"110100100",
  26373=>"000000101",
  26374=>"000010110",
  26375=>"011001010",
  26376=>"000000001",
  26377=>"011110000",
  26378=>"111001100",
  26379=>"011001101",
  26380=>"000100001",
  26381=>"110001110",
  26382=>"101111101",
  26383=>"010011110",
  26384=>"001001000",
  26385=>"001010111",
  26386=>"000011000",
  26387=>"111000100",
  26388=>"010010000",
  26389=>"011100101",
  26390=>"111011011",
  26391=>"000010101",
  26392=>"001001010",
  26393=>"110000010",
  26394=>"001010101",
  26395=>"111101100",
  26396=>"110111000",
  26397=>"011110010",
  26398=>"100011010",
  26399=>"000010001",
  26400=>"100011001",
  26401=>"100010100",
  26402=>"111111110",
  26403=>"110111110",
  26404=>"100111101",
  26405=>"000010101",
  26406=>"101111110",
  26407=>"000000011",
  26408=>"010100000",
  26409=>"000000101",
  26410=>"110011111",
  26411=>"101101101",
  26412=>"000010100",
  26413=>"110111101",
  26414=>"110000111",
  26415=>"110010100",
  26416=>"011001011",
  26417=>"010101111",
  26418=>"001100101",
  26419=>"010111011",
  26420=>"001011001",
  26421=>"111101001",
  26422=>"100011011",
  26423=>"001010011",
  26424=>"101111000",
  26425=>"010010001",
  26426=>"101001011",
  26427=>"000100110",
  26428=>"000001010",
  26429=>"101000100",
  26430=>"111010010",
  26431=>"111010101",
  26432=>"010100011",
  26433=>"000010011",
  26434=>"101101111",
  26435=>"101000001",
  26436=>"101010100",
  26437=>"110101001",
  26438=>"000100001",
  26439=>"101010111",
  26440=>"010010001",
  26441=>"111110011",
  26442=>"000110111",
  26443=>"111010101",
  26444=>"110110000",
  26445=>"111110111",
  26446=>"101110000",
  26447=>"111110001",
  26448=>"000001100",
  26449=>"001101111",
  26450=>"101000110",
  26451=>"000000000",
  26452=>"101101100",
  26453=>"110010110",
  26454=>"010000101",
  26455=>"000000010",
  26456=>"011010001",
  26457=>"011101001",
  26458=>"101000100",
  26459=>"010111011",
  26460=>"000000110",
  26461=>"001000101",
  26462=>"001001111",
  26463=>"100101101",
  26464=>"011101100",
  26465=>"101000001",
  26466=>"110111000",
  26467=>"001001101",
  26468=>"101011011",
  26469=>"000000001",
  26470=>"110010100",
  26471=>"010110110",
  26472=>"001010101",
  26473=>"100110010",
  26474=>"110100101",
  26475=>"011111010",
  26476=>"111101001",
  26477=>"011001011",
  26478=>"110001110",
  26479=>"100001110",
  26480=>"100001100",
  26481=>"011001011",
  26482=>"001101110",
  26483=>"001011100",
  26484=>"111101110",
  26485=>"001000100",
  26486=>"111101101",
  26487=>"111101100",
  26488=>"011001110",
  26489=>"100001110",
  26490=>"110001111",
  26491=>"001011000",
  26492=>"111010001",
  26493=>"011001100",
  26494=>"111000000",
  26495=>"110000000",
  26496=>"110011100",
  26497=>"110000000",
  26498=>"110111011",
  26499=>"010000011",
  26500=>"001011100",
  26501=>"111110111",
  26502=>"001011011",
  26503=>"000000010",
  26504=>"000001110",
  26505=>"011011111",
  26506=>"100111110",
  26507=>"000011111",
  26508=>"011110011",
  26509=>"011101000",
  26510=>"101001000",
  26511=>"111110100",
  26512=>"100111001",
  26513=>"100000100",
  26514=>"111101111",
  26515=>"100111110",
  26516=>"011111001",
  26517=>"110001011",
  26518=>"000101101",
  26519=>"110100001",
  26520=>"101101001",
  26521=>"111001100",
  26522=>"100110010",
  26523=>"010011011",
  26524=>"101100011",
  26525=>"001010110",
  26526=>"001101111",
  26527=>"011111111",
  26528=>"110001011",
  26529=>"000001011",
  26530=>"010011010",
  26531=>"111000111",
  26532=>"110001110",
  26533=>"000000110",
  26534=>"010110000",
  26535=>"101101010",
  26536=>"001110011",
  26537=>"000010001",
  26538=>"100110101",
  26539=>"111110101",
  26540=>"000001010",
  26541=>"010011010",
  26542=>"111000110",
  26543=>"001110001",
  26544=>"010000110",
  26545=>"011000111",
  26546=>"010011111",
  26547=>"111010100",
  26548=>"111011011",
  26549=>"100010110",
  26550=>"011011001",
  26551=>"111011010",
  26552=>"011000111",
  26553=>"001001110",
  26554=>"100010000",
  26555=>"101001010",
  26556=>"011010011",
  26557=>"110000010",
  26558=>"111111110",
  26559=>"101101110",
  26560=>"100000001",
  26561=>"111010110",
  26562=>"000010001",
  26563=>"111001101",
  26564=>"110110011",
  26565=>"111111001",
  26566=>"000001101",
  26567=>"110110001",
  26568=>"011001100",
  26569=>"101011101",
  26570=>"001011110",
  26571=>"111110101",
  26572=>"011110010",
  26573=>"110101010",
  26574=>"000100011",
  26575=>"010001011",
  26576=>"011010101",
  26577=>"010101011",
  26578=>"011001011",
  26579=>"000010000",
  26580=>"101010100",
  26581=>"111011010",
  26582=>"101100011",
  26583=>"101110001",
  26584=>"110000011",
  26585=>"110011101",
  26586=>"101100111",
  26587=>"000001110",
  26588=>"100000011",
  26589=>"100101111",
  26590=>"111100100",
  26591=>"101101010",
  26592=>"111111100",
  26593=>"101111011",
  26594=>"101001000",
  26595=>"001001011",
  26596=>"111111001",
  26597=>"000101100",
  26598=>"000110011",
  26599=>"011001011",
  26600=>"011110110",
  26601=>"111111111",
  26602=>"111001101",
  26603=>"110110010",
  26604=>"000101010",
  26605=>"011001000",
  26606=>"100010110",
  26607=>"100100100",
  26608=>"110111111",
  26609=>"110110011",
  26610=>"010000101",
  26611=>"000011110",
  26612=>"000000010",
  26613=>"110000101",
  26614=>"001000011",
  26615=>"101010100",
  26616=>"111001101",
  26617=>"100111111",
  26618=>"011011101",
  26619=>"011110011",
  26620=>"110011000",
  26621=>"111101111",
  26622=>"001001100",
  26623=>"000111011",
  26624=>"101111110",
  26625=>"011100001",
  26626=>"001110111",
  26627=>"111000110",
  26628=>"101011111",
  26629=>"100101011",
  26630=>"000011110",
  26631=>"110001010",
  26632=>"001001000",
  26633=>"111001011",
  26634=>"011001010",
  26635=>"000011001",
  26636=>"001000011",
  26637=>"010100011",
  26638=>"111001110",
  26639=>"011000111",
  26640=>"010010000",
  26641=>"101001111",
  26642=>"101011111",
  26643=>"000110010",
  26644=>"001110101",
  26645=>"000011110",
  26646=>"110011110",
  26647=>"111001111",
  26648=>"101111001",
  26649=>"000100010",
  26650=>"101011111",
  26651=>"011110100",
  26652=>"101011010",
  26653=>"010011011",
  26654=>"100101000",
  26655=>"010111111",
  26656=>"001101010",
  26657=>"111011101",
  26658=>"000011100",
  26659=>"010100101",
  26660=>"000001010",
  26661=>"000111001",
  26662=>"101101010",
  26663=>"000111101",
  26664=>"000011100",
  26665=>"100101000",
  26666=>"001100011",
  26667=>"100000100",
  26668=>"110001110",
  26669=>"100100000",
  26670=>"100111101",
  26671=>"000001100",
  26672=>"110100011",
  26673=>"100100010",
  26674=>"110101111",
  26675=>"111001001",
  26676=>"101001100",
  26677=>"001000001",
  26678=>"000111110",
  26679=>"000011010",
  26680=>"001000110",
  26681=>"011101001",
  26682=>"110100011",
  26683=>"111011110",
  26684=>"011001101",
  26685=>"000111110",
  26686=>"110111010",
  26687=>"011001011",
  26688=>"100110100",
  26689=>"000010010",
  26690=>"100101010",
  26691=>"111100100",
  26692=>"011011111",
  26693=>"010011101",
  26694=>"010011000",
  26695=>"000000001",
  26696=>"101010101",
  26697=>"110101100",
  26698=>"001100010",
  26699=>"010000010",
  26700=>"000000010",
  26701=>"101010010",
  26702=>"011101110",
  26703=>"011001101",
  26704=>"100101110",
  26705=>"110001010",
  26706=>"111101011",
  26707=>"001000110",
  26708=>"000101101",
  26709=>"101111101",
  26710=>"101001001",
  26711=>"001000000",
  26712=>"001011011",
  26713=>"110100011",
  26714=>"001010010",
  26715=>"001001101",
  26716=>"101000110",
  26717=>"000010011",
  26718=>"000110011",
  26719=>"110000100",
  26720=>"010000000",
  26721=>"101010101",
  26722=>"001100111",
  26723=>"010111101",
  26724=>"110101000",
  26725=>"101001100",
  26726=>"101010000",
  26727=>"101110000",
  26728=>"011101011",
  26729=>"001011110",
  26730=>"001011110",
  26731=>"001000010",
  26732=>"001000000",
  26733=>"000110000",
  26734=>"001101000",
  26735=>"111111100",
  26736=>"000001001",
  26737=>"111101000",
  26738=>"101100101",
  26739=>"100101111",
  26740=>"111001010",
  26741=>"010000001",
  26742=>"110000100",
  26743=>"111010010",
  26744=>"110111010",
  26745=>"100001110",
  26746=>"001001100",
  26747=>"110101101",
  26748=>"101111000",
  26749=>"101010010",
  26750=>"001100111",
  26751=>"001000111",
  26752=>"100111100",
  26753=>"110110000",
  26754=>"100011111",
  26755=>"110100010",
  26756=>"101111111",
  26757=>"001111001",
  26758=>"111001000",
  26759=>"101000111",
  26760=>"011110100",
  26761=>"110111000",
  26762=>"100111111",
  26763=>"111100101",
  26764=>"101010011",
  26765=>"010110101",
  26766=>"101001111",
  26767=>"111111011",
  26768=>"000000111",
  26769=>"100100100",
  26770=>"000100111",
  26771=>"001000000",
  26772=>"010100101",
  26773=>"000101010",
  26774=>"011101010",
  26775=>"110000111",
  26776=>"110000011",
  26777=>"011000100",
  26778=>"100001111",
  26779=>"011001001",
  26780=>"101011011",
  26781=>"110111111",
  26782=>"111101000",
  26783=>"010011110",
  26784=>"111101111",
  26785=>"011001111",
  26786=>"101100000",
  26787=>"000000001",
  26788=>"111100101",
  26789=>"000111010",
  26790=>"110011101",
  26791=>"110001000",
  26792=>"010101000",
  26793=>"001001011",
  26794=>"001010001",
  26795=>"010010110",
  26796=>"000000010",
  26797=>"011111111",
  26798=>"000000001",
  26799=>"010111000",
  26800=>"000101100",
  26801=>"111101000",
  26802=>"011001010",
  26803=>"100011010",
  26804=>"110010100",
  26805=>"110001101",
  26806=>"101010110",
  26807=>"011011010",
  26808=>"010011111",
  26809=>"100001110",
  26810=>"001011011",
  26811=>"010100010",
  26812=>"011111001",
  26813=>"001001000",
  26814=>"001001110",
  26815=>"111110111",
  26816=>"000010111",
  26817=>"101100110",
  26818=>"100100001",
  26819=>"011001000",
  26820=>"101010101",
  26821=>"100001011",
  26822=>"001011011",
  26823=>"011010011",
  26824=>"000001001",
  26825=>"011110101",
  26826=>"000100000",
  26827=>"101111111",
  26828=>"101001000",
  26829=>"010111010",
  26830=>"001101010",
  26831=>"010100101",
  26832=>"011110110",
  26833=>"111110110",
  26834=>"111000000",
  26835=>"101000011",
  26836=>"110111001",
  26837=>"001010011",
  26838=>"000100111",
  26839=>"100010101",
  26840=>"100000010",
  26841=>"100110000",
  26842=>"011100000",
  26843=>"111100110",
  26844=>"000000101",
  26845=>"100000101",
  26846=>"001101101",
  26847=>"011000000",
  26848=>"101001110",
  26849=>"110100101",
  26850=>"010000000",
  26851=>"101111011",
  26852=>"000000100",
  26853=>"011000001",
  26854=>"011000010",
  26855=>"000100001",
  26856=>"001101110",
  26857=>"011011111",
  26858=>"001101100",
  26859=>"001111100",
  26860=>"101000010",
  26861=>"000000100",
  26862=>"111101000",
  26863=>"011100111",
  26864=>"110100110",
  26865=>"011101011",
  26866=>"101001001",
  26867=>"000100010",
  26868=>"011110001",
  26869=>"001101010",
  26870=>"100001001",
  26871=>"000000001",
  26872=>"101000111",
  26873=>"101011101",
  26874=>"010101110",
  26875=>"001011101",
  26876=>"001111001",
  26877=>"110101001",
  26878=>"110000000",
  26879=>"111111001",
  26880=>"011111111",
  26881=>"001000110",
  26882=>"011001000",
  26883=>"110110111",
  26884=>"010100101",
  26885=>"000101110",
  26886=>"010110000",
  26887=>"011011111",
  26888=>"111011100",
  26889=>"001011100",
  26890=>"011011011",
  26891=>"100001010",
  26892=>"111110100",
  26893=>"111000000",
  26894=>"100111010",
  26895=>"011110111",
  26896=>"010000110",
  26897=>"010001001",
  26898=>"010111011",
  26899=>"100001110",
  26900=>"111110001",
  26901=>"101010011",
  26902=>"010100011",
  26903=>"110101110",
  26904=>"010110111",
  26905=>"001011110",
  26906=>"101100100",
  26907=>"010010111",
  26908=>"101100001",
  26909=>"100101110",
  26910=>"010100011",
  26911=>"000001010",
  26912=>"010110011",
  26913=>"111010111",
  26914=>"110111101",
  26915=>"000100000",
  26916=>"001101000",
  26917=>"110001101",
  26918=>"000100011",
  26919=>"110111101",
  26920=>"010101010",
  26921=>"011110010",
  26922=>"000010000",
  26923=>"001110011",
  26924=>"011110010",
  26925=>"010000000",
  26926=>"000101001",
  26927=>"000011101",
  26928=>"111000001",
  26929=>"001011101",
  26930=>"110111111",
  26931=>"101001101",
  26932=>"001010101",
  26933=>"010010001",
  26934=>"010100000",
  26935=>"000111110",
  26936=>"000100101",
  26937=>"010111110",
  26938=>"111001000",
  26939=>"011011000",
  26940=>"000000110",
  26941=>"101100010",
  26942=>"001101010",
  26943=>"110111111",
  26944=>"110101100",
  26945=>"001110011",
  26946=>"010010101",
  26947=>"000110110",
  26948=>"010111111",
  26949=>"101101100",
  26950=>"100101011",
  26951=>"011110110",
  26952=>"101001011",
  26953=>"010010001",
  26954=>"111010100",
  26955=>"001010101",
  26956=>"111110000",
  26957=>"100111010",
  26958=>"101001011",
  26959=>"110011100",
  26960=>"001001100",
  26961=>"000111100",
  26962=>"000011010",
  26963=>"000000011",
  26964=>"000110110",
  26965=>"010100111",
  26966=>"111011110",
  26967=>"111011100",
  26968=>"101011010",
  26969=>"111111011",
  26970=>"000000001",
  26971=>"010111111",
  26972=>"000110110",
  26973=>"101000111",
  26974=>"111101110",
  26975=>"001011111",
  26976=>"100111111",
  26977=>"000001001",
  26978=>"010101110",
  26979=>"101111110",
  26980=>"110111010",
  26981=>"110110010",
  26982=>"111101001",
  26983=>"111000000",
  26984=>"110010001",
  26985=>"000110010",
  26986=>"101001001",
  26987=>"110100101",
  26988=>"000000100",
  26989=>"110010000",
  26990=>"101010100",
  26991=>"111100111",
  26992=>"000100101",
  26993=>"011101011",
  26994=>"011101100",
  26995=>"100001001",
  26996=>"110000111",
  26997=>"100010001",
  26998=>"001010100",
  26999=>"000011111",
  27000=>"011111001",
  27001=>"010100110",
  27002=>"101011101",
  27003=>"011100010",
  27004=>"010100010",
  27005=>"011100111",
  27006=>"001001101",
  27007=>"011011001",
  27008=>"111101110",
  27009=>"111001000",
  27010=>"110011011",
  27011=>"100001111",
  27012=>"101110100",
  27013=>"100110000",
  27014=>"010111011",
  27015=>"001111001",
  27016=>"101011101",
  27017=>"000000100",
  27018=>"000010100",
  27019=>"001000110",
  27020=>"110110010",
  27021=>"001100100",
  27022=>"000110111",
  27023=>"110011001",
  27024=>"000110111",
  27025=>"000000001",
  27026=>"011110011",
  27027=>"100011010",
  27028=>"100001010",
  27029=>"000000011",
  27030=>"010001010",
  27031=>"001110111",
  27032=>"000011100",
  27033=>"011110000",
  27034=>"011111100",
  27035=>"111010001",
  27036=>"000101111",
  27037=>"001000101",
  27038=>"011000000",
  27039=>"110010000",
  27040=>"001100001",
  27041=>"101000111",
  27042=>"100001001",
  27043=>"000000000",
  27044=>"011001010",
  27045=>"000000000",
  27046=>"010010111",
  27047=>"100000111",
  27048=>"010101100",
  27049=>"100010100",
  27050=>"111110100",
  27051=>"111111101",
  27052=>"101000100",
  27053=>"011000011",
  27054=>"010100110",
  27055=>"011100111",
  27056=>"110110101",
  27057=>"000011000",
  27058=>"000100010",
  27059=>"100001011",
  27060=>"111010111",
  27061=>"010100001",
  27062=>"010011110",
  27063=>"101010010",
  27064=>"001001000",
  27065=>"000110011",
  27066=>"111101000",
  27067=>"110111100",
  27068=>"010111100",
  27069=>"000101101",
  27070=>"010101011",
  27071=>"110101011",
  27072=>"011110101",
  27073=>"101111111",
  27074=>"111100110",
  27075=>"000001100",
  27076=>"001011110",
  27077=>"101110001",
  27078=>"110001001",
  27079=>"000011111",
  27080=>"011001100",
  27081=>"001101000",
  27082=>"111111001",
  27083=>"110111000",
  27084=>"100111110",
  27085=>"000010110",
  27086=>"000110000",
  27087=>"100010011",
  27088=>"111101101",
  27089=>"000010111",
  27090=>"111110010",
  27091=>"110101001",
  27092=>"010000110",
  27093=>"100100001",
  27094=>"111101101",
  27095=>"011010000",
  27096=>"011010001",
  27097=>"000001010",
  27098=>"010101000",
  27099=>"101110100",
  27100=>"000111100",
  27101=>"111111111",
  27102=>"101011111",
  27103=>"111110110",
  27104=>"100100100",
  27105=>"100011101",
  27106=>"110100010",
  27107=>"100100111",
  27108=>"110010110",
  27109=>"010110011",
  27110=>"000110011",
  27111=>"000111111",
  27112=>"001000111",
  27113=>"100001101",
  27114=>"100100101",
  27115=>"001100010",
  27116=>"100000011",
  27117=>"001000101",
  27118=>"101101101",
  27119=>"110000000",
  27120=>"110110000",
  27121=>"011010010",
  27122=>"000101111",
  27123=>"000011000",
  27124=>"100000000",
  27125=>"010111110",
  27126=>"001001011",
  27127=>"000001011",
  27128=>"100111100",
  27129=>"001010000",
  27130=>"010011111",
  27131=>"010001110",
  27132=>"111100011",
  27133=>"011101101",
  27134=>"010101001",
  27135=>"101000100",
  27136=>"111101111",
  27137=>"000011001",
  27138=>"101101110",
  27139=>"001100100",
  27140=>"110001100",
  27141=>"111001100",
  27142=>"100101010",
  27143=>"010101100",
  27144=>"010001010",
  27145=>"110100001",
  27146=>"000000010",
  27147=>"001001100",
  27148=>"001111110",
  27149=>"000101001",
  27150=>"000101100",
  27151=>"111100111",
  27152=>"000001101",
  27153=>"001010010",
  27154=>"010000101",
  27155=>"101100111",
  27156=>"001110011",
  27157=>"101101110",
  27158=>"001001110",
  27159=>"001100000",
  27160=>"110000001",
  27161=>"110101001",
  27162=>"101100100",
  27163=>"111001001",
  27164=>"100000101",
  27165=>"001110110",
  27166=>"101010101",
  27167=>"110101110",
  27168=>"010110010",
  27169=>"000101101",
  27170=>"001000100",
  27171=>"000001110",
  27172=>"110110010",
  27173=>"011111000",
  27174=>"101001001",
  27175=>"011000000",
  27176=>"110011101",
  27177=>"011101101",
  27178=>"011010001",
  27179=>"110100110",
  27180=>"100010011",
  27181=>"000110011",
  27182=>"100111010",
  27183=>"011001110",
  27184=>"011110001",
  27185=>"011001001",
  27186=>"001000111",
  27187=>"101111100",
  27188=>"101100100",
  27189=>"111011001",
  27190=>"110101111",
  27191=>"000100001",
  27192=>"111101010",
  27193=>"110101011",
  27194=>"110100100",
  27195=>"100010011",
  27196=>"110111111",
  27197=>"011010001",
  27198=>"101000111",
  27199=>"101110010",
  27200=>"110111111",
  27201=>"000001001",
  27202=>"111011001",
  27203=>"100010011",
  27204=>"011100010",
  27205=>"101111011",
  27206=>"010000001",
  27207=>"111111111",
  27208=>"011101011",
  27209=>"010110111",
  27210=>"010001001",
  27211=>"100101011",
  27212=>"011111011",
  27213=>"100010101",
  27214=>"101111101",
  27215=>"001001100",
  27216=>"000010000",
  27217=>"011111111",
  27218=>"101000011",
  27219=>"111000010",
  27220=>"101010101",
  27221=>"011001000",
  27222=>"100011111",
  27223=>"001001100",
  27224=>"011001110",
  27225=>"100010000",
  27226=>"100001011",
  27227=>"000101001",
  27228=>"101011010",
  27229=>"100011000",
  27230=>"001110101",
  27231=>"101001011",
  27232=>"111110010",
  27233=>"001101000",
  27234=>"000111101",
  27235=>"101100011",
  27236=>"001110111",
  27237=>"001001101",
  27238=>"001001110",
  27239=>"111100001",
  27240=>"100100000",
  27241=>"000110101",
  27242=>"100111110",
  27243=>"000010000",
  27244=>"110111100",
  27245=>"000011111",
  27246=>"000100110",
  27247=>"001101100",
  27248=>"110110000",
  27249=>"111110111",
  27250=>"000111011",
  27251=>"000111010",
  27252=>"110110101",
  27253=>"100010010",
  27254=>"111101101",
  27255=>"000010110",
  27256=>"001100010",
  27257=>"111111000",
  27258=>"100111000",
  27259=>"010110111",
  27260=>"100110101",
  27261=>"011000100",
  27262=>"000110000",
  27263=>"110110100",
  27264=>"100000010",
  27265=>"111110001",
  27266=>"111111111",
  27267=>"000000101",
  27268=>"111000000",
  27269=>"011110011",
  27270=>"000011010",
  27271=>"110010010",
  27272=>"011110010",
  27273=>"011000101",
  27274=>"111110101",
  27275=>"000100111",
  27276=>"111001101",
  27277=>"000111111",
  27278=>"111100110",
  27279=>"010110110",
  27280=>"011010011",
  27281=>"101001111",
  27282=>"011010010",
  27283=>"111110100",
  27284=>"001000010",
  27285=>"100001010",
  27286=>"010111011",
  27287=>"101000100",
  27288=>"110001010",
  27289=>"100010100",
  27290=>"010100101",
  27291=>"100001010",
  27292=>"010010001",
  27293=>"101000001",
  27294=>"110011100",
  27295=>"001100010",
  27296=>"001011010",
  27297=>"001010011",
  27298=>"001010100",
  27299=>"101010100",
  27300=>"100110011",
  27301=>"000000010",
  27302=>"111100100",
  27303=>"010000000",
  27304=>"110000001",
  27305=>"011001010",
  27306=>"000010101",
  27307=>"010000000",
  27308=>"111000000",
  27309=>"010010101",
  27310=>"100111100",
  27311=>"111001101",
  27312=>"010101110",
  27313=>"011000010",
  27314=>"010011101",
  27315=>"010101110",
  27316=>"010101011",
  27317=>"111111000",
  27318=>"110110100",
  27319=>"101010001",
  27320=>"110001001",
  27321=>"101001010",
  27322=>"110000100",
  27323=>"111000010",
  27324=>"000010011",
  27325=>"101000011",
  27326=>"100111011",
  27327=>"101101001",
  27328=>"100101100",
  27329=>"111000000",
  27330=>"010000111",
  27331=>"100000111",
  27332=>"100001110",
  27333=>"000001111",
  27334=>"101000110",
  27335=>"010100011",
  27336=>"100001101",
  27337=>"110011001",
  27338=>"010101100",
  27339=>"101100011",
  27340=>"010101110",
  27341=>"100101111",
  27342=>"001101110",
  27343=>"101100111",
  27344=>"000000111",
  27345=>"111000100",
  27346=>"110111011",
  27347=>"011011101",
  27348=>"011100100",
  27349=>"001110011",
  27350=>"110001100",
  27351=>"101001011",
  27352=>"001010111",
  27353=>"001110001",
  27354=>"100000100",
  27355=>"000011110",
  27356=>"000110100",
  27357=>"010110110",
  27358=>"010001111",
  27359=>"101000001",
  27360=>"010000111",
  27361=>"011001000",
  27362=>"111110010",
  27363=>"101111101",
  27364=>"011001111",
  27365=>"110010101",
  27366=>"111101000",
  27367=>"000000000",
  27368=>"100100110",
  27369=>"101100011",
  27370=>"100111011",
  27371=>"000001111",
  27372=>"111101011",
  27373=>"110001100",
  27374=>"100100111",
  27375=>"110101111",
  27376=>"000000110",
  27377=>"001001110",
  27378=>"000000100",
  27379=>"010000000",
  27380=>"110100010",
  27381=>"000111100",
  27382=>"111100011",
  27383=>"111100111",
  27384=>"000111100",
  27385=>"001111010",
  27386=>"101010010",
  27387=>"010110000",
  27388=>"011100111",
  27389=>"110111011",
  27390=>"000111101",
  27391=>"010010110",
  27392=>"001111000",
  27393=>"111000100",
  27394=>"100000111",
  27395=>"100101101",
  27396=>"111001011",
  27397=>"000110001",
  27398=>"010001101",
  27399=>"000110000",
  27400=>"001110000",
  27401=>"111110111",
  27402=>"001011101",
  27403=>"001001100",
  27404=>"011000111",
  27405=>"100011110",
  27406=>"101000000",
  27407=>"001100001",
  27408=>"011110001",
  27409=>"101001010",
  27410=>"011000000",
  27411=>"111001000",
  27412=>"001010110",
  27413=>"101101101",
  27414=>"111100111",
  27415=>"101101011",
  27416=>"001001001",
  27417=>"111100001",
  27418=>"110001100",
  27419=>"101001111",
  27420=>"010011011",
  27421=>"010010111",
  27422=>"111101110",
  27423=>"000010011",
  27424=>"111101010",
  27425=>"000000011",
  27426=>"100011000",
  27427=>"001000101",
  27428=>"100110010",
  27429=>"000000101",
  27430=>"010010101",
  27431=>"000010110",
  27432=>"010011110",
  27433=>"101110111",
  27434=>"010001010",
  27435=>"110111011",
  27436=>"110001000",
  27437=>"011000001",
  27438=>"001110111",
  27439=>"111010111",
  27440=>"000011000",
  27441=>"000001111",
  27442=>"111000111",
  27443=>"010111111",
  27444=>"101000110",
  27445=>"000000000",
  27446=>"110010010",
  27447=>"001010010",
  27448=>"000010101",
  27449=>"101000000",
  27450=>"101011010",
  27451=>"011110100",
  27452=>"011100000",
  27453=>"001010110",
  27454=>"010000011",
  27455=>"111001101",
  27456=>"110011010",
  27457=>"010000011",
  27458=>"000000000",
  27459=>"010111000",
  27460=>"111010111",
  27461=>"100011111",
  27462=>"101001001",
  27463=>"001001110",
  27464=>"100001100",
  27465=>"001111101",
  27466=>"011110110",
  27467=>"001000100",
  27468=>"001111101",
  27469=>"011010100",
  27470=>"100001011",
  27471=>"110111101",
  27472=>"110001001",
  27473=>"100100001",
  27474=>"011101110",
  27475=>"000010001",
  27476=>"100110100",
  27477=>"010110010",
  27478=>"100011100",
  27479=>"111011010",
  27480=>"000011100",
  27481=>"110000010",
  27482=>"111000100",
  27483=>"000011000",
  27484=>"101000001",
  27485=>"110000000",
  27486=>"011100100",
  27487=>"000001011",
  27488=>"000001010",
  27489=>"111100110",
  27490=>"110001010",
  27491=>"000011111",
  27492=>"010000100",
  27493=>"000010110",
  27494=>"100010101",
  27495=>"010100111",
  27496=>"110000001",
  27497=>"101000001",
  27498=>"010111011",
  27499=>"001100101",
  27500=>"000100100",
  27501=>"001001001",
  27502=>"101100010",
  27503=>"110111111",
  27504=>"100011011",
  27505=>"011110100",
  27506=>"100001111",
  27507=>"100110111",
  27508=>"010110010",
  27509=>"111101101",
  27510=>"101101011",
  27511=>"010100000",
  27512=>"000110100",
  27513=>"001000010",
  27514=>"001100001",
  27515=>"011001000",
  27516=>"110110101",
  27517=>"111011010",
  27518=>"110010100",
  27519=>"110011001",
  27520=>"111110110",
  27521=>"011110010",
  27522=>"000010011",
  27523=>"001111111",
  27524=>"101111100",
  27525=>"001000010",
  27526=>"100100100",
  27527=>"001010101",
  27528=>"000111010",
  27529=>"101100110",
  27530=>"000000010",
  27531=>"001111100",
  27532=>"010000000",
  27533=>"011110100",
  27534=>"001001001",
  27535=>"100010001",
  27536=>"110011000",
  27537=>"000011100",
  27538=>"100101011",
  27539=>"000001011",
  27540=>"010001100",
  27541=>"001101110",
  27542=>"101100110",
  27543=>"000100110",
  27544=>"110111001",
  27545=>"001000010",
  27546=>"110010010",
  27547=>"000001101",
  27548=>"110111111",
  27549=>"101010000",
  27550=>"101010001",
  27551=>"000110100",
  27552=>"011101110",
  27553=>"100111101",
  27554=>"011011011",
  27555=>"011111110",
  27556=>"001101001",
  27557=>"011110100",
  27558=>"010001011",
  27559=>"011000011",
  27560=>"100101001",
  27561=>"100000000",
  27562=>"111111001",
  27563=>"101111101",
  27564=>"010011101",
  27565=>"111010000",
  27566=>"000010100",
  27567=>"010010010",
  27568=>"111110111",
  27569=>"010001100",
  27570=>"110000100",
  27571=>"011110010",
  27572=>"011001001",
  27573=>"010010111",
  27574=>"010011001",
  27575=>"110010101",
  27576=>"100100100",
  27577=>"011100110",
  27578=>"111110110",
  27579=>"110101010",
  27580=>"111000011",
  27581=>"110011100",
  27582=>"001001010",
  27583=>"111101111",
  27584=>"001101111",
  27585=>"101001001",
  27586=>"111110101",
  27587=>"000001001",
  27588=>"010010100",
  27589=>"001010101",
  27590=>"001111000",
  27591=>"010000001",
  27592=>"011001000",
  27593=>"100000101",
  27594=>"010000100",
  27595=>"100000000",
  27596=>"000111000",
  27597=>"010000010",
  27598=>"001111100",
  27599=>"110011110",
  27600=>"010100010",
  27601=>"000000010",
  27602=>"000000100",
  27603=>"001001001",
  27604=>"101010000",
  27605=>"110011110",
  27606=>"001001110",
  27607=>"000001000",
  27608=>"001010101",
  27609=>"111110011",
  27610=>"011001000",
  27611=>"111111001",
  27612=>"011001101",
  27613=>"011111011",
  27614=>"000001110",
  27615=>"100010011",
  27616=>"010001110",
  27617=>"000100101",
  27618=>"000111000",
  27619=>"101111111",
  27620=>"000000100",
  27621=>"111011101",
  27622=>"001001111",
  27623=>"000101000",
  27624=>"111001000",
  27625=>"010100110",
  27626=>"000011010",
  27627=>"001110011",
  27628=>"111010111",
  27629=>"101010111",
  27630=>"001101011",
  27631=>"111010010",
  27632=>"001000101",
  27633=>"011011100",
  27634=>"111001101",
  27635=>"010101001",
  27636=>"001100000",
  27637=>"101010010",
  27638=>"011100100",
  27639=>"111110011",
  27640=>"101111101",
  27641=>"101111101",
  27642=>"000111001",
  27643=>"000100111",
  27644=>"111000100",
  27645=>"111010001",
  27646=>"110101011",
  27647=>"011100111",
  27648=>"100010010",
  27649=>"001010011",
  27650=>"110111011",
  27651=>"010101111",
  27652=>"000000000",
  27653=>"010111001",
  27654=>"100101110",
  27655=>"110100000",
  27656=>"110001101",
  27657=>"000100110",
  27658=>"111001011",
  27659=>"010100110",
  27660=>"000001011",
  27661=>"111110100",
  27662=>"111010101",
  27663=>"111001111",
  27664=>"001010010",
  27665=>"110000111",
  27666=>"000101010",
  27667=>"101111111",
  27668=>"000010100",
  27669=>"110101111",
  27670=>"001101000",
  27671=>"011110010",
  27672=>"000110100",
  27673=>"010001111",
  27674=>"101000001",
  27675=>"111111111",
  27676=>"101001001",
  27677=>"101110000",
  27678=>"111010011",
  27679=>"100001011",
  27680=>"000010010",
  27681=>"010101011",
  27682=>"010011001",
  27683=>"110111101",
  27684=>"000101111",
  27685=>"110000110",
  27686=>"010111101",
  27687=>"101100110",
  27688=>"000001110",
  27689=>"010010110",
  27690=>"001000010",
  27691=>"000111101",
  27692=>"110100010",
  27693=>"100010111",
  27694=>"100001001",
  27695=>"011001101",
  27696=>"111101100",
  27697=>"001110100",
  27698=>"111010001",
  27699=>"110101000",
  27700=>"100000100",
  27701=>"010000011",
  27702=>"110011010",
  27703=>"110110011",
  27704=>"110011100",
  27705=>"010001001",
  27706=>"100100000",
  27707=>"101001101",
  27708=>"000100101",
  27709=>"101000101",
  27710=>"000000011",
  27711=>"100110110",
  27712=>"111101011",
  27713=>"000010010",
  27714=>"010010000",
  27715=>"001100000",
  27716=>"010111101",
  27717=>"001111010",
  27718=>"110001010",
  27719=>"101101000",
  27720=>"100111000",
  27721=>"101011011",
  27722=>"011001000",
  27723=>"100000111",
  27724=>"010110010",
  27725=>"000101110",
  27726=>"010111101",
  27727=>"010011011",
  27728=>"100001001",
  27729=>"011101111",
  27730=>"001111110",
  27731=>"110011110",
  27732=>"000010110",
  27733=>"110111100",
  27734=>"101111110",
  27735=>"110110011",
  27736=>"011110000",
  27737=>"011101110",
  27738=>"110011000",
  27739=>"000111000",
  27740=>"100100110",
  27741=>"000010001",
  27742=>"100000010",
  27743=>"000010011",
  27744=>"111111111",
  27745=>"101101110",
  27746=>"011101001",
  27747=>"110111011",
  27748=>"100001100",
  27749=>"110101110",
  27750=>"011110000",
  27751=>"001110000",
  27752=>"011001011",
  27753=>"100100001",
  27754=>"000000000",
  27755=>"010111100",
  27756=>"110000111",
  27757=>"111100111",
  27758=>"011000001",
  27759=>"100011010",
  27760=>"001101010",
  27761=>"110010110",
  27762=>"011011010",
  27763=>"110101100",
  27764=>"010110011",
  27765=>"111110000",
  27766=>"100000100",
  27767=>"010110101",
  27768=>"001010010",
  27769=>"110110000",
  27770=>"001000100",
  27771=>"000100010",
  27772=>"110101001",
  27773=>"110010000",
  27774=>"010100110",
  27775=>"001000101",
  27776=>"100001111",
  27777=>"111000110",
  27778=>"110011100",
  27779=>"000011001",
  27780=>"010001000",
  27781=>"000011111",
  27782=>"000110110",
  27783=>"001100010",
  27784=>"010111111",
  27785=>"000001010",
  27786=>"100000000",
  27787=>"010010101",
  27788=>"101100010",
  27789=>"101010000",
  27790=>"111011101",
  27791=>"111111010",
  27792=>"100000110",
  27793=>"100101111",
  27794=>"101000010",
  27795=>"111101111",
  27796=>"100000011",
  27797=>"010110100",
  27798=>"110101110",
  27799=>"000101011",
  27800=>"000000000",
  27801=>"011101101",
  27802=>"001110001",
  27803=>"011001111",
  27804=>"011100111",
  27805=>"000010001",
  27806=>"000000100",
  27807=>"011000001",
  27808=>"010001000",
  27809=>"110110001",
  27810=>"011111000",
  27811=>"100011000",
  27812=>"010001001",
  27813=>"101100110",
  27814=>"010110111",
  27815=>"110001010",
  27816=>"110010001",
  27817=>"010110110",
  27818=>"011001011",
  27819=>"110010000",
  27820=>"101111001",
  27821=>"001000000",
  27822=>"101101000",
  27823=>"110110101",
  27824=>"000010000",
  27825=>"100001000",
  27826=>"000110110",
  27827=>"001001000",
  27828=>"111100011",
  27829=>"011000110",
  27830=>"111010010",
  27831=>"100011100",
  27832=>"011100011",
  27833=>"010110011",
  27834=>"011011010",
  27835=>"111111110",
  27836=>"111101110",
  27837=>"011001010",
  27838=>"110000110",
  27839=>"001000011",
  27840=>"000000011",
  27841=>"100000101",
  27842=>"000011001",
  27843=>"100011111",
  27844=>"011011001",
  27845=>"010010110",
  27846=>"001110001",
  27847=>"000100101",
  27848=>"111011111",
  27849=>"100010110",
  27850=>"101001001",
  27851=>"111100001",
  27852=>"001010010",
  27853=>"111111100",
  27854=>"010111000",
  27855=>"001011111",
  27856=>"111000100",
  27857=>"110110011",
  27858=>"101000100",
  27859=>"101001000",
  27860=>"101001101",
  27861=>"100001001",
  27862=>"101101110",
  27863=>"100001100",
  27864=>"000111000",
  27865=>"111100000",
  27866=>"110010110",
  27867=>"111101011",
  27868=>"011010001",
  27869=>"101101100",
  27870=>"000111011",
  27871=>"111111000",
  27872=>"100101110",
  27873=>"011100000",
  27874=>"100101111",
  27875=>"111101111",
  27876=>"000011100",
  27877=>"001111000",
  27878=>"001011000",
  27879=>"111011100",
  27880=>"101010111",
  27881=>"110110101",
  27882=>"000100010",
  27883=>"011101111",
  27884=>"010001000",
  27885=>"100101011",
  27886=>"001010110",
  27887=>"000100110",
  27888=>"101101101",
  27889=>"011011101",
  27890=>"000111110",
  27891=>"000100011",
  27892=>"010011001",
  27893=>"000100110",
  27894=>"111100010",
  27895=>"110011101",
  27896=>"001000110",
  27897=>"010001100",
  27898=>"000111000",
  27899=>"101111100",
  27900=>"100001010",
  27901=>"010111110",
  27902=>"111111001",
  27903=>"001010100",
  27904=>"001011101",
  27905=>"000111000",
  27906=>"011101111",
  27907=>"110000001",
  27908=>"100010001",
  27909=>"110101111",
  27910=>"011100100",
  27911=>"111100110",
  27912=>"001100100",
  27913=>"110101010",
  27914=>"111100110",
  27915=>"010010111",
  27916=>"111011101",
  27917=>"001110000",
  27918=>"000001000",
  27919=>"000001010",
  27920=>"101111000",
  27921=>"001110110",
  27922=>"101011011",
  27923=>"000011100",
  27924=>"111110111",
  27925=>"101010011",
  27926=>"000001101",
  27927=>"101000100",
  27928=>"110111101",
  27929=>"110011001",
  27930=>"110100111",
  27931=>"101111111",
  27932=>"001111011",
  27933=>"101000111",
  27934=>"100110110",
  27935=>"001001101",
  27936=>"000111101",
  27937=>"011111001",
  27938=>"001101000",
  27939=>"000010010",
  27940=>"101111011",
  27941=>"110100001",
  27942=>"010111110",
  27943=>"100011100",
  27944=>"000000011",
  27945=>"101000010",
  27946=>"110110101",
  27947=>"101110000",
  27948=>"110100000",
  27949=>"010100001",
  27950=>"000000010",
  27951=>"000100110",
  27952=>"010111101",
  27953=>"011100101",
  27954=>"011001101",
  27955=>"110010000",
  27956=>"001100000",
  27957=>"101000011",
  27958=>"011111010",
  27959=>"100010111",
  27960=>"000100111",
  27961=>"011110111",
  27962=>"001111010",
  27963=>"111010000",
  27964=>"001101010",
  27965=>"100110011",
  27966=>"110001011",
  27967=>"001001100",
  27968=>"001111000",
  27969=>"100101001",
  27970=>"000111111",
  27971=>"101010100",
  27972=>"010011011",
  27973=>"110110101",
  27974=>"010010011",
  27975=>"010001101",
  27976=>"101010000",
  27977=>"111010001",
  27978=>"101110100",
  27979=>"000011101",
  27980=>"011110110",
  27981=>"010000110",
  27982=>"000000000",
  27983=>"100010010",
  27984=>"110101101",
  27985=>"001101001",
  27986=>"000100011",
  27987=>"000011100",
  27988=>"100111100",
  27989=>"011000111",
  27990=>"100000011",
  27991=>"010001000",
  27992=>"011100100",
  27993=>"110100111",
  27994=>"010110001",
  27995=>"011111010",
  27996=>"101000011",
  27997=>"010110010",
  27998=>"000001011",
  27999=>"111010111",
  28000=>"010000101",
  28001=>"111111111",
  28002=>"010110001",
  28003=>"010100011",
  28004=>"001010100",
  28005=>"011001001",
  28006=>"000000010",
  28007=>"110101111",
  28008=>"001011010",
  28009=>"000100111",
  28010=>"001001110",
  28011=>"000101110",
  28012=>"010010100",
  28013=>"010101010",
  28014=>"101101000",
  28015=>"011010100",
  28016=>"111100001",
  28017=>"011101000",
  28018=>"010010000",
  28019=>"101110000",
  28020=>"011100110",
  28021=>"000110011",
  28022=>"001010001",
  28023=>"011011111",
  28024=>"100011100",
  28025=>"110110000",
  28026=>"111010011",
  28027=>"110100101",
  28028=>"100001001",
  28029=>"000010000",
  28030=>"000000001",
  28031=>"111011111",
  28032=>"000001000",
  28033=>"001010011",
  28034=>"001011000",
  28035=>"011101001",
  28036=>"100001111",
  28037=>"010011010",
  28038=>"101111100",
  28039=>"000001001",
  28040=>"000111010",
  28041=>"100011011",
  28042=>"000011111",
  28043=>"100100000",
  28044=>"100110101",
  28045=>"000001000",
  28046=>"010101101",
  28047=>"000110101",
  28048=>"100100011",
  28049=>"000000001",
  28050=>"101100111",
  28051=>"011000001",
  28052=>"000011010",
  28053=>"101000010",
  28054=>"111110111",
  28055=>"101011111",
  28056=>"011011010",
  28057=>"001111011",
  28058=>"010100001",
  28059=>"111110110",
  28060=>"011111011",
  28061=>"100010111",
  28062=>"000011111",
  28063=>"010001000",
  28064=>"010011001",
  28065=>"100100100",
  28066=>"110100000",
  28067=>"111111111",
  28068=>"011011000",
  28069=>"001010010",
  28070=>"110011000",
  28071=>"110010011",
  28072=>"101111011",
  28073=>"111101111",
  28074=>"011100000",
  28075=>"010011001",
  28076=>"000111010",
  28077=>"001010010",
  28078=>"110001100",
  28079=>"011001011",
  28080=>"110111111",
  28081=>"010000110",
  28082=>"000011100",
  28083=>"111111101",
  28084=>"000101110",
  28085=>"110000000",
  28086=>"000011011",
  28087=>"111010110",
  28088=>"100101111",
  28089=>"000100011",
  28090=>"011110000",
  28091=>"101010010",
  28092=>"110100010",
  28093=>"000001101",
  28094=>"001110101",
  28095=>"111000000",
  28096=>"100100100",
  28097=>"100010010",
  28098=>"000001100",
  28099=>"111001000",
  28100=>"001010000",
  28101=>"011101001",
  28102=>"100001111",
  28103=>"101101101",
  28104=>"110011100",
  28105=>"100101110",
  28106=>"100001101",
  28107=>"110011111",
  28108=>"110101100",
  28109=>"111110001",
  28110=>"111101110",
  28111=>"100101110",
  28112=>"110110101",
  28113=>"100101000",
  28114=>"001011111",
  28115=>"000000011",
  28116=>"101111100",
  28117=>"010110000",
  28118=>"011110001",
  28119=>"010100100",
  28120=>"011000101",
  28121=>"011001010",
  28122=>"010010111",
  28123=>"111001111",
  28124=>"111100010",
  28125=>"111101000",
  28126=>"110101110",
  28127=>"001110001",
  28128=>"000110110",
  28129=>"000101110",
  28130=>"101111111",
  28131=>"110000100",
  28132=>"100100010",
  28133=>"000001110",
  28134=>"001100110",
  28135=>"010000001",
  28136=>"000111011",
  28137=>"111111110",
  28138=>"001000100",
  28139=>"110101101",
  28140=>"000001000",
  28141=>"110100000",
  28142=>"001110001",
  28143=>"100111001",
  28144=>"100001101",
  28145=>"110001001",
  28146=>"100110110",
  28147=>"100111111",
  28148=>"011010000",
  28149=>"001000000",
  28150=>"100110001",
  28151=>"110001000",
  28152=>"001011000",
  28153=>"011001110",
  28154=>"111100110",
  28155=>"001110000",
  28156=>"111101111",
  28157=>"000000101",
  28158=>"010001111",
  28159=>"101111000",
  28160=>"100011010",
  28161=>"100001010",
  28162=>"110110011",
  28163=>"111100100",
  28164=>"110001110",
  28165=>"000111100",
  28166=>"011000001",
  28167=>"001111000",
  28168=>"010000000",
  28169=>"101100101",
  28170=>"101100101",
  28171=>"001101010",
  28172=>"101111001",
  28173=>"010110011",
  28174=>"001000010",
  28175=>"100011101",
  28176=>"001001001",
  28177=>"111101010",
  28178=>"001010010",
  28179=>"010111101",
  28180=>"000000111",
  28181=>"001101000",
  28182=>"111100010",
  28183=>"111000100",
  28184=>"111111001",
  28185=>"010010000",
  28186=>"101000110",
  28187=>"001010100",
  28188=>"110100011",
  28189=>"011000011",
  28190=>"100001010",
  28191=>"111110011",
  28192=>"010100110",
  28193=>"101010100",
  28194=>"010111110",
  28195=>"010001011",
  28196=>"110010110",
  28197=>"100010100",
  28198=>"100010110",
  28199=>"010010110",
  28200=>"001000001",
  28201=>"001000001",
  28202=>"000110010",
  28203=>"011110001",
  28204=>"000010010",
  28205=>"000100000",
  28206=>"001000000",
  28207=>"000001011",
  28208=>"111100010",
  28209=>"111101110",
  28210=>"010101010",
  28211=>"000010100",
  28212=>"110111000",
  28213=>"001011010",
  28214=>"101001001",
  28215=>"000111111",
  28216=>"101000000",
  28217=>"100111100",
  28218=>"100011000",
  28219=>"000110111",
  28220=>"110010111",
  28221=>"101101011",
  28222=>"010011101",
  28223=>"000110001",
  28224=>"100011111",
  28225=>"010100010",
  28226=>"000110000",
  28227=>"011111001",
  28228=>"111101101",
  28229=>"111101001",
  28230=>"010001010",
  28231=>"001011100",
  28232=>"001110111",
  28233=>"000101100",
  28234=>"101011011",
  28235=>"001000101",
  28236=>"011100110",
  28237=>"100101111",
  28238=>"100101010",
  28239=>"110110000",
  28240=>"000000101",
  28241=>"110111111",
  28242=>"101010101",
  28243=>"001110100",
  28244=>"100010100",
  28245=>"101011110",
  28246=>"110111000",
  28247=>"000110101",
  28248=>"000000110",
  28249=>"110111000",
  28250=>"111011001",
  28251=>"000100111",
  28252=>"011100110",
  28253=>"010111011",
  28254=>"000000101",
  28255=>"110001011",
  28256=>"011001110",
  28257=>"110000001",
  28258=>"111001011",
  28259=>"011100110",
  28260=>"010111111",
  28261=>"000100101",
  28262=>"010000010",
  28263=>"100011000",
  28264=>"011100000",
  28265=>"110000111",
  28266=>"010110111",
  28267=>"110111111",
  28268=>"001010001",
  28269=>"100000101",
  28270=>"110110101",
  28271=>"101111100",
  28272=>"001000101",
  28273=>"001001110",
  28274=>"111110011",
  28275=>"010111111",
  28276=>"110100100",
  28277=>"100011111",
  28278=>"101111011",
  28279=>"100000000",
  28280=>"001011010",
  28281=>"010111011",
  28282=>"111000110",
  28283=>"001000111",
  28284=>"011110000",
  28285=>"000001100",
  28286=>"101100010",
  28287=>"010011010",
  28288=>"110001011",
  28289=>"100101110",
  28290=>"101010100",
  28291=>"001101001",
  28292=>"010101110",
  28293=>"100101011",
  28294=>"101100110",
  28295=>"001000110",
  28296=>"001110100",
  28297=>"010111011",
  28298=>"111111111",
  28299=>"000000110",
  28300=>"111001010",
  28301=>"000011111",
  28302=>"100101110",
  28303=>"100001111",
  28304=>"101000000",
  28305=>"001010110",
  28306=>"000100000",
  28307=>"000010111",
  28308=>"100000110",
  28309=>"001100110",
  28310=>"000111100",
  28311=>"001100101",
  28312=>"000001011",
  28313=>"011110110",
  28314=>"001111000",
  28315=>"000010001",
  28316=>"000010100",
  28317=>"111010101",
  28318=>"110000000",
  28319=>"110011110",
  28320=>"111110100",
  28321=>"111111011",
  28322=>"100101011",
  28323=>"111011010",
  28324=>"100100110",
  28325=>"101110011",
  28326=>"111111011",
  28327=>"110001111",
  28328=>"001101101",
  28329=>"011100111",
  28330=>"101000101",
  28331=>"000000000",
  28332=>"001110000",
  28333=>"000010100",
  28334=>"111100100",
  28335=>"011100111",
  28336=>"110000000",
  28337=>"110010010",
  28338=>"011011001",
  28339=>"011010011",
  28340=>"101111000",
  28341=>"000101110",
  28342=>"101110010",
  28343=>"101010110",
  28344=>"100001000",
  28345=>"111010101",
  28346=>"001011011",
  28347=>"111100111",
  28348=>"010100111",
  28349=>"110000000",
  28350=>"110010110",
  28351=>"011011001",
  28352=>"110100110",
  28353=>"011010101",
  28354=>"111001011",
  28355=>"110101100",
  28356=>"000001011",
  28357=>"111001100",
  28358=>"011010001",
  28359=>"000100110",
  28360=>"111000100",
  28361=>"110110001",
  28362=>"101100110",
  28363=>"101010001",
  28364=>"011011100",
  28365=>"010001000",
  28366=>"010011011",
  28367=>"101000101",
  28368=>"010001010",
  28369=>"110010001",
  28370=>"011101010",
  28371=>"110110101",
  28372=>"101000110",
  28373=>"010000011",
  28374=>"000011010",
  28375=>"100001111",
  28376=>"000110000",
  28377=>"100000000",
  28378=>"011101110",
  28379=>"011011101",
  28380=>"111101011",
  28381=>"000010011",
  28382=>"111100011",
  28383=>"100010110",
  28384=>"111010111",
  28385=>"110000001",
  28386=>"001001001",
  28387=>"100100110",
  28388=>"111111100",
  28389=>"000100111",
  28390=>"100010111",
  28391=>"000000011",
  28392=>"101111000",
  28393=>"100010110",
  28394=>"110111011",
  28395=>"010111010",
  28396=>"011010111",
  28397=>"100001000",
  28398=>"011000110",
  28399=>"000110101",
  28400=>"011010111",
  28401=>"011001011",
  28402=>"101011011",
  28403=>"001111010",
  28404=>"110011000",
  28405=>"101000101",
  28406=>"100000000",
  28407=>"010011011",
  28408=>"001010000",
  28409=>"100001110",
  28410=>"001101110",
  28411=>"010100100",
  28412=>"111111010",
  28413=>"111111101",
  28414=>"000000000",
  28415=>"101010111",
  28416=>"111110000",
  28417=>"011001100",
  28418=>"101011111",
  28419=>"000000011",
  28420=>"100110010",
  28421=>"001001001",
  28422=>"111000110",
  28423=>"010111100",
  28424=>"010001111",
  28425=>"111001110",
  28426=>"011111010",
  28427=>"100010110",
  28428=>"010111110",
  28429=>"000111000",
  28430=>"001001110",
  28431=>"001101100",
  28432=>"111100001",
  28433=>"110011001",
  28434=>"111101110",
  28435=>"110100000",
  28436=>"001001011",
  28437=>"101111011",
  28438=>"011000100",
  28439=>"100011000",
  28440=>"110111010",
  28441=>"011111101",
  28442=>"001000110",
  28443=>"110101110",
  28444=>"011000110",
  28445=>"000001001",
  28446=>"000011100",
  28447=>"110100000",
  28448=>"010001101",
  28449=>"000001110",
  28450=>"111000000",
  28451=>"001000011",
  28452=>"110100010",
  28453=>"100001100",
  28454=>"100001100",
  28455=>"010111010",
  28456=>"011111111",
  28457=>"101100000",
  28458=>"101011101",
  28459=>"000111000",
  28460=>"000010111",
  28461=>"011110111",
  28462=>"010100101",
  28463=>"100010011",
  28464=>"011111101",
  28465=>"111001110",
  28466=>"111001000",
  28467=>"110011011",
  28468=>"101011001",
  28469=>"110101010",
  28470=>"111001011",
  28471=>"010110110",
  28472=>"010110000",
  28473=>"010111001",
  28474=>"000010011",
  28475=>"111111011",
  28476=>"000101100",
  28477=>"111010101",
  28478=>"011001100",
  28479=>"101011001",
  28480=>"000111001",
  28481=>"011000100",
  28482=>"000101100",
  28483=>"111011100",
  28484=>"000110000",
  28485=>"111000100",
  28486=>"010100011",
  28487=>"111010000",
  28488=>"110000010",
  28489=>"101110000",
  28490=>"011110111",
  28491=>"000111000",
  28492=>"001110001",
  28493=>"110010111",
  28494=>"010100101",
  28495=>"100111111",
  28496=>"101101001",
  28497=>"000100000",
  28498=>"001010001",
  28499=>"110001000",
  28500=>"100010011",
  28501=>"110000001",
  28502=>"000001111",
  28503=>"000101000",
  28504=>"100110100",
  28505=>"101111111",
  28506=>"000011110",
  28507=>"000100010",
  28508=>"000111000",
  28509=>"101100011",
  28510=>"000011110",
  28511=>"101010110",
  28512=>"110111110",
  28513=>"110110100",
  28514=>"111000011",
  28515=>"011100100",
  28516=>"011100110",
  28517=>"010010011",
  28518=>"111101000",
  28519=>"110101010",
  28520=>"100001000",
  28521=>"011001011",
  28522=>"101100010",
  28523=>"101000010",
  28524=>"011100101",
  28525=>"000001110",
  28526=>"110000110",
  28527=>"010001011",
  28528=>"111011111",
  28529=>"011011100",
  28530=>"010110100",
  28531=>"010011110",
  28532=>"100110110",
  28533=>"111010101",
  28534=>"111001110",
  28535=>"011000100",
  28536=>"011100011",
  28537=>"000011000",
  28538=>"011000011",
  28539=>"011100001",
  28540=>"010000000",
  28541=>"000100011",
  28542=>"111010100",
  28543=>"011110001",
  28544=>"000110000",
  28545=>"111010111",
  28546=>"100011111",
  28547=>"011100110",
  28548=>"111000110",
  28549=>"001000011",
  28550=>"010011010",
  28551=>"011111110",
  28552=>"011010101",
  28553=>"000000111",
  28554=>"010110001",
  28555=>"110110100",
  28556=>"110010000",
  28557=>"111100001",
  28558=>"011011110",
  28559=>"011101101",
  28560=>"011010001",
  28561=>"000011011",
  28562=>"111001100",
  28563=>"001000011",
  28564=>"110001110",
  28565=>"110001110",
  28566=>"110110001",
  28567=>"000001000",
  28568=>"111110011",
  28569=>"000000101",
  28570=>"000110000",
  28571=>"011011000",
  28572=>"010011010",
  28573=>"110010110",
  28574=>"110000100",
  28575=>"111110111",
  28576=>"001110101",
  28577=>"011011111",
  28578=>"010001110",
  28579=>"110100000",
  28580=>"000010000",
  28581=>"100101101",
  28582=>"101000010",
  28583=>"100011101",
  28584=>"010110101",
  28585=>"000011011",
  28586=>"101111101",
  28587=>"110001111",
  28588=>"001111010",
  28589=>"111101001",
  28590=>"011011000",
  28591=>"011110011",
  28592=>"111111100",
  28593=>"110010011",
  28594=>"001001110",
  28595=>"011101100",
  28596=>"001110100",
  28597=>"010010111",
  28598=>"010110110",
  28599=>"111111001",
  28600=>"101000000",
  28601=>"100011111",
  28602=>"011001111",
  28603=>"100000001",
  28604=>"110011010",
  28605=>"010001100",
  28606=>"100111001",
  28607=>"010000111",
  28608=>"010110000",
  28609=>"001000010",
  28610=>"110101111",
  28611=>"010010111",
  28612=>"010010000",
  28613=>"000000011",
  28614=>"011010100",
  28615=>"100111101",
  28616=>"000010101",
  28617=>"011100100",
  28618=>"111010000",
  28619=>"000001010",
  28620=>"110110010",
  28621=>"101000000",
  28622=>"001001000",
  28623=>"011111000",
  28624=>"101000100",
  28625=>"111111100",
  28626=>"011000010",
  28627=>"000111001",
  28628=>"111111111",
  28629=>"110110101",
  28630=>"100000000",
  28631=>"111101110",
  28632=>"000110000",
  28633=>"100001100",
  28634=>"000100000",
  28635=>"100100000",
  28636=>"010001110",
  28637=>"011100011",
  28638=>"011101101",
  28639=>"010000110",
  28640=>"110000111",
  28641=>"000100111",
  28642=>"111111101",
  28643=>"111000100",
  28644=>"000110011",
  28645=>"001010110",
  28646=>"000000011",
  28647=>"111010101",
  28648=>"011111000",
  28649=>"100001110",
  28650=>"001000110",
  28651=>"000101000",
  28652=>"011110010",
  28653=>"111000101",
  28654=>"001000100",
  28655=>"101011000",
  28656=>"000100010",
  28657=>"000111001",
  28658=>"101110101",
  28659=>"010100101",
  28660=>"100101011",
  28661=>"111001001",
  28662=>"110101010",
  28663=>"100000000",
  28664=>"010110000",
  28665=>"011000011",
  28666=>"000011000",
  28667=>"111010000",
  28668=>"010100001",
  28669=>"110000000",
  28670=>"110000010",
  28671=>"010000111",
  28672=>"000010000",
  28673=>"001100001",
  28674=>"011011001",
  28675=>"101100110",
  28676=>"010001011",
  28677=>"100101011",
  28678=>"110100010",
  28679=>"010111100",
  28680=>"000010000",
  28681=>"000001010",
  28682=>"000111101",
  28683=>"001110110",
  28684=>"111000000",
  28685=>"000011000",
  28686=>"111101110",
  28687=>"111011110",
  28688=>"110111000",
  28689=>"101000111",
  28690=>"101100101",
  28691=>"010011101",
  28692=>"011100010",
  28693=>"000010011",
  28694=>"001111101",
  28695=>"100111000",
  28696=>"101110110",
  28697=>"001100110",
  28698=>"111011000",
  28699=>"111011101",
  28700=>"101010110",
  28701=>"110110001",
  28702=>"000000101",
  28703=>"100001000",
  28704=>"110110010",
  28705=>"101001100",
  28706=>"100111101",
  28707=>"000100101",
  28708=>"001111101",
  28709=>"010010000",
  28710=>"001010010",
  28711=>"010001011",
  28712=>"101101001",
  28713=>"110100101",
  28714=>"100110000",
  28715=>"000100111",
  28716=>"010011011",
  28717=>"100011110",
  28718=>"101101001",
  28719=>"111001000",
  28720=>"000101000",
  28721=>"101011110",
  28722=>"010111110",
  28723=>"010010111",
  28724=>"010000000",
  28725=>"000000000",
  28726=>"001011110",
  28727=>"010001110",
  28728=>"001111100",
  28729=>"110000001",
  28730=>"001000111",
  28731=>"000111100",
  28732=>"110011001",
  28733=>"000010001",
  28734=>"110001000",
  28735=>"011010110",
  28736=>"111100011",
  28737=>"110010100",
  28738=>"111101010",
  28739=>"101101011",
  28740=>"101111111",
  28741=>"111000101",
  28742=>"010100001",
  28743=>"001011100",
  28744=>"000110001",
  28745=>"010101110",
  28746=>"000001101",
  28747=>"101110000",
  28748=>"010000001",
  28749=>"100111010",
  28750=>"111001000",
  28751=>"111101100",
  28752=>"100001001",
  28753=>"000000100",
  28754=>"101000110",
  28755=>"110101001",
  28756=>"010111101",
  28757=>"011001110",
  28758=>"110101001",
  28759=>"100100110",
  28760=>"110100001",
  28761=>"101100101",
  28762=>"111101110",
  28763=>"110100100",
  28764=>"010111000",
  28765=>"110001110",
  28766=>"111100001",
  28767=>"000001110",
  28768=>"101100101",
  28769=>"001010111",
  28770=>"001100010",
  28771=>"011000000",
  28772=>"111111011",
  28773=>"011101100",
  28774=>"101010111",
  28775=>"001000111",
  28776=>"111001101",
  28777=>"110111110",
  28778=>"110011110",
  28779=>"110101111",
  28780=>"001101010",
  28781=>"111000000",
  28782=>"101001001",
  28783=>"000000011",
  28784=>"111110101",
  28785=>"000000001",
  28786=>"111101011",
  28787=>"100100100",
  28788=>"010101101",
  28789=>"111010001",
  28790=>"001001111",
  28791=>"111011001",
  28792=>"100111010",
  28793=>"010101101",
  28794=>"000101000",
  28795=>"101001010",
  28796=>"010101100",
  28797=>"110000100",
  28798=>"110000111",
  28799=>"101011011",
  28800=>"011011001",
  28801=>"101011101",
  28802=>"001010010",
  28803=>"101100000",
  28804=>"000100000",
  28805=>"100110100",
  28806=>"110010100",
  28807=>"110111110",
  28808=>"101100011",
  28809=>"000100111",
  28810=>"110111001",
  28811=>"110011101",
  28812=>"111100011",
  28813=>"000001011",
  28814=>"000110011",
  28815=>"010111101",
  28816=>"111010110",
  28817=>"000000010",
  28818=>"000001000",
  28819=>"011000010",
  28820=>"000000000",
  28821=>"110101101",
  28822=>"111001100",
  28823=>"001100111",
  28824=>"000100000",
  28825=>"110101001",
  28826=>"100111100",
  28827=>"101111000",
  28828=>"000001000",
  28829=>"010111000",
  28830=>"100100010",
  28831=>"011011101",
  28832=>"000101000",
  28833=>"001101110",
  28834=>"111111111",
  28835=>"111010110",
  28836=>"011100010",
  28837=>"010000011",
  28838=>"011000110",
  28839=>"001011011",
  28840=>"001101111",
  28841=>"011000000",
  28842=>"100111111",
  28843=>"100010001",
  28844=>"000010100",
  28845=>"111001100",
  28846=>"110000000",
  28847=>"101000000",
  28848=>"101000111",
  28849=>"101000000",
  28850=>"100100101",
  28851=>"010000001",
  28852=>"110011111",
  28853=>"010011011",
  28854=>"101010001",
  28855=>"101111101",
  28856=>"100001000",
  28857=>"110111111",
  28858=>"000101110",
  28859=>"111111000",
  28860=>"101001010",
  28861=>"011110011",
  28862=>"100010100",
  28863=>"011011010",
  28864=>"110111110",
  28865=>"010000111",
  28866=>"000110011",
  28867=>"011000010",
  28868=>"101001000",
  28869=>"111110001",
  28870=>"000111010",
  28871=>"110111100",
  28872=>"110111111",
  28873=>"111110101",
  28874=>"110111100",
  28875=>"101110001",
  28876=>"001100111",
  28877=>"110100101",
  28878=>"110010000",
  28879=>"001001100",
  28880=>"111111101",
  28881=>"111001010",
  28882=>"110101010",
  28883=>"000001010",
  28884=>"110100011",
  28885=>"100000101",
  28886=>"010011000",
  28887=>"010011000",
  28888=>"111011111",
  28889=>"001101010",
  28890=>"101001001",
  28891=>"000001100",
  28892=>"101000010",
  28893=>"110110110",
  28894=>"001001001",
  28895=>"101001111",
  28896=>"000110011",
  28897=>"111101000",
  28898=>"110111001",
  28899=>"101010010",
  28900=>"111000011",
  28901=>"000000100",
  28902=>"000111101",
  28903=>"001110001",
  28904=>"000111010",
  28905=>"000010110",
  28906=>"110111000",
  28907=>"010111110",
  28908=>"000011001",
  28909=>"100011011",
  28910=>"100011110",
  28911=>"101010110",
  28912=>"100011010",
  28913=>"001000000",
  28914=>"100000010",
  28915=>"001001101",
  28916=>"111001101",
  28917=>"000111110",
  28918=>"111101110",
  28919=>"000001110",
  28920=>"101011101",
  28921=>"110010110",
  28922=>"111000101",
  28923=>"011100010",
  28924=>"011100100",
  28925=>"000000000",
  28926=>"101011100",
  28927=>"010001010",
  28928=>"010001111",
  28929=>"010100001",
  28930=>"001111100",
  28931=>"010010110",
  28932=>"010010011",
  28933=>"001110101",
  28934=>"111100011",
  28935=>"000011111",
  28936=>"100011110",
  28937=>"000010010",
  28938=>"010010001",
  28939=>"111110001",
  28940=>"011111011",
  28941=>"111011000",
  28942=>"011010101",
  28943=>"111110110",
  28944=>"100111011",
  28945=>"110101000",
  28946=>"000011101",
  28947=>"100111000",
  28948=>"111111110",
  28949=>"001111110",
  28950=>"101010110",
  28951=>"111111001",
  28952=>"011001100",
  28953=>"000110110",
  28954=>"110101011",
  28955=>"011101000",
  28956=>"101011011",
  28957=>"111000010",
  28958=>"011111111",
  28959=>"000001111",
  28960=>"110000111",
  28961=>"001000000",
  28962=>"010111111",
  28963=>"000111000",
  28964=>"110110001",
  28965=>"101111011",
  28966=>"110100101",
  28967=>"000100101",
  28968=>"100011000",
  28969=>"111001100",
  28970=>"010011110",
  28971=>"110101010",
  28972=>"010011100",
  28973=>"010010000",
  28974=>"001000111",
  28975=>"100000011",
  28976=>"001101010",
  28977=>"001001101",
  28978=>"111010000",
  28979=>"010000011",
  28980=>"100101101",
  28981=>"000000110",
  28982=>"101010010",
  28983=>"110000000",
  28984=>"011000110",
  28985=>"100100001",
  28986=>"111011110",
  28987=>"101011011",
  28988=>"000111001",
  28989=>"110111010",
  28990=>"000111000",
  28991=>"100100011",
  28992=>"111000010",
  28993=>"010110110",
  28994=>"000100100",
  28995=>"000000101",
  28996=>"010001010",
  28997=>"000010001",
  28998=>"101110100",
  28999=>"000100001",
  29000=>"010001111",
  29001=>"100101000",
  29002=>"001001001",
  29003=>"110010000",
  29004=>"010000001",
  29005=>"111101000",
  29006=>"110110011",
  29007=>"000011010",
  29008=>"110010000",
  29009=>"110011000",
  29010=>"100001110",
  29011=>"001100010",
  29012=>"111111110",
  29013=>"100011110",
  29014=>"000011011",
  29015=>"110001010",
  29016=>"100000111",
  29017=>"000100111",
  29018=>"010100001",
  29019=>"000100101",
  29020=>"011101010",
  29021=>"110101001",
  29022=>"111111011",
  29023=>"101000101",
  29024=>"111010000",
  29025=>"011111110",
  29026=>"010000111",
  29027=>"011011000",
  29028=>"111000110",
  29029=>"000110111",
  29030=>"000100100",
  29031=>"010100000",
  29032=>"101100001",
  29033=>"010100110",
  29034=>"110111010",
  29035=>"111010000",
  29036=>"100000100",
  29037=>"110100000",
  29038=>"011010001",
  29039=>"100011110",
  29040=>"000010110",
  29041=>"101101001",
  29042=>"110100001",
  29043=>"100000110",
  29044=>"000101000",
  29045=>"010111000",
  29046=>"111001111",
  29047=>"000111111",
  29048=>"111101111",
  29049=>"000111000",
  29050=>"001100011",
  29051=>"110100100",
  29052=>"000001000",
  29053=>"011111000",
  29054=>"111000010",
  29055=>"110110011",
  29056=>"110001110",
  29057=>"001110111",
  29058=>"101001011",
  29059=>"000010000",
  29060=>"011110001",
  29061=>"011000010",
  29062=>"100010010",
  29063=>"000000110",
  29064=>"000010011",
  29065=>"101111111",
  29066=>"011001110",
  29067=>"100100001",
  29068=>"100011110",
  29069=>"111011000",
  29070=>"011010010",
  29071=>"101010101",
  29072=>"001010011",
  29073=>"001101111",
  29074=>"101011011",
  29075=>"011111001",
  29076=>"110101011",
  29077=>"001001100",
  29078=>"000110111",
  29079=>"110001110",
  29080=>"101010010",
  29081=>"100001100",
  29082=>"100110001",
  29083=>"001011100",
  29084=>"100000111",
  29085=>"000100000",
  29086=>"111011111",
  29087=>"111000001",
  29088=>"110111010",
  29089=>"011000000",
  29090=>"010101001",
  29091=>"100001111",
  29092=>"011111001",
  29093=>"010001011",
  29094=>"101000000",
  29095=>"011000110",
  29096=>"101011111",
  29097=>"111110101",
  29098=>"100111111",
  29099=>"011101110",
  29100=>"011001100",
  29101=>"111001100",
  29102=>"100111001",
  29103=>"000001001",
  29104=>"000100110",
  29105=>"101111110",
  29106=>"100000010",
  29107=>"101100011",
  29108=>"110000100",
  29109=>"000111010",
  29110=>"110111111",
  29111=>"111001001",
  29112=>"000111000",
  29113=>"010011110",
  29114=>"010110111",
  29115=>"100110000",
  29116=>"111000000",
  29117=>"011001010",
  29118=>"001001010",
  29119=>"001011000",
  29120=>"110101000",
  29121=>"110000000",
  29122=>"000110110",
  29123=>"001010000",
  29124=>"011100110",
  29125=>"101111100",
  29126=>"010010111",
  29127=>"000101001",
  29128=>"111001101",
  29129=>"000100111",
  29130=>"111100111",
  29131=>"100101000",
  29132=>"001111100",
  29133=>"010010000",
  29134=>"101001111",
  29135=>"100010110",
  29136=>"100011011",
  29137=>"011010010",
  29138=>"110100101",
  29139=>"000011110",
  29140=>"100000011",
  29141=>"011010000",
  29142=>"101111000",
  29143=>"110000000",
  29144=>"010010001",
  29145=>"100010010",
  29146=>"111010011",
  29147=>"100010010",
  29148=>"011001011",
  29149=>"110100010",
  29150=>"001110001",
  29151=>"110010101",
  29152=>"000000111",
  29153=>"000011011",
  29154=>"011100101",
  29155=>"100010100",
  29156=>"100001101",
  29157=>"000100111",
  29158=>"001010000",
  29159=>"110010100",
  29160=>"011101000",
  29161=>"011111101",
  29162=>"111111011",
  29163=>"001110001",
  29164=>"000111001",
  29165=>"111110101",
  29166=>"011010111",
  29167=>"000001110",
  29168=>"001101010",
  29169=>"101000010",
  29170=>"011001010",
  29171=>"100000111",
  29172=>"110100110",
  29173=>"001011011",
  29174=>"110110110",
  29175=>"010000101",
  29176=>"011011100",
  29177=>"001100001",
  29178=>"100000010",
  29179=>"111110100",
  29180=>"010011111",
  29181=>"111111110",
  29182=>"111111111",
  29183=>"100001111",
  29184=>"001101110",
  29185=>"001111111",
  29186=>"000101101",
  29187=>"101111011",
  29188=>"101101100",
  29189=>"110001111",
  29190=>"011010101",
  29191=>"110000001",
  29192=>"110001111",
  29193=>"011000100",
  29194=>"100111100",
  29195=>"001000011",
  29196=>"111111011",
  29197=>"100001101",
  29198=>"001100111",
  29199=>"000010000",
  29200=>"100001010",
  29201=>"000110001",
  29202=>"001111011",
  29203=>"001110001",
  29204=>"110110001",
  29205=>"010000010",
  29206=>"000110100",
  29207=>"000101101",
  29208=>"001011011",
  29209=>"011111110",
  29210=>"101110000",
  29211=>"100101001",
  29212=>"101101011",
  29213=>"010011000",
  29214=>"001101011",
  29215=>"100101010",
  29216=>"001110001",
  29217=>"110001010",
  29218=>"110100101",
  29219=>"111001000",
  29220=>"000101111",
  29221=>"011011010",
  29222=>"100001010",
  29223=>"000101101",
  29224=>"010010101",
  29225=>"110111101",
  29226=>"100101010",
  29227=>"010001001",
  29228=>"000011011",
  29229=>"000101001",
  29230=>"111111011",
  29231=>"000001011",
  29232=>"110010101",
  29233=>"110111111",
  29234=>"010110011",
  29235=>"100000101",
  29236=>"001000011",
  29237=>"000100000",
  29238=>"100000010",
  29239=>"101111010",
  29240=>"001010100",
  29241=>"111101010",
  29242=>"011110111",
  29243=>"110100101",
  29244=>"100011011",
  29245=>"110101110",
  29246=>"101000001",
  29247=>"100010010",
  29248=>"001111011",
  29249=>"101010100",
  29250=>"111001010",
  29251=>"000001000",
  29252=>"101100100",
  29253=>"000111111",
  29254=>"100100011",
  29255=>"111110110",
  29256=>"001011111",
  29257=>"001111000",
  29258=>"011000010",
  29259=>"011111101",
  29260=>"000011100",
  29261=>"101110010",
  29262=>"010100010",
  29263=>"000111010",
  29264=>"111101110",
  29265=>"110000110",
  29266=>"110100010",
  29267=>"110001001",
  29268=>"110010010",
  29269=>"011101111",
  29270=>"011111100",
  29271=>"011011110",
  29272=>"110001011",
  29273=>"111100111",
  29274=>"000111010",
  29275=>"110000010",
  29276=>"010110001",
  29277=>"000111011",
  29278=>"111111011",
  29279=>"101100111",
  29280=>"010001111",
  29281=>"000011011",
  29282=>"010010000",
  29283=>"000010010",
  29284=>"110100110",
  29285=>"111000010",
  29286=>"010000111",
  29287=>"111111001",
  29288=>"001111010",
  29289=>"100110111",
  29290=>"000001001",
  29291=>"100110100",
  29292=>"010110110",
  29293=>"010101011",
  29294=>"111011111",
  29295=>"100011111",
  29296=>"011001000",
  29297=>"011101001",
  29298=>"000011000",
  29299=>"111010001",
  29300=>"010001010",
  29301=>"001111001",
  29302=>"100100111",
  29303=>"010000010",
  29304=>"010101000",
  29305=>"101111111",
  29306=>"110100100",
  29307=>"011011001",
  29308=>"011100010",
  29309=>"100001011",
  29310=>"110101100",
  29311=>"011011010",
  29312=>"001100110",
  29313=>"100100110",
  29314=>"001111110",
  29315=>"010011000",
  29316=>"111010110",
  29317=>"111000110",
  29318=>"110010001",
  29319=>"011000111",
  29320=>"001001011",
  29321=>"001101101",
  29322=>"110010000",
  29323=>"010010001",
  29324=>"100011101",
  29325=>"110111101",
  29326=>"001111101",
  29327=>"111001110",
  29328=>"001011010",
  29329=>"000100100",
  29330=>"001111110",
  29331=>"111111011",
  29332=>"100011000",
  29333=>"111001101",
  29334=>"100100011",
  29335=>"001000100",
  29336=>"111011011",
  29337=>"110001001",
  29338=>"011010100",
  29339=>"100001000",
  29340=>"100101011",
  29341=>"101111100",
  29342=>"101000000",
  29343=>"001101000",
  29344=>"000000001",
  29345=>"111010010",
  29346=>"010101100",
  29347=>"001101110",
  29348=>"010011000",
  29349=>"101111101",
  29350=>"110000111",
  29351=>"110111000",
  29352=>"110011011",
  29353=>"100100100",
  29354=>"011100101",
  29355=>"001000000",
  29356=>"111011111",
  29357=>"110111100",
  29358=>"001001110",
  29359=>"000110000",
  29360=>"010001001",
  29361=>"000001111",
  29362=>"000111000",
  29363=>"011100100",
  29364=>"111011110",
  29365=>"011110100",
  29366=>"001011101",
  29367=>"000111101",
  29368=>"111011111",
  29369=>"010101100",
  29370=>"011001010",
  29371=>"010000100",
  29372=>"000010010",
  29373=>"011010101",
  29374=>"000011010",
  29375=>"100111001",
  29376=>"101001101",
  29377=>"111010010",
  29378=>"010001001",
  29379=>"001101100",
  29380=>"000011001",
  29381=>"001110110",
  29382=>"111010110",
  29383=>"100010100",
  29384=>"000100011",
  29385=>"011101001",
  29386=>"100001000",
  29387=>"111111110",
  29388=>"111101001",
  29389=>"010001011",
  29390=>"000111111",
  29391=>"010000010",
  29392=>"101100101",
  29393=>"011001100",
  29394=>"110010011",
  29395=>"000110011",
  29396=>"100110100",
  29397=>"110001110",
  29398=>"100010100",
  29399=>"011010110",
  29400=>"101100001",
  29401=>"111010101",
  29402=>"010100111",
  29403=>"101010010",
  29404=>"111110000",
  29405=>"110000110",
  29406=>"100101001",
  29407=>"010110000",
  29408=>"100100010",
  29409=>"000001011",
  29410=>"111101010",
  29411=>"000011110",
  29412=>"101001001",
  29413=>"110100100",
  29414=>"000110110",
  29415=>"001101010",
  29416=>"011011101",
  29417=>"110010011",
  29418=>"000011001",
  29419=>"010001001",
  29420=>"110111110",
  29421=>"000110011",
  29422=>"100000010",
  29423=>"010111010",
  29424=>"010010111",
  29425=>"111101010",
  29426=>"011101001",
  29427=>"101100010",
  29428=>"000000101",
  29429=>"101010101",
  29430=>"011000100",
  29431=>"001010011",
  29432=>"111110010",
  29433=>"111000010",
  29434=>"011010001",
  29435=>"100100011",
  29436=>"101110000",
  29437=>"111011110",
  29438=>"110101011",
  29439=>"001101010",
  29440=>"101110110",
  29441=>"010111010",
  29442=>"100110101",
  29443=>"010101000",
  29444=>"011111100",
  29445=>"111101000",
  29446=>"101011110",
  29447=>"100001011",
  29448=>"100110011",
  29449=>"010100111",
  29450=>"010000111",
  29451=>"111110100",
  29452=>"110101110",
  29453=>"000111010",
  29454=>"100100011",
  29455=>"100100110",
  29456=>"110010110",
  29457=>"011101111",
  29458=>"100101100",
  29459=>"000011001",
  29460=>"101010101",
  29461=>"011010000",
  29462=>"100100110",
  29463=>"100101100",
  29464=>"110100111",
  29465=>"010001000",
  29466=>"101010100",
  29467=>"010000100",
  29468=>"010011111",
  29469=>"010011100",
  29470=>"100011110",
  29471=>"000101100",
  29472=>"111101101",
  29473=>"001001101",
  29474=>"111110111",
  29475=>"110110100",
  29476=>"010000010",
  29477=>"101110111",
  29478=>"011000000",
  29479=>"010000010",
  29480=>"101000101",
  29481=>"001110010",
  29482=>"100100101",
  29483=>"011000000",
  29484=>"001110010",
  29485=>"010100000",
  29486=>"100000001",
  29487=>"110010010",
  29488=>"111101111",
  29489=>"011010100",
  29490=>"000100010",
  29491=>"001111111",
  29492=>"000100111",
  29493=>"010111110",
  29494=>"110001110",
  29495=>"001010111",
  29496=>"111111100",
  29497=>"100000100",
  29498=>"010000001",
  29499=>"100011000",
  29500=>"101001000",
  29501=>"000111100",
  29502=>"000101011",
  29503=>"010101111",
  29504=>"011001111",
  29505=>"101111000",
  29506=>"011101110",
  29507=>"100000010",
  29508=>"101110000",
  29509=>"111011011",
  29510=>"100101101",
  29511=>"111110101",
  29512=>"000000001",
  29513=>"111100100",
  29514=>"011000011",
  29515=>"011010101",
  29516=>"001000001",
  29517=>"000011111",
  29518=>"000100110",
  29519=>"011100001",
  29520=>"101101110",
  29521=>"010101101",
  29522=>"011101010",
  29523=>"000010011",
  29524=>"001101001",
  29525=>"111101011",
  29526=>"111101111",
  29527=>"000000011",
  29528=>"111111101",
  29529=>"100010101",
  29530=>"000000011",
  29531=>"111110101",
  29532=>"001010011",
  29533=>"110000100",
  29534=>"010101001",
  29535=>"110100101",
  29536=>"011000011",
  29537=>"000101000",
  29538=>"111100111",
  29539=>"110111010",
  29540=>"101011110",
  29541=>"011110001",
  29542=>"111000000",
  29543=>"000000001",
  29544=>"110110101",
  29545=>"011101000",
  29546=>"010100100",
  29547=>"101111011",
  29548=>"001111100",
  29549=>"010000010",
  29550=>"110001010",
  29551=>"100001100",
  29552=>"110101010",
  29553=>"001100001",
  29554=>"011111011",
  29555=>"010100100",
  29556=>"100110110",
  29557=>"110011000",
  29558=>"101011101",
  29559=>"110001000",
  29560=>"010011000",
  29561=>"100011010",
  29562=>"100110111",
  29563=>"100000010",
  29564=>"000011101",
  29565=>"111101000",
  29566=>"000010101",
  29567=>"101101011",
  29568=>"000011001",
  29569=>"000010100",
  29570=>"010111001",
  29571=>"000010010",
  29572=>"110111111",
  29573=>"011010111",
  29574=>"101110110",
  29575=>"010011110",
  29576=>"100011001",
  29577=>"010000111",
  29578=>"110100010",
  29579=>"111010111",
  29580=>"110000101",
  29581=>"111111110",
  29582=>"010011100",
  29583=>"110110101",
  29584=>"100000010",
  29585=>"010000001",
  29586=>"000100011",
  29587=>"101010001",
  29588=>"101001011",
  29589=>"000000000",
  29590=>"100111010",
  29591=>"110000001",
  29592=>"011101000",
  29593=>"000001011",
  29594=>"000011110",
  29595=>"101101001",
  29596=>"000111000",
  29597=>"000110100",
  29598=>"110000000",
  29599=>"001011010",
  29600=>"000001110",
  29601=>"010100000",
  29602=>"011001110",
  29603=>"110100000",
  29604=>"100010110",
  29605=>"110101000",
  29606=>"101010100",
  29607=>"101001110",
  29608=>"100010100",
  29609=>"000001100",
  29610=>"011110101",
  29611=>"000100101",
  29612=>"001000110",
  29613=>"001111011",
  29614=>"111110000",
  29615=>"001101110",
  29616=>"001111110",
  29617=>"000110110",
  29618=>"100100100",
  29619=>"011001000",
  29620=>"111111111",
  29621=>"010000001",
  29622=>"101001111",
  29623=>"110001001",
  29624=>"111100101",
  29625=>"010010011",
  29626=>"111100101",
  29627=>"011011100",
  29628=>"101101100",
  29629=>"010100110",
  29630=>"011100101",
  29631=>"110110100",
  29632=>"000100001",
  29633=>"011110111",
  29634=>"101101001",
  29635=>"011001000",
  29636=>"111111101",
  29637=>"010111001",
  29638=>"011101000",
  29639=>"011101100",
  29640=>"101010100",
  29641=>"011000011",
  29642=>"111100010",
  29643=>"111010101",
  29644=>"010100001",
  29645=>"100110100",
  29646=>"101001100",
  29647=>"100111110",
  29648=>"000101111",
  29649=>"111011011",
  29650=>"110011000",
  29651=>"000010010",
  29652=>"111111011",
  29653=>"001010011",
  29654=>"100001000",
  29655=>"010111101",
  29656=>"110001101",
  29657=>"011011010",
  29658=>"001011000",
  29659=>"001100011",
  29660=>"010000101",
  29661=>"101111010",
  29662=>"001001110",
  29663=>"000110010",
  29664=>"110011001",
  29665=>"011011001",
  29666=>"101100001",
  29667=>"001000111",
  29668=>"110010000",
  29669=>"100110011",
  29670=>"111000101",
  29671=>"011010010",
  29672=>"010111100",
  29673=>"010100100",
  29674=>"001111100",
  29675=>"000000100",
  29676=>"101010000",
  29677=>"100001100",
  29678=>"111011000",
  29679=>"000111010",
  29680=>"110011111",
  29681=>"010100101",
  29682=>"110110001",
  29683=>"110100011",
  29684=>"111110011",
  29685=>"000011000",
  29686=>"011011100",
  29687=>"111110111",
  29688=>"111111100",
  29689=>"111001000",
  29690=>"110100111",
  29691=>"101101000",
  29692=>"001111101",
  29693=>"001011101",
  29694=>"101011010",
  29695=>"101001011",
  29696=>"101101101",
  29697=>"000010110",
  29698=>"110110011",
  29699=>"000101111",
  29700=>"110010100",
  29701=>"111111110",
  29702=>"110010110",
  29703=>"010000110",
  29704=>"000100111",
  29705=>"010110101",
  29706=>"011100011",
  29707=>"010011111",
  29708=>"101000100",
  29709=>"110110000",
  29710=>"110101101",
  29711=>"000010101",
  29712=>"011011000",
  29713=>"010111101",
  29714=>"100010101",
  29715=>"000000001",
  29716=>"001001010",
  29717=>"111100110",
  29718=>"010010010",
  29719=>"011100110",
  29720=>"110011100",
  29721=>"000001000",
  29722=>"100010011",
  29723=>"001101100",
  29724=>"100011011",
  29725=>"000100000",
  29726=>"001011011",
  29727=>"100101010",
  29728=>"101000000",
  29729=>"100010001",
  29730=>"111011000",
  29731=>"000000011",
  29732=>"011110000",
  29733=>"001111111",
  29734=>"100001011",
  29735=>"100010000",
  29736=>"110110000",
  29737=>"000101000",
  29738=>"111101110",
  29739=>"101100000",
  29740=>"000011011",
  29741=>"010011101",
  29742=>"110010100",
  29743=>"111100000",
  29744=>"001001001",
  29745=>"101000101",
  29746=>"100011001",
  29747=>"010101011",
  29748=>"000000010",
  29749=>"111001011",
  29750=>"011001110",
  29751=>"001101010",
  29752=>"001100111",
  29753=>"111111111",
  29754=>"000110001",
  29755=>"100111110",
  29756=>"110001000",
  29757=>"010011000",
  29758=>"111111000",
  29759=>"100001010",
  29760=>"010101000",
  29761=>"100010001",
  29762=>"110001001",
  29763=>"111101101",
  29764=>"100100111",
  29765=>"110111010",
  29766=>"100000010",
  29767=>"110101011",
  29768=>"011011000",
  29769=>"101010111",
  29770=>"110011101",
  29771=>"001011110",
  29772=>"010000010",
  29773=>"111001110",
  29774=>"100101110",
  29775=>"011001110",
  29776=>"100101101",
  29777=>"000111110",
  29778=>"110111100",
  29779=>"101000000",
  29780=>"101111001",
  29781=>"001010001",
  29782=>"010000001",
  29783=>"000101001",
  29784=>"100100010",
  29785=>"001000010",
  29786=>"100011111",
  29787=>"001000011",
  29788=>"100100011",
  29789=>"100101010",
  29790=>"110101101",
  29791=>"111001010",
  29792=>"000010111",
  29793=>"111100000",
  29794=>"100100000",
  29795=>"110100000",
  29796=>"001110111",
  29797=>"111011111",
  29798=>"101011011",
  29799=>"111101000",
  29800=>"110111011",
  29801=>"100011111",
  29802=>"011000000",
  29803=>"111000011",
  29804=>"000110011",
  29805=>"111000101",
  29806=>"000101001",
  29807=>"011111111",
  29808=>"110000010",
  29809=>"010011000",
  29810=>"000001110",
  29811=>"100101000",
  29812=>"011101111",
  29813=>"101000111",
  29814=>"100111011",
  29815=>"000000010",
  29816=>"110010011",
  29817=>"000010010",
  29818=>"100100000",
  29819=>"011110110",
  29820=>"011100000",
  29821=>"110110100",
  29822=>"101010011",
  29823=>"011011010",
  29824=>"110000001",
  29825=>"010011000",
  29826=>"000111101",
  29827=>"011010011",
  29828=>"101001011",
  29829=>"110111111",
  29830=>"100101101",
  29831=>"011001101",
  29832=>"110111101",
  29833=>"001111100",
  29834=>"100010111",
  29835=>"010001111",
  29836=>"011111111",
  29837=>"110111010",
  29838=>"111010111",
  29839=>"000101001",
  29840=>"010011000",
  29841=>"110101111",
  29842=>"100101100",
  29843=>"111001100",
  29844=>"010100000",
  29845=>"110110111",
  29846=>"101000110",
  29847=>"100110011",
  29848=>"000100111",
  29849=>"000001010",
  29850=>"011000101",
  29851=>"110000000",
  29852=>"001100111",
  29853=>"110010100",
  29854=>"011110101",
  29855=>"111001010",
  29856=>"000100010",
  29857=>"010110111",
  29858=>"000101110",
  29859=>"000101111",
  29860=>"010000101",
  29861=>"011101001",
  29862=>"110010000",
  29863=>"111011111",
  29864=>"110011010",
  29865=>"010011010",
  29866=>"000001111",
  29867=>"011000010",
  29868=>"001001011",
  29869=>"000111111",
  29870=>"111111010",
  29871=>"001101000",
  29872=>"001110001",
  29873=>"100100010",
  29874=>"000010000",
  29875=>"010000111",
  29876=>"100101010",
  29877=>"001101100",
  29878=>"011110100",
  29879=>"110110010",
  29880=>"110111100",
  29881=>"101001011",
  29882=>"011111011",
  29883=>"010010001",
  29884=>"001000001",
  29885=>"101011010",
  29886=>"111001100",
  29887=>"111001001",
  29888=>"010011100",
  29889=>"000101000",
  29890=>"001011001",
  29891=>"111110001",
  29892=>"110000010",
  29893=>"001110011",
  29894=>"010111110",
  29895=>"110100110",
  29896=>"000111100",
  29897=>"110100101",
  29898=>"111110111",
  29899=>"011101011",
  29900=>"001001001",
  29901=>"111111100",
  29902=>"000011111",
  29903=>"110010101",
  29904=>"001110100",
  29905=>"001100110",
  29906=>"100000100",
  29907=>"000111011",
  29908=>"100110101",
  29909=>"010001011",
  29910=>"010111011",
  29911=>"011010000",
  29912=>"101011010",
  29913=>"101111100",
  29914=>"110110011",
  29915=>"000111010",
  29916=>"000010011",
  29917=>"110001011",
  29918=>"011001011",
  29919=>"100000010",
  29920=>"111100111",
  29921=>"100000011",
  29922=>"010111110",
  29923=>"001111000",
  29924=>"110010111",
  29925=>"000100011",
  29926=>"110110110",
  29927=>"100110001",
  29928=>"010100011",
  29929=>"011110010",
  29930=>"101111111",
  29931=>"110001111",
  29932=>"011110011",
  29933=>"000101011",
  29934=>"000100010",
  29935=>"100111111",
  29936=>"011000100",
  29937=>"000110000",
  29938=>"011111101",
  29939=>"100001010",
  29940=>"000101001",
  29941=>"100101000",
  29942=>"011011000",
  29943=>"100010111",
  29944=>"011010011",
  29945=>"101011010",
  29946=>"011011001",
  29947=>"111001000",
  29948=>"010100010",
  29949=>"001001111",
  29950=>"110011100",
  29951=>"000100001",
  29952=>"001011101",
  29953=>"010010010",
  29954=>"010000101",
  29955=>"100110001",
  29956=>"010000111",
  29957=>"111011000",
  29958=>"000001110",
  29959=>"101100000",
  29960=>"011111111",
  29961=>"001011111",
  29962=>"001101001",
  29963=>"000100101",
  29964=>"011011000",
  29965=>"101110000",
  29966=>"100111001",
  29967=>"000111101",
  29968=>"001100111",
  29969=>"101000101",
  29970=>"001100100",
  29971=>"010000101",
  29972=>"110111001",
  29973=>"011000000",
  29974=>"000011000",
  29975=>"100010000",
  29976=>"000111110",
  29977=>"111011000",
  29978=>"011001111",
  29979=>"100000001",
  29980=>"010010111",
  29981=>"110100100",
  29982=>"001100100",
  29983=>"000100001",
  29984=>"001001011",
  29985=>"011111001",
  29986=>"000100101",
  29987=>"110100010",
  29988=>"000101010",
  29989=>"111010011",
  29990=>"110110100",
  29991=>"111111100",
  29992=>"010100001",
  29993=>"110011010",
  29994=>"101001111",
  29995=>"101110001",
  29996=>"111001000",
  29997=>"000111011",
  29998=>"100001100",
  29999=>"001100100",
  30000=>"011111001",
  30001=>"100100000",
  30002=>"101010110",
  30003=>"101010111",
  30004=>"110000110",
  30005=>"101101110",
  30006=>"010000110",
  30007=>"111111110",
  30008=>"100110111",
  30009=>"101000011",
  30010=>"100101110",
  30011=>"111101110",
  30012=>"111010011",
  30013=>"000101000",
  30014=>"010011100",
  30015=>"111101011",
  30016=>"111000000",
  30017=>"100000011",
  30018=>"001011101",
  30019=>"011011001",
  30020=>"001000100",
  30021=>"010010111",
  30022=>"110110001",
  30023=>"101100010",
  30024=>"111011000",
  30025=>"010011101",
  30026=>"111001010",
  30027=>"001011010",
  30028=>"101111000",
  30029=>"010101110",
  30030=>"101100111",
  30031=>"011001100",
  30032=>"000000001",
  30033=>"111011101",
  30034=>"000100111",
  30035=>"111011000",
  30036=>"100001101",
  30037=>"111011000",
  30038=>"111010110",
  30039=>"101100110",
  30040=>"110000101",
  30041=>"110111101",
  30042=>"010000000",
  30043=>"000101101",
  30044=>"000011111",
  30045=>"111011100",
  30046=>"111011010",
  30047=>"110101111",
  30048=>"111110000",
  30049=>"011010110",
  30050=>"010001010",
  30051=>"111110100",
  30052=>"100000111",
  30053=>"000010111",
  30054=>"011110001",
  30055=>"110011101",
  30056=>"001101111",
  30057=>"101000001",
  30058=>"010110110",
  30059=>"000111011",
  30060=>"001011100",
  30061=>"011100011",
  30062=>"101000101",
  30063=>"011011100",
  30064=>"001100000",
  30065=>"011000111",
  30066=>"001111111",
  30067=>"101101111",
  30068=>"110101101",
  30069=>"000100100",
  30070=>"011001100",
  30071=>"110110100",
  30072=>"001111001",
  30073=>"000111110",
  30074=>"101100111",
  30075=>"010110011",
  30076=>"111101000",
  30077=>"111000101",
  30078=>"001001010",
  30079=>"110110000",
  30080=>"111010011",
  30081=>"001011100",
  30082=>"001110100",
  30083=>"001110011",
  30084=>"111000011",
  30085=>"001011100",
  30086=>"000001110",
  30087=>"000101010",
  30088=>"101100110",
  30089=>"000011111",
  30090=>"011010010",
  30091=>"001010000",
  30092=>"101000111",
  30093=>"001001010",
  30094=>"110101111",
  30095=>"100010101",
  30096=>"110110001",
  30097=>"000011011",
  30098=>"101001101",
  30099=>"101101110",
  30100=>"100011001",
  30101=>"000000111",
  30102=>"101011101",
  30103=>"011111111",
  30104=>"001000010",
  30105=>"010000100",
  30106=>"100100011",
  30107=>"000101100",
  30108=>"101011010",
  30109=>"010011100",
  30110=>"111100110",
  30111=>"111111110",
  30112=>"000001101",
  30113=>"000101010",
  30114=>"101110000",
  30115=>"110000000",
  30116=>"011100110",
  30117=>"110111100",
  30118=>"011011011",
  30119=>"000000000",
  30120=>"000100111",
  30121=>"010110001",
  30122=>"100101100",
  30123=>"100010000",
  30124=>"100000010",
  30125=>"000001110",
  30126=>"000101100",
  30127=>"011111110",
  30128=>"000000000",
  30129=>"000011100",
  30130=>"000100010",
  30131=>"011100101",
  30132=>"010110001",
  30133=>"110000011",
  30134=>"100101101",
  30135=>"101011001",
  30136=>"101001100",
  30137=>"010101010",
  30138=>"011101110",
  30139=>"010110000",
  30140=>"110011010",
  30141=>"100001101",
  30142=>"010000011",
  30143=>"101111001",
  30144=>"000000000",
  30145=>"101010100",
  30146=>"010001101",
  30147=>"111011000",
  30148=>"011001100",
  30149=>"101000001",
  30150=>"101010110",
  30151=>"111000111",
  30152=>"101010110",
  30153=>"000101110",
  30154=>"111001101",
  30155=>"000010000",
  30156=>"001010110",
  30157=>"001000001",
  30158=>"010011011",
  30159=>"111110101",
  30160=>"110111101",
  30161=>"111111110",
  30162=>"001011101",
  30163=>"111101100",
  30164=>"011010101",
  30165=>"111101000",
  30166=>"111011000",
  30167=>"100000100",
  30168=>"101110110",
  30169=>"000100111",
  30170=>"010100011",
  30171=>"110111000",
  30172=>"010100100",
  30173=>"111111111",
  30174=>"110111101",
  30175=>"000010111",
  30176=>"101101100",
  30177=>"111010101",
  30178=>"100100110",
  30179=>"001100101",
  30180=>"011001100",
  30181=>"001011000",
  30182=>"111010100",
  30183=>"010110000",
  30184=>"001011010",
  30185=>"001010110",
  30186=>"000010110",
  30187=>"101101010",
  30188=>"010010000",
  30189=>"110101001",
  30190=>"110000100",
  30191=>"100110000",
  30192=>"000001010",
  30193=>"011011001",
  30194=>"010101000",
  30195=>"010111001",
  30196=>"011111110",
  30197=>"011010001",
  30198=>"101010111",
  30199=>"010001001",
  30200=>"111001100",
  30201=>"001001111",
  30202=>"010001110",
  30203=>"010110010",
  30204=>"110111010",
  30205=>"111101111",
  30206=>"001110111",
  30207=>"000010110",
  30208=>"001111011",
  30209=>"110101011",
  30210=>"010010000",
  30211=>"001010101",
  30212=>"001100011",
  30213=>"010100100",
  30214=>"100111011",
  30215=>"100001101",
  30216=>"010110011",
  30217=>"000100000",
  30218=>"000100001",
  30219=>"100011111",
  30220=>"010001010",
  30221=>"110111011",
  30222=>"000011000",
  30223=>"001101010",
  30224=>"010011111",
  30225=>"111011000",
  30226=>"011110111",
  30227=>"000100011",
  30228=>"101110001",
  30229=>"010101110",
  30230=>"101001000",
  30231=>"100101011",
  30232=>"001001000",
  30233=>"010101010",
  30234=>"001001000",
  30235=>"001100110",
  30236=>"111110011",
  30237=>"011010101",
  30238=>"101100101",
  30239=>"110111000",
  30240=>"010001001",
  30241=>"111100011",
  30242=>"001101001",
  30243=>"001101110",
  30244=>"101110110",
  30245=>"011100000",
  30246=>"101001010",
  30247=>"001001110",
  30248=>"100010011",
  30249=>"101101010",
  30250=>"010011001",
  30251=>"101000100",
  30252=>"111001111",
  30253=>"101100110",
  30254=>"111111001",
  30255=>"010101011",
  30256=>"101111010",
  30257=>"001100010",
  30258=>"010111000",
  30259=>"000101110",
  30260=>"001101000",
  30261=>"110010011",
  30262=>"110101100",
  30263=>"010100111",
  30264=>"100001111",
  30265=>"110110110",
  30266=>"110101101",
  30267=>"011110010",
  30268=>"111011101",
  30269=>"000100011",
  30270=>"111101101",
  30271=>"100000000",
  30272=>"001011101",
  30273=>"011011101",
  30274=>"000110011",
  30275=>"100100100",
  30276=>"001001010",
  30277=>"001011010",
  30278=>"010110011",
  30279=>"001111000",
  30280=>"111011111",
  30281=>"011101101",
  30282=>"101110101",
  30283=>"010110010",
  30284=>"001110000",
  30285=>"100100010",
  30286=>"101010000",
  30287=>"111011110",
  30288=>"100010101",
  30289=>"010101011",
  30290=>"100101000",
  30291=>"010011100",
  30292=>"010000101",
  30293=>"000010001",
  30294=>"000100010",
  30295=>"110010100",
  30296=>"010100100",
  30297=>"010111011",
  30298=>"110111111",
  30299=>"111001011",
  30300=>"011101010",
  30301=>"101101110",
  30302=>"110000010",
  30303=>"000111111",
  30304=>"001100010",
  30305=>"000001000",
  30306=>"010111110",
  30307=>"111101011",
  30308=>"000101101",
  30309=>"100101111",
  30310=>"110100111",
  30311=>"100010101",
  30312=>"100010111",
  30313=>"011100010",
  30314=>"100010011",
  30315=>"110000001",
  30316=>"100110000",
  30317=>"010111111",
  30318=>"011110101",
  30319=>"101101010",
  30320=>"111100011",
  30321=>"111110000",
  30322=>"101101001",
  30323=>"010111101",
  30324=>"001111010",
  30325=>"111110000",
  30326=>"000100010",
  30327=>"111101111",
  30328=>"000110111",
  30329=>"110100011",
  30330=>"011110010",
  30331=>"111111011",
  30332=>"000000110",
  30333=>"110111011",
  30334=>"111100100",
  30335=>"101011000",
  30336=>"001010010",
  30337=>"011010001",
  30338=>"001110010",
  30339=>"111101111",
  30340=>"010001011",
  30341=>"010100111",
  30342=>"010000100",
  30343=>"111010010",
  30344=>"101011001",
  30345=>"100001101",
  30346=>"111111101",
  30347=>"010000001",
  30348=>"100010000",
  30349=>"001101100",
  30350=>"010000010",
  30351=>"110000010",
  30352=>"110011111",
  30353=>"000110000",
  30354=>"011101010",
  30355=>"100111100",
  30356=>"010001011",
  30357=>"001010001",
  30358=>"010000000",
  30359=>"001000000",
  30360=>"100110100",
  30361=>"010111001",
  30362=>"010110101",
  30363=>"101011010",
  30364=>"101111001",
  30365=>"011010001",
  30366=>"001101111",
  30367=>"001111110",
  30368=>"000001101",
  30369=>"010111110",
  30370=>"101101001",
  30371=>"011111111",
  30372=>"000010010",
  30373=>"001000110",
  30374=>"101011000",
  30375=>"101111110",
  30376=>"101000101",
  30377=>"101000000",
  30378=>"111000011",
  30379=>"001111110",
  30380=>"111011011",
  30381=>"000100100",
  30382=>"100101001",
  30383=>"000001110",
  30384=>"111011100",
  30385=>"101010010",
  30386=>"010100101",
  30387=>"000110000",
  30388=>"111011111",
  30389=>"001000010",
  30390=>"111101000",
  30391=>"111101010",
  30392=>"000011011",
  30393=>"111100111",
  30394=>"001100010",
  30395=>"101000110",
  30396=>"010010100",
  30397=>"001001001",
  30398=>"001000001",
  30399=>"101101100",
  30400=>"011101010",
  30401=>"011110100",
  30402=>"101101100",
  30403=>"000100101",
  30404=>"010111011",
  30405=>"111111101",
  30406=>"111101010",
  30407=>"000010010",
  30408=>"000111100",
  30409=>"000110100",
  30410=>"111100100",
  30411=>"001011000",
  30412=>"011001110",
  30413=>"010001000",
  30414=>"111111001",
  30415=>"001111001",
  30416=>"001110011",
  30417=>"111001110",
  30418=>"100001100",
  30419=>"011010111",
  30420=>"010111000",
  30421=>"111010010",
  30422=>"001110010",
  30423=>"001101101",
  30424=>"000001000",
  30425=>"110010101",
  30426=>"101010011",
  30427=>"001111000",
  30428=>"000010001",
  30429=>"110110010",
  30430=>"100000010",
  30431=>"101101001",
  30432=>"110110110",
  30433=>"100010000",
  30434=>"110100100",
  30435=>"111111100",
  30436=>"100010001",
  30437=>"010001000",
  30438=>"101110000",
  30439=>"101001001",
  30440=>"100001110",
  30441=>"000010100",
  30442=>"111111001",
  30443=>"010001011",
  30444=>"001000110",
  30445=>"010001010",
  30446=>"101111110",
  30447=>"011001100",
  30448=>"000001110",
  30449=>"010110001",
  30450=>"000100010",
  30451=>"000001100",
  30452=>"111100110",
  30453=>"010101010",
  30454=>"000100101",
  30455=>"100110101",
  30456=>"001001010",
  30457=>"000010110",
  30458=>"001011111",
  30459=>"101001001",
  30460=>"011011001",
  30461=>"110001110",
  30462=>"100001011",
  30463=>"100100110",
  30464=>"000000100",
  30465=>"110011001",
  30466=>"100110001",
  30467=>"010101111",
  30468=>"101011001",
  30469=>"111010110",
  30470=>"011110001",
  30471=>"100000000",
  30472=>"011101010",
  30473=>"110010111",
  30474=>"011100110",
  30475=>"001100011",
  30476=>"100000000",
  30477=>"101001010",
  30478=>"011000110",
  30479=>"101010100",
  30480=>"100101101",
  30481=>"011110111",
  30482=>"110100100",
  30483=>"010011011",
  30484=>"100011100",
  30485=>"001011100",
  30486=>"100110011",
  30487=>"110111010",
  30488=>"011001001",
  30489=>"111001000",
  30490=>"001001000",
  30491=>"111111110",
  30492=>"110101001",
  30493=>"110101100",
  30494=>"100010101",
  30495=>"110011001",
  30496=>"000001101",
  30497=>"011000101",
  30498=>"001110000",
  30499=>"111001000",
  30500=>"000001000",
  30501=>"001001011",
  30502=>"110111010",
  30503=>"010100110",
  30504=>"001110101",
  30505=>"110111010",
  30506=>"001110010",
  30507=>"000110110",
  30508=>"101101010",
  30509=>"000100111",
  30510=>"101010011",
  30511=>"101000110",
  30512=>"001100111",
  30513=>"000101000",
  30514=>"011000100",
  30515=>"100110101",
  30516=>"100000110",
  30517=>"001110011",
  30518=>"001000001",
  30519=>"100000010",
  30520=>"100000010",
  30521=>"001100100",
  30522=>"101100010",
  30523=>"101100011",
  30524=>"111101111",
  30525=>"111001010",
  30526=>"001110111",
  30527=>"111010110",
  30528=>"000100111",
  30529=>"010001111",
  30530=>"101010011",
  30531=>"000111000",
  30532=>"001110000",
  30533=>"011111101",
  30534=>"101100001",
  30535=>"001001100",
  30536=>"111110011",
  30537=>"000110111",
  30538=>"111101011",
  30539=>"000110011",
  30540=>"101111101",
  30541=>"110111100",
  30542=>"101111000",
  30543=>"110000001",
  30544=>"100100111",
  30545=>"101101010",
  30546=>"000111001",
  30547=>"101101001",
  30548=>"010011111",
  30549=>"000001101",
  30550=>"011000101",
  30551=>"101111111",
  30552=>"010110001",
  30553=>"100011000",
  30554=>"100011110",
  30555=>"101010010",
  30556=>"111111100",
  30557=>"111011100",
  30558=>"101110111",
  30559=>"100010110",
  30560=>"011101011",
  30561=>"010010010",
  30562=>"000000100",
  30563=>"010101000",
  30564=>"000010111",
  30565=>"100011011",
  30566=>"111001010",
  30567=>"000111110",
  30568=>"000100011",
  30569=>"011110100",
  30570=>"110111100",
  30571=>"110111110",
  30572=>"001100100",
  30573=>"010001100",
  30574=>"010100100",
  30575=>"001010001",
  30576=>"000000101",
  30577=>"010011101",
  30578=>"111100111",
  30579=>"111000110",
  30580=>"011011001",
  30581=>"111111001",
  30582=>"001010101",
  30583=>"001001111",
  30584=>"101011100",
  30585=>"011000101",
  30586=>"000100001",
  30587=>"000111000",
  30588=>"011100101",
  30589=>"111100010",
  30590=>"010111011",
  30591=>"101010001",
  30592=>"101011011",
  30593=>"010100010",
  30594=>"001111000",
  30595=>"100011011",
  30596=>"000101011",
  30597=>"101101011",
  30598=>"100010100",
  30599=>"001111110",
  30600=>"111011001",
  30601=>"011111110",
  30602=>"001010011",
  30603=>"000010001",
  30604=>"010010101",
  30605=>"111010111",
  30606=>"010100000",
  30607=>"110111100",
  30608=>"110111010",
  30609=>"000110011",
  30610=>"110100110",
  30611=>"000000111",
  30612=>"101001001",
  30613=>"101011101",
  30614=>"001000001",
  30615=>"000011001",
  30616=>"010100101",
  30617=>"000101101",
  30618=>"010101001",
  30619=>"011010001",
  30620=>"111011110",
  30621=>"000011000",
  30622=>"010001000",
  30623=>"001011000",
  30624=>"011000001",
  30625=>"010010100",
  30626=>"010101100",
  30627=>"010010010",
  30628=>"100011101",
  30629=>"011110110",
  30630=>"001000110",
  30631=>"111000001",
  30632=>"011000110",
  30633=>"000011000",
  30634=>"101101101",
  30635=>"111001001",
  30636=>"101001111",
  30637=>"001001110",
  30638=>"110100110",
  30639=>"100001000",
  30640=>"111010010",
  30641=>"010001000",
  30642=>"110001101",
  30643=>"000001011",
  30644=>"111110000",
  30645=>"000001100",
  30646=>"010000011",
  30647=>"001110010",
  30648=>"110011101",
  30649=>"010000000",
  30650=>"100000100",
  30651=>"011000000",
  30652=>"000000000",
  30653=>"100011000",
  30654=>"101100011",
  30655=>"110111100",
  30656=>"110001101",
  30657=>"011000101",
  30658=>"011010000",
  30659=>"100001101",
  30660=>"000000001",
  30661=>"010110101",
  30662=>"111110010",
  30663=>"000010010",
  30664=>"101000100",
  30665=>"010010011",
  30666=>"000001101",
  30667=>"101111010",
  30668=>"101111010",
  30669=>"100000110",
  30670=>"110001011",
  30671=>"111011110",
  30672=>"100010001",
  30673=>"101011101",
  30674=>"001101000",
  30675=>"011010101",
  30676=>"010000001",
  30677=>"110100101",
  30678=>"000110100",
  30679=>"100011111",
  30680=>"111111110",
  30681=>"000111000",
  30682=>"011000001",
  30683=>"011111100",
  30684=>"010010110",
  30685=>"010111100",
  30686=>"001001100",
  30687=>"010000110",
  30688=>"101101011",
  30689=>"110001011",
  30690=>"001001111",
  30691=>"001001001",
  30692=>"001011100",
  30693=>"111011000",
  30694=>"110100001",
  30695=>"100110100",
  30696=>"001000000",
  30697=>"011011001",
  30698=>"110100110",
  30699=>"100000111",
  30700=>"110110001",
  30701=>"000011001",
  30702=>"011100000",
  30703=>"001111001",
  30704=>"001111111",
  30705=>"100111010",
  30706=>"010110110",
  30707=>"001010100",
  30708=>"101110101",
  30709=>"111011011",
  30710=>"000111000",
  30711=>"111111101",
  30712=>"111010111",
  30713=>"101110000",
  30714=>"110111000",
  30715=>"010001011",
  30716=>"000001110",
  30717=>"111110101",
  30718=>"100111101",
  30719=>"101011110",
  30720=>"011001111",
  30721=>"101110110",
  30722=>"010011101",
  30723=>"111110101",
  30724=>"000111101",
  30725=>"010011100",
  30726=>"110010111",
  30727=>"100110000",
  30728=>"100101111",
  30729=>"001111010",
  30730=>"001000001",
  30731=>"111101010",
  30732=>"101111011",
  30733=>"111011011",
  30734=>"111100110",
  30735=>"110110111",
  30736=>"011110011",
  30737=>"111001101",
  30738=>"111011011",
  30739=>"000001100",
  30740=>"000000000",
  30741=>"110110110",
  30742=>"111001110",
  30743=>"011000010",
  30744=>"110110001",
  30745=>"000000010",
  30746=>"000101111",
  30747=>"000110001",
  30748=>"111101111",
  30749=>"011101110",
  30750=>"000011110",
  30751=>"101110100",
  30752=>"000001111",
  30753=>"011101001",
  30754=>"100000010",
  30755=>"101000000",
  30756=>"100110010",
  30757=>"001111100",
  30758=>"111101100",
  30759=>"110010101",
  30760=>"110110000",
  30761=>"001010101",
  30762=>"100111010",
  30763=>"111000110",
  30764=>"000100110",
  30765=>"011111000",
  30766=>"100111101",
  30767=>"101100001",
  30768=>"101011111",
  30769=>"001100100",
  30770=>"010011000",
  30771=>"010011010",
  30772=>"100111001",
  30773=>"010001010",
  30774=>"110100111",
  30775=>"011010111",
  30776=>"111111100",
  30777=>"011011110",
  30778=>"001001111",
  30779=>"100001010",
  30780=>"101110101",
  30781=>"000000001",
  30782=>"000101110",
  30783=>"111100000",
  30784=>"110001010",
  30785=>"100001101",
  30786=>"110100001",
  30787=>"110000110",
  30788=>"000010100",
  30789=>"100100011",
  30790=>"100000101",
  30791=>"100100010",
  30792=>"011110000",
  30793=>"111100110",
  30794=>"000111011",
  30795=>"001110111",
  30796=>"100000011",
  30797=>"010010101",
  30798=>"010011111",
  30799=>"010110110",
  30800=>"111010101",
  30801=>"010001100",
  30802=>"110101000",
  30803=>"001110010",
  30804=>"100011111",
  30805=>"010100110",
  30806=>"000100111",
  30807=>"001010000",
  30808=>"111111110",
  30809=>"100000101",
  30810=>"110111101",
  30811=>"100111001",
  30812=>"001111101",
  30813=>"111001101",
  30814=>"010100001",
  30815=>"110110000",
  30816=>"010000001",
  30817=>"111001001",
  30818=>"001000000",
  30819=>"101100100",
  30820=>"011001010",
  30821=>"100111001",
  30822=>"101100011",
  30823=>"000100101",
  30824=>"111101101",
  30825=>"010001101",
  30826=>"111110110",
  30827=>"001110101",
  30828=>"001110011",
  30829=>"111110100",
  30830=>"111010110",
  30831=>"100111100",
  30832=>"100001010",
  30833=>"001100100",
  30834=>"101000111",
  30835=>"001100010",
  30836=>"010101100",
  30837=>"011011011",
  30838=>"010011011",
  30839=>"010100110",
  30840=>"001100010",
  30841=>"110100010",
  30842=>"111011101",
  30843=>"111000101",
  30844=>"001000011",
  30845=>"110001011",
  30846=>"101101110",
  30847=>"111011111",
  30848=>"001100001",
  30849=>"001110101",
  30850=>"110001110",
  30851=>"010011111",
  30852=>"010111000",
  30853=>"000000101",
  30854=>"110000111",
  30855=>"000001101",
  30856=>"100001110",
  30857=>"110101000",
  30858=>"000101111",
  30859=>"101111111",
  30860=>"111100011",
  30861=>"000000111",
  30862=>"011001111",
  30863=>"110011000",
  30864=>"000000000",
  30865=>"100111010",
  30866=>"001011000",
  30867=>"101100011",
  30868=>"010100111",
  30869=>"001001001",
  30870=>"011001001",
  30871=>"001100111",
  30872=>"100111000",
  30873=>"010010110",
  30874=>"101001010",
  30875=>"000001101",
  30876=>"001110010",
  30877=>"110110010",
  30878=>"010011101",
  30879=>"111010010",
  30880=>"110101111",
  30881=>"010010001",
  30882=>"011101100",
  30883=>"010100100",
  30884=>"000100011",
  30885=>"100110111",
  30886=>"000010001",
  30887=>"100101101",
  30888=>"111100011",
  30889=>"001110000",
  30890=>"011001000",
  30891=>"000000011",
  30892=>"000101101",
  30893=>"101010111",
  30894=>"000010010",
  30895=>"000101011",
  30896=>"100101011",
  30897=>"000011000",
  30898=>"100110100",
  30899=>"000000011",
  30900=>"101101001",
  30901=>"101110011",
  30902=>"011101100",
  30903=>"001100000",
  30904=>"001100100",
  30905=>"001101011",
  30906=>"001000101",
  30907=>"110010010",
  30908=>"010111011",
  30909=>"001101101",
  30910=>"010011001",
  30911=>"001100010",
  30912=>"111011111",
  30913=>"001011101",
  30914=>"001011110",
  30915=>"000111001",
  30916=>"110101111",
  30917=>"101011111",
  30918=>"111111010",
  30919=>"100000111",
  30920=>"011101000",
  30921=>"000011110",
  30922=>"110000110",
  30923=>"000001001",
  30924=>"110010001",
  30925=>"000111110",
  30926=>"010100100",
  30927=>"101100110",
  30928=>"111111000",
  30929=>"000001101",
  30930=>"000011111",
  30931=>"100001101",
  30932=>"001001110",
  30933=>"001011111",
  30934=>"110011010",
  30935=>"100001011",
  30936=>"101011101",
  30937=>"100000101",
  30938=>"111101111",
  30939=>"111010011",
  30940=>"111101011",
  30941=>"001110101",
  30942=>"101110101",
  30943=>"001000110",
  30944=>"101000001",
  30945=>"001100000",
  30946=>"010011100",
  30947=>"001111100",
  30948=>"100101100",
  30949=>"000101000",
  30950=>"101101101",
  30951=>"101000011",
  30952=>"000111010",
  30953=>"001101010",
  30954=>"011011011",
  30955=>"000101100",
  30956=>"110110010",
  30957=>"101000111",
  30958=>"111111010",
  30959=>"100001111",
  30960=>"011111000",
  30961=>"110010000",
  30962=>"101100010",
  30963=>"010011001",
  30964=>"011011001",
  30965=>"101000101",
  30966=>"001000001",
  30967=>"010000111",
  30968=>"100010010",
  30969=>"111011000",
  30970=>"010101001",
  30971=>"101001001",
  30972=>"111000100",
  30973=>"110110011",
  30974=>"110111010",
  30975=>"000101001",
  30976=>"001110000",
  30977=>"011011110",
  30978=>"000101111",
  30979=>"100100000",
  30980=>"101110100",
  30981=>"011101110",
  30982=>"110000000",
  30983=>"111100000",
  30984=>"111001001",
  30985=>"001010000",
  30986=>"110000001",
  30987=>"100100001",
  30988=>"001011110",
  30989=>"000011100",
  30990=>"000101011",
  30991=>"000111010",
  30992=>"110010001",
  30993=>"001000100",
  30994=>"000001010",
  30995=>"000011011",
  30996=>"100010110",
  30997=>"001111111",
  30998=>"011111101",
  30999=>"011001010",
  31000=>"110101001",
  31001=>"001101101",
  31002=>"111001111",
  31003=>"111110101",
  31004=>"110110111",
  31005=>"001001100",
  31006=>"001001011",
  31007=>"100001100",
  31008=>"100000001",
  31009=>"100110001",
  31010=>"010101000",
  31011=>"111011000",
  31012=>"100111111",
  31013=>"101100100",
  31014=>"000010001",
  31015=>"111101001",
  31016=>"010111101",
  31017=>"000000110",
  31018=>"100011010",
  31019=>"001010101",
  31020=>"000000010",
  31021=>"000110111",
  31022=>"110001100",
  31023=>"010010001",
  31024=>"101000010",
  31025=>"111010100",
  31026=>"001100110",
  31027=>"110010011",
  31028=>"001010100",
  31029=>"100000111",
  31030=>"100111100",
  31031=>"001101001",
  31032=>"010010110",
  31033=>"001100100",
  31034=>"110010111",
  31035=>"101101110",
  31036=>"100011000",
  31037=>"100110000",
  31038=>"101010100",
  31039=>"001110101",
  31040=>"001101111",
  31041=>"100000100",
  31042=>"100011111",
  31043=>"001000010",
  31044=>"000000001",
  31045=>"100001001",
  31046=>"100001111",
  31047=>"100011110",
  31048=>"101011111",
  31049=>"000000100",
  31050=>"001001000",
  31051=>"010101001",
  31052=>"000111000",
  31053=>"010001001",
  31054=>"010110100",
  31055=>"011111111",
  31056=>"111110001",
  31057=>"101100010",
  31058=>"001010010",
  31059=>"111101000",
  31060=>"000101100",
  31061=>"101000100",
  31062=>"000101110",
  31063=>"100010010",
  31064=>"000001000",
  31065=>"100000010",
  31066=>"101110100",
  31067=>"001010110",
  31068=>"100110011",
  31069=>"011111111",
  31070=>"101010100",
  31071=>"110010100",
  31072=>"111101111",
  31073=>"001100111",
  31074=>"010100111",
  31075=>"010011111",
  31076=>"011110111",
  31077=>"010100011",
  31078=>"010100111",
  31079=>"010101011",
  31080=>"111110010",
  31081=>"000111101",
  31082=>"011100001",
  31083=>"011000111",
  31084=>"110011010",
  31085=>"001000111",
  31086=>"111000101",
  31087=>"110100010",
  31088=>"111100011",
  31089=>"100010010",
  31090=>"110010101",
  31091=>"000000010",
  31092=>"111100001",
  31093=>"011100001",
  31094=>"000101000",
  31095=>"001100111",
  31096=>"110111010",
  31097=>"110000100",
  31098=>"101110000",
  31099=>"101100110",
  31100=>"100111000",
  31101=>"000100101",
  31102=>"100101111",
  31103=>"010000000",
  31104=>"000010011",
  31105=>"101000101",
  31106=>"011110000",
  31107=>"101111101",
  31108=>"010011101",
  31109=>"011000000",
  31110=>"100011111",
  31111=>"111111110",
  31112=>"111100001",
  31113=>"111100110",
  31114=>"001000111",
  31115=>"001100011",
  31116=>"001000111",
  31117=>"111000000",
  31118=>"100111100",
  31119=>"001010010",
  31120=>"110111010",
  31121=>"000100000",
  31122=>"010011100",
  31123=>"110011100",
  31124=>"100111011",
  31125=>"110100000",
  31126=>"101001111",
  31127=>"001110100",
  31128=>"011011001",
  31129=>"000000011",
  31130=>"101000011",
  31131=>"000011010",
  31132=>"101010101",
  31133=>"000111111",
  31134=>"101001111",
  31135=>"111111010",
  31136=>"100101000",
  31137=>"010010110",
  31138=>"111011101",
  31139=>"000010101",
  31140=>"101011000",
  31141=>"010111011",
  31142=>"000000010",
  31143=>"100001001",
  31144=>"001101111",
  31145=>"011001011",
  31146=>"001101111",
  31147=>"111001000",
  31148=>"101011110",
  31149=>"111100010",
  31150=>"001101111",
  31151=>"101111111",
  31152=>"100101010",
  31153=>"100101100",
  31154=>"100100000",
  31155=>"111001011",
  31156=>"001110111",
  31157=>"100000010",
  31158=>"100100100",
  31159=>"000010000",
  31160=>"101111110",
  31161=>"000111011",
  31162=>"000110001",
  31163=>"111111011",
  31164=>"111111111",
  31165=>"011100001",
  31166=>"000001011",
  31167=>"100110000",
  31168=>"011010011",
  31169=>"111100111",
  31170=>"110001100",
  31171=>"100001101",
  31172=>"000001011",
  31173=>"100011000",
  31174=>"010010010",
  31175=>"010001111",
  31176=>"000011111",
  31177=>"111111100",
  31178=>"110100100",
  31179=>"100010101",
  31180=>"001000110",
  31181=>"011100100",
  31182=>"111010000",
  31183=>"011000000",
  31184=>"100101110",
  31185=>"110010101",
  31186=>"001011000",
  31187=>"001011111",
  31188=>"011111111",
  31189=>"010011101",
  31190=>"101001001",
  31191=>"110100111",
  31192=>"010111111",
  31193=>"011000101",
  31194=>"101101111",
  31195=>"100011111",
  31196=>"101011010",
  31197=>"010011001",
  31198=>"111010010",
  31199=>"001000111",
  31200=>"110100011",
  31201=>"110101101",
  31202=>"110111110",
  31203=>"111111111",
  31204=>"100101100",
  31205=>"111000100",
  31206=>"011001010",
  31207=>"000011000",
  31208=>"010000010",
  31209=>"000110101",
  31210=>"000001110",
  31211=>"000000111",
  31212=>"000110001",
  31213=>"011100000",
  31214=>"011101111",
  31215=>"011110001",
  31216=>"100011001",
  31217=>"010111000",
  31218=>"101100000",
  31219=>"000001000",
  31220=>"011110110",
  31221=>"110001110",
  31222=>"001110100",
  31223=>"101100100",
  31224=>"001101000",
  31225=>"101110000",
  31226=>"100111110",
  31227=>"100001011",
  31228=>"000110111",
  31229=>"101011010",
  31230=>"100100001",
  31231=>"101101110",
  31232=>"100101001",
  31233=>"110000000",
  31234=>"101001001",
  31235=>"111011100",
  31236=>"110011000",
  31237=>"110101110",
  31238=>"000000010",
  31239=>"011000110",
  31240=>"110100000",
  31241=>"110000011",
  31242=>"010010011",
  31243=>"000111000",
  31244=>"000100000",
  31245=>"110101010",
  31246=>"010100100",
  31247=>"101110000",
  31248=>"111001011",
  31249=>"111001001",
  31250=>"100111110",
  31251=>"101010101",
  31252=>"001001101",
  31253=>"011001011",
  31254=>"111011101",
  31255=>"011100010",
  31256=>"011101101",
  31257=>"110011011",
  31258=>"111111010",
  31259=>"101001001",
  31260=>"100001111",
  31261=>"010010101",
  31262=>"000001000",
  31263=>"011011011",
  31264=>"011101000",
  31265=>"010001011",
  31266=>"100001110",
  31267=>"110100100",
  31268=>"111110101",
  31269=>"000001011",
  31270=>"111000011",
  31271=>"000000111",
  31272=>"010101011",
  31273=>"000011010",
  31274=>"000110110",
  31275=>"101110111",
  31276=>"111000101",
  31277=>"011100101",
  31278=>"110001110",
  31279=>"011011100",
  31280=>"110100010",
  31281=>"100100110",
  31282=>"000011001",
  31283=>"111111011",
  31284=>"000111000",
  31285=>"010100110",
  31286=>"100101101",
  31287=>"000110010",
  31288=>"000000001",
  31289=>"001011001",
  31290=>"011000110",
  31291=>"000010101",
  31292=>"011101011",
  31293=>"100010010",
  31294=>"100111101",
  31295=>"110001010",
  31296=>"001111101",
  31297=>"110001110",
  31298=>"011010010",
  31299=>"010100110",
  31300=>"101001101",
  31301=>"011100001",
  31302=>"011101101",
  31303=>"001100010",
  31304=>"001011101",
  31305=>"000110010",
  31306=>"001010100",
  31307=>"000110001",
  31308=>"101001111",
  31309=>"101000101",
  31310=>"001110110",
  31311=>"100010101",
  31312=>"000001101",
  31313=>"000100111",
  31314=>"001001001",
  31315=>"000010010",
  31316=>"011011010",
  31317=>"110011011",
  31318=>"100110111",
  31319=>"001001000",
  31320=>"011101110",
  31321=>"010010001",
  31322=>"000101001",
  31323=>"100011001",
  31324=>"101010000",
  31325=>"110101010",
  31326=>"100011101",
  31327=>"000011110",
  31328=>"001010000",
  31329=>"010100010",
  31330=>"001111110",
  31331=>"010110010",
  31332=>"110011010",
  31333=>"111000111",
  31334=>"011100010",
  31335=>"010011111",
  31336=>"001101001",
  31337=>"100011111",
  31338=>"001101010",
  31339=>"011001100",
  31340=>"010101011",
  31341=>"111101111",
  31342=>"001111011",
  31343=>"000001100",
  31344=>"101000100",
  31345=>"011001111",
  31346=>"101111110",
  31347=>"110101000",
  31348=>"100110110",
  31349=>"001001100",
  31350=>"100011110",
  31351=>"001001110",
  31352=>"101110100",
  31353=>"111111010",
  31354=>"100010101",
  31355=>"010000110",
  31356=>"100100001",
  31357=>"001101101",
  31358=>"010110100",
  31359=>"000011110",
  31360=>"100100000",
  31361=>"010100110",
  31362=>"110010000",
  31363=>"010011001",
  31364=>"110101000",
  31365=>"010001000",
  31366=>"111001010",
  31367=>"111101111",
  31368=>"110111100",
  31369=>"001001100",
  31370=>"111100101",
  31371=>"000010010",
  31372=>"010111100",
  31373=>"000110011",
  31374=>"110010101",
  31375=>"010111111",
  31376=>"001111001",
  31377=>"000011001",
  31378=>"010111001",
  31379=>"110110100",
  31380=>"001010100",
  31381=>"000001001",
  31382=>"101001100",
  31383=>"011000000",
  31384=>"010000101",
  31385=>"101000001",
  31386=>"000101001",
  31387=>"100111001",
  31388=>"011000010",
  31389=>"111111101",
  31390=>"010001000",
  31391=>"100100010",
  31392=>"111101101",
  31393=>"011100111",
  31394=>"010111010",
  31395=>"010111100",
  31396=>"010100000",
  31397=>"101011010",
  31398=>"111001010",
  31399=>"000010100",
  31400=>"110110001",
  31401=>"001100001",
  31402=>"011110010",
  31403=>"111111100",
  31404=>"111111101",
  31405=>"010001110",
  31406=>"111101000",
  31407=>"110001111",
  31408=>"000110010",
  31409=>"101001101",
  31410=>"011110111",
  31411=>"110111110",
  31412=>"110111111",
  31413=>"000111111",
  31414=>"110100111",
  31415=>"011101100",
  31416=>"010001001",
  31417=>"010111101",
  31418=>"101110001",
  31419=>"001101110",
  31420=>"110010101",
  31421=>"001000111",
  31422=>"001000101",
  31423=>"110101000",
  31424=>"001111110",
  31425=>"101010011",
  31426=>"111011010",
  31427=>"101001000",
  31428=>"000011001",
  31429=>"000000000",
  31430=>"100100100",
  31431=>"000110110",
  31432=>"101011100",
  31433=>"100001001",
  31434=>"110010011",
  31435=>"111000001",
  31436=>"101110010",
  31437=>"000000101",
  31438=>"110111111",
  31439=>"001000001",
  31440=>"001011111",
  31441=>"010101100",
  31442=>"010010001",
  31443=>"011000110",
  31444=>"000001000",
  31445=>"000010111",
  31446=>"010100100",
  31447=>"011000101",
  31448=>"010101100",
  31449=>"100101000",
  31450=>"000100110",
  31451=>"101111001",
  31452=>"000100101",
  31453=>"101111000",
  31454=>"010111000",
  31455=>"100100111",
  31456=>"000111101",
  31457=>"101101110",
  31458=>"001110000",
  31459=>"000001110",
  31460=>"000110101",
  31461=>"101101100",
  31462=>"001110110",
  31463=>"001010100",
  31464=>"001111110",
  31465=>"000100111",
  31466=>"100111100",
  31467=>"010001000",
  31468=>"010000011",
  31469=>"011001001",
  31470=>"001001100",
  31471=>"000100110",
  31472=>"011101111",
  31473=>"000000101",
  31474=>"110000011",
  31475=>"010010011",
  31476=>"100100110",
  31477=>"001101101",
  31478=>"111111100",
  31479=>"011100100",
  31480=>"011110011",
  31481=>"100101110",
  31482=>"111010001",
  31483=>"001100100",
  31484=>"000100111",
  31485=>"100000001",
  31486=>"110001110",
  31487=>"000111101",
  31488=>"001100000",
  31489=>"001011011",
  31490=>"111000000",
  31491=>"010001111",
  31492=>"100000000",
  31493=>"110111110",
  31494=>"010010100",
  31495=>"000000000",
  31496=>"101011111",
  31497=>"000100101",
  31498=>"100010011",
  31499=>"001000000",
  31500=>"011101011",
  31501=>"011010011",
  31502=>"111011100",
  31503=>"011101011",
  31504=>"001110000",
  31505=>"101010100",
  31506=>"111010101",
  31507=>"010010111",
  31508=>"101010010",
  31509=>"110110011",
  31510=>"101111011",
  31511=>"110000010",
  31512=>"011011010",
  31513=>"001000110",
  31514=>"110001010",
  31515=>"011000010",
  31516=>"010000000",
  31517=>"100111110",
  31518=>"011100101",
  31519=>"111110100",
  31520=>"001101111",
  31521=>"110010110",
  31522=>"111000101",
  31523=>"111000110",
  31524=>"111011011",
  31525=>"011100010",
  31526=>"101011101",
  31527=>"001010010",
  31528=>"100100100",
  31529=>"010100011",
  31530=>"110010111",
  31531=>"011011110",
  31532=>"100000010",
  31533=>"010001001",
  31534=>"001000110",
  31535=>"111100010",
  31536=>"000111000",
  31537=>"011100011",
  31538=>"101100011",
  31539=>"111101001",
  31540=>"001011001",
  31541=>"000011111",
  31542=>"000010010",
  31543=>"111001000",
  31544=>"110001101",
  31545=>"101101011",
  31546=>"001001111",
  31547=>"010010100",
  31548=>"101100111",
  31549=>"100111101",
  31550=>"010110000",
  31551=>"000011001",
  31552=>"001110111",
  31553=>"010111011",
  31554=>"110111000",
  31555=>"100111101",
  31556=>"110100100",
  31557=>"001001010",
  31558=>"110010111",
  31559=>"001001011",
  31560=>"000010000",
  31561=>"100100100",
  31562=>"111010010",
  31563=>"100111100",
  31564=>"000111011",
  31565=>"011100000",
  31566=>"100101000",
  31567=>"000101001",
  31568=>"011000110",
  31569=>"011110011",
  31570=>"111001100",
  31571=>"001011111",
  31572=>"110000111",
  31573=>"110001111",
  31574=>"111000101",
  31575=>"000110000",
  31576=>"010110011",
  31577=>"110000010",
  31578=>"110110010",
  31579=>"010100001",
  31580=>"000110001",
  31581=>"000000111",
  31582=>"011011110",
  31583=>"000010111",
  31584=>"010001111",
  31585=>"111111110",
  31586=>"000010101",
  31587=>"101111111",
  31588=>"001000000",
  31589=>"110101011",
  31590=>"001011000",
  31591=>"100111011",
  31592=>"110101111",
  31593=>"001111001",
  31594=>"000110100",
  31595=>"001000000",
  31596=>"010000101",
  31597=>"110110111",
  31598=>"101010100",
  31599=>"111111101",
  31600=>"011010010",
  31601=>"011000101",
  31602=>"001111000",
  31603=>"001111110",
  31604=>"010101001",
  31605=>"100000000",
  31606=>"110011111",
  31607=>"000011000",
  31608=>"010011111",
  31609=>"100001000",
  31610=>"011100111",
  31611=>"110110011",
  31612=>"100100100",
  31613=>"011101011",
  31614=>"111111111",
  31615=>"110011111",
  31616=>"100000110",
  31617=>"000011001",
  31618=>"101001110",
  31619=>"000001101",
  31620=>"100000110",
  31621=>"110010101",
  31622=>"101010000",
  31623=>"111000111",
  31624=>"001001101",
  31625=>"000010000",
  31626=>"010001110",
  31627=>"010010000",
  31628=>"100111111",
  31629=>"011000001",
  31630=>"101100010",
  31631=>"011111101",
  31632=>"011101100",
  31633=>"111000001",
  31634=>"000111000",
  31635=>"010100001",
  31636=>"110110100",
  31637=>"000011000",
  31638=>"100010111",
  31639=>"101011100",
  31640=>"111000001",
  31641=>"100001101",
  31642=>"111111001",
  31643=>"111011010",
  31644=>"010011001",
  31645=>"011111000",
  31646=>"000100101",
  31647=>"010010110",
  31648=>"010010011",
  31649=>"101100011",
  31650=>"001010001",
  31651=>"101001101",
  31652=>"100100101",
  31653=>"101000000",
  31654=>"010011110",
  31655=>"001100010",
  31656=>"111111110",
  31657=>"111111000",
  31658=>"000000000",
  31659=>"110011100",
  31660=>"010101001",
  31661=>"111011010",
  31662=>"100001101",
  31663=>"100111100",
  31664=>"111010010",
  31665=>"011110111",
  31666=>"101000011",
  31667=>"011000111",
  31668=>"011111010",
  31669=>"100010000",
  31670=>"001001110",
  31671=>"011001011",
  31672=>"110111011",
  31673=>"111000100",
  31674=>"000011000",
  31675=>"101110111",
  31676=>"111000011",
  31677=>"001110011",
  31678=>"011011111",
  31679=>"100101100",
  31680=>"000011110",
  31681=>"000110111",
  31682=>"100000000",
  31683=>"011011110",
  31684=>"111000001",
  31685=>"010000111",
  31686=>"101010110",
  31687=>"110000110",
  31688=>"000001010",
  31689=>"100000001",
  31690=>"101100101",
  31691=>"100000011",
  31692=>"011110101",
  31693=>"000010000",
  31694=>"111001100",
  31695=>"011011000",
  31696=>"001110010",
  31697=>"101110001",
  31698=>"000101001",
  31699=>"101010110",
  31700=>"010010100",
  31701=>"010001101",
  31702=>"010111111",
  31703=>"010110111",
  31704=>"010000101",
  31705=>"000010111",
  31706=>"001101100",
  31707=>"110110000",
  31708=>"010101110",
  31709=>"100110111",
  31710=>"010101001",
  31711=>"001111100",
  31712=>"110011000",
  31713=>"110101110",
  31714=>"110100011",
  31715=>"011000000",
  31716=>"010100110",
  31717=>"100110101",
  31718=>"100110001",
  31719=>"110101011",
  31720=>"000100110",
  31721=>"000001001",
  31722=>"010110100",
  31723=>"110000110",
  31724=>"010011101",
  31725=>"000010110",
  31726=>"111100011",
  31727=>"000100101",
  31728=>"101010101",
  31729=>"111001001",
  31730=>"101001111",
  31731=>"110101010",
  31732=>"001001101",
  31733=>"001001101",
  31734=>"011000111",
  31735=>"000101001",
  31736=>"100001101",
  31737=>"100101010",
  31738=>"100000111",
  31739=>"001011001",
  31740=>"100111111",
  31741=>"011111000",
  31742=>"010100000",
  31743=>"010010000",
  31744=>"111101000",
  31745=>"000000101",
  31746=>"110010011",
  31747=>"001111010",
  31748=>"110010101",
  31749=>"111100110",
  31750=>"111101111",
  31751=>"000000100",
  31752=>"011110101",
  31753=>"101101110",
  31754=>"001000110",
  31755=>"111011111",
  31756=>"111011010",
  31757=>"001011010",
  31758=>"000101110",
  31759=>"001101010",
  31760=>"001000101",
  31761=>"101111100",
  31762=>"011100010",
  31763=>"111000110",
  31764=>"010100000",
  31765=>"011000110",
  31766=>"101001000",
  31767=>"001000101",
  31768=>"011011111",
  31769=>"111010110",
  31770=>"110100011",
  31771=>"100001110",
  31772=>"100101000",
  31773=>"001111100",
  31774=>"011100010",
  31775=>"010000111",
  31776=>"011001010",
  31777=>"111111111",
  31778=>"111010001",
  31779=>"100110001",
  31780=>"110110001",
  31781=>"101110000",
  31782=>"101110111",
  31783=>"100001110",
  31784=>"111111011",
  31785=>"101011101",
  31786=>"001110100",
  31787=>"111111001",
  31788=>"000011010",
  31789=>"111101111",
  31790=>"111111111",
  31791=>"011000001",
  31792=>"101101111",
  31793=>"001101011",
  31794=>"111101001",
  31795=>"000000000",
  31796=>"110101111",
  31797=>"001010001",
  31798=>"111110101",
  31799=>"001001011",
  31800=>"101011010",
  31801=>"001110110",
  31802=>"100101001",
  31803=>"000110001",
  31804=>"101011001",
  31805=>"110010101",
  31806=>"011001110",
  31807=>"111100011",
  31808=>"001011011",
  31809=>"100111010",
  31810=>"010100111",
  31811=>"100100110",
  31812=>"001000010",
  31813=>"000001001",
  31814=>"101101110",
  31815=>"001010010",
  31816=>"001101100",
  31817=>"011101111",
  31818=>"000101000",
  31819=>"110010001",
  31820=>"000101000",
  31821=>"110100010",
  31822=>"100011110",
  31823=>"001101110",
  31824=>"100001010",
  31825=>"101010000",
  31826=>"111011110",
  31827=>"111110010",
  31828=>"000010110",
  31829=>"000110110",
  31830=>"011000010",
  31831=>"110110011",
  31832=>"111111010",
  31833=>"010000000",
  31834=>"110011000",
  31835=>"110000111",
  31836=>"111000011",
  31837=>"010010001",
  31838=>"100111110",
  31839=>"111101110",
  31840=>"010100000",
  31841=>"011101110",
  31842=>"100100110",
  31843=>"000110011",
  31844=>"001110011",
  31845=>"010001101",
  31846=>"101000011",
  31847=>"111101111",
  31848=>"100100011",
  31849=>"001000100",
  31850=>"010110011",
  31851=>"011111010",
  31852=>"001101101",
  31853=>"110011010",
  31854=>"111101001",
  31855=>"011111101",
  31856=>"100101111",
  31857=>"000110100",
  31858=>"010111000",
  31859=>"100111111",
  31860=>"010100000",
  31861=>"111100010",
  31862=>"100100010",
  31863=>"100101100",
  31864=>"111100010",
  31865=>"110111001",
  31866=>"111111000",
  31867=>"001111010",
  31868=>"101111011",
  31869=>"101101001",
  31870=>"101101010",
  31871=>"010000010",
  31872=>"101110111",
  31873=>"100101111",
  31874=>"100101011",
  31875=>"111111101",
  31876=>"001100010",
  31877=>"101011110",
  31878=>"111111110",
  31879=>"000000111",
  31880=>"011010001",
  31881=>"011010001",
  31882=>"110101010",
  31883=>"101001011",
  31884=>"010010101",
  31885=>"000000101",
  31886=>"000010001",
  31887=>"000101001",
  31888=>"101110110",
  31889=>"000110100",
  31890=>"000011000",
  31891=>"000101010",
  31892=>"110011000",
  31893=>"100111010",
  31894=>"110101100",
  31895=>"111000001",
  31896=>"110010111",
  31897=>"010000111",
  31898=>"101110001",
  31899=>"111000110",
  31900=>"101110011",
  31901=>"010011111",
  31902=>"001010101",
  31903=>"000001110",
  31904=>"000100001",
  31905=>"101111011",
  31906=>"110011100",
  31907=>"010010111",
  31908=>"100000001",
  31909=>"111011010",
  31910=>"010000011",
  31911=>"101001011",
  31912=>"110000001",
  31913=>"101101111",
  31914=>"110101001",
  31915=>"010110000",
  31916=>"011000101",
  31917=>"000001111",
  31918=>"110011111",
  31919=>"110011000",
  31920=>"000010111",
  31921=>"110101100",
  31922=>"110011001",
  31923=>"101001001",
  31924=>"100000110",
  31925=>"110000000",
  31926=>"010010111",
  31927=>"110010110",
  31928=>"010000010",
  31929=>"111110011",
  31930=>"010000101",
  31931=>"001101000",
  31932=>"010101000",
  31933=>"100111110",
  31934=>"011011011",
  31935=>"110101010",
  31936=>"101101010",
  31937=>"110001101",
  31938=>"100100001",
  31939=>"101011110",
  31940=>"111111111",
  31941=>"111110110",
  31942=>"010101010",
  31943=>"001010010",
  31944=>"100101001",
  31945=>"100000001",
  31946=>"011000010",
  31947=>"111110100",
  31948=>"111011010",
  31949=>"111101111",
  31950=>"111101100",
  31951=>"100010100",
  31952=>"111010001",
  31953=>"000010111",
  31954=>"111001101",
  31955=>"001111101",
  31956=>"100010000",
  31957=>"010100101",
  31958=>"111000011",
  31959=>"001010111",
  31960=>"000001000",
  31961=>"100110011",
  31962=>"000001010",
  31963=>"110010001",
  31964=>"010010101",
  31965=>"111001110",
  31966=>"111111110",
  31967=>"000111111",
  31968=>"011111100",
  31969=>"000011000",
  31970=>"110110011",
  31971=>"111010010",
  31972=>"000011010",
  31973=>"101110011",
  31974=>"110111010",
  31975=>"111010101",
  31976=>"100001100",
  31977=>"100110100",
  31978=>"100000100",
  31979=>"010110011",
  31980=>"111011100",
  31981=>"100011111",
  31982=>"010010011",
  31983=>"101001100",
  31984=>"111110000",
  31985=>"111010000",
  31986=>"101110110",
  31987=>"001011110",
  31988=>"010010000",
  31989=>"010110011",
  31990=>"100001110",
  31991=>"101011110",
  31992=>"001101110",
  31993=>"100100111",
  31994=>"100011000",
  31995=>"110111101",
  31996=>"011110101",
  31997=>"000111010",
  31998=>"011111110",
  31999=>"001011000",
  32000=>"011111111",
  32001=>"000111001",
  32002=>"101000111",
  32003=>"101111011",
  32004=>"011101010",
  32005=>"111111011",
  32006=>"001111100",
  32007=>"101100000",
  32008=>"100111011",
  32009=>"011101101",
  32010=>"100111001",
  32011=>"001101111",
  32012=>"001000111",
  32013=>"111011111",
  32014=>"111110011",
  32015=>"001001111",
  32016=>"000001001",
  32017=>"110011101",
  32018=>"010001100",
  32019=>"111110000",
  32020=>"111101101",
  32021=>"101101111",
  32022=>"010001001",
  32023=>"100001111",
  32024=>"110111100",
  32025=>"100111000",
  32026=>"010010111",
  32027=>"011000100",
  32028=>"010101111",
  32029=>"101101111",
  32030=>"100111100",
  32031=>"110100111",
  32032=>"011000010",
  32033=>"111011000",
  32034=>"111100111",
  32035=>"010100000",
  32036=>"001101010",
  32037=>"000110000",
  32038=>"100001111",
  32039=>"100010101",
  32040=>"000100100",
  32041=>"011101110",
  32042=>"101100100",
  32043=>"000110001",
  32044=>"000001110",
  32045=>"010000010",
  32046=>"110110010",
  32047=>"010101010",
  32048=>"010101111",
  32049=>"011000001",
  32050=>"000011011",
  32051=>"111101110",
  32052=>"111110001",
  32053=>"100011100",
  32054=>"110100000",
  32055=>"001010010",
  32056=>"010000011",
  32057=>"101000011",
  32058=>"110110000",
  32059=>"101010110",
  32060=>"101110001",
  32061=>"010000010",
  32062=>"000101100",
  32063=>"000010101",
  32064=>"010101010",
  32065=>"111001100",
  32066=>"000010010",
  32067=>"111101100",
  32068=>"110100111",
  32069=>"101100111",
  32070=>"001011100",
  32071=>"000011000",
  32072=>"000000101",
  32073=>"111110001",
  32074=>"010000110",
  32075=>"111001100",
  32076=>"110010110",
  32077=>"000000011",
  32078=>"110000110",
  32079=>"111111000",
  32080=>"101101111",
  32081=>"010111011",
  32082=>"000101001",
  32083=>"101010100",
  32084=>"111110101",
  32085=>"111010100",
  32086=>"110011011",
  32087=>"110110110",
  32088=>"001100111",
  32089=>"100000110",
  32090=>"001110110",
  32091=>"111111011",
  32092=>"000011101",
  32093=>"001011111",
  32094=>"001010001",
  32095=>"100010010",
  32096=>"110011011",
  32097=>"110011010",
  32098=>"001110001",
  32099=>"101101111",
  32100=>"010111100",
  32101=>"000110010",
  32102=>"010000001",
  32103=>"100001010",
  32104=>"111011000",
  32105=>"111101101",
  32106=>"011110000",
  32107=>"100101001",
  32108=>"010100000",
  32109=>"111101000",
  32110=>"000011010",
  32111=>"001000011",
  32112=>"001001010",
  32113=>"100011111",
  32114=>"100100011",
  32115=>"101011011",
  32116=>"111111000",
  32117=>"000110001",
  32118=>"100000000",
  32119=>"101101001",
  32120=>"000000101",
  32121=>"000001011",
  32122=>"110111010",
  32123=>"010110000",
  32124=>"011101101",
  32125=>"010010111",
  32126=>"100100000",
  32127=>"000011001",
  32128=>"000000111",
  32129=>"101001100",
  32130=>"000011010",
  32131=>"001011011",
  32132=>"100001111",
  32133=>"111110011",
  32134=>"011001001",
  32135=>"010101011",
  32136=>"101000011",
  32137=>"101000110",
  32138=>"101000101",
  32139=>"000010000",
  32140=>"010101000",
  32141=>"101110001",
  32142=>"111111111",
  32143=>"100001101",
  32144=>"010010011",
  32145=>"100001111",
  32146=>"100100100",
  32147=>"101100110",
  32148=>"111111110",
  32149=>"110000001",
  32150=>"110010000",
  32151=>"010010011",
  32152=>"010010101",
  32153=>"111101010",
  32154=>"011011101",
  32155=>"000010110",
  32156=>"110011011",
  32157=>"110011000",
  32158=>"111010111",
  32159=>"001010000",
  32160=>"100100010",
  32161=>"000100101",
  32162=>"101101010",
  32163=>"111110011",
  32164=>"010010011",
  32165=>"100100011",
  32166=>"100010110",
  32167=>"011011011",
  32168=>"100001000",
  32169=>"100000110",
  32170=>"110001100",
  32171=>"000010100",
  32172=>"110011100",
  32173=>"000100100",
  32174=>"000111001",
  32175=>"101111010",
  32176=>"001111001",
  32177=>"001110101",
  32178=>"000000100",
  32179=>"111111000",
  32180=>"001011000",
  32181=>"010101011",
  32182=>"101010010",
  32183=>"100111011",
  32184=>"001001110",
  32185=>"011111101",
  32186=>"011011100",
  32187=>"101000010",
  32188=>"101000100",
  32189=>"111110000",
  32190=>"110001010",
  32191=>"111111000",
  32192=>"110011101",
  32193=>"010110110",
  32194=>"110100100",
  32195=>"010010111",
  32196=>"010001110",
  32197=>"000001110",
  32198=>"111100000",
  32199=>"000111001",
  32200=>"110001001",
  32201=>"011010000",
  32202=>"010110110",
  32203=>"010001111",
  32204=>"011101100",
  32205=>"001110100",
  32206=>"000001010",
  32207=>"001101101",
  32208=>"010001010",
  32209=>"011110101",
  32210=>"110100011",
  32211=>"111010101",
  32212=>"001101101",
  32213=>"101010000",
  32214=>"000101110",
  32215=>"011011111",
  32216=>"011110011",
  32217=>"111101001",
  32218=>"111010100",
  32219=>"110100111",
  32220=>"111000001",
  32221=>"110101011",
  32222=>"011011111",
  32223=>"000010101",
  32224=>"000001001",
  32225=>"110100001",
  32226=>"000111010",
  32227=>"000011011",
  32228=>"010111001",
  32229=>"010011100",
  32230=>"111000000",
  32231=>"111111110",
  32232=>"111100001",
  32233=>"100111100",
  32234=>"000000010",
  32235=>"011101011",
  32236=>"000010110",
  32237=>"110101011",
  32238=>"101110101",
  32239=>"001001000",
  32240=>"010101101",
  32241=>"011101110",
  32242=>"111010100",
  32243=>"110111001",
  32244=>"110111000",
  32245=>"010001001",
  32246=>"111111110",
  32247=>"111111101",
  32248=>"111011000",
  32249=>"101010010",
  32250=>"111000111",
  32251=>"010101111",
  32252=>"111010101",
  32253=>"001000101",
  32254=>"011000010",
  32255=>"011101111",
  32256=>"001001100",
  32257=>"000000000",
  32258=>"111001010",
  32259=>"101000011",
  32260=>"111111110",
  32261=>"111101101",
  32262=>"000101001",
  32263=>"111010000",
  32264=>"000101001",
  32265=>"110000000",
  32266=>"000000000",
  32267=>"010001011",
  32268=>"111101100",
  32269=>"011110010",
  32270=>"011001101",
  32271=>"111111111",
  32272=>"000100011",
  32273=>"010100011",
  32274=>"100001111",
  32275=>"000000101",
  32276=>"110000010",
  32277=>"111010001",
  32278=>"000000011",
  32279=>"100001111",
  32280=>"111001011",
  32281=>"100000111",
  32282=>"110111111",
  32283=>"000001110",
  32284=>"111000111",
  32285=>"100010001",
  32286=>"111001110",
  32287=>"011011100",
  32288=>"111100101",
  32289=>"000000000",
  32290=>"010000010",
  32291=>"101110110",
  32292=>"100111111",
  32293=>"001111110",
  32294=>"011000100",
  32295=>"000011011",
  32296=>"100000001",
  32297=>"001010101",
  32298=>"000000100",
  32299=>"111000011",
  32300=>"111110001",
  32301=>"111101100",
  32302=>"001011110",
  32303=>"001100110",
  32304=>"000010000",
  32305=>"111001000",
  32306=>"001101010",
  32307=>"101011101",
  32308=>"101101001",
  32309=>"110011101",
  32310=>"110101101",
  32311=>"100001001",
  32312=>"100100110",
  32313=>"010000000",
  32314=>"011101010",
  32315=>"110100100",
  32316=>"100100000",
  32317=>"110100100",
  32318=>"100100011",
  32319=>"011111010",
  32320=>"111101001",
  32321=>"011111011",
  32322=>"011100101",
  32323=>"110111111",
  32324=>"111001010",
  32325=>"010010110",
  32326=>"100001101",
  32327=>"000011001",
  32328=>"101000100",
  32329=>"101000001",
  32330=>"111000100",
  32331=>"000001010",
  32332=>"111101111",
  32333=>"110110001",
  32334=>"011000010",
  32335=>"010110001",
  32336=>"100000110",
  32337=>"010100111",
  32338=>"011111110",
  32339=>"101000110",
  32340=>"011011110",
  32341=>"111110101",
  32342=>"101101100",
  32343=>"100001011",
  32344=>"101001001",
  32345=>"011000100",
  32346=>"111101100",
  32347=>"000010111",
  32348=>"111010110",
  32349=>"111110111",
  32350=>"001100111",
  32351=>"000111011",
  32352=>"010100000",
  32353=>"010100110",
  32354=>"011111010",
  32355=>"111100011",
  32356=>"000001101",
  32357=>"011010110",
  32358=>"111011101",
  32359=>"101001000",
  32360=>"100100010",
  32361=>"010101110",
  32362=>"010011110",
  32363=>"010011100",
  32364=>"000101110",
  32365=>"011100000",
  32366=>"011001110",
  32367=>"111100010",
  32368=>"100111101",
  32369=>"110110101",
  32370=>"110110000",
  32371=>"001101101",
  32372=>"011001101",
  32373=>"111001110",
  32374=>"111110100",
  32375=>"111000001",
  32376=>"101110000",
  32377=>"010111110",
  32378=>"100000000",
  32379=>"111001101",
  32380=>"111101011",
  32381=>"100111001",
  32382=>"110111010",
  32383=>"010110110",
  32384=>"010111011",
  32385=>"111111001",
  32386=>"111000110",
  32387=>"101111010",
  32388=>"101101000",
  32389=>"101101001",
  32390=>"011101001",
  32391=>"001000010",
  32392=>"101001111",
  32393=>"011000110",
  32394=>"000100101",
  32395=>"101000100",
  32396=>"000110111",
  32397=>"010010110",
  32398=>"001000000",
  32399=>"010111110",
  32400=>"110011111",
  32401=>"011101000",
  32402=>"110001011",
  32403=>"111101110",
  32404=>"110001110",
  32405=>"101110010",
  32406=>"000011110",
  32407=>"011100101",
  32408=>"101101111",
  32409=>"101001111",
  32410=>"010001000",
  32411=>"001011111",
  32412=>"101100010",
  32413=>"001011010",
  32414=>"010100000",
  32415=>"000011110",
  32416=>"011100000",
  32417=>"110100000",
  32418=>"101101011",
  32419=>"100100100",
  32420=>"111101110",
  32421=>"000011011",
  32422=>"000100001",
  32423=>"010010101",
  32424=>"101111100",
  32425=>"001000000",
  32426=>"011001000",
  32427=>"101010011",
  32428=>"001111000",
  32429=>"110011111",
  32430=>"110110010",
  32431=>"011110001",
  32432=>"000001100",
  32433=>"001010011",
  32434=>"000000000",
  32435=>"011010100",
  32436=>"110011101",
  32437=>"101111111",
  32438=>"111001101",
  32439=>"111110110",
  32440=>"010000110",
  32441=>"100000000",
  32442=>"111010110",
  32443=>"100101101",
  32444=>"001000101",
  32445=>"111001101",
  32446=>"010100101",
  32447=>"011011101",
  32448=>"010001011",
  32449=>"101010101",
  32450=>"111001001",
  32451=>"001100010",
  32452=>"101010000",
  32453=>"010000000",
  32454=>"111101000",
  32455=>"101110000",
  32456=>"101110110",
  32457=>"001101101",
  32458=>"111101011",
  32459=>"101111100",
  32460=>"000111001",
  32461=>"010000010",
  32462=>"000111000",
  32463=>"001110001",
  32464=>"110010001",
  32465=>"101101011",
  32466=>"001001100",
  32467=>"001011010",
  32468=>"100010001",
  32469=>"011101001",
  32470=>"001101101",
  32471=>"011011101",
  32472=>"000001101",
  32473=>"110010110",
  32474=>"100100111",
  32475=>"000010100",
  32476=>"110101011",
  32477=>"010010010",
  32478=>"000011011",
  32479=>"111101011",
  32480=>"110110100",
  32481=>"101000111",
  32482=>"011010001",
  32483=>"110000110",
  32484=>"000101110",
  32485=>"001010000",
  32486=>"000001000",
  32487=>"000101010",
  32488=>"001001101",
  32489=>"111011111",
  32490=>"100000101",
  32491=>"111111011",
  32492=>"010101011",
  32493=>"000101010",
  32494=>"000111110",
  32495=>"100101111",
  32496=>"101000111",
  32497=>"110101101",
  32498=>"110100011",
  32499=>"111110000",
  32500=>"001110001",
  32501=>"100011110",
  32502=>"011110000",
  32503=>"110000111",
  32504=>"010010000",
  32505=>"000000000",
  32506=>"010110100",
  32507=>"001001011",
  32508=>"111111000",
  32509=>"111101010",
  32510=>"000110111",
  32511=>"000111111",
  32512=>"100011110",
  32513=>"111100111",
  32514=>"011101101",
  32515=>"111100000",
  32516=>"001000110",
  32517=>"110110111",
  32518=>"011110001",
  32519=>"000000001",
  32520=>"101000110",
  32521=>"001100001",
  32522=>"111000010",
  32523=>"010001101",
  32524=>"101101000",
  32525=>"100101101",
  32526=>"010100001",
  32527=>"111111010",
  32528=>"101100110",
  32529=>"101010011",
  32530=>"010010001",
  32531=>"011010110",
  32532=>"110001100",
  32533=>"011001000",
  32534=>"001000010",
  32535=>"010111010",
  32536=>"100100100",
  32537=>"111000011",
  32538=>"101111000",
  32539=>"011001111",
  32540=>"110011000",
  32541=>"001011110",
  32542=>"011010011",
  32543=>"111000010",
  32544=>"000011111",
  32545=>"111101000",
  32546=>"001000010",
  32547=>"110000101",
  32548=>"111001111",
  32549=>"101010000",
  32550=>"110000000",
  32551=>"110101101",
  32552=>"111100100",
  32553=>"000011110",
  32554=>"111110100",
  32555=>"011000000",
  32556=>"011110111",
  32557=>"101100111",
  32558=>"100010101",
  32559=>"011011011",
  32560=>"010000100",
  32561=>"001111011",
  32562=>"110011001",
  32563=>"100001000",
  32564=>"000100000",
  32565=>"000010001",
  32566=>"000110011",
  32567=>"000011010",
  32568=>"110000000",
  32569=>"010011011",
  32570=>"110011000",
  32571=>"001000001",
  32572=>"101111110",
  32573=>"101100000",
  32574=>"101001111",
  32575=>"101010001",
  32576=>"001110000",
  32577=>"011011010",
  32578=>"011001111",
  32579=>"011001110",
  32580=>"000010101",
  32581=>"001101100",
  32582=>"111010010",
  32583=>"000111111",
  32584=>"111100111",
  32585=>"011100011",
  32586=>"011010001",
  32587=>"100100110",
  32588=>"010111100",
  32589=>"001110110",
  32590=>"001000100",
  32591=>"010011010",
  32592=>"101101001",
  32593=>"110001011",
  32594=>"011011101",
  32595=>"100010111",
  32596=>"101001110",
  32597=>"011011101",
  32598=>"111011111",
  32599=>"011111110",
  32600=>"001000010",
  32601=>"011011110",
  32602=>"001001000",
  32603=>"110001110",
  32604=>"001100001",
  32605=>"001010001",
  32606=>"100100100",
  32607=>"110110010",
  32608=>"101101111",
  32609=>"111110011",
  32610=>"101010001",
  32611=>"111010111",
  32612=>"100010011",
  32613=>"100011100",
  32614=>"111100110",
  32615=>"101011101",
  32616=>"111100100",
  32617=>"100101010",
  32618=>"100100100",
  32619=>"101101010",
  32620=>"011101111",
  32621=>"101000000",
  32622=>"111000110",
  32623=>"100101111",
  32624=>"011000110",
  32625=>"011000011",
  32626=>"000110101",
  32627=>"001010101",
  32628=>"111000011",
  32629=>"010001111",
  32630=>"101100001",
  32631=>"101111101",
  32632=>"110100000",
  32633=>"111011000",
  32634=>"111111111",
  32635=>"100111111",
  32636=>"010111001",
  32637=>"010101101",
  32638=>"010000011",
  32639=>"110111001",
  32640=>"111010001",
  32641=>"110101000",
  32642=>"101101111",
  32643=>"111010010",
  32644=>"111111111",
  32645=>"110111000",
  32646=>"000110100",
  32647=>"000111001",
  32648=>"010000001",
  32649=>"010000100",
  32650=>"110010010",
  32651=>"010100000",
  32652=>"000001011",
  32653=>"101101001",
  32654=>"010110000",
  32655=>"011011111",
  32656=>"000011010",
  32657=>"111000010",
  32658=>"101100001",
  32659=>"011100111",
  32660=>"011100011",
  32661=>"101111111",
  32662=>"111101011",
  32663=>"100001000",
  32664=>"010001100",
  32665=>"010000010",
  32666=>"101010011",
  32667=>"001010011",
  32668=>"001010111",
  32669=>"111101110",
  32670=>"100110001",
  32671=>"110111000",
  32672=>"110000101",
  32673=>"010011001",
  32674=>"111010001",
  32675=>"100001100",
  32676=>"100000110",
  32677=>"111101001",
  32678=>"001010110",
  32679=>"111111011",
  32680=>"110110100",
  32681=>"000100111",
  32682=>"101110011",
  32683=>"011110011",
  32684=>"000011111",
  32685=>"000111010",
  32686=>"111011011",
  32687=>"100100110",
  32688=>"111110110",
  32689=>"010000000",
  32690=>"011101110",
  32691=>"111100100",
  32692=>"101001101",
  32693=>"110101110",
  32694=>"111001111",
  32695=>"000100001",
  32696=>"111110110",
  32697=>"000001001",
  32698=>"101110101",
  32699=>"011101011",
  32700=>"101101111",
  32701=>"111110101",
  32702=>"011000001",
  32703=>"000111011",
  32704=>"100110111",
  32705=>"001011001",
  32706=>"101110111",
  32707=>"010100010",
  32708=>"000111000",
  32709=>"100011001",
  32710=>"100101101",
  32711=>"001110111",
  32712=>"011110000",
  32713=>"111101101",
  32714=>"000001010",
  32715=>"011011111",
  32716=>"111010000",
  32717=>"011100100",
  32718=>"010111111",
  32719=>"110011010",
  32720=>"100001001",
  32721=>"000011001",
  32722=>"001000000",
  32723=>"101000001",
  32724=>"101111111",
  32725=>"100011010",
  32726=>"101100101",
  32727=>"100001000",
  32728=>"000111100",
  32729=>"000100110",
  32730=>"100101010",
  32731=>"100011100",
  32732=>"010010000",
  32733=>"101000110",
  32734=>"011010111",
  32735=>"101001111",
  32736=>"111101101",
  32737=>"100000010",
  32738=>"011001001",
  32739=>"100111111",
  32740=>"100101010",
  32741=>"010101000",
  32742=>"101101111",
  32743=>"110000011",
  32744=>"110000010",
  32745=>"100001111",
  32746=>"011111111",
  32747=>"001111011",
  32748=>"101101001",
  32749=>"011010111",
  32750=>"001011111",
  32751=>"001000100",
  32752=>"110010010",
  32753=>"001010011",
  32754=>"100110001",
  32755=>"110101011",
  32756=>"010001111",
  32757=>"010111011",
  32758=>"101111110",
  32759=>"111001100",
  32760=>"001111100",
  32761=>"111101001",
  32762=>"011010111",
  32763=>"001100011",
  32764=>"111101111",
  32765=>"001001101",
  32766=>"000001100",
  32767=>"110001000",
  32768=>"101110000",
  32769=>"010111010",
  32770=>"011000011",
  32771=>"001000111",
  32772=>"001001100",
  32773=>"110010101",
  32774=>"111111111",
  32775=>"011011000",
  32776=>"100010010",
  32777=>"010101100",
  32778=>"100101011",
  32779=>"111001100",
  32780=>"110011111",
  32781=>"111100010",
  32782=>"111010001",
  32783=>"110011111",
  32784=>"101010110",
  32785=>"111011101",
  32786=>"001010000",
  32787=>"001010101",
  32788=>"001100001",
  32789=>"100010100",
  32790=>"111101101",
  32791=>"111100001",
  32792=>"010000110",
  32793=>"100110000",
  32794=>"111110000",
  32795=>"101010001",
  32796=>"111100010",
  32797=>"101001110",
  32798=>"110011111",
  32799=>"011000001",
  32800=>"111001101",
  32801=>"111111010",
  32802=>"011111000",
  32803=>"001100001",
  32804=>"000011001",
  32805=>"110110111",
  32806=>"101100101",
  32807=>"111101110",
  32808=>"111001101",
  32809=>"100111010",
  32810=>"001000101",
  32811=>"110110001",
  32812=>"111110111",
  32813=>"011001100",
  32814=>"000010100",
  32815=>"100000010",
  32816=>"111100000",
  32817=>"001111101",
  32818=>"010011111",
  32819=>"101100010",
  32820=>"011010100",
  32821=>"100111110",
  32822=>"010001101",
  32823=>"111110110",
  32824=>"100001010",
  32825=>"000010101",
  32826=>"101001100",
  32827=>"010011110",
  32828=>"000000110",
  32829=>"011100111",
  32830=>"001001011",
  32831=>"101011010",
  32832=>"111111010",
  32833=>"011000010",
  32834=>"110110010",
  32835=>"100111001",
  32836=>"011000000",
  32837=>"100000010",
  32838=>"010010110",
  32839=>"100000010",
  32840=>"001011010",
  32841=>"101100010",
  32842=>"010011101",
  32843=>"111101001",
  32844=>"010011111",
  32845=>"011001110",
  32846=>"111110001",
  32847=>"111011100",
  32848=>"000001010",
  32849=>"111110010",
  32850=>"110010100",
  32851=>"100110011",
  32852=>"000001101",
  32853=>"010000101",
  32854=>"011011100",
  32855=>"000011111",
  32856=>"011010101",
  32857=>"010010101",
  32858=>"100001111",
  32859=>"111000100",
  32860=>"010100010",
  32861=>"000101011",
  32862=>"010110011",
  32863=>"111101011",
  32864=>"001000110",
  32865=>"001001001",
  32866=>"111100101",
  32867=>"000011101",
  32868=>"111001000",
  32869=>"110111010",
  32870=>"000101000",
  32871=>"111110010",
  32872=>"001000100",
  32873=>"101011000",
  32874=>"000100010",
  32875=>"001010100",
  32876=>"101101100",
  32877=>"101110101",
  32878=>"001010010",
  32879=>"111011111",
  32880=>"000110111",
  32881=>"000101111",
  32882=>"111110011",
  32883=>"000111101",
  32884=>"110111011",
  32885=>"001100100",
  32886=>"101101000",
  32887=>"100010011",
  32888=>"101101000",
  32889=>"110110001",
  32890=>"011000001",
  32891=>"001001010",
  32892=>"101110110",
  32893=>"011100111",
  32894=>"111100000",
  32895=>"010011000",
  32896=>"101011111",
  32897=>"001101101",
  32898=>"000100001",
  32899=>"100111010",
  32900=>"111100111",
  32901=>"000011010",
  32902=>"001011001",
  32903=>"111010100",
  32904=>"010000100",
  32905=>"110110001",
  32906=>"110001110",
  32907=>"110010001",
  32908=>"001110101",
  32909=>"000110110",
  32910=>"100101001",
  32911=>"101011100",
  32912=>"101101101",
  32913=>"000110110",
  32914=>"111011110",
  32915=>"110100100",
  32916=>"000011010",
  32917=>"011111110",
  32918=>"100101100",
  32919=>"010111010",
  32920=>"100001110",
  32921=>"111000011",
  32922=>"010000011",
  32923=>"010011110",
  32924=>"010000010",
  32925=>"000100010",
  32926=>"110011001",
  32927=>"000010101",
  32928=>"100011110",
  32929=>"100010000",
  32930=>"000111001",
  32931=>"111001111",
  32932=>"101111101",
  32933=>"111100100",
  32934=>"100010110",
  32935=>"000010000",
  32936=>"100010001",
  32937=>"111010111",
  32938=>"101010110",
  32939=>"101100000",
  32940=>"101000010",
  32941=>"111000011",
  32942=>"101100100",
  32943=>"101010100",
  32944=>"001010000",
  32945=>"001101101",
  32946=>"101101111",
  32947=>"110111000",
  32948=>"101001000",
  32949=>"001111111",
  32950=>"000011011",
  32951=>"011001110",
  32952=>"001001110",
  32953=>"110111101",
  32954=>"010110101",
  32955=>"000101011",
  32956=>"100001111",
  32957=>"000011010",
  32958=>"110000110",
  32959=>"011110001",
  32960=>"100100110",
  32961=>"100111101",
  32962=>"101101110",
  32963=>"010110100",
  32964=>"001010110",
  32965=>"010000100",
  32966=>"000100011",
  32967=>"111111111",
  32968=>"111111100",
  32969=>"111001110",
  32970=>"000001110",
  32971=>"000111101",
  32972=>"001111111",
  32973=>"100110000",
  32974=>"100011110",
  32975=>"011000010",
  32976=>"011100100",
  32977=>"111101111",
  32978=>"001100011",
  32979=>"110110011",
  32980=>"001010011",
  32981=>"100111111",
  32982=>"010100111",
  32983=>"000111000",
  32984=>"101000010",
  32985=>"000101000",
  32986=>"001000011",
  32987=>"000011011",
  32988=>"111010011",
  32989=>"011001001",
  32990=>"010001011",
  32991=>"100111010",
  32992=>"001101111",
  32993=>"110101101",
  32994=>"000110000",
  32995=>"010010011",
  32996=>"100110100",
  32997=>"000111111",
  32998=>"011010010",
  32999=>"011110000",
  33000=>"000010101",
  33001=>"100001101",
  33002=>"111111110",
  33003=>"111000110",
  33004=>"100111011",
  33005=>"010100010",
  33006=>"101000011",
  33007=>"000001101",
  33008=>"111000001",
  33009=>"100101100",
  33010=>"110011100",
  33011=>"000111000",
  33012=>"000101011",
  33013=>"010111101",
  33014=>"110110110",
  33015=>"000001101",
  33016=>"111010100",
  33017=>"000010001",
  33018=>"100110010",
  33019=>"000011100",
  33020=>"011001100",
  33021=>"001100011",
  33022=>"000011111",
  33023=>"001100001",
  33024=>"111011010",
  33025=>"001110111",
  33026=>"010001010",
  33027=>"010010110",
  33028=>"101100101",
  33029=>"111100001",
  33030=>"101011000",
  33031=>"010100000",
  33032=>"010110110",
  33033=>"010101111",
  33034=>"111100001",
  33035=>"111101100",
  33036=>"011001100",
  33037=>"011000100",
  33038=>"011101101",
  33039=>"011001010",
  33040=>"101111110",
  33041=>"010110110",
  33042=>"001100110",
  33043=>"011101001",
  33044=>"111110010",
  33045=>"101101101",
  33046=>"000100011",
  33047=>"001011110",
  33048=>"000010100",
  33049=>"111000101",
  33050=>"101011111",
  33051=>"001011010",
  33052=>"111101111",
  33053=>"001000101",
  33054=>"101110010",
  33055=>"000111010",
  33056=>"101100000",
  33057=>"110101110",
  33058=>"000000000",
  33059=>"001100101",
  33060=>"110001001",
  33061=>"001100101",
  33062=>"011000110",
  33063=>"011100101",
  33064=>"010000011",
  33065=>"110010111",
  33066=>"111001110",
  33067=>"101001101",
  33068=>"111000100",
  33069=>"010110010",
  33070=>"001010000",
  33071=>"111100000",
  33072=>"111100101",
  33073=>"111111101",
  33074=>"110101101",
  33075=>"110000101",
  33076=>"001110110",
  33077=>"011000001",
  33078=>"101110001",
  33079=>"011101111",
  33080=>"101010111",
  33081=>"110000000",
  33082=>"100010100",
  33083=>"110111010",
  33084=>"011011000",
  33085=>"110101110",
  33086=>"101011000",
  33087=>"110010111",
  33088=>"001110011",
  33089=>"111010111",
  33090=>"000111011",
  33091=>"010101110",
  33092=>"000111111",
  33093=>"010010110",
  33094=>"011001101",
  33095=>"111000010",
  33096=>"000010001",
  33097=>"010110011",
  33098=>"011001011",
  33099=>"001011011",
  33100=>"101001110",
  33101=>"001000101",
  33102=>"000011110",
  33103=>"010110001",
  33104=>"000101000",
  33105=>"100111000",
  33106=>"110001000",
  33107=>"111101001",
  33108=>"000011000",
  33109=>"111100111",
  33110=>"111000000",
  33111=>"010110001",
  33112=>"011100000",
  33113=>"000010001",
  33114=>"110011011",
  33115=>"010000110",
  33116=>"101110111",
  33117=>"101100101",
  33118=>"100110110",
  33119=>"110000001",
  33120=>"011011000",
  33121=>"100001111",
  33122=>"010010000",
  33123=>"101001010",
  33124=>"000111101",
  33125=>"111010111",
  33126=>"101010011",
  33127=>"100000000",
  33128=>"011111010",
  33129=>"100000010",
  33130=>"101111101",
  33131=>"100000101",
  33132=>"111000011",
  33133=>"000010000",
  33134=>"100011110",
  33135=>"110101010",
  33136=>"001111111",
  33137=>"000000000",
  33138=>"010000001",
  33139=>"110010101",
  33140=>"101000110",
  33141=>"000100011",
  33142=>"011110000",
  33143=>"110111101",
  33144=>"000110111",
  33145=>"001111110",
  33146=>"100110001",
  33147=>"100010101",
  33148=>"000111111",
  33149=>"111111111",
  33150=>"010010000",
  33151=>"111110111",
  33152=>"110011111",
  33153=>"101010010",
  33154=>"100001111",
  33155=>"000110000",
  33156=>"101010011",
  33157=>"001000100",
  33158=>"101000111",
  33159=>"010010000",
  33160=>"010010001",
  33161=>"011010010",
  33162=>"010010001",
  33163=>"100001111",
  33164=>"011100111",
  33165=>"111110010",
  33166=>"000011000",
  33167=>"010100010",
  33168=>"111110010",
  33169=>"110110001",
  33170=>"100000010",
  33171=>"001011000",
  33172=>"111110100",
  33173=>"001101100",
  33174=>"010010000",
  33175=>"101111110",
  33176=>"000010000",
  33177=>"011000000",
  33178=>"110101101",
  33179=>"001000111",
  33180=>"110011100",
  33181=>"111100111",
  33182=>"101101010",
  33183=>"001001001",
  33184=>"001000111",
  33185=>"011100101",
  33186=>"110110101",
  33187=>"011101110",
  33188=>"110111010",
  33189=>"001111111",
  33190=>"011110111",
  33191=>"100101111",
  33192=>"110110001",
  33193=>"001100001",
  33194=>"101011110",
  33195=>"011000000",
  33196=>"110110010",
  33197=>"101011011",
  33198=>"101010110",
  33199=>"000010000",
  33200=>"101011101",
  33201=>"100001000",
  33202=>"101100001",
  33203=>"001000000",
  33204=>"110100010",
  33205=>"111111000",
  33206=>"100000010",
  33207=>"111111111",
  33208=>"011111000",
  33209=>"110100111",
  33210=>"011101010",
  33211=>"110110001",
  33212=>"100111110",
  33213=>"011000111",
  33214=>"111110001",
  33215=>"000000010",
  33216=>"110101111",
  33217=>"000100000",
  33218=>"100111111",
  33219=>"011001000",
  33220=>"111000111",
  33221=>"011101101",
  33222=>"100001111",
  33223=>"001000011",
  33224=>"101010100",
  33225=>"101011111",
  33226=>"011101111",
  33227=>"000011000",
  33228=>"000110101",
  33229=>"010001010",
  33230=>"111010000",
  33231=>"000100100",
  33232=>"010100010",
  33233=>"000001011",
  33234=>"001111100",
  33235=>"101000010",
  33236=>"111100001",
  33237=>"011111100",
  33238=>"111111011",
  33239=>"010000100",
  33240=>"010010101",
  33241=>"011001101",
  33242=>"000110011",
  33243=>"010100001",
  33244=>"000010101",
  33245=>"011001101",
  33246=>"001110000",
  33247=>"010000001",
  33248=>"000001110",
  33249=>"100001100",
  33250=>"011111101",
  33251=>"000110010",
  33252=>"101100000",
  33253=>"101000000",
  33254=>"100101111",
  33255=>"100011011",
  33256=>"000110001",
  33257=>"001001110",
  33258=>"111001111",
  33259=>"011001011",
  33260=>"010010100",
  33261=>"110111111",
  33262=>"111111001",
  33263=>"011100000",
  33264=>"000111010",
  33265=>"101011100",
  33266=>"101011100",
  33267=>"010010011",
  33268=>"110001001",
  33269=>"111100111",
  33270=>"000000110",
  33271=>"111110011",
  33272=>"010100100",
  33273=>"110011000",
  33274=>"111011101",
  33275=>"010111000",
  33276=>"110011011",
  33277=>"100000001",
  33278=>"100011101",
  33279=>"011001100",
  33280=>"101111110",
  33281=>"010010011",
  33282=>"000111111",
  33283=>"000001110",
  33284=>"111111110",
  33285=>"000001011",
  33286=>"011100101",
  33287=>"101111110",
  33288=>"111101001",
  33289=>"111010000",
  33290=>"111111111",
  33291=>"011100101",
  33292=>"101110111",
  33293=>"111000010",
  33294=>"010101000",
  33295=>"000100000",
  33296=>"011111100",
  33297=>"001101101",
  33298=>"001000000",
  33299=>"110100100",
  33300=>"110100101",
  33301=>"011010111",
  33302=>"101010010",
  33303=>"000000110",
  33304=>"011100101",
  33305=>"111011001",
  33306=>"111110100",
  33307=>"010001111",
  33308=>"001101011",
  33309=>"000010100",
  33310=>"100111011",
  33311=>"110110111",
  33312=>"000011010",
  33313=>"010100001",
  33314=>"110000100",
  33315=>"111000111",
  33316=>"111101101",
  33317=>"011111000",
  33318=>"111110111",
  33319=>"100100100",
  33320=>"000001101",
  33321=>"000110111",
  33322=>"001000110",
  33323=>"111010010",
  33324=>"110111111",
  33325=>"010111011",
  33326=>"101001010",
  33327=>"110111101",
  33328=>"100001000",
  33329=>"110011011",
  33330=>"110001010",
  33331=>"111100111",
  33332=>"101001010",
  33333=>"000110010",
  33334=>"101001011",
  33335=>"010001110",
  33336=>"100000000",
  33337=>"000110101",
  33338=>"010011010",
  33339=>"111000011",
  33340=>"111001001",
  33341=>"111000000",
  33342=>"011001000",
  33343=>"111010111",
  33344=>"111110111",
  33345=>"001010001",
  33346=>"111000110",
  33347=>"011101100",
  33348=>"010101101",
  33349=>"001101000",
  33350=>"100101001",
  33351=>"000000000",
  33352=>"010111111",
  33353=>"100110010",
  33354=>"101101100",
  33355=>"000001101",
  33356=>"010110100",
  33357=>"101101100",
  33358=>"001001111",
  33359=>"110010111",
  33360=>"001100010",
  33361=>"001001101",
  33362=>"100000001",
  33363=>"111100001",
  33364=>"100011001",
  33365=>"111100011",
  33366=>"001000111",
  33367=>"111000111",
  33368=>"111011010",
  33369=>"001110001",
  33370=>"110011100",
  33371=>"000100111",
  33372=>"000111101",
  33373=>"100000001",
  33374=>"010100101",
  33375=>"000100001",
  33376=>"010001010",
  33377=>"000011000",
  33378=>"001101010",
  33379=>"101000101",
  33380=>"100001000",
  33381=>"100011001",
  33382=>"001101011",
  33383=>"000110000",
  33384=>"100101010",
  33385=>"011110100",
  33386=>"101110110",
  33387=>"010111110",
  33388=>"001101101",
  33389=>"001111110",
  33390=>"100100001",
  33391=>"011000000",
  33392=>"111001011",
  33393=>"110001000",
  33394=>"000010011",
  33395=>"011110010",
  33396=>"000110011",
  33397=>"101110001",
  33398=>"001111000",
  33399=>"110010011",
  33400=>"101000011",
  33401=>"111100111",
  33402=>"010001101",
  33403=>"100101011",
  33404=>"001011001",
  33405=>"011010000",
  33406=>"111001010",
  33407=>"111101010",
  33408=>"111101001",
  33409=>"111000110",
  33410=>"101101010",
  33411=>"011010000",
  33412=>"011101000",
  33413=>"100010101",
  33414=>"110111001",
  33415=>"110011010",
  33416=>"101111001",
  33417=>"011111000",
  33418=>"100110100",
  33419=>"111001101",
  33420=>"111001001",
  33421=>"100000110",
  33422=>"111101100",
  33423=>"001000011",
  33424=>"000100001",
  33425=>"011000101",
  33426=>"110111011",
  33427=>"100001100",
  33428=>"000101110",
  33429=>"001101000",
  33430=>"111000011",
  33431=>"101010000",
  33432=>"100001100",
  33433=>"000001010",
  33434=>"011111110",
  33435=>"001100101",
  33436=>"100101011",
  33437=>"000110100",
  33438=>"111101100",
  33439=>"101011011",
  33440=>"110100001",
  33441=>"110110110",
  33442=>"010000010",
  33443=>"111010100",
  33444=>"110100100",
  33445=>"011101110",
  33446=>"011000010",
  33447=>"011011000",
  33448=>"111110000",
  33449=>"101100111",
  33450=>"101000100",
  33451=>"000011100",
  33452=>"010010001",
  33453=>"101001000",
  33454=>"101110100",
  33455=>"101000100",
  33456=>"011010000",
  33457=>"101011101",
  33458=>"001001100",
  33459=>"001100010",
  33460=>"110001110",
  33461=>"111010110",
  33462=>"100110001",
  33463=>"000010111",
  33464=>"110001000",
  33465=>"000011111",
  33466=>"001011100",
  33467=>"000011000",
  33468=>"111011001",
  33469=>"001011110",
  33470=>"111101101",
  33471=>"111100100",
  33472=>"111011111",
  33473=>"001111000",
  33474=>"000101100",
  33475=>"010001000",
  33476=>"101110001",
  33477=>"000001001",
  33478=>"110011100",
  33479=>"000100011",
  33480=>"100001010",
  33481=>"000100110",
  33482=>"100111011",
  33483=>"100001111",
  33484=>"011011110",
  33485=>"010111100",
  33486=>"000000111",
  33487=>"000010110",
  33488=>"001111111",
  33489=>"011101011",
  33490=>"101011101",
  33491=>"111101110",
  33492=>"100100100",
  33493=>"000111101",
  33494=>"011010001",
  33495=>"000101010",
  33496=>"010110011",
  33497=>"100010111",
  33498=>"000000000",
  33499=>"011000010",
  33500=>"001011000",
  33501=>"101110011",
  33502=>"100010000",
  33503=>"101100000",
  33504=>"110011010",
  33505=>"001010101",
  33506=>"101010110",
  33507=>"110010010",
  33508=>"000010011",
  33509=>"000001100",
  33510=>"011011110",
  33511=>"000000011",
  33512=>"111111100",
  33513=>"000100100",
  33514=>"000010011",
  33515=>"101100010",
  33516=>"010000100",
  33517=>"001010011",
  33518=>"101100010",
  33519=>"000111100",
  33520=>"000100011",
  33521=>"011011101",
  33522=>"011000110",
  33523=>"010010101",
  33524=>"010011111",
  33525=>"001000001",
  33526=>"110100011",
  33527=>"011111000",
  33528=>"111110000",
  33529=>"010100000",
  33530=>"001011111",
  33531=>"011000000",
  33532=>"111110111",
  33533=>"111100101",
  33534=>"000000010",
  33535=>"100111011",
  33536=>"000010011",
  33537=>"011101100",
  33538=>"110101110",
  33539=>"000000110",
  33540=>"100000101",
  33541=>"101010111",
  33542=>"111001110",
  33543=>"001001100",
  33544=>"001010100",
  33545=>"001110001",
  33546=>"111010000",
  33547=>"100110110",
  33548=>"100001101",
  33549=>"011110110",
  33550=>"011101100",
  33551=>"010011110",
  33552=>"111010101",
  33553=>"000100011",
  33554=>"011101110",
  33555=>"100011110",
  33556=>"101010010",
  33557=>"111000111",
  33558=>"000101000",
  33559=>"111001110",
  33560=>"100010010",
  33561=>"110001111",
  33562=>"001111110",
  33563=>"111101010",
  33564=>"100011001",
  33565=>"111001010",
  33566=>"100111110",
  33567=>"010100110",
  33568=>"110000111",
  33569=>"101011011",
  33570=>"000101100",
  33571=>"001010111",
  33572=>"010100010",
  33573=>"010100110",
  33574=>"111001110",
  33575=>"010011110",
  33576=>"000101110",
  33577=>"010100010",
  33578=>"100111001",
  33579=>"011011111",
  33580=>"011100011",
  33581=>"010111111",
  33582=>"101100000",
  33583=>"010001101",
  33584=>"101000111",
  33585=>"010001000",
  33586=>"011000001",
  33587=>"010111001",
  33588=>"111000111",
  33589=>"010110010",
  33590=>"111100011",
  33591=>"001101110",
  33592=>"101111000",
  33593=>"001011111",
  33594=>"111000000",
  33595=>"010010010",
  33596=>"010111001",
  33597=>"011000001",
  33598=>"010110101",
  33599=>"010001101",
  33600=>"101000001",
  33601=>"111010010",
  33602=>"000010000",
  33603=>"101011100",
  33604=>"000011101",
  33605=>"000011101",
  33606=>"110100111",
  33607=>"000000100",
  33608=>"101000111",
  33609=>"100101101",
  33610=>"100110001",
  33611=>"100110001",
  33612=>"000001011",
  33613=>"001001001",
  33614=>"101111111",
  33615=>"110000111",
  33616=>"100101000",
  33617=>"010011011",
  33618=>"011100100",
  33619=>"011101110",
  33620=>"101101011",
  33621=>"000001001",
  33622=>"011101110",
  33623=>"111101000",
  33624=>"111011100",
  33625=>"000110110",
  33626=>"100110101",
  33627=>"011011000",
  33628=>"000011010",
  33629=>"011101111",
  33630=>"001111100",
  33631=>"111110011",
  33632=>"100111101",
  33633=>"111101111",
  33634=>"010001111",
  33635=>"111011110",
  33636=>"000100110",
  33637=>"000101001",
  33638=>"111111000",
  33639=>"001111010",
  33640=>"011001001",
  33641=>"000010100",
  33642=>"000101101",
  33643=>"100001110",
  33644=>"100000000",
  33645=>"101010011",
  33646=>"001100110",
  33647=>"100100110",
  33648=>"111111011",
  33649=>"000000010",
  33650=>"010000001",
  33651=>"100110111",
  33652=>"001011101",
  33653=>"101011010",
  33654=>"100010010",
  33655=>"100000010",
  33656=>"101111001",
  33657=>"001110101",
  33658=>"011100110",
  33659=>"001111011",
  33660=>"101111101",
  33661=>"001001000",
  33662=>"000100010",
  33663=>"001110111",
  33664=>"101011000",
  33665=>"100110011",
  33666=>"000001001",
  33667=>"010101111",
  33668=>"111010111",
  33669=>"011001001",
  33670=>"101100001",
  33671=>"100010110",
  33672=>"100111100",
  33673=>"100011110",
  33674=>"011111100",
  33675=>"000001011",
  33676=>"011001000",
  33677=>"000001110",
  33678=>"111110000",
  33679=>"101111011",
  33680=>"100110110",
  33681=>"010101011",
  33682=>"101111110",
  33683=>"010000011",
  33684=>"101110010",
  33685=>"110010100",
  33686=>"111000011",
  33687=>"101010010",
  33688=>"011111000",
  33689=>"010110101",
  33690=>"000001000",
  33691=>"110100111",
  33692=>"011001101",
  33693=>"001000110",
  33694=>"111001001",
  33695=>"110010001",
  33696=>"001111010",
  33697=>"011100110",
  33698=>"110001111",
  33699=>"110010011",
  33700=>"001010011",
  33701=>"011100100",
  33702=>"111110101",
  33703=>"010010100",
  33704=>"001011011",
  33705=>"010011001",
  33706=>"101011110",
  33707=>"010001001",
  33708=>"110000011",
  33709=>"110011010",
  33710=>"101011111",
  33711=>"011110000",
  33712=>"001111100",
  33713=>"000001000",
  33714=>"011101110",
  33715=>"001001000",
  33716=>"110001110",
  33717=>"000000010",
  33718=>"110010111",
  33719=>"111011101",
  33720=>"111101000",
  33721=>"000101110",
  33722=>"101101001",
  33723=>"001100110",
  33724=>"001110111",
  33725=>"100111111",
  33726=>"110010110",
  33727=>"010101110",
  33728=>"011001011",
  33729=>"100110110",
  33730=>"001010100",
  33731=>"000110011",
  33732=>"010111010",
  33733=>"001001010",
  33734=>"111100111",
  33735=>"010010111",
  33736=>"011001011",
  33737=>"010110100",
  33738=>"111001111",
  33739=>"100110011",
  33740=>"100110111",
  33741=>"111101110",
  33742=>"101100001",
  33743=>"101001000",
  33744=>"110010011",
  33745=>"100001011",
  33746=>"000010011",
  33747=>"101011010",
  33748=>"010011111",
  33749=>"011000011",
  33750=>"101001000",
  33751=>"111001000",
  33752=>"110010110",
  33753=>"001010101",
  33754=>"010111011",
  33755=>"000001101",
  33756=>"101001101",
  33757=>"001011000",
  33758=>"100100110",
  33759=>"111111011",
  33760=>"010111110",
  33761=>"101101111",
  33762=>"011100101",
  33763=>"111110110",
  33764=>"000010110",
  33765=>"010001101",
  33766=>"011000101",
  33767=>"101100000",
  33768=>"001100111",
  33769=>"001111111",
  33770=>"100100101",
  33771=>"100100011",
  33772=>"011101101",
  33773=>"010011011",
  33774=>"100010011",
  33775=>"111010110",
  33776=>"010000001",
  33777=>"001011011",
  33778=>"000001101",
  33779=>"011110010",
  33780=>"011001100",
  33781=>"000110000",
  33782=>"011101110",
  33783=>"011101101",
  33784=>"111010111",
  33785=>"000100000",
  33786=>"110111001",
  33787=>"101111001",
  33788=>"100011101",
  33789=>"001100110",
  33790=>"101111111",
  33791=>"011100001",
  33792=>"100010100",
  33793=>"100110100",
  33794=>"110010010",
  33795=>"011100110",
  33796=>"010100111",
  33797=>"010000101",
  33798=>"111010011",
  33799=>"011110110",
  33800=>"011110110",
  33801=>"001000101",
  33802=>"001100101",
  33803=>"000001000",
  33804=>"111010100",
  33805=>"010011110",
  33806=>"110111001",
  33807=>"000101000",
  33808=>"101000000",
  33809=>"000000111",
  33810=>"001010000",
  33811=>"000110101",
  33812=>"010010000",
  33813=>"011111111",
  33814=>"101011111",
  33815=>"101101110",
  33816=>"010100011",
  33817=>"111000111",
  33818=>"110001111",
  33819=>"101111001",
  33820=>"001010100",
  33821=>"010101110",
  33822=>"011001110",
  33823=>"000100010",
  33824=>"010010000",
  33825=>"100111011",
  33826=>"000011110",
  33827=>"000111101",
  33828=>"001110111",
  33829=>"000010101",
  33830=>"011101111",
  33831=>"111110100",
  33832=>"011000100",
  33833=>"010100010",
  33834=>"011010111",
  33835=>"110001110",
  33836=>"001000001",
  33837=>"010100100",
  33838=>"000001000",
  33839=>"001001000",
  33840=>"011001101",
  33841=>"100100110",
  33842=>"100101001",
  33843=>"000011010",
  33844=>"101111110",
  33845=>"001001110",
  33846=>"000001010",
  33847=>"111110001",
  33848=>"011011001",
  33849=>"001111010",
  33850=>"100111111",
  33851=>"111101001",
  33852=>"101111100",
  33853=>"000101101",
  33854=>"011101001",
  33855=>"000001000",
  33856=>"110110001",
  33857=>"101111100",
  33858=>"101000111",
  33859=>"011011101",
  33860=>"010100101",
  33861=>"000000001",
  33862=>"110000000",
  33863=>"000101110",
  33864=>"000100100",
  33865=>"100001110",
  33866=>"111010011",
  33867=>"011011100",
  33868=>"011010100",
  33869=>"011101111",
  33870=>"111110011",
  33871=>"111011101",
  33872=>"111000011",
  33873=>"000100100",
  33874=>"110011110",
  33875=>"111011110",
  33876=>"011001110",
  33877=>"010001001",
  33878=>"100011110",
  33879=>"110101111",
  33880=>"001000110",
  33881=>"111011011",
  33882=>"011101101",
  33883=>"110101110",
  33884=>"001011010",
  33885=>"001010010",
  33886=>"100000100",
  33887=>"111011011",
  33888=>"000100111",
  33889=>"001110100",
  33890=>"111010101",
  33891=>"100101000",
  33892=>"010000110",
  33893=>"100000110",
  33894=>"100100010",
  33895=>"100010001",
  33896=>"000000000",
  33897=>"111010001",
  33898=>"101001100",
  33899=>"011110110",
  33900=>"101001000",
  33901=>"000000110",
  33902=>"101100100",
  33903=>"111101010",
  33904=>"110011100",
  33905=>"111001100",
  33906=>"001101010",
  33907=>"010110110",
  33908=>"010000011",
  33909=>"000010011",
  33910=>"100110011",
  33911=>"110110110",
  33912=>"001000010",
  33913=>"101100111",
  33914=>"001011100",
  33915=>"011010111",
  33916=>"000011001",
  33917=>"001010110",
  33918=>"111111000",
  33919=>"101001011",
  33920=>"111111111",
  33921=>"111100010",
  33922=>"000111100",
  33923=>"001000110",
  33924=>"100001010",
  33925=>"001111011",
  33926=>"001110110",
  33927=>"011000000",
  33928=>"100111100",
  33929=>"001011000",
  33930=>"000000001",
  33931=>"101101000",
  33932=>"111010100",
  33933=>"101011011",
  33934=>"100110011",
  33935=>"001111010",
  33936=>"010111000",
  33937=>"010101110",
  33938=>"000100011",
  33939=>"111111111",
  33940=>"111110011",
  33941=>"111111111",
  33942=>"101100000",
  33943=>"010110111",
  33944=>"001110010",
  33945=>"111100111",
  33946=>"101101010",
  33947=>"000011000",
  33948=>"110101111",
  33949=>"001100000",
  33950=>"100000000",
  33951=>"011100000",
  33952=>"100100000",
  33953=>"101100100",
  33954=>"111101111",
  33955=>"100110111",
  33956=>"001010010",
  33957=>"010101001",
  33958=>"111001111",
  33959=>"110010000",
  33960=>"101010001",
  33961=>"001010101",
  33962=>"111100111",
  33963=>"001010011",
  33964=>"110010000",
  33965=>"100110010",
  33966=>"010011010",
  33967=>"001011010",
  33968=>"000111000",
  33969=>"010110100",
  33970=>"000000001",
  33971=>"111011100",
  33972=>"001100100",
  33973=>"101111111",
  33974=>"110001110",
  33975=>"000111100",
  33976=>"001111010",
  33977=>"100110101",
  33978=>"100110010",
  33979=>"000111101",
  33980=>"001011111",
  33981=>"001001010",
  33982=>"101111000",
  33983=>"010000000",
  33984=>"010111111",
  33985=>"111011101",
  33986=>"110011000",
  33987=>"000000010",
  33988=>"111100001",
  33989=>"010111100",
  33990=>"111110010",
  33991=>"100101011",
  33992=>"111111111",
  33993=>"101100111",
  33994=>"101011010",
  33995=>"101000010",
  33996=>"010101001",
  33997=>"111111101",
  33998=>"011001111",
  33999=>"011010111",
  34000=>"101011010",
  34001=>"000000110",
  34002=>"110111101",
  34003=>"010001011",
  34004=>"100101111",
  34005=>"101010010",
  34006=>"111010111",
  34007=>"111001000",
  34008=>"110100000",
  34009=>"100011111",
  34010=>"010100111",
  34011=>"100101110",
  34012=>"101001110",
  34013=>"001111011",
  34014=>"000010000",
  34015=>"100011100",
  34016=>"101110101",
  34017=>"010001100",
  34018=>"111000101",
  34019=>"001000001",
  34020=>"000010110",
  34021=>"101000111",
  34022=>"000111101",
  34023=>"000010101",
  34024=>"111110010",
  34025=>"110110110",
  34026=>"110010111",
  34027=>"111011010",
  34028=>"010100110",
  34029=>"011000010",
  34030=>"000011101",
  34031=>"000111000",
  34032=>"111110010",
  34033=>"100000010",
  34034=>"100111110",
  34035=>"100100011",
  34036=>"101000101",
  34037=>"000101010",
  34038=>"111110101",
  34039=>"000001001",
  34040=>"101011111",
  34041=>"001001011",
  34042=>"001100011",
  34043=>"110111110",
  34044=>"001010111",
  34045=>"101100101",
  34046=>"101101110",
  34047=>"110110001",
  34048=>"101111101",
  34049=>"111110010",
  34050=>"111000011",
  34051=>"100110001",
  34052=>"100100100",
  34053=>"101000100",
  34054=>"110100100",
  34055=>"101000010",
  34056=>"010101011",
  34057=>"110101000",
  34058=>"000001101",
  34059=>"001111110",
  34060=>"010001000",
  34061=>"000111111",
  34062=>"010001000",
  34063=>"100110111",
  34064=>"101111000",
  34065=>"110110110",
  34066=>"001110011",
  34067=>"011100011",
  34068=>"001001000",
  34069=>"100110010",
  34070=>"110011001",
  34071=>"001101100",
  34072=>"001011001",
  34073=>"110000011",
  34074=>"010101111",
  34075=>"100110000",
  34076=>"011111010",
  34077=>"001001001",
  34078=>"110111110",
  34079=>"011000001",
  34080=>"000001001",
  34081=>"110010111",
  34082=>"000010100",
  34083=>"100011111",
  34084=>"000001001",
  34085=>"101010111",
  34086=>"101011000",
  34087=>"010100111",
  34088=>"101011010",
  34089=>"011111111",
  34090=>"001001011",
  34091=>"011101010",
  34092=>"010001000",
  34093=>"111110100",
  34094=>"100001010",
  34095=>"000010111",
  34096=>"110111110",
  34097=>"110011001",
  34098=>"011111000",
  34099=>"010000001",
  34100=>"110010010",
  34101=>"000100010",
  34102=>"000110110",
  34103=>"111111011",
  34104=>"000100010",
  34105=>"001101110",
  34106=>"101001100",
  34107=>"100110001",
  34108=>"100010100",
  34109=>"110111100",
  34110=>"110100001",
  34111=>"000110101",
  34112=>"110101101",
  34113=>"011100101",
  34114=>"100111000",
  34115=>"000010001",
  34116=>"011100111",
  34117=>"001100001",
  34118=>"001111001",
  34119=>"000100000",
  34120=>"100100001",
  34121=>"001100101",
  34122=>"101010101",
  34123=>"000100111",
  34124=>"001111101",
  34125=>"111101100",
  34126=>"111100001",
  34127=>"010001110",
  34128=>"100001000",
  34129=>"111111011",
  34130=>"010101101",
  34131=>"000010001",
  34132=>"001001001",
  34133=>"000110110",
  34134=>"001001001",
  34135=>"011110110",
  34136=>"111110010",
  34137=>"011100111",
  34138=>"111111011",
  34139=>"110110000",
  34140=>"101011011",
  34141=>"011100110",
  34142=>"000110001",
  34143=>"111110111",
  34144=>"100001111",
  34145=>"011111110",
  34146=>"110010001",
  34147=>"001001010",
  34148=>"010001101",
  34149=>"111001110",
  34150=>"101100001",
  34151=>"111111100",
  34152=>"101111001",
  34153=>"010010000",
  34154=>"010001111",
  34155=>"011001001",
  34156=>"000100011",
  34157=>"000011100",
  34158=>"000111110",
  34159=>"111110111",
  34160=>"100100110",
  34161=>"110100111",
  34162=>"111001010",
  34163=>"111001101",
  34164=>"000010100",
  34165=>"100101110",
  34166=>"101000110",
  34167=>"011001101",
  34168=>"000111010",
  34169=>"000000001",
  34170=>"001111001",
  34171=>"000000100",
  34172=>"010110101",
  34173=>"001001101",
  34174=>"010111110",
  34175=>"001110000",
  34176=>"000000101",
  34177=>"100000101",
  34178=>"100101110",
  34179=>"011011110",
  34180=>"111110010",
  34181=>"001000100",
  34182=>"111010101",
  34183=>"000100000",
  34184=>"101110111",
  34185=>"000101001",
  34186=>"110001110",
  34187=>"001010010",
  34188=>"100101101",
  34189=>"110010110",
  34190=>"000110011",
  34191=>"100101011",
  34192=>"111110100",
  34193=>"110001001",
  34194=>"011011110",
  34195=>"110011000",
  34196=>"100110000",
  34197=>"001101100",
  34198=>"111111110",
  34199=>"100110010",
  34200=>"010001001",
  34201=>"011100100",
  34202=>"010000111",
  34203=>"111100111",
  34204=>"101001010",
  34205=>"100010111",
  34206=>"100110010",
  34207=>"101001010",
  34208=>"111110100",
  34209=>"011101100",
  34210=>"101000001",
  34211=>"111000100",
  34212=>"000001111",
  34213=>"010010000",
  34214=>"001001001",
  34215=>"111100100",
  34216=>"010000011",
  34217=>"100000010",
  34218=>"110110000",
  34219=>"001111110",
  34220=>"101111110",
  34221=>"001111100",
  34222=>"011100101",
  34223=>"110110010",
  34224=>"000010000",
  34225=>"101011000",
  34226=>"000110010",
  34227=>"111011111",
  34228=>"111010111",
  34229=>"110110010",
  34230=>"101110001",
  34231=>"100001100",
  34232=>"100100110",
  34233=>"101011101",
  34234=>"111011111",
  34235=>"001100010",
  34236=>"000000000",
  34237=>"000101110",
  34238=>"101010000",
  34239=>"011010100",
  34240=>"000000101",
  34241=>"110010101",
  34242=>"100011001",
  34243=>"001001000",
  34244=>"101011111",
  34245=>"110111010",
  34246=>"011101101",
  34247=>"000100010",
  34248=>"100001001",
  34249=>"010110111",
  34250=>"001000101",
  34251=>"001000100",
  34252=>"111100111",
  34253=>"000111010",
  34254=>"100111001",
  34255=>"101111001",
  34256=>"111100011",
  34257=>"101111011",
  34258=>"101001000",
  34259=>"100101001",
  34260=>"101101001",
  34261=>"000111101",
  34262=>"000101001",
  34263=>"010000001",
  34264=>"011000101",
  34265=>"001010000",
  34266=>"110110001",
  34267=>"010100100",
  34268=>"110110110",
  34269=>"101001100",
  34270=>"101100100",
  34271=>"000110110",
  34272=>"000000011",
  34273=>"101001110",
  34274=>"000011111",
  34275=>"000000110",
  34276=>"010100011",
  34277=>"010011111",
  34278=>"010101110",
  34279=>"001101100",
  34280=>"011111110",
  34281=>"110011101",
  34282=>"000101100",
  34283=>"100111110",
  34284=>"001000001",
  34285=>"000010011",
  34286=>"010001010",
  34287=>"010010000",
  34288=>"010000100",
  34289=>"110111001",
  34290=>"101100110",
  34291=>"001000011",
  34292=>"101001010",
  34293=>"011101110",
  34294=>"011001001",
  34295=>"010001111",
  34296=>"011110010",
  34297=>"000000011",
  34298=>"010101100",
  34299=>"011000010",
  34300=>"101100000",
  34301=>"011011011",
  34302=>"001100111",
  34303=>"010000001",
  34304=>"011011010",
  34305=>"000000101",
  34306=>"001101010",
  34307=>"010100100",
  34308=>"110111111",
  34309=>"101000000",
  34310=>"001111011",
  34311=>"110111010",
  34312=>"001000001",
  34313=>"111111100",
  34314=>"010001101",
  34315=>"111111101",
  34316=>"011000000",
  34317=>"011101110",
  34318=>"101111101",
  34319=>"111101001",
  34320=>"001111111",
  34321=>"011001111",
  34322=>"111000010",
  34323=>"111100011",
  34324=>"100110011",
  34325=>"010001010",
  34326=>"000110001",
  34327=>"010011011",
  34328=>"000100010",
  34329=>"110000010",
  34330=>"101111111",
  34331=>"010100011",
  34332=>"010110000",
  34333=>"101101000",
  34334=>"000011100",
  34335=>"000110101",
  34336=>"100010110",
  34337=>"000110111",
  34338=>"000100101",
  34339=>"100101001",
  34340=>"011110001",
  34341=>"001000011",
  34342=>"110110010",
  34343=>"111101000",
  34344=>"000010001",
  34345=>"011000000",
  34346=>"100000100",
  34347=>"011010101",
  34348=>"000100111",
  34349=>"011010010",
  34350=>"100011111",
  34351=>"010001111",
  34352=>"000100110",
  34353=>"111000111",
  34354=>"101101011",
  34355=>"111100001",
  34356=>"001100000",
  34357=>"100001000",
  34358=>"101101011",
  34359=>"011000110",
  34360=>"111001010",
  34361=>"100000110",
  34362=>"010001000",
  34363=>"011010101",
  34364=>"111111111",
  34365=>"001110111",
  34366=>"111111110",
  34367=>"100111000",
  34368=>"001010101",
  34369=>"100000001",
  34370=>"011010000",
  34371=>"011000001",
  34372=>"111110000",
  34373=>"111011100",
  34374=>"011001111",
  34375=>"100111011",
  34376=>"010100000",
  34377=>"000100000",
  34378=>"000000001",
  34379=>"100111100",
  34380=>"010000000",
  34381=>"100011111",
  34382=>"101100101",
  34383=>"110101011",
  34384=>"011011011",
  34385=>"000001011",
  34386=>"110111111",
  34387=>"000010111",
  34388=>"011001110",
  34389=>"111101110",
  34390=>"010001110",
  34391=>"110101011",
  34392=>"001001001",
  34393=>"110100011",
  34394=>"100011010",
  34395=>"011110000",
  34396=>"011001110",
  34397=>"111011111",
  34398=>"110100111",
  34399=>"100000000",
  34400=>"110110111",
  34401=>"001011111",
  34402=>"111001000",
  34403=>"110000100",
  34404=>"110110110",
  34405=>"000011100",
  34406=>"111110011",
  34407=>"101110110",
  34408=>"001100010",
  34409=>"111100001",
  34410=>"111001111",
  34411=>"111001100",
  34412=>"000010111",
  34413=>"001110110",
  34414=>"000010010",
  34415=>"001011101",
  34416=>"000000001",
  34417=>"001010111",
  34418=>"101010111",
  34419=>"010000010",
  34420=>"111110011",
  34421=>"111100001",
  34422=>"101010110",
  34423=>"100010111",
  34424=>"111110110",
  34425=>"011001011",
  34426=>"111111011",
  34427=>"011001000",
  34428=>"110100000",
  34429=>"001000111",
  34430=>"000100111",
  34431=>"100000101",
  34432=>"101010111",
  34433=>"100111011",
  34434=>"001001100",
  34435=>"001011010",
  34436=>"010111000",
  34437=>"100111101",
  34438=>"010100001",
  34439=>"101010111",
  34440=>"010110111",
  34441=>"001011011",
  34442=>"110110101",
  34443=>"101110100",
  34444=>"101111111",
  34445=>"100100110",
  34446=>"101101110",
  34447=>"000000000",
  34448=>"000110001",
  34449=>"111001101",
  34450=>"001010101",
  34451=>"010010010",
  34452=>"100001101",
  34453=>"110101001",
  34454=>"110111101",
  34455=>"110101011",
  34456=>"011000100",
  34457=>"110011111",
  34458=>"000101101",
  34459=>"111011101",
  34460=>"010010001",
  34461=>"011010000",
  34462=>"111111100",
  34463=>"000010011",
  34464=>"100011111",
  34465=>"101000001",
  34466=>"111111110",
  34467=>"000011010",
  34468=>"101010100",
  34469=>"100101111",
  34470=>"110010001",
  34471=>"001010000",
  34472=>"111110010",
  34473=>"111011110",
  34474=>"001011101",
  34475=>"011101000",
  34476=>"001001010",
  34477=>"101011111",
  34478=>"101010101",
  34479=>"111110000",
  34480=>"101100010",
  34481=>"011100111",
  34482=>"101111001",
  34483=>"011100100",
  34484=>"001010011",
  34485=>"000101010",
  34486=>"011101100",
  34487=>"110001001",
  34488=>"000001001",
  34489=>"100000001",
  34490=>"110110010",
  34491=>"101110111",
  34492=>"111100011",
  34493=>"101101101",
  34494=>"001101010",
  34495=>"010100110",
  34496=>"101010011",
  34497=>"101101011",
  34498=>"110110111",
  34499=>"000001010",
  34500=>"011110000",
  34501=>"011011110",
  34502=>"100010101",
  34503=>"101101100",
  34504=>"101000100",
  34505=>"000001000",
  34506=>"001111011",
  34507=>"110101100",
  34508=>"000011101",
  34509=>"010100111",
  34510=>"000001010",
  34511=>"110011010",
  34512=>"101011011",
  34513=>"101001111",
  34514=>"111010011",
  34515=>"011110011",
  34516=>"101001110",
  34517=>"010010011",
  34518=>"110100011",
  34519=>"001010001",
  34520=>"111111000",
  34521=>"101011001",
  34522=>"110000000",
  34523=>"000000101",
  34524=>"110010110",
  34525=>"101010100",
  34526=>"011000101",
  34527=>"000010001",
  34528=>"100111110",
  34529=>"110000110",
  34530=>"011010000",
  34531=>"110100101",
  34532=>"011000111",
  34533=>"101001010",
  34534=>"001111101",
  34535=>"100101010",
  34536=>"000001001",
  34537=>"111010101",
  34538=>"101010110",
  34539=>"010110100",
  34540=>"000000001",
  34541=>"000011100",
  34542=>"111011010",
  34543=>"110011101",
  34544=>"001011011",
  34545=>"111011110",
  34546=>"100010100",
  34547=>"011101000",
  34548=>"000101100",
  34549=>"000000100",
  34550=>"011111011",
  34551=>"100001101",
  34552=>"011011101",
  34553=>"010010011",
  34554=>"100100111",
  34555=>"001011100",
  34556=>"111110000",
  34557=>"001110011",
  34558=>"100111110",
  34559=>"010010111",
  34560=>"111010110",
  34561=>"111110101",
  34562=>"111011110",
  34563=>"101101111",
  34564=>"001001010",
  34565=>"000000011",
  34566=>"101000101",
  34567=>"010000100",
  34568=>"000110000",
  34569=>"000000100",
  34570=>"011101001",
  34571=>"011000000",
  34572=>"010001001",
  34573=>"001111100",
  34574=>"111100101",
  34575=>"001010100",
  34576=>"001110111",
  34577=>"000001110",
  34578=>"101001101",
  34579=>"100010110",
  34580=>"101101101",
  34581=>"101101010",
  34582=>"011001000",
  34583=>"101100011",
  34584=>"000000000",
  34585=>"110101101",
  34586=>"110001101",
  34587=>"100111010",
  34588=>"011001011",
  34589=>"110101100",
  34590=>"101001111",
  34591=>"010011001",
  34592=>"111000010",
  34593=>"001101011",
  34594=>"010101011",
  34595=>"101100111",
  34596=>"010111011",
  34597=>"000010010",
  34598=>"011000100",
  34599=>"000110110",
  34600=>"111110110",
  34601=>"000101100",
  34602=>"001110000",
  34603=>"001011000",
  34604=>"000110111",
  34605=>"101111111",
  34606=>"010001001",
  34607=>"110011111",
  34608=>"111000100",
  34609=>"100100000",
  34610=>"011100110",
  34611=>"000011001",
  34612=>"100000000",
  34613=>"010110011",
  34614=>"111011011",
  34615=>"110000000",
  34616=>"101111101",
  34617=>"100100111",
  34618=>"000100101",
  34619=>"011111110",
  34620=>"001110100",
  34621=>"111000111",
  34622=>"011010111",
  34623=>"100010100",
  34624=>"101101101",
  34625=>"111001001",
  34626=>"010001100",
  34627=>"100111111",
  34628=>"000000000",
  34629=>"100010101",
  34630=>"000110010",
  34631=>"100001101",
  34632=>"011001011",
  34633=>"110101100",
  34634=>"001000100",
  34635=>"101100001",
  34636=>"001001010",
  34637=>"100001110",
  34638=>"010100001",
  34639=>"100111111",
  34640=>"000001000",
  34641=>"001000101",
  34642=>"011010111",
  34643=>"000001110",
  34644=>"001001000",
  34645=>"111100010",
  34646=>"011111011",
  34647=>"101011100",
  34648=>"110000111",
  34649=>"010001110",
  34650=>"000000010",
  34651=>"100101111",
  34652=>"011110001",
  34653=>"101011100",
  34654=>"001000100",
  34655=>"000000100",
  34656=>"010100010",
  34657=>"000001111",
  34658=>"001000100",
  34659=>"101000001",
  34660=>"111011000",
  34661=>"001101100",
  34662=>"101001011",
  34663=>"111111010",
  34664=>"001111101",
  34665=>"000101110",
  34666=>"100010110",
  34667=>"101010111",
  34668=>"010011111",
  34669=>"010001111",
  34670=>"010001000",
  34671=>"010000100",
  34672=>"010010100",
  34673=>"100001101",
  34674=>"000111101",
  34675=>"011101001",
  34676=>"001110110",
  34677=>"000111111",
  34678=>"110110111",
  34679=>"111010000",
  34680=>"010000001",
  34681=>"011100101",
  34682=>"011100101",
  34683=>"101101110",
  34684=>"000101010",
  34685=>"110111000",
  34686=>"001101111",
  34687=>"010100101",
  34688=>"111100110",
  34689=>"101110100",
  34690=>"010101010",
  34691=>"010000111",
  34692=>"110001101",
  34693=>"111001001",
  34694=>"001000101",
  34695=>"101011110",
  34696=>"010010011",
  34697=>"011100011",
  34698=>"000100100",
  34699=>"000011010",
  34700=>"010010100",
  34701=>"011111111",
  34702=>"011001001",
  34703=>"000110011",
  34704=>"110011000",
  34705=>"100111001",
  34706=>"111010001",
  34707=>"111101000",
  34708=>"100100010",
  34709=>"110101011",
  34710=>"000011010",
  34711=>"111110100",
  34712=>"011101100",
  34713=>"101110010",
  34714=>"001001110",
  34715=>"001000000",
  34716=>"001011000",
  34717=>"001011111",
  34718=>"010110001",
  34719=>"001111011",
  34720=>"010110011",
  34721=>"011100011",
  34722=>"110101110",
  34723=>"001000010",
  34724=>"100101001",
  34725=>"001011101",
  34726=>"011001101",
  34727=>"101100010",
  34728=>"010101111",
  34729=>"000101001",
  34730=>"010000101",
  34731=>"000000001",
  34732=>"011110011",
  34733=>"100101101",
  34734=>"000100010",
  34735=>"100100001",
  34736=>"000100011",
  34737=>"110110111",
  34738=>"101011111",
  34739=>"110000111",
  34740=>"011110011",
  34741=>"001111011",
  34742=>"000010000",
  34743=>"101101101",
  34744=>"000101000",
  34745=>"110000100",
  34746=>"111101111",
  34747=>"110011110",
  34748=>"101011001",
  34749=>"100110001",
  34750=>"011110011",
  34751=>"110011011",
  34752=>"100110110",
  34753=>"001000111",
  34754=>"000000111",
  34755=>"110111100",
  34756=>"001001011",
  34757=>"101010110",
  34758=>"101000000",
  34759=>"001100001",
  34760=>"001101110",
  34761=>"100001110",
  34762=>"110111001",
  34763=>"010010011",
  34764=>"110001001",
  34765=>"111001010",
  34766=>"100111111",
  34767=>"100010011",
  34768=>"011101100",
  34769=>"110100000",
  34770=>"100010111",
  34771=>"101001001",
  34772=>"110001000",
  34773=>"100110111",
  34774=>"101101011",
  34775=>"110111010",
  34776=>"000010110",
  34777=>"011011100",
  34778=>"110111111",
  34779=>"010110100",
  34780=>"011100001",
  34781=>"101001000",
  34782=>"011101010",
  34783=>"010010000",
  34784=>"101001010",
  34785=>"100000000",
  34786=>"000011101",
  34787=>"100010111",
  34788=>"010011110",
  34789=>"110101011",
  34790=>"111101110",
  34791=>"000000111",
  34792=>"001011111",
  34793=>"111111010",
  34794=>"101010110",
  34795=>"110100010",
  34796=>"111111111",
  34797=>"010111101",
  34798=>"111010000",
  34799=>"111110111",
  34800=>"001110010",
  34801=>"100011010",
  34802=>"001100001",
  34803=>"010011110",
  34804=>"011010001",
  34805=>"111110111",
  34806=>"001000010",
  34807=>"100011011",
  34808=>"001010000",
  34809=>"010001011",
  34810=>"101100101",
  34811=>"111000001",
  34812=>"110100000",
  34813=>"000010110",
  34814=>"111001011",
  34815=>"001010001",
  34816=>"101000000",
  34817=>"111011100",
  34818=>"001010110",
  34819=>"100010000",
  34820=>"110100101",
  34821=>"001010111",
  34822=>"110111111",
  34823=>"001100001",
  34824=>"010011100",
  34825=>"010101000",
  34826=>"010101000",
  34827=>"000111010",
  34828=>"111011100",
  34829=>"111010000",
  34830=>"011000011",
  34831=>"000000011",
  34832=>"000111111",
  34833=>"001100111",
  34834=>"001101011",
  34835=>"010000000",
  34836=>"000110001",
  34837=>"101001111",
  34838=>"100010110",
  34839=>"001000000",
  34840=>"000010110",
  34841=>"010001000",
  34842=>"100100101",
  34843=>"100010001",
  34844=>"101111111",
  34845=>"010001101",
  34846=>"000010010",
  34847=>"000000101",
  34848=>"010000111",
  34849=>"111111100",
  34850=>"010011111",
  34851=>"011011101",
  34852=>"101111110",
  34853=>"010110100",
  34854=>"111011001",
  34855=>"011011111",
  34856=>"000001011",
  34857=>"111100111",
  34858=>"110010101",
  34859=>"010000111",
  34860=>"000010110",
  34861=>"000110100",
  34862=>"000111000",
  34863=>"111101000",
  34864=>"111000010",
  34865=>"010010001",
  34866=>"001001111",
  34867=>"101111111",
  34868=>"101111110",
  34869=>"001011010",
  34870=>"110100101",
  34871=>"011001100",
  34872=>"101101000",
  34873=>"011101111",
  34874=>"111110111",
  34875=>"000010010",
  34876=>"011001011",
  34877=>"100101110",
  34878=>"000010000",
  34879=>"001101111",
  34880=>"010111011",
  34881=>"001110111",
  34882=>"110000101",
  34883=>"110010011",
  34884=>"100111100",
  34885=>"111111100",
  34886=>"000110000",
  34887=>"000111010",
  34888=>"000000000",
  34889=>"000110011",
  34890=>"000010110",
  34891=>"110000101",
  34892=>"110010001",
  34893=>"110111100",
  34894=>"011011111",
  34895=>"000101011",
  34896=>"010000010",
  34897=>"010110011",
  34898=>"011110110",
  34899=>"111000000",
  34900=>"110000110",
  34901=>"010010110",
  34902=>"100001110",
  34903=>"110011101",
  34904=>"101101000",
  34905=>"101100101",
  34906=>"100110100",
  34907=>"110010011",
  34908=>"111000111",
  34909=>"011001111",
  34910=>"111100010",
  34911=>"100000001",
  34912=>"110101111",
  34913=>"001111010",
  34914=>"010100011",
  34915=>"101111001",
  34916=>"110010000",
  34917=>"111011010",
  34918=>"110000011",
  34919=>"110111111",
  34920=>"011110110",
  34921=>"001101001",
  34922=>"111011001",
  34923=>"101011100",
  34924=>"010001001",
  34925=>"001111001",
  34926=>"011010011",
  34927=>"110011100",
  34928=>"010110110",
  34929=>"001110111",
  34930=>"000100010",
  34931=>"110111000",
  34932=>"111110101",
  34933=>"001001001",
  34934=>"101101111",
  34935=>"101101000",
  34936=>"011001010",
  34937=>"110010100",
  34938=>"000001010",
  34939=>"101010101",
  34940=>"110110110",
  34941=>"010101011",
  34942=>"011000100",
  34943=>"000001010",
  34944=>"010010010",
  34945=>"000110010",
  34946=>"111101010",
  34947=>"110011011",
  34948=>"101110001",
  34949=>"111111100",
  34950=>"100001000",
  34951=>"011001100",
  34952=>"011001100",
  34953=>"100011010",
  34954=>"000101010",
  34955=>"111110111",
  34956=>"011001101",
  34957=>"110111000",
  34958=>"001100000",
  34959=>"011110001",
  34960=>"000101101",
  34961=>"101010000",
  34962=>"000010010",
  34963=>"000001000",
  34964=>"100011010",
  34965=>"011000001",
  34966=>"000001100",
  34967=>"000101000",
  34968=>"111111111",
  34969=>"110011101",
  34970=>"000110111",
  34971=>"110001000",
  34972=>"110001111",
  34973=>"010100111",
  34974=>"010001101",
  34975=>"001100111",
  34976=>"010000001",
  34977=>"100100011",
  34978=>"101001011",
  34979=>"010001010",
  34980=>"111001111",
  34981=>"000000011",
  34982=>"011101110",
  34983=>"110000011",
  34984=>"011001101",
  34985=>"010011000",
  34986=>"111111000",
  34987=>"110111010",
  34988=>"010000101",
  34989=>"101100100",
  34990=>"000111000",
  34991=>"011010101",
  34992=>"011110000",
  34993=>"110110010",
  34994=>"011100110",
  34995=>"110110001",
  34996=>"000100000",
  34997=>"001101000",
  34998=>"101000110",
  34999=>"110001100",
  35000=>"000011000",
  35001=>"111001111",
  35002=>"110100101",
  35003=>"100100010",
  35004=>"101001101",
  35005=>"111001110",
  35006=>"011001001",
  35007=>"001001001",
  35008=>"101011101",
  35009=>"101101000",
  35010=>"100011110",
  35011=>"010010101",
  35012=>"110110100",
  35013=>"101000110",
  35014=>"000000100",
  35015=>"100110101",
  35016=>"000101101",
  35017=>"110101101",
  35018=>"100010010",
  35019=>"111001111",
  35020=>"000101011",
  35021=>"100101101",
  35022=>"110000110",
  35023=>"111100110",
  35024=>"100110011",
  35025=>"111010010",
  35026=>"111100101",
  35027=>"100011010",
  35028=>"001100000",
  35029=>"010100001",
  35030=>"011011111",
  35031=>"000101100",
  35032=>"011100111",
  35033=>"010111010",
  35034=>"010100111",
  35035=>"100111000",
  35036=>"001101010",
  35037=>"100001100",
  35038=>"001011110",
  35039=>"101100101",
  35040=>"000101000",
  35041=>"010010000",
  35042=>"101010100",
  35043=>"011101101",
  35044=>"001110110",
  35045=>"000001111",
  35046=>"110010100",
  35047=>"000001000",
  35048=>"111001100",
  35049=>"101111110",
  35050=>"100010101",
  35051=>"101111101",
  35052=>"010100110",
  35053=>"011000111",
  35054=>"010100101",
  35055=>"111011100",
  35056=>"110111100",
  35057=>"111010001",
  35058=>"010010101",
  35059=>"111110100",
  35060=>"110110100",
  35061=>"011000000",
  35062=>"110100000",
  35063=>"101111011",
  35064=>"001101011",
  35065=>"101011110",
  35066=>"100000010",
  35067=>"000100101",
  35068=>"000001000",
  35069=>"110010000",
  35070=>"110010010",
  35071=>"010000101",
  35072=>"100001010",
  35073=>"100011001",
  35074=>"101011010",
  35075=>"111010011",
  35076=>"000010100",
  35077=>"010100000",
  35078=>"110101100",
  35079=>"110010100",
  35080=>"110001011",
  35081=>"110101010",
  35082=>"100000101",
  35083=>"010111001",
  35084=>"011110111",
  35085=>"100001101",
  35086=>"110100101",
  35087=>"101100010",
  35088=>"011110110",
  35089=>"111010101",
  35090=>"101110000",
  35091=>"100011001",
  35092=>"010110010",
  35093=>"100110000",
  35094=>"110101110",
  35095=>"101010101",
  35096=>"101001100",
  35097=>"101111101",
  35098=>"001111000",
  35099=>"000011101",
  35100=>"000110111",
  35101=>"000000100",
  35102=>"101101011",
  35103=>"101011011",
  35104=>"010010110",
  35105=>"110000101",
  35106=>"101001111",
  35107=>"110000111",
  35108=>"001100100",
  35109=>"010100111",
  35110=>"000000000",
  35111=>"110110000",
  35112=>"101100010",
  35113=>"100001101",
  35114=>"001111111",
  35115=>"011101010",
  35116=>"101110001",
  35117=>"100101001",
  35118=>"010110100",
  35119=>"100110100",
  35120=>"010100001",
  35121=>"110111101",
  35122=>"000111111",
  35123=>"000101110",
  35124=>"011000011",
  35125=>"010110000",
  35126=>"101000000",
  35127=>"101011110",
  35128=>"111111111",
  35129=>"001011100",
  35130=>"100001100",
  35131=>"001101111",
  35132=>"001111111",
  35133=>"011110000",
  35134=>"001001001",
  35135=>"011100101",
  35136=>"011011010",
  35137=>"011101010",
  35138=>"000001000",
  35139=>"110100111",
  35140=>"110000010",
  35141=>"110010010",
  35142=>"100100001",
  35143=>"000000100",
  35144=>"101000001",
  35145=>"100100000",
  35146=>"100000100",
  35147=>"101000100",
  35148=>"011100001",
  35149=>"010101011",
  35150=>"110011111",
  35151=>"000010001",
  35152=>"110011010",
  35153=>"111101000",
  35154=>"101100011",
  35155=>"100011000",
  35156=>"111111111",
  35157=>"011000011",
  35158=>"111111111",
  35159=>"110001100",
  35160=>"101000010",
  35161=>"111100101",
  35162=>"000011001",
  35163=>"100011010",
  35164=>"000010010",
  35165=>"100111111",
  35166=>"111011101",
  35167=>"000011111",
  35168=>"100111000",
  35169=>"101011100",
  35170=>"111101001",
  35171=>"110010110",
  35172=>"011001011",
  35173=>"110100100",
  35174=>"101011000",
  35175=>"101101011",
  35176=>"010011011",
  35177=>"010000010",
  35178=>"100110111",
  35179=>"010101000",
  35180=>"110111100",
  35181=>"000000100",
  35182=>"011110011",
  35183=>"101001110",
  35184=>"111110000",
  35185=>"010010110",
  35186=>"010110100",
  35187=>"111100010",
  35188=>"010101111",
  35189=>"011011010",
  35190=>"000111010",
  35191=>"111101110",
  35192=>"111110111",
  35193=>"001011111",
  35194=>"111101101",
  35195=>"111111001",
  35196=>"000000110",
  35197=>"111011000",
  35198=>"110000011",
  35199=>"001110111",
  35200=>"110100101",
  35201=>"101001010",
  35202=>"000010011",
  35203=>"010100000",
  35204=>"000101101",
  35205=>"000111110",
  35206=>"000100011",
  35207=>"110100111",
  35208=>"011000110",
  35209=>"011010110",
  35210=>"100010000",
  35211=>"110001001",
  35212=>"011100111",
  35213=>"100001000",
  35214=>"010100111",
  35215=>"111111111",
  35216=>"111110010",
  35217=>"100001000",
  35218=>"101111000",
  35219=>"111011111",
  35220=>"000001000",
  35221=>"110101100",
  35222=>"001011010",
  35223=>"011111101",
  35224=>"011000001",
  35225=>"011111110",
  35226=>"010010111",
  35227=>"000001110",
  35228=>"010001101",
  35229=>"010000000",
  35230=>"111111110",
  35231=>"110101110",
  35232=>"101001001",
  35233=>"010100001",
  35234=>"111111000",
  35235=>"001111001",
  35236=>"001000011",
  35237=>"000001010",
  35238=>"111111001",
  35239=>"011110010",
  35240=>"111010101",
  35241=>"101110011",
  35242=>"100001110",
  35243=>"111100110",
  35244=>"000110010",
  35245=>"010010100",
  35246=>"111111110",
  35247=>"010010000",
  35248=>"111101011",
  35249=>"011101011",
  35250=>"100001001",
  35251=>"000111110",
  35252=>"010100000",
  35253=>"110010011",
  35254=>"000100000",
  35255=>"111011100",
  35256=>"111000111",
  35257=>"101010111",
  35258=>"010110111",
  35259=>"110101000",
  35260=>"010010000",
  35261=>"101001110",
  35262=>"110001110",
  35263=>"010100101",
  35264=>"001000000",
  35265=>"100111101",
  35266=>"111100010",
  35267=>"100000011",
  35268=>"110010110",
  35269=>"010000100",
  35270=>"000110001",
  35271=>"101011110",
  35272=>"101010111",
  35273=>"001110111",
  35274=>"111100000",
  35275=>"110011010",
  35276=>"111010101",
  35277=>"110110100",
  35278=>"011000011",
  35279=>"100001000",
  35280=>"011110010",
  35281=>"001100001",
  35282=>"010110110",
  35283=>"011111110",
  35284=>"001000100",
  35285=>"001101000",
  35286=>"111100000",
  35287=>"110111000",
  35288=>"110110111",
  35289=>"001011101",
  35290=>"001111011",
  35291=>"110100010",
  35292=>"001101111",
  35293=>"001010011",
  35294=>"110110011",
  35295=>"100111110",
  35296=>"100011011",
  35297=>"000010111",
  35298=>"110011111",
  35299=>"001000111",
  35300=>"101101101",
  35301=>"000100001",
  35302=>"110000100",
  35303=>"001101111",
  35304=>"111010110",
  35305=>"010010010",
  35306=>"111010110",
  35307=>"101001000",
  35308=>"010000111",
  35309=>"000100111",
  35310=>"100010000",
  35311=>"110110111",
  35312=>"101111011",
  35313=>"100100000",
  35314=>"011000110",
  35315=>"010111001",
  35316=>"010111001",
  35317=>"111100111",
  35318=>"100110011",
  35319=>"010110111",
  35320=>"100111010",
  35321=>"001100010",
  35322=>"101101111",
  35323=>"110101110",
  35324=>"110100100",
  35325=>"100001101",
  35326=>"001111110",
  35327=>"010000111",
  35328=>"100001101",
  35329=>"100100000",
  35330=>"010011100",
  35331=>"111001110",
  35332=>"110010100",
  35333=>"000111101",
  35334=>"011110001",
  35335=>"011000011",
  35336=>"110001010",
  35337=>"000110011",
  35338=>"111010111",
  35339=>"001010000",
  35340=>"100101001",
  35341=>"001010100",
  35342=>"001000111",
  35343=>"000110011",
  35344=>"100000000",
  35345=>"001001000",
  35346=>"001110101",
  35347=>"001001001",
  35348=>"110010101",
  35349=>"000110101",
  35350=>"100101000",
  35351=>"011010100",
  35352=>"111011111",
  35353=>"101001100",
  35354=>"010100101",
  35355=>"111101010",
  35356=>"000110001",
  35357=>"000111101",
  35358=>"110101100",
  35359=>"110010000",
  35360=>"110100110",
  35361=>"110110100",
  35362=>"111110110",
  35363=>"010000110",
  35364=>"010001110",
  35365=>"010000101",
  35366=>"101110011",
  35367=>"111110111",
  35368=>"011000101",
  35369=>"011011010",
  35370=>"110001111",
  35371=>"001110010",
  35372=>"000111111",
  35373=>"000101000",
  35374=>"010111110",
  35375=>"100011111",
  35376=>"001110110",
  35377=>"101000000",
  35378=>"110100000",
  35379=>"100110010",
  35380=>"011110010",
  35381=>"011110011",
  35382=>"110100000",
  35383=>"111010110",
  35384=>"111001010",
  35385=>"101011101",
  35386=>"000010000",
  35387=>"100011000",
  35388=>"101010011",
  35389=>"100100111",
  35390=>"000110100",
  35391=>"100111100",
  35392=>"111110001",
  35393=>"000100100",
  35394=>"110000000",
  35395=>"100110110",
  35396=>"101101000",
  35397=>"110010111",
  35398=>"110000000",
  35399=>"111011110",
  35400=>"110110111",
  35401=>"010111000",
  35402=>"111111110",
  35403=>"001110001",
  35404=>"000111011",
  35405=>"101100011",
  35406=>"100111111",
  35407=>"011110011",
  35408=>"111101100",
  35409=>"101110011",
  35410=>"100101000",
  35411=>"001001110",
  35412=>"000001010",
  35413=>"011001001",
  35414=>"010111111",
  35415=>"011101110",
  35416=>"110001001",
  35417=>"111110101",
  35418=>"010100110",
  35419=>"110101101",
  35420=>"111000011",
  35421=>"000000101",
  35422=>"101011101",
  35423=>"000001001",
  35424=>"100111100",
  35425=>"011001011",
  35426=>"000010000",
  35427=>"111100110",
  35428=>"110110101",
  35429=>"111011000",
  35430=>"101010001",
  35431=>"001101010",
  35432=>"010000111",
  35433=>"100000000",
  35434=>"011000100",
  35435=>"011001010",
  35436=>"011000010",
  35437=>"001010010",
  35438=>"010000011",
  35439=>"010000100",
  35440=>"010011110",
  35441=>"111101101",
  35442=>"010110001",
  35443=>"001100000",
  35444=>"101111110",
  35445=>"111011110",
  35446=>"000100000",
  35447=>"101000011",
  35448=>"000011101",
  35449=>"111100011",
  35450=>"110001011",
  35451=>"011010100",
  35452=>"000010111",
  35453=>"000001000",
  35454=>"001111111",
  35455=>"101111010",
  35456=>"110011010",
  35457=>"000101000",
  35458=>"010110011",
  35459=>"001011110",
  35460=>"101111100",
  35461=>"010110100",
  35462=>"111111001",
  35463=>"100011111",
  35464=>"101111100",
  35465=>"001000010",
  35466=>"111111101",
  35467=>"001111001",
  35468=>"000100010",
  35469=>"111000000",
  35470=>"100110001",
  35471=>"000100111",
  35472=>"010110000",
  35473=>"000101111",
  35474=>"001101000",
  35475=>"001111011",
  35476=>"000101111",
  35477=>"110011110",
  35478=>"111001110",
  35479=>"100001110",
  35480=>"011110010",
  35481=>"100000100",
  35482=>"000000001",
  35483=>"011010011",
  35484=>"110111010",
  35485=>"101110010",
  35486=>"000000111",
  35487=>"011100011",
  35488=>"001011011",
  35489=>"011101011",
  35490=>"000001101",
  35491=>"110110111",
  35492=>"010100010",
  35493=>"011100100",
  35494=>"111001100",
  35495=>"101111111",
  35496=>"001110101",
  35497=>"000100001",
  35498=>"111000110",
  35499=>"011010111",
  35500=>"010110000",
  35501=>"011010111",
  35502=>"000010001",
  35503=>"000110101",
  35504=>"010101000",
  35505=>"100001111",
  35506=>"111101000",
  35507=>"001001110",
  35508=>"110011110",
  35509=>"001101110",
  35510=>"110000010",
  35511=>"000010101",
  35512=>"010111111",
  35513=>"101101011",
  35514=>"011101001",
  35515=>"000011100",
  35516=>"010000100",
  35517=>"001011101",
  35518=>"100110111",
  35519=>"110011111",
  35520=>"111001010",
  35521=>"000101000",
  35522=>"111011011",
  35523=>"001100011",
  35524=>"010111010",
  35525=>"110000101",
  35526=>"101010100",
  35527=>"001010110",
  35528=>"000010010",
  35529=>"010001110",
  35530=>"011000000",
  35531=>"110011101",
  35532=>"100110001",
  35533=>"000100011",
  35534=>"111110100",
  35535=>"110000100",
  35536=>"000100011",
  35537=>"100110001",
  35538=>"100001010",
  35539=>"100011111",
  35540=>"001101101",
  35541=>"111110110",
  35542=>"010101100",
  35543=>"000010010",
  35544=>"010001010",
  35545=>"111110001",
  35546=>"011111101",
  35547=>"101101010",
  35548=>"101111110",
  35549=>"111111001",
  35550=>"001110111",
  35551=>"001011011",
  35552=>"101001000",
  35553=>"111011100",
  35554=>"101000010",
  35555=>"000111101",
  35556=>"100011110",
  35557=>"110010111",
  35558=>"111101010",
  35559=>"100001111",
  35560=>"010110011",
  35561=>"011101011",
  35562=>"001100010",
  35563=>"000110111",
  35564=>"110000101",
  35565=>"110011111",
  35566=>"101101110",
  35567=>"001110001",
  35568=>"000010110",
  35569=>"010010100",
  35570=>"111111000",
  35571=>"101011001",
  35572=>"010100000",
  35573=>"010001110",
  35574=>"000111011",
  35575=>"100011101",
  35576=>"000010110",
  35577=>"110010110",
  35578=>"000010000",
  35579=>"010011101",
  35580=>"000110000",
  35581=>"111111110",
  35582=>"001010110",
  35583=>"110001101",
  35584=>"100000111",
  35585=>"011011000",
  35586=>"110100111",
  35587=>"111001100",
  35588=>"011011100",
  35589=>"111111010",
  35590=>"111111010",
  35591=>"010000000",
  35592=>"000100011",
  35593=>"010001111",
  35594=>"000000010",
  35595=>"100011011",
  35596=>"001001001",
  35597=>"011110001",
  35598=>"001011000",
  35599=>"100010010",
  35600=>"101111110",
  35601=>"111000001",
  35602=>"111011001",
  35603=>"011101100",
  35604=>"011000011",
  35605=>"010000111",
  35606=>"100011100",
  35607=>"111000111",
  35608=>"110101111",
  35609=>"000110001",
  35610=>"110110010",
  35611=>"111101110",
  35612=>"101010111",
  35613=>"100000001",
  35614=>"011110000",
  35615=>"001000011",
  35616=>"011010011",
  35617=>"001110000",
  35618=>"101000100",
  35619=>"010100000",
  35620=>"101100001",
  35621=>"111100111",
  35622=>"000000000",
  35623=>"111011110",
  35624=>"010100011",
  35625=>"110011100",
  35626=>"010100010",
  35627=>"101000101",
  35628=>"110001101",
  35629=>"010011101",
  35630=>"100001100",
  35631=>"000000110",
  35632=>"100000110",
  35633=>"000000101",
  35634=>"101111111",
  35635=>"100011000",
  35636=>"111101011",
  35637=>"000001110",
  35638=>"000010010",
  35639=>"001010011",
  35640=>"110100011",
  35641=>"101011011",
  35642=>"010011101",
  35643=>"111111111",
  35644=>"111111010",
  35645=>"110011110",
  35646=>"110101010",
  35647=>"101010100",
  35648=>"111111001",
  35649=>"110010001",
  35650=>"000010000",
  35651=>"101111111",
  35652=>"010110011",
  35653=>"001000010",
  35654=>"110011100",
  35655=>"001111010",
  35656=>"110000001",
  35657=>"000000001",
  35658=>"100011001",
  35659=>"100011010",
  35660=>"010001110",
  35661=>"000101000",
  35662=>"101101101",
  35663=>"100110010",
  35664=>"110010111",
  35665=>"010001100",
  35666=>"110001100",
  35667=>"110011111",
  35668=>"100001111",
  35669=>"101111110",
  35670=>"001000101",
  35671=>"011001110",
  35672=>"110000000",
  35673=>"101100011",
  35674=>"101100000",
  35675=>"011001111",
  35676=>"010010101",
  35677=>"010011100",
  35678=>"010000001",
  35679=>"111101101",
  35680=>"110001101",
  35681=>"000111100",
  35682=>"110111001",
  35683=>"000000101",
  35684=>"101000011",
  35685=>"011010100",
  35686=>"001011101",
  35687=>"010110111",
  35688=>"101111111",
  35689=>"100001111",
  35690=>"110010010",
  35691=>"110000011",
  35692=>"100100111",
  35693=>"010101000",
  35694=>"000111001",
  35695=>"100001100",
  35696=>"110111111",
  35697=>"011100110",
  35698=>"000111000",
  35699=>"110011101",
  35700=>"010100100",
  35701=>"111111010",
  35702=>"011010011",
  35703=>"001100000",
  35704=>"010011000",
  35705=>"000101010",
  35706=>"000001001",
  35707=>"110110000",
  35708=>"010101110",
  35709=>"000111101",
  35710=>"100100101",
  35711=>"110011001",
  35712=>"001110011",
  35713=>"100111101",
  35714=>"110101011",
  35715=>"011000111",
  35716=>"000110100",
  35717=>"000001100",
  35718=>"001111111",
  35719=>"011111010",
  35720=>"111101010",
  35721=>"100111000",
  35722=>"010110011",
  35723=>"111111111",
  35724=>"000001101",
  35725=>"010110001",
  35726=>"011000000",
  35727=>"001010100",
  35728=>"101101000",
  35729=>"000000010",
  35730=>"011001111",
  35731=>"010110001",
  35732=>"010111011",
  35733=>"000101110",
  35734=>"100101101",
  35735=>"011010100",
  35736=>"000000000",
  35737=>"000010111",
  35738=>"011110101",
  35739=>"010010011",
  35740=>"001010010",
  35741=>"111110111",
  35742=>"101000111",
  35743=>"001100111",
  35744=>"011000101",
  35745=>"000100001",
  35746=>"011011110",
  35747=>"111111011",
  35748=>"010101001",
  35749=>"001101111",
  35750=>"111100110",
  35751=>"000001000",
  35752=>"111111110",
  35753=>"100000101",
  35754=>"111000001",
  35755=>"010111101",
  35756=>"100100111",
  35757=>"100000000",
  35758=>"011110001",
  35759=>"110000101",
  35760=>"100111010",
  35761=>"001010000",
  35762=>"000000011",
  35763=>"000100000",
  35764=>"000100011",
  35765=>"010101101",
  35766=>"100111110",
  35767=>"000001010",
  35768=>"110011000",
  35769=>"000001010",
  35770=>"001110110",
  35771=>"100111110",
  35772=>"111100011",
  35773=>"100001000",
  35774=>"000010010",
  35775=>"010101000",
  35776=>"100000100",
  35777=>"101100000",
  35778=>"011100111",
  35779=>"001010000",
  35780=>"000000000",
  35781=>"101101011",
  35782=>"110111011",
  35783=>"010101101",
  35784=>"000110000",
  35785=>"011110001",
  35786=>"101011001",
  35787=>"000111001",
  35788=>"010010011",
  35789=>"100001001",
  35790=>"110111010",
  35791=>"110100100",
  35792=>"010110000",
  35793=>"111111001",
  35794=>"101000110",
  35795=>"111011011",
  35796=>"111111110",
  35797=>"010110010",
  35798=>"000111111",
  35799=>"010101011",
  35800=>"000010001",
  35801=>"111101011",
  35802=>"110110111",
  35803=>"110010000",
  35804=>"001000000",
  35805=>"000001011",
  35806=>"010100111",
  35807=>"011000111",
  35808=>"011101101",
  35809=>"001001011",
  35810=>"000000010",
  35811=>"100011110",
  35812=>"110010010",
  35813=>"100110110",
  35814=>"000111100",
  35815=>"100111001",
  35816=>"111011011",
  35817=>"111011000",
  35818=>"101101011",
  35819=>"100010101",
  35820=>"000101000",
  35821=>"110011111",
  35822=>"111001001",
  35823=>"111010010",
  35824=>"101111010",
  35825=>"100101010",
  35826=>"111000000",
  35827=>"010010001",
  35828=>"111000010",
  35829=>"001000000",
  35830=>"011110111",
  35831=>"011011100",
  35832=>"000110010",
  35833=>"101011000",
  35834=>"110100110",
  35835=>"110011001",
  35836=>"010000010",
  35837=>"011100011",
  35838=>"110110011",
  35839=>"000011110",
  35840=>"011001100",
  35841=>"100001000",
  35842=>"100010101",
  35843=>"100101111",
  35844=>"111000000",
  35845=>"111101010",
  35846=>"010010011",
  35847=>"011110110",
  35848=>"000110111",
  35849=>"000101101",
  35850=>"001001000",
  35851=>"110010101",
  35852=>"100010000",
  35853=>"000111111",
  35854=>"001101101",
  35855=>"111100001",
  35856=>"001000001",
  35857=>"110011001",
  35858=>"110011000",
  35859=>"000110111",
  35860=>"101110001",
  35861=>"100110111",
  35862=>"010101111",
  35863=>"010110000",
  35864=>"000100110",
  35865=>"111101011",
  35866=>"011110100",
  35867=>"000011001",
  35868=>"101101101",
  35869=>"000011100",
  35870=>"011010101",
  35871=>"000101111",
  35872=>"011110001",
  35873=>"010011001",
  35874=>"010011011",
  35875=>"001111111",
  35876=>"010010000",
  35877=>"001000001",
  35878=>"011010011",
  35879=>"110111000",
  35880=>"111111001",
  35881=>"010000000",
  35882=>"110001100",
  35883=>"111000100",
  35884=>"000011011",
  35885=>"000101110",
  35886=>"011100001",
  35887=>"101110101",
  35888=>"010001010",
  35889=>"011110011",
  35890=>"001000101",
  35891=>"010111111",
  35892=>"101100110",
  35893=>"001111110",
  35894=>"110110111",
  35895=>"001111011",
  35896=>"001100001",
  35897=>"001000110",
  35898=>"000001111",
  35899=>"001011000",
  35900=>"010111001",
  35901=>"101001010",
  35902=>"001000111",
  35903=>"011111011",
  35904=>"101001110",
  35905=>"011110111",
  35906=>"100000010",
  35907=>"111000011",
  35908=>"000011001",
  35909=>"011000110",
  35910=>"110011101",
  35911=>"000100111",
  35912=>"100110000",
  35913=>"000101101",
  35914=>"001000011",
  35915=>"011001101",
  35916=>"100000010",
  35917=>"000000101",
  35918=>"011101111",
  35919=>"000101001",
  35920=>"010100000",
  35921=>"100101000",
  35922=>"101110000",
  35923=>"101010100",
  35924=>"011110101",
  35925=>"011010001",
  35926=>"000001010",
  35927=>"011110101",
  35928=>"110001000",
  35929=>"000111101",
  35930=>"001010011",
  35931=>"110111101",
  35932=>"000001101",
  35933=>"110000000",
  35934=>"110111100",
  35935=>"011001111",
  35936=>"010001010",
  35937=>"101111000",
  35938=>"110000101",
  35939=>"011000000",
  35940=>"000010111",
  35941=>"001010101",
  35942=>"011000001",
  35943=>"011101101",
  35944=>"101111001",
  35945=>"100000000",
  35946=>"101011101",
  35947=>"100101110",
  35948=>"100100111",
  35949=>"110000001",
  35950=>"000000010",
  35951=>"101000010",
  35952=>"111010011",
  35953=>"111011011",
  35954=>"101100101",
  35955=>"110101100",
  35956=>"110100011",
  35957=>"101111010",
  35958=>"010000000",
  35959=>"101100011",
  35960=>"010010000",
  35961=>"110001100",
  35962=>"111100000",
  35963=>"001011000",
  35964=>"101000001",
  35965=>"110011101",
  35966=>"110000100",
  35967=>"111111111",
  35968=>"110100111",
  35969=>"010010010",
  35970=>"111001010",
  35971=>"001001110",
  35972=>"101111110",
  35973=>"011100000",
  35974=>"000011011",
  35975=>"000011010",
  35976=>"111001010",
  35977=>"001100011",
  35978=>"101000111",
  35979=>"111010110",
  35980=>"010100100",
  35981=>"101010100",
  35982=>"001011111",
  35983=>"111001000",
  35984=>"010000000",
  35985=>"001011011",
  35986=>"000000001",
  35987=>"111110001",
  35988=>"000011101",
  35989=>"010001111",
  35990=>"010011111",
  35991=>"110100010",
  35992=>"010101010",
  35993=>"101111111",
  35994=>"110001000",
  35995=>"011010100",
  35996=>"001001010",
  35997=>"110101111",
  35998=>"000100111",
  35999=>"100101100",
  36000=>"100001011",
  36001=>"101100000",
  36002=>"010000101",
  36003=>"110111110",
  36004=>"101101010",
  36005=>"011000010",
  36006=>"101011110",
  36007=>"000000010",
  36008=>"100010110",
  36009=>"101011101",
  36010=>"111111111",
  36011=>"011011000",
  36012=>"110110111",
  36013=>"110001100",
  36014=>"000000010",
  36015=>"110000011",
  36016=>"001010001",
  36017=>"010000001",
  36018=>"111010010",
  36019=>"011001100",
  36020=>"101001111",
  36021=>"100001000",
  36022=>"010000011",
  36023=>"101010100",
  36024=>"010101100",
  36025=>"101000111",
  36026=>"010111010",
  36027=>"111010111",
  36028=>"001000110",
  36029=>"000000001",
  36030=>"111110011",
  36031=>"101001011",
  36032=>"010101100",
  36033=>"100100011",
  36034=>"001011101",
  36035=>"000011001",
  36036=>"000011011",
  36037=>"011011100",
  36038=>"101010011",
  36039=>"000000001",
  36040=>"111000010",
  36041=>"000101110",
  36042=>"111000001",
  36043=>"000011100",
  36044=>"101110000",
  36045=>"110110100",
  36046=>"011111100",
  36047=>"101101000",
  36048=>"011101101",
  36049=>"001011101",
  36050=>"000000010",
  36051=>"000011011",
  36052=>"010110011",
  36053=>"010011001",
  36054=>"011111001",
  36055=>"110111011",
  36056=>"101000100",
  36057=>"010110010",
  36058=>"011110110",
  36059=>"111111010",
  36060=>"001000110",
  36061=>"101001110",
  36062=>"110110001",
  36063=>"000010111",
  36064=>"001001100",
  36065=>"110000001",
  36066=>"000111000",
  36067=>"001000011",
  36068=>"100000000",
  36069=>"001000100",
  36070=>"111111101",
  36071=>"100101101",
  36072=>"011101010",
  36073=>"100110000",
  36074=>"011010100",
  36075=>"001100111",
  36076=>"000101000",
  36077=>"000110111",
  36078=>"000100101",
  36079=>"000111111",
  36080=>"011100001",
  36081=>"101111110",
  36082=>"000101110",
  36083=>"111100111",
  36084=>"100010101",
  36085=>"000101010",
  36086=>"111101011",
  36087=>"111110001",
  36088=>"110100000",
  36089=>"101100101",
  36090=>"100011000",
  36091=>"011010001",
  36092=>"001100001",
  36093=>"011110010",
  36094=>"111111010",
  36095=>"000100111",
  36096=>"011101110",
  36097=>"010001100",
  36098=>"000010111",
  36099=>"000111110",
  36100=>"001001010",
  36101=>"100111100",
  36102=>"001110010",
  36103=>"001010000",
  36104=>"100101010",
  36105=>"110000010",
  36106=>"101100110",
  36107=>"100100000",
  36108=>"110000110",
  36109=>"110100101",
  36110=>"011000011",
  36111=>"101010001",
  36112=>"110010001",
  36113=>"110001001",
  36114=>"100011011",
  36115=>"001111011",
  36116=>"000100110",
  36117=>"000011101",
  36118=>"111010001",
  36119=>"101110110",
  36120=>"110000010",
  36121=>"001001100",
  36122=>"110100110",
  36123=>"111000111",
  36124=>"010101001",
  36125=>"001100111",
  36126=>"011111010",
  36127=>"110001000",
  36128=>"100111001",
  36129=>"111001111",
  36130=>"100010101",
  36131=>"111111000",
  36132=>"111001111",
  36133=>"110011010",
  36134=>"001100000",
  36135=>"101110110",
  36136=>"011101001",
  36137=>"111010010",
  36138=>"110101000",
  36139=>"110111110",
  36140=>"001010100",
  36141=>"110000001",
  36142=>"011001110",
  36143=>"110110000",
  36144=>"111111010",
  36145=>"000101110",
  36146=>"111101010",
  36147=>"000010101",
  36148=>"111100101",
  36149=>"111100101",
  36150=>"110011100",
  36151=>"111111111",
  36152=>"101001000",
  36153=>"001011110",
  36154=>"000111100",
  36155=>"101011001",
  36156=>"101011010",
  36157=>"000110110",
  36158=>"111001101",
  36159=>"111011010",
  36160=>"010100100",
  36161=>"011010010",
  36162=>"010101000",
  36163=>"010000011",
  36164=>"011011000",
  36165=>"010111001",
  36166=>"100000001",
  36167=>"000000100",
  36168=>"000010111",
  36169=>"110111011",
  36170=>"110010101",
  36171=>"100111001",
  36172=>"000010011",
  36173=>"000100100",
  36174=>"011101101",
  36175=>"111000100",
  36176=>"011010010",
  36177=>"111110001",
  36178=>"001111001",
  36179=>"100001001",
  36180=>"011101010",
  36181=>"101001001",
  36182=>"110100111",
  36183=>"110000101",
  36184=>"100011100",
  36185=>"110100010",
  36186=>"000001100",
  36187=>"100011000",
  36188=>"111011110",
  36189=>"101000000",
  36190=>"101011001",
  36191=>"100001001",
  36192=>"001000100",
  36193=>"001011101",
  36194=>"111100111",
  36195=>"111010001",
  36196=>"110100100",
  36197=>"110001000",
  36198=>"000101101",
  36199=>"011001000",
  36200=>"110101010",
  36201=>"001111011",
  36202=>"000001111",
  36203=>"101111010",
  36204=>"001001001",
  36205=>"111110110",
  36206=>"011110111",
  36207=>"101101111",
  36208=>"110001001",
  36209=>"011010110",
  36210=>"110110001",
  36211=>"100110000",
  36212=>"100100001",
  36213=>"101001000",
  36214=>"010001101",
  36215=>"001001110",
  36216=>"000111001",
  36217=>"100011010",
  36218=>"111011101",
  36219=>"110001111",
  36220=>"001000101",
  36221=>"011101010",
  36222=>"111100001",
  36223=>"111101010",
  36224=>"001011000",
  36225=>"111000111",
  36226=>"110110011",
  36227=>"000011010",
  36228=>"111010000",
  36229=>"111111100",
  36230=>"000110001",
  36231=>"001111001",
  36232=>"011110100",
  36233=>"000101001",
  36234=>"101110001",
  36235=>"100010000",
  36236=>"101111000",
  36237=>"000100101",
  36238=>"111101000",
  36239=>"001111010",
  36240=>"001000100",
  36241=>"111100001",
  36242=>"110010100",
  36243=>"111001100",
  36244=>"011110001",
  36245=>"000000011",
  36246=>"110101100",
  36247=>"111000000",
  36248=>"010000111",
  36249=>"010011101",
  36250=>"101111011",
  36251=>"100111011",
  36252=>"010101110",
  36253=>"101011000",
  36254=>"100111110",
  36255=>"100011000",
  36256=>"001001110",
  36257=>"011110100",
  36258=>"111101000",
  36259=>"010111010",
  36260=>"011111101",
  36261=>"101011011",
  36262=>"111000110",
  36263=>"000011010",
  36264=>"000100101",
  36265=>"001100111",
  36266=>"001001011",
  36267=>"100000011",
  36268=>"000010111",
  36269=>"101101010",
  36270=>"001100000",
  36271=>"001110111",
  36272=>"110010101",
  36273=>"000000110",
  36274=>"001100001",
  36275=>"001100001",
  36276=>"001100000",
  36277=>"010000111",
  36278=>"110000011",
  36279=>"110001000",
  36280=>"110111111",
  36281=>"111101011",
  36282=>"001011011",
  36283=>"000110110",
  36284=>"000001101",
  36285=>"101011110",
  36286=>"100110111",
  36287=>"101011010",
  36288=>"110100000",
  36289=>"101110001",
  36290=>"111010111",
  36291=>"111111010",
  36292=>"001010011",
  36293=>"011001000",
  36294=>"001010100",
  36295=>"011101111",
  36296=>"010011111",
  36297=>"110100101",
  36298=>"111000010",
  36299=>"001111000",
  36300=>"000001101",
  36301=>"100100010",
  36302=>"011000000",
  36303=>"100011010",
  36304=>"001001010",
  36305=>"001011111",
  36306=>"011011001",
  36307=>"000100000",
  36308=>"010011111",
  36309=>"111011001",
  36310=>"011110111",
  36311=>"111000100",
  36312=>"000000111",
  36313=>"000001010",
  36314=>"000101110",
  36315=>"000010011",
  36316=>"110000010",
  36317=>"110001011",
  36318=>"001000111",
  36319=>"001001110",
  36320=>"101101011",
  36321=>"101101010",
  36322=>"110100000",
  36323=>"000011011",
  36324=>"111111001",
  36325=>"011110100",
  36326=>"110001100",
  36327=>"000000101",
  36328=>"010010001",
  36329=>"000011101",
  36330=>"110101000",
  36331=>"000111010",
  36332=>"000100010",
  36333=>"100110011",
  36334=>"011010011",
  36335=>"011101101",
  36336=>"000101010",
  36337=>"101001100",
  36338=>"100010100",
  36339=>"000010000",
  36340=>"100010111",
  36341=>"010011000",
  36342=>"011100111",
  36343=>"010111100",
  36344=>"010110001",
  36345=>"111001001",
  36346=>"010010000",
  36347=>"100000000",
  36348=>"101000101",
  36349=>"001000101",
  36350=>"001000100",
  36351=>"111010110",
  36352=>"100110001",
  36353=>"010111100",
  36354=>"111011110",
  36355=>"001101001",
  36356=>"001001000",
  36357=>"111111110",
  36358=>"000001110",
  36359=>"100111010",
  36360=>"110000111",
  36361=>"100101011",
  36362=>"101101110",
  36363=>"010110000",
  36364=>"100110011",
  36365=>"100001001",
  36366=>"101110000",
  36367=>"000010011",
  36368=>"110001011",
  36369=>"010010110",
  36370=>"000001010",
  36371=>"101001000",
  36372=>"100101111",
  36373=>"101100111",
  36374=>"011111111",
  36375=>"000000010",
  36376=>"111010100",
  36377=>"000110000",
  36378=>"110101111",
  36379=>"001110100",
  36380=>"101111111",
  36381=>"111011111",
  36382=>"001110001",
  36383=>"100110001",
  36384=>"111000100",
  36385=>"001000010",
  36386=>"011101101",
  36387=>"101010111",
  36388=>"010110100",
  36389=>"000010100",
  36390=>"111101110",
  36391=>"010001011",
  36392=>"111110000",
  36393=>"000011111",
  36394=>"001110100",
  36395=>"110000000",
  36396=>"000100111",
  36397=>"010001100",
  36398=>"111110111",
  36399=>"000011001",
  36400=>"111001101",
  36401=>"011011100",
  36402=>"000101000",
  36403=>"000010000",
  36404=>"110011001",
  36405=>"111001101",
  36406=>"001010100",
  36407=>"000111001",
  36408=>"111101011",
  36409=>"000000011",
  36410=>"101110110",
  36411=>"110111100",
  36412=>"010000000",
  36413=>"101000000",
  36414=>"111111001",
  36415=>"010000110",
  36416=>"011001010",
  36417=>"000000001",
  36418=>"011111010",
  36419=>"100101011",
  36420=>"111111101",
  36421=>"101100000",
  36422=>"011111110",
  36423=>"110101001",
  36424=>"101010010",
  36425=>"001100000",
  36426=>"011110111",
  36427=>"000000100",
  36428=>"101011100",
  36429=>"110110101",
  36430=>"001010010",
  36431=>"111111010",
  36432=>"001000000",
  36433=>"101011110",
  36434=>"111000001",
  36435=>"010111100",
  36436=>"001010101",
  36437=>"010010110",
  36438=>"000110011",
  36439=>"100001001",
  36440=>"010101100",
  36441=>"010011010",
  36442=>"110110111",
  36443=>"101111101",
  36444=>"010011111",
  36445=>"010110100",
  36446=>"011110111",
  36447=>"101101111",
  36448=>"110111011",
  36449=>"011101001",
  36450=>"110010011",
  36451=>"010111001",
  36452=>"010010011",
  36453=>"100010000",
  36454=>"110001100",
  36455=>"101010100",
  36456=>"010100000",
  36457=>"110000000",
  36458=>"000111010",
  36459=>"111010000",
  36460=>"111111010",
  36461=>"101101010",
  36462=>"011001010",
  36463=>"001001110",
  36464=>"100110111",
  36465=>"101101110",
  36466=>"010101111",
  36467=>"111110101",
  36468=>"011111001",
  36469=>"101110011",
  36470=>"111110111",
  36471=>"001000100",
  36472=>"011011111",
  36473=>"011110000",
  36474=>"111101110",
  36475=>"101111011",
  36476=>"110011111",
  36477=>"111000001",
  36478=>"000010000",
  36479=>"101000010",
  36480=>"001101011",
  36481=>"110110100",
  36482=>"001001000",
  36483=>"101100001",
  36484=>"110100111",
  36485=>"010011101",
  36486=>"100111100",
  36487=>"110101100",
  36488=>"001000011",
  36489=>"010000101",
  36490=>"010001110",
  36491=>"000010011",
  36492=>"101110111",
  36493=>"111100101",
  36494=>"110100001",
  36495=>"100011001",
  36496=>"000111000",
  36497=>"001101001",
  36498=>"010001111",
  36499=>"011010101",
  36500=>"010000011",
  36501=>"000101011",
  36502=>"011100000",
  36503=>"011010000",
  36504=>"111111011",
  36505=>"110110101",
  36506=>"111010101",
  36507=>"011110011",
  36508=>"111111010",
  36509=>"101000110",
  36510=>"110110110",
  36511=>"110110011",
  36512=>"101010111",
  36513=>"111000110",
  36514=>"101101010",
  36515=>"010010010",
  36516=>"000101100",
  36517=>"101000100",
  36518=>"010000111",
  36519=>"111110011",
  36520=>"100100101",
  36521=>"001111111",
  36522=>"100100000",
  36523=>"101101000",
  36524=>"101001010",
  36525=>"110100000",
  36526=>"010101011",
  36527=>"111001111",
  36528=>"011100000",
  36529=>"001100010",
  36530=>"010111000",
  36531=>"010001110",
  36532=>"010101010",
  36533=>"010110110",
  36534=>"100011011",
  36535=>"111011100",
  36536=>"011010100",
  36537=>"100110101",
  36538=>"100101001",
  36539=>"011000000",
  36540=>"101111111",
  36541=>"011110000",
  36542=>"011111001",
  36543=>"000010010",
  36544=>"111111010",
  36545=>"010011011",
  36546=>"100010000",
  36547=>"000100111",
  36548=>"001110100",
  36549=>"101101110",
  36550=>"100111110",
  36551=>"101100011",
  36552=>"100111100",
  36553=>"011100000",
  36554=>"100101111",
  36555=>"100111011",
  36556=>"101001011",
  36557=>"011010111",
  36558=>"101001101",
  36559=>"000100101",
  36560=>"001011010",
  36561=>"111000011",
  36562=>"011110110",
  36563=>"011110001",
  36564=>"001111001",
  36565=>"101000000",
  36566=>"100001111",
  36567=>"101011011",
  36568=>"101101111",
  36569=>"100010010",
  36570=>"100011000",
  36571=>"110011001",
  36572=>"101011100",
  36573=>"100000111",
  36574=>"010101110",
  36575=>"010001111",
  36576=>"111000100",
  36577=>"011101110",
  36578=>"001111000",
  36579=>"110010001",
  36580=>"011001011",
  36581=>"010000011",
  36582=>"001111101",
  36583=>"101001001",
  36584=>"011010101",
  36585=>"101111000",
  36586=>"010111011",
  36587=>"110010010",
  36588=>"000001111",
  36589=>"011111000",
  36590=>"110110100",
  36591=>"010001001",
  36592=>"001110100",
  36593=>"011011100",
  36594=>"101000010",
  36595=>"100100000",
  36596=>"010100111",
  36597=>"110111010",
  36598=>"111111101",
  36599=>"010011011",
  36600=>"100010100",
  36601=>"110111100",
  36602=>"011110110",
  36603=>"101110001",
  36604=>"001111111",
  36605=>"010101011",
  36606=>"111001011",
  36607=>"000101111",
  36608=>"011010010",
  36609=>"010101110",
  36610=>"110110110",
  36611=>"000111011",
  36612=>"001100101",
  36613=>"110001011",
  36614=>"000101001",
  36615=>"001011110",
  36616=>"011111011",
  36617=>"111001100",
  36618=>"111110010",
  36619=>"010101000",
  36620=>"000001110",
  36621=>"100001010",
  36622=>"100001010",
  36623=>"110001000",
  36624=>"001110111",
  36625=>"101001110",
  36626=>"110110000",
  36627=>"011010001",
  36628=>"000000110",
  36629=>"101001010",
  36630=>"101010011",
  36631=>"110001101",
  36632=>"001011001",
  36633=>"111000111",
  36634=>"000100110",
  36635=>"101001010",
  36636=>"011000101",
  36637=>"100010100",
  36638=>"101010110",
  36639=>"000111010",
  36640=>"101001011",
  36641=>"111110111",
  36642=>"111100101",
  36643=>"001100001",
  36644=>"110011101",
  36645=>"100110100",
  36646=>"110010000",
  36647=>"000101100",
  36648=>"101101101",
  36649=>"111111010",
  36650=>"011000100",
  36651=>"101011001",
  36652=>"111110100",
  36653=>"001000010",
  36654=>"000100010",
  36655=>"110100101",
  36656=>"010000011",
  36657=>"101100100",
  36658=>"001000101",
  36659=>"111111101",
  36660=>"001011111",
  36661=>"110010101",
  36662=>"011100100",
  36663=>"111101001",
  36664=>"110110110",
  36665=>"100111010",
  36666=>"110100110",
  36667=>"111011100",
  36668=>"011010000",
  36669=>"010011111",
  36670=>"111001110",
  36671=>"000100101",
  36672=>"010011001",
  36673=>"010010110",
  36674=>"111110000",
  36675=>"011001000",
  36676=>"011111111",
  36677=>"010101001",
  36678=>"101111111",
  36679=>"001100100",
  36680=>"011101000",
  36681=>"110101100",
  36682=>"011101110",
  36683=>"001011011",
  36684=>"110111001",
  36685=>"111101011",
  36686=>"111110110",
  36687=>"001011010",
  36688=>"111101010",
  36689=>"001101100",
  36690=>"010010110",
  36691=>"101111101",
  36692=>"111110111",
  36693=>"101101101",
  36694=>"001001000",
  36695=>"100111000",
  36696=>"101000000",
  36697=>"111011000",
  36698=>"101010111",
  36699=>"100011110",
  36700=>"010110001",
  36701=>"001100110",
  36702=>"111111111",
  36703=>"011111000",
  36704=>"101011000",
  36705=>"100110001",
  36706=>"000010100",
  36707=>"111101010",
  36708=>"001010000",
  36709=>"111101011",
  36710=>"101111011",
  36711=>"110010111",
  36712=>"000000111",
  36713=>"100010000",
  36714=>"111111011",
  36715=>"010010010",
  36716=>"000100100",
  36717=>"001110111",
  36718=>"110001110",
  36719=>"010000111",
  36720=>"011100000",
  36721=>"111011110",
  36722=>"011110101",
  36723=>"011000011",
  36724=>"101111010",
  36725=>"000110110",
  36726=>"000110011",
  36727=>"110110111",
  36728=>"011000011",
  36729=>"110101000",
  36730=>"110000000",
  36731=>"010101100",
  36732=>"111000101",
  36733=>"110101000",
  36734=>"000110010",
  36735=>"101100111",
  36736=>"010001000",
  36737=>"000111001",
  36738=>"000101101",
  36739=>"100100111",
  36740=>"000011100",
  36741=>"101111110",
  36742=>"110011101",
  36743=>"011101110",
  36744=>"111111010",
  36745=>"001000100",
  36746=>"000000101",
  36747=>"110100001",
  36748=>"001011001",
  36749=>"010100101",
  36750=>"101111101",
  36751=>"010110101",
  36752=>"101111101",
  36753=>"100000010",
  36754=>"111100101",
  36755=>"111000011",
  36756=>"111101111",
  36757=>"010011100",
  36758=>"011110111",
  36759=>"111110001",
  36760=>"000010001",
  36761=>"001100011",
  36762=>"011011100",
  36763=>"111100100",
  36764=>"010100010",
  36765=>"110100001",
  36766=>"010010000",
  36767=>"101100101",
  36768=>"110110000",
  36769=>"000000011",
  36770=>"100110011",
  36771=>"111111110",
  36772=>"010011001",
  36773=>"111110000",
  36774=>"101011011",
  36775=>"100100011",
  36776=>"110110101",
  36777=>"101110100",
  36778=>"101001100",
  36779=>"100111100",
  36780=>"111111011",
  36781=>"111100000",
  36782=>"001111111",
  36783=>"000100101",
  36784=>"000001111",
  36785=>"000011010",
  36786=>"011100010",
  36787=>"001101001",
  36788=>"101111011",
  36789=>"110010010",
  36790=>"011100100",
  36791=>"001010100",
  36792=>"110010010",
  36793=>"100101000",
  36794=>"110000010",
  36795=>"001010110",
  36796=>"100010001",
  36797=>"011001010",
  36798=>"010111010",
  36799=>"101001000",
  36800=>"111000111",
  36801=>"101111001",
  36802=>"110101001",
  36803=>"010101000",
  36804=>"101100011",
  36805=>"011101001",
  36806=>"000001010",
  36807=>"010101101",
  36808=>"100010001",
  36809=>"101110100",
  36810=>"100110011",
  36811=>"110000110",
  36812=>"000001111",
  36813=>"000111011",
  36814=>"111110111",
  36815=>"010001101",
  36816=>"011000011",
  36817=>"010011111",
  36818=>"010110010",
  36819=>"000000100",
  36820=>"011011010",
  36821=>"010111000",
  36822=>"000111010",
  36823=>"000110110",
  36824=>"011100010",
  36825=>"100011001",
  36826=>"000011010",
  36827=>"001011110",
  36828=>"110100001",
  36829=>"000111010",
  36830=>"111100101",
  36831=>"101110110",
  36832=>"101110111",
  36833=>"000100000",
  36834=>"110010100",
  36835=>"101000011",
  36836=>"001111001",
  36837=>"011101110",
  36838=>"000001111",
  36839=>"000111100",
  36840=>"000111010",
  36841=>"111110011",
  36842=>"111011100",
  36843=>"001000111",
  36844=>"000110011",
  36845=>"001011000",
  36846=>"001101110",
  36847=>"100110001",
  36848=>"111001011",
  36849=>"011101110",
  36850=>"100100110",
  36851=>"111100000",
  36852=>"100010010",
  36853=>"000001001",
  36854=>"110010110",
  36855=>"001100101",
  36856=>"111010000",
  36857=>"011111000",
  36858=>"010100010",
  36859=>"001011011",
  36860=>"011001100",
  36861=>"000110110",
  36862=>"010101101",
  36863=>"100010011",
  36864=>"101110000",
  36865=>"101111001",
  36866=>"111110000",
  36867=>"101011010",
  36868=>"110101100",
  36869=>"111000010",
  36870=>"010100111",
  36871=>"111111100",
  36872=>"001110010",
  36873=>"010001100",
  36874=>"110110011",
  36875=>"110100011",
  36876=>"010100000",
  36877=>"000101010",
  36878=>"111011001",
  36879=>"000010111",
  36880=>"100111111",
  36881=>"010100101",
  36882=>"010111001",
  36883=>"101010111",
  36884=>"100001101",
  36885=>"111100110",
  36886=>"001101111",
  36887=>"110010001",
  36888=>"010110111",
  36889=>"100010001",
  36890=>"011100011",
  36891=>"000101001",
  36892=>"010111100",
  36893=>"011000101",
  36894=>"100101100",
  36895=>"101001110",
  36896=>"011000101",
  36897=>"110010011",
  36898=>"110010101",
  36899=>"011100110",
  36900=>"101011100",
  36901=>"000001100",
  36902=>"001101101",
  36903=>"010111110",
  36904=>"010101111",
  36905=>"100000101",
  36906=>"010110011",
  36907=>"101100011",
  36908=>"111101110",
  36909=>"100100100",
  36910=>"101001010",
  36911=>"110011000",
  36912=>"000001110",
  36913=>"000100010",
  36914=>"001011001",
  36915=>"100000010",
  36916=>"000110011",
  36917=>"011011001",
  36918=>"111110101",
  36919=>"000001101",
  36920=>"000100110",
  36921=>"010011111",
  36922=>"000100011",
  36923=>"101100101",
  36924=>"010001011",
  36925=>"011110010",
  36926=>"111000010",
  36927=>"010110110",
  36928=>"101011010",
  36929=>"111100100",
  36930=>"100000100",
  36931=>"001000010",
  36932=>"101111010",
  36933=>"111111010",
  36934=>"011000001",
  36935=>"000100011",
  36936=>"101010001",
  36937=>"010111111",
  36938=>"100011011",
  36939=>"101111000",
  36940=>"001100111",
  36941=>"101100000",
  36942=>"111101101",
  36943=>"001110001",
  36944=>"111100000",
  36945=>"000000010",
  36946=>"101001111",
  36947=>"100001010",
  36948=>"100110100",
  36949=>"100001100",
  36950=>"111000100",
  36951=>"110110111",
  36952=>"001100110",
  36953=>"101001100",
  36954=>"000111101",
  36955=>"100011110",
  36956=>"111110100",
  36957=>"100100000",
  36958=>"010010001",
  36959=>"010011011",
  36960=>"011110011",
  36961=>"011001100",
  36962=>"101111010",
  36963=>"011000000",
  36964=>"001011101",
  36965=>"000101110",
  36966=>"011111010",
  36967=>"100000000",
  36968=>"100110110",
  36969=>"110101111",
  36970=>"000000101",
  36971=>"000011111",
  36972=>"111000000",
  36973=>"011110000",
  36974=>"110000110",
  36975=>"000111100",
  36976=>"100111101",
  36977=>"101010010",
  36978=>"001110110",
  36979=>"100010111",
  36980=>"010110010",
  36981=>"110001010",
  36982=>"010000100",
  36983=>"010000011",
  36984=>"000100111",
  36985=>"111001011",
  36986=>"110010110",
  36987=>"010001100",
  36988=>"011101100",
  36989=>"110101000",
  36990=>"001001010",
  36991=>"110110111",
  36992=>"000001100",
  36993=>"000110101",
  36994=>"101100100",
  36995=>"110101111",
  36996=>"100010011",
  36997=>"010101111",
  36998=>"100000000",
  36999=>"110101101",
  37000=>"010010010",
  37001=>"101111000",
  37002=>"000110011",
  37003=>"101110010",
  37004=>"001010010",
  37005=>"110010110",
  37006=>"111110001",
  37007=>"000001011",
  37008=>"011010010",
  37009=>"010000010",
  37010=>"010001000",
  37011=>"100011001",
  37012=>"011011000",
  37013=>"100101011",
  37014=>"100000000",
  37015=>"011111111",
  37016=>"001100110",
  37017=>"101101101",
  37018=>"011110010",
  37019=>"101010000",
  37020=>"000010000",
  37021=>"100110101",
  37022=>"111110101",
  37023=>"101001011",
  37024=>"000000111",
  37025=>"100110111",
  37026=>"101100000",
  37027=>"001111101",
  37028=>"010010010",
  37029=>"000000001",
  37030=>"011010101",
  37031=>"001001111",
  37032=>"010111100",
  37033=>"001110111",
  37034=>"100110011",
  37035=>"010101011",
  37036=>"011111011",
  37037=>"000000110",
  37038=>"101011001",
  37039=>"011110100",
  37040=>"011100100",
  37041=>"010011000",
  37042=>"111110010",
  37043=>"001001001",
  37044=>"001010010",
  37045=>"001011001",
  37046=>"110001010",
  37047=>"111111000",
  37048=>"100110000",
  37049=>"011001011",
  37050=>"110011111",
  37051=>"001110010",
  37052=>"001100101",
  37053=>"010110011",
  37054=>"101011111",
  37055=>"000111011",
  37056=>"000100001",
  37057=>"001011100",
  37058=>"101001100",
  37059=>"000000011",
  37060=>"011001101",
  37061=>"100010000",
  37062=>"110011000",
  37063=>"001011101",
  37064=>"110110110",
  37065=>"110101111",
  37066=>"011100101",
  37067=>"101111110",
  37068=>"111101110",
  37069=>"101011011",
  37070=>"100010010",
  37071=>"101000000",
  37072=>"100010000",
  37073=>"100100100",
  37074=>"111110110",
  37075=>"110010010",
  37076=>"100001010",
  37077=>"101100001",
  37078=>"101101110",
  37079=>"110010101",
  37080=>"100111000",
  37081=>"100111011",
  37082=>"100000101",
  37083=>"110000010",
  37084=>"101001110",
  37085=>"000001001",
  37086=>"011010111",
  37087=>"001000100",
  37088=>"011110011",
  37089=>"101011110",
  37090=>"010010110",
  37091=>"100000101",
  37092=>"001110101",
  37093=>"011100100",
  37094=>"001000101",
  37095=>"101101101",
  37096=>"111001011",
  37097=>"000011001",
  37098=>"111010100",
  37099=>"100110100",
  37100=>"001010100",
  37101=>"000111111",
  37102=>"110001111",
  37103=>"000010000",
  37104=>"110110110",
  37105=>"100111100",
  37106=>"110011000",
  37107=>"110100001",
  37108=>"000011110",
  37109=>"000000100",
  37110=>"010010100",
  37111=>"101111001",
  37112=>"110111110",
  37113=>"001010110",
  37114=>"111010000",
  37115=>"111101011",
  37116=>"001010111",
  37117=>"001000101",
  37118=>"000101000",
  37119=>"101110011",
  37120=>"011011111",
  37121=>"010001010",
  37122=>"010000011",
  37123=>"001011111",
  37124=>"100110111",
  37125=>"100110111",
  37126=>"001001000",
  37127=>"101010101",
  37128=>"111101010",
  37129=>"010010111",
  37130=>"000111110",
  37131=>"100010000",
  37132=>"000010101",
  37133=>"001011000",
  37134=>"100101000",
  37135=>"000011000",
  37136=>"001000001",
  37137=>"011100000",
  37138=>"000111101",
  37139=>"110110111",
  37140=>"110000101",
  37141=>"010011101",
  37142=>"100010000",
  37143=>"100100010",
  37144=>"110011101",
  37145=>"011011001",
  37146=>"110111101",
  37147=>"101110111",
  37148=>"001101000",
  37149=>"010100001",
  37150=>"111010101",
  37151=>"100011000",
  37152=>"001101010",
  37153=>"010100001",
  37154=>"110111001",
  37155=>"110010000",
  37156=>"011010000",
  37157=>"010110111",
  37158=>"100001101",
  37159=>"011010011",
  37160=>"000011110",
  37161=>"100000110",
  37162=>"111100000",
  37163=>"110010101",
  37164=>"011010001",
  37165=>"100111011",
  37166=>"000110001",
  37167=>"010000011",
  37168=>"100010110",
  37169=>"010010110",
  37170=>"100101111",
  37171=>"010000000",
  37172=>"011101000",
  37173=>"001011111",
  37174=>"101101100",
  37175=>"110101100",
  37176=>"001101101",
  37177=>"010101110",
  37178=>"000100011",
  37179=>"001010011",
  37180=>"001100001",
  37181=>"111110000",
  37182=>"110100000",
  37183=>"010011011",
  37184=>"111111010",
  37185=>"000101101",
  37186=>"011000110",
  37187=>"010110101",
  37188=>"000111101",
  37189=>"100100010",
  37190=>"010111111",
  37191=>"001110011",
  37192=>"000101010",
  37193=>"010101101",
  37194=>"101000000",
  37195=>"011010110",
  37196=>"010111100",
  37197=>"001111001",
  37198=>"000111000",
  37199=>"111000010",
  37200=>"101011111",
  37201=>"111111111",
  37202=>"001010011",
  37203=>"100101000",
  37204=>"101011101",
  37205=>"111010000",
  37206=>"110000110",
  37207=>"001111001",
  37208=>"000011101",
  37209=>"011101110",
  37210=>"000010100",
  37211=>"110110110",
  37212=>"110101110",
  37213=>"000101110",
  37214=>"011011010",
  37215=>"001001111",
  37216=>"100101001",
  37217=>"101100001",
  37218=>"100110101",
  37219=>"010000101",
  37220=>"010010100",
  37221=>"100001111",
  37222=>"011011001",
  37223=>"111101101",
  37224=>"001100011",
  37225=>"010111111",
  37226=>"001111111",
  37227=>"000110000",
  37228=>"011010111",
  37229=>"101111111",
  37230=>"000011011",
  37231=>"110111111",
  37232=>"000110010",
  37233=>"111010001",
  37234=>"011100001",
  37235=>"000101001",
  37236=>"100101111",
  37237=>"010011111",
  37238=>"100100101",
  37239=>"100011110",
  37240=>"000010010",
  37241=>"110110111",
  37242=>"010001111",
  37243=>"101111011",
  37244=>"100110001",
  37245=>"011111001",
  37246=>"111001001",
  37247=>"000111011",
  37248=>"010000111",
  37249=>"000011000",
  37250=>"000100010",
  37251=>"110001101",
  37252=>"101100010",
  37253=>"110111001",
  37254=>"011111101",
  37255=>"110110110",
  37256=>"110100111",
  37257=>"111000000",
  37258=>"110100000",
  37259=>"011100010",
  37260=>"011101011",
  37261=>"110101000",
  37262=>"111110000",
  37263=>"111010010",
  37264=>"100111110",
  37265=>"101010100",
  37266=>"011100001",
  37267=>"000100110",
  37268=>"110100101",
  37269=>"100001110",
  37270=>"100001100",
  37271=>"010111111",
  37272=>"100100111",
  37273=>"100100010",
  37274=>"011011001",
  37275=>"111110001",
  37276=>"100001111",
  37277=>"011110000",
  37278=>"000100000",
  37279=>"111100110",
  37280=>"101101011",
  37281=>"011010010",
  37282=>"001100010",
  37283=>"001000000",
  37284=>"111101001",
  37285=>"000101111",
  37286=>"101100111",
  37287=>"100000011",
  37288=>"111011100",
  37289=>"010010111",
  37290=>"001001101",
  37291=>"001000001",
  37292=>"000010100",
  37293=>"111100010",
  37294=>"110111011",
  37295=>"001000001",
  37296=>"100100110",
  37297=>"101000000",
  37298=>"000010110",
  37299=>"100101110",
  37300=>"110010010",
  37301=>"100101011",
  37302=>"101111110",
  37303=>"110111010",
  37304=>"110111000",
  37305=>"000011111",
  37306=>"100100101",
  37307=>"101110011",
  37308=>"100110010",
  37309=>"001110010",
  37310=>"111111000",
  37311=>"100010011",
  37312=>"110011000",
  37313=>"010111000",
  37314=>"101011111",
  37315=>"101101100",
  37316=>"001011000",
  37317=>"010111110",
  37318=>"110100110",
  37319=>"111101000",
  37320=>"111000111",
  37321=>"111000001",
  37322=>"100000101",
  37323=>"100010001",
  37324=>"100011011",
  37325=>"100110001",
  37326=>"101110001",
  37327=>"000110101",
  37328=>"111101010",
  37329=>"011011000",
  37330=>"000001001",
  37331=>"111000110",
  37332=>"001011111",
  37333=>"011101001",
  37334=>"111011100",
  37335=>"001011011",
  37336=>"000110110",
  37337=>"001011011",
  37338=>"110110100",
  37339=>"111011110",
  37340=>"101001011",
  37341=>"001010010",
  37342=>"010110111",
  37343=>"101001100",
  37344=>"110000100",
  37345=>"010011100",
  37346=>"110110010",
  37347=>"111011101",
  37348=>"100001010",
  37349=>"001101110",
  37350=>"110010001",
  37351=>"110000001",
  37352=>"110001011",
  37353=>"101001011",
  37354=>"111010101",
  37355=>"110111010",
  37356=>"111111010",
  37357=>"001101010",
  37358=>"111100111",
  37359=>"110100001",
  37360=>"001001000",
  37361=>"010110001",
  37362=>"110000111",
  37363=>"000000100",
  37364=>"011111110",
  37365=>"010111011",
  37366=>"001011010",
  37367=>"111000110",
  37368=>"101011000",
  37369=>"000011010",
  37370=>"000011011",
  37371=>"111000111",
  37372=>"100010010",
  37373=>"101101100",
  37374=>"000000000",
  37375=>"000001001",
  37376=>"101111111",
  37377=>"010101010",
  37378=>"000111001",
  37379=>"010100000",
  37380=>"011000000",
  37381=>"001011010",
  37382=>"001000010",
  37383=>"110110111",
  37384=>"011011011",
  37385=>"100001010",
  37386=>"001011110",
  37387=>"110011101",
  37388=>"101100010",
  37389=>"001000010",
  37390=>"000101010",
  37391=>"110011010",
  37392=>"111101100",
  37393=>"111010001",
  37394=>"101010100",
  37395=>"011010001",
  37396=>"011111010",
  37397=>"000010100",
  37398=>"111110001",
  37399=>"001111110",
  37400=>"101111011",
  37401=>"110111001",
  37402=>"111000011",
  37403=>"001111010",
  37404=>"001011011",
  37405=>"100110000",
  37406=>"101010101",
  37407=>"011101101",
  37408=>"001101001",
  37409=>"111011001",
  37410=>"011001111",
  37411=>"101100001",
  37412=>"011100100",
  37413=>"000010010",
  37414=>"110001011",
  37415=>"000001101",
  37416=>"010111111",
  37417=>"010101011",
  37418=>"111000000",
  37419=>"101100011",
  37420=>"011000111",
  37421=>"010000110",
  37422=>"100000001",
  37423=>"100100111",
  37424=>"011110011",
  37425=>"011001110",
  37426=>"110000011",
  37427=>"011100001",
  37428=>"101110011",
  37429=>"000000010",
  37430=>"011001110",
  37431=>"000001110",
  37432=>"000101011",
  37433=>"111110110",
  37434=>"111111001",
  37435=>"100101011",
  37436=>"001010111",
  37437=>"000100010",
  37438=>"010110010",
  37439=>"111101111",
  37440=>"100110010",
  37441=>"010110111",
  37442=>"000111011",
  37443=>"101001010",
  37444=>"100111011",
  37445=>"001111011",
  37446=>"111111010",
  37447=>"110000100",
  37448=>"111010010",
  37449=>"111101001",
  37450=>"000000011",
  37451=>"100011000",
  37452=>"100101110",
  37453=>"110000001",
  37454=>"110111110",
  37455=>"111001000",
  37456=>"001111111",
  37457=>"100000111",
  37458=>"111100101",
  37459=>"110110101",
  37460=>"001010100",
  37461=>"101110010",
  37462=>"001000010",
  37463=>"100011001",
  37464=>"110001110",
  37465=>"111000110",
  37466=>"100010100",
  37467=>"000111100",
  37468=>"001011010",
  37469=>"101000001",
  37470=>"101111100",
  37471=>"111101111",
  37472=>"011001000",
  37473=>"011001110",
  37474=>"011101111",
  37475=>"001100010",
  37476=>"011111011",
  37477=>"101110111",
  37478=>"000100101",
  37479=>"101010100",
  37480=>"010101111",
  37481=>"110011001",
  37482=>"101110011",
  37483=>"010111111",
  37484=>"101000101",
  37485=>"011011100",
  37486=>"010111011",
  37487=>"110110110",
  37488=>"011001000",
  37489=>"101000000",
  37490=>"101101010",
  37491=>"010011010",
  37492=>"100000001",
  37493=>"001100100",
  37494=>"000011101",
  37495=>"000000000",
  37496=>"111101101",
  37497=>"111100011",
  37498=>"101110110",
  37499=>"000101010",
  37500=>"000000111",
  37501=>"101001010",
  37502=>"100010000",
  37503=>"010001101",
  37504=>"011010000",
  37505=>"011110011",
  37506=>"111011101",
  37507=>"001011000",
  37508=>"001001011",
  37509=>"000010111",
  37510=>"000111100",
  37511=>"111111101",
  37512=>"001111101",
  37513=>"110101001",
  37514=>"100011101",
  37515=>"000111000",
  37516=>"001000110",
  37517=>"111111111",
  37518=>"111001000",
  37519=>"011111110",
  37520=>"010100011",
  37521=>"110111001",
  37522=>"110111100",
  37523=>"000101100",
  37524=>"100000010",
  37525=>"000010011",
  37526=>"100010000",
  37527=>"010011010",
  37528=>"101111011",
  37529=>"010011110",
  37530=>"011011100",
  37531=>"000001011",
  37532=>"000110010",
  37533=>"111011001",
  37534=>"111100100",
  37535=>"110010100",
  37536=>"110101110",
  37537=>"101010101",
  37538=>"001001010",
  37539=>"101100101",
  37540=>"101111011",
  37541=>"110010001",
  37542=>"110011100",
  37543=>"000111010",
  37544=>"000101101",
  37545=>"011101000",
  37546=>"100001011",
  37547=>"000111111",
  37548=>"101111010",
  37549=>"011010111",
  37550=>"110111101",
  37551=>"000110100",
  37552=>"001101000",
  37553=>"111000111",
  37554=>"011000100",
  37555=>"011001111",
  37556=>"001011011",
  37557=>"111011001",
  37558=>"011111111",
  37559=>"111001111",
  37560=>"100110100",
  37561=>"000111100",
  37562=>"000011110",
  37563=>"111011100",
  37564=>"100011001",
  37565=>"000101000",
  37566=>"000001100",
  37567=>"001100000",
  37568=>"011111101",
  37569=>"000101111",
  37570=>"000011101",
  37571=>"010011010",
  37572=>"101110001",
  37573=>"100111010",
  37574=>"010101000",
  37575=>"111000110",
  37576=>"011010111",
  37577=>"101001001",
  37578=>"100001001",
  37579=>"011101001",
  37580=>"101011000",
  37581=>"101110100",
  37582=>"100110000",
  37583=>"101010000",
  37584=>"000000000",
  37585=>"000011000",
  37586=>"101101110",
  37587=>"010011000",
  37588=>"111111000",
  37589=>"100001101",
  37590=>"011100000",
  37591=>"111000110",
  37592=>"000111011",
  37593=>"111111011",
  37594=>"110011111",
  37595=>"010001011",
  37596=>"001110101",
  37597=>"111010011",
  37598=>"111000101",
  37599=>"000101000",
  37600=>"110101001",
  37601=>"011100110",
  37602=>"000110010",
  37603=>"001110101",
  37604=>"000001100",
  37605=>"011110111",
  37606=>"101000000",
  37607=>"001000011",
  37608=>"001011101",
  37609=>"110111111",
  37610=>"110111101",
  37611=>"100001000",
  37612=>"000010101",
  37613=>"001110100",
  37614=>"110001111",
  37615=>"000001101",
  37616=>"110010001",
  37617=>"000110101",
  37618=>"111011101",
  37619=>"010001011",
  37620=>"110110110",
  37621=>"100110101",
  37622=>"101000111",
  37623=>"110011101",
  37624=>"010011111",
  37625=>"110100001",
  37626=>"110100011",
  37627=>"001111011",
  37628=>"000101001",
  37629=>"010110011",
  37630=>"011110100",
  37631=>"010010010",
  37632=>"010001001",
  37633=>"100111000",
  37634=>"011101100",
  37635=>"010000001",
  37636=>"011110000",
  37637=>"001011010",
  37638=>"001110011",
  37639=>"111010110",
  37640=>"010111100",
  37641=>"011100010",
  37642=>"110000000",
  37643=>"101101011",
  37644=>"100110100",
  37645=>"011111100",
  37646=>"100100101",
  37647=>"101011011",
  37648=>"111111100",
  37649=>"010010101",
  37650=>"001111011",
  37651=>"000111101",
  37652=>"001001010",
  37653=>"011011111",
  37654=>"110000011",
  37655=>"000100111",
  37656=>"101100101",
  37657=>"110000001",
  37658=>"010111110",
  37659=>"001011111",
  37660=>"100001101",
  37661=>"000111101",
  37662=>"101011111",
  37663=>"101011100",
  37664=>"000011110",
  37665=>"011011110",
  37666=>"110100010",
  37667=>"001011010",
  37668=>"100110111",
  37669=>"111000010",
  37670=>"100100101",
  37671=>"011101100",
  37672=>"101110011",
  37673=>"111001000",
  37674=>"111101011",
  37675=>"010010001",
  37676=>"011001100",
  37677=>"011110001",
  37678=>"111110011",
  37679=>"110001001",
  37680=>"110101001",
  37681=>"111101000",
  37682=>"100110100",
  37683=>"001010011",
  37684=>"010111001",
  37685=>"010111110",
  37686=>"000011110",
  37687=>"101001011",
  37688=>"000010000",
  37689=>"111111011",
  37690=>"111011011",
  37691=>"001110011",
  37692=>"011110011",
  37693=>"010100011",
  37694=>"111010011",
  37695=>"011001110",
  37696=>"101000100",
  37697=>"001001011",
  37698=>"010010110",
  37699=>"010000100",
  37700=>"001001110",
  37701=>"110101001",
  37702=>"011110101",
  37703=>"011001111",
  37704=>"110111011",
  37705=>"110101111",
  37706=>"011101000",
  37707=>"010111111",
  37708=>"111011101",
  37709=>"101000010",
  37710=>"001000100",
  37711=>"011000110",
  37712=>"101011001",
  37713=>"011111010",
  37714=>"111000101",
  37715=>"000010110",
  37716=>"110111111",
  37717=>"000101000",
  37718=>"000110100",
  37719=>"010001000",
  37720=>"011111001",
  37721=>"010010100",
  37722=>"000010011",
  37723=>"001110110",
  37724=>"001000110",
  37725=>"100101010",
  37726=>"010111101",
  37727=>"100000101",
  37728=>"010011110",
  37729=>"111011101",
  37730=>"010010001",
  37731=>"000101011",
  37732=>"100101000",
  37733=>"001101101",
  37734=>"111101110",
  37735=>"011010011",
  37736=>"000100010",
  37737=>"011111101",
  37738=>"101111110",
  37739=>"000100110",
  37740=>"101000100",
  37741=>"110100101",
  37742=>"001000111",
  37743=>"100111011",
  37744=>"111111110",
  37745=>"001001011",
  37746=>"000101110",
  37747=>"110000011",
  37748=>"010100001",
  37749=>"000000101",
  37750=>"000000111",
  37751=>"101101011",
  37752=>"110111111",
  37753=>"010010001",
  37754=>"101101110",
  37755=>"001001000",
  37756=>"000011010",
  37757=>"101001111",
  37758=>"001000000",
  37759=>"111000011",
  37760=>"101011011",
  37761=>"000011101",
  37762=>"000001000",
  37763=>"101101000",
  37764=>"110111010",
  37765=>"010010000",
  37766=>"001010100",
  37767=>"101000110",
  37768=>"111111011",
  37769=>"111010010",
  37770=>"010000011",
  37771=>"000010000",
  37772=>"010111101",
  37773=>"111110101",
  37774=>"001010100",
  37775=>"101111100",
  37776=>"111000110",
  37777=>"001011101",
  37778=>"011010000",
  37779=>"001010001",
  37780=>"001001101",
  37781=>"101011001",
  37782=>"010011101",
  37783=>"001111010",
  37784=>"110001010",
  37785=>"110101101",
  37786=>"101000001",
  37787=>"111110011",
  37788=>"100100010",
  37789=>"011101100",
  37790=>"000000101",
  37791=>"001001001",
  37792=>"111010011",
  37793=>"111010110",
  37794=>"111010110",
  37795=>"111000011",
  37796=>"000010101",
  37797=>"001101010",
  37798=>"000110001",
  37799=>"000000100",
  37800=>"111101110",
  37801=>"111011101",
  37802=>"101000101",
  37803=>"011011101",
  37804=>"110111011",
  37805=>"111011001",
  37806=>"111111000",
  37807=>"111100100",
  37808=>"000001011",
  37809=>"101110010",
  37810=>"110010001",
  37811=>"101110100",
  37812=>"101011101",
  37813=>"001000111",
  37814=>"010000110",
  37815=>"100010000",
  37816=>"010001110",
  37817=>"111110010",
  37818=>"010110100",
  37819=>"001001101",
  37820=>"100010110",
  37821=>"010101111",
  37822=>"011110000",
  37823=>"101001101",
  37824=>"010000010",
  37825=>"000011000",
  37826=>"011110100",
  37827=>"001001111",
  37828=>"100011010",
  37829=>"110001011",
  37830=>"000110011",
  37831=>"100001100",
  37832=>"001111101",
  37833=>"101001110",
  37834=>"011010110",
  37835=>"010011011",
  37836=>"010101001",
  37837=>"000000000",
  37838=>"000001111",
  37839=>"010100111",
  37840=>"000010111",
  37841=>"000100111",
  37842=>"011001001",
  37843=>"101010011",
  37844=>"011011000",
  37845=>"100111010",
  37846=>"100101001",
  37847=>"000001101",
  37848=>"000101100",
  37849=>"100101011",
  37850=>"111000101",
  37851=>"101110111",
  37852=>"111101000",
  37853=>"101001000",
  37854=>"101001111",
  37855=>"000111011",
  37856=>"010010010",
  37857=>"101000100",
  37858=>"001000010",
  37859=>"101101101",
  37860=>"000001001",
  37861=>"000010111",
  37862=>"000010010",
  37863=>"011110011",
  37864=>"101100100",
  37865=>"001110010",
  37866=>"111100010",
  37867=>"010110100",
  37868=>"001000001",
  37869=>"000000010",
  37870=>"100111110",
  37871=>"110101101",
  37872=>"100000101",
  37873=>"001110110",
  37874=>"001111111",
  37875=>"010010000",
  37876=>"100101001",
  37877=>"110111101",
  37878=>"111110101",
  37879=>"101110010",
  37880=>"000001110",
  37881=>"010110100",
  37882=>"100111111",
  37883=>"100010110",
  37884=>"000010101",
  37885=>"001001111",
  37886=>"011100101",
  37887=>"000011110",
  37888=>"111111101",
  37889=>"011000110",
  37890=>"010110011",
  37891=>"100000110",
  37892=>"100111010",
  37893=>"111011001",
  37894=>"010000101",
  37895=>"000001010",
  37896=>"001011010",
  37897=>"101110111",
  37898=>"010101001",
  37899=>"010011000",
  37900=>"100100001",
  37901=>"111100100",
  37902=>"011011111",
  37903=>"111010010",
  37904=>"111010001",
  37905=>"011000001",
  37906=>"011111011",
  37907=>"111001010",
  37908=>"110000000",
  37909=>"001011010",
  37910=>"100000001",
  37911=>"000101010",
  37912=>"100111001",
  37913=>"001000110",
  37914=>"110011001",
  37915=>"001000111",
  37916=>"100100000",
  37917=>"100111011",
  37918=>"101100010",
  37919=>"010000000",
  37920=>"111000001",
  37921=>"101010011",
  37922=>"010110111",
  37923=>"001011011",
  37924=>"001010001",
  37925=>"011100010",
  37926=>"110110101",
  37927=>"011111101",
  37928=>"100101001",
  37929=>"111111111",
  37930=>"110111111",
  37931=>"101001000",
  37932=>"011100111",
  37933=>"101000011",
  37934=>"110000001",
  37935=>"011111011",
  37936=>"111000000",
  37937=>"110001101",
  37938=>"000111101",
  37939=>"110000000",
  37940=>"010001100",
  37941=>"010011010",
  37942=>"011010110",
  37943=>"101101010",
  37944=>"000010000",
  37945=>"000111000",
  37946=>"111111111",
  37947=>"011110101",
  37948=>"011001001",
  37949=>"011110111",
  37950=>"001000010",
  37951=>"000010010",
  37952=>"100000011",
  37953=>"111100000",
  37954=>"011010110",
  37955=>"111011110",
  37956=>"101110101",
  37957=>"100011000",
  37958=>"010110111",
  37959=>"000000000",
  37960=>"111010001",
  37961=>"000001110",
  37962=>"101110100",
  37963=>"000100110",
  37964=>"100100111",
  37965=>"000111000",
  37966=>"100111011",
  37967=>"101111101",
  37968=>"010101110",
  37969=>"001001010",
  37970=>"110100000",
  37971=>"000000001",
  37972=>"011000110",
  37973=>"111011000",
  37974=>"100101010",
  37975=>"010010000",
  37976=>"101111000",
  37977=>"000110011",
  37978=>"000011011",
  37979=>"010000001",
  37980=>"010001101",
  37981=>"000100100",
  37982=>"110100100",
  37983=>"011011010",
  37984=>"100101000",
  37985=>"011111001",
  37986=>"000100110",
  37987=>"000011010",
  37988=>"110010001",
  37989=>"000010000",
  37990=>"101111000",
  37991=>"011010110",
  37992=>"100101100",
  37993=>"111011101",
  37994=>"000101110",
  37995=>"100101001",
  37996=>"100000101",
  37997=>"001110001",
  37998=>"111110010",
  37999=>"111011111",
  38000=>"000110111",
  38001=>"010111011",
  38002=>"010110100",
  38003=>"110001011",
  38004=>"110110111",
  38005=>"101010101",
  38006=>"011011101",
  38007=>"011111000",
  38008=>"110100010",
  38009=>"001011100",
  38010=>"111011000",
  38011=>"111000011",
  38012=>"010101101",
  38013=>"001100100",
  38014=>"000010100",
  38015=>"101011111",
  38016=>"100010011",
  38017=>"001100010",
  38018=>"000100110",
  38019=>"011010001",
  38020=>"001011000",
  38021=>"011010000",
  38022=>"010001001",
  38023=>"001010101",
  38024=>"110111101",
  38025=>"110010000",
  38026=>"001001101",
  38027=>"101110010",
  38028=>"001001010",
  38029=>"001101000",
  38030=>"000001000",
  38031=>"000101001",
  38032=>"010001000",
  38033=>"011010100",
  38034=>"000101100",
  38035=>"011111111",
  38036=>"111110111",
  38037=>"000111010",
  38038=>"100010000",
  38039=>"001011010",
  38040=>"010001011",
  38041=>"010001000",
  38042=>"111111001",
  38043=>"100110010",
  38044=>"101111110",
  38045=>"001110010",
  38046=>"000010010",
  38047=>"110111111",
  38048=>"000000100",
  38049=>"011011001",
  38050=>"111100010",
  38051=>"101011010",
  38052=>"110010110",
  38053=>"100111010",
  38054=>"001100000",
  38055=>"011011110",
  38056=>"110110000",
  38057=>"010010010",
  38058=>"001101010",
  38059=>"001001100",
  38060=>"011010110",
  38061=>"111101010",
  38062=>"101101100",
  38063=>"101000111",
  38064=>"001000000",
  38065=>"000000000",
  38066=>"100110010",
  38067=>"000001111",
  38068=>"011110101",
  38069=>"010000000",
  38070=>"110001110",
  38071=>"010010110",
  38072=>"000001010",
  38073=>"001100011",
  38074=>"101000110",
  38075=>"101111110",
  38076=>"100011011",
  38077=>"010110010",
  38078=>"101010100",
  38079=>"100011010",
  38080=>"110010011",
  38081=>"001111111",
  38082=>"011001001",
  38083=>"111001010",
  38084=>"111001011",
  38085=>"111010001",
  38086=>"000001101",
  38087=>"000111000",
  38088=>"110001010",
  38089=>"101001100",
  38090=>"111011110",
  38091=>"001111111",
  38092=>"001111001",
  38093=>"010001001",
  38094=>"110110001",
  38095=>"011001101",
  38096=>"101100010",
  38097=>"111111100",
  38098=>"000101111",
  38099=>"111000111",
  38100=>"110011001",
  38101=>"001100000",
  38102=>"011000100",
  38103=>"010110111",
  38104=>"100000000",
  38105=>"010010111",
  38106=>"010010100",
  38107=>"100100111",
  38108=>"011010010",
  38109=>"011111000",
  38110=>"011010100",
  38111=>"111110000",
  38112=>"101001011",
  38113=>"101001000",
  38114=>"001010000",
  38115=>"010000011",
  38116=>"011110010",
  38117=>"010000010",
  38118=>"001101000",
  38119=>"110110001",
  38120=>"010110100",
  38121=>"101011110",
  38122=>"010111010",
  38123=>"001110000",
  38124=>"100101101",
  38125=>"000010010",
  38126=>"110001100",
  38127=>"100111011",
  38128=>"100101110",
  38129=>"110110011",
  38130=>"001001011",
  38131=>"110110001",
  38132=>"100100101",
  38133=>"001101110",
  38134=>"111011111",
  38135=>"100111111",
  38136=>"101101101",
  38137=>"010100111",
  38138=>"101001101",
  38139=>"010111010",
  38140=>"001111110",
  38141=>"101110001",
  38142=>"001011001",
  38143=>"100111111",
  38144=>"010011001",
  38145=>"010000101",
  38146=>"010110111",
  38147=>"111010101",
  38148=>"000010010",
  38149=>"100001111",
  38150=>"010100011",
  38151=>"000000101",
  38152=>"110110101",
  38153=>"101111101",
  38154=>"001110100",
  38155=>"101001100",
  38156=>"011111100",
  38157=>"110101101",
  38158=>"011111000",
  38159=>"000001011",
  38160=>"001000101",
  38161=>"111011110",
  38162=>"011011001",
  38163=>"111011100",
  38164=>"000110100",
  38165=>"001000110",
  38166=>"001000011",
  38167=>"000000100",
  38168=>"111001110",
  38169=>"010100101",
  38170=>"100110101",
  38171=>"010010110",
  38172=>"111011001",
  38173=>"011010010",
  38174=>"100100110",
  38175=>"000001110",
  38176=>"100110000",
  38177=>"101100001",
  38178=>"010101100",
  38179=>"111010100",
  38180=>"010000001",
  38181=>"101101011",
  38182=>"010001100",
  38183=>"010001010",
  38184=>"101110010",
  38185=>"010011000",
  38186=>"101000110",
  38187=>"110110000",
  38188=>"111001000",
  38189=>"000000011",
  38190=>"100010011",
  38191=>"100110110",
  38192=>"001101000",
  38193=>"111101111",
  38194=>"010011111",
  38195=>"100011111",
  38196=>"001010011",
  38197=>"011010101",
  38198=>"000110110",
  38199=>"001111100",
  38200=>"010001100",
  38201=>"010000000",
  38202=>"001110000",
  38203=>"100000110",
  38204=>"101001001",
  38205=>"111101111",
  38206=>"001100110",
  38207=>"011000101",
  38208=>"010000001",
  38209=>"010101101",
  38210=>"101100110",
  38211=>"010011000",
  38212=>"100000100",
  38213=>"111111011",
  38214=>"000110011",
  38215=>"000001110",
  38216=>"011111000",
  38217=>"011000101",
  38218=>"101100111",
  38219=>"111010001",
  38220=>"110001100",
  38221=>"010011101",
  38222=>"001110000",
  38223=>"001011001",
  38224=>"101001111",
  38225=>"000010111",
  38226=>"010100010",
  38227=>"100000011",
  38228=>"000000000",
  38229=>"101111101",
  38230=>"000001010",
  38231=>"111110001",
  38232=>"110110110",
  38233=>"000110110",
  38234=>"000101011",
  38235=>"011110111",
  38236=>"001101010",
  38237=>"010101111",
  38238=>"110000111",
  38239=>"010001111",
  38240=>"101001001",
  38241=>"000110000",
  38242=>"010001101",
  38243=>"000000001",
  38244=>"100110110",
  38245=>"010010001",
  38246=>"011000110",
  38247=>"101111111",
  38248=>"010011110",
  38249=>"000110001",
  38250=>"010110010",
  38251=>"011111110",
  38252=>"000110000",
  38253=>"111000111",
  38254=>"110000011",
  38255=>"111110111",
  38256=>"010100111",
  38257=>"100000100",
  38258=>"011010111",
  38259=>"100110001",
  38260=>"111111100",
  38261=>"111100101",
  38262=>"110110010",
  38263=>"100000100",
  38264=>"110110110",
  38265=>"100100110",
  38266=>"000000111",
  38267=>"011011100",
  38268=>"111010100",
  38269=>"000100111",
  38270=>"000110001",
  38271=>"011001110",
  38272=>"101010000",
  38273=>"001100000",
  38274=>"110011100",
  38275=>"100001001",
  38276=>"011010010",
  38277=>"101011011",
  38278=>"011111111",
  38279=>"101000100",
  38280=>"101010011",
  38281=>"011001110",
  38282=>"011101000",
  38283=>"010111010",
  38284=>"100110110",
  38285=>"001001001",
  38286=>"101110101",
  38287=>"011111100",
  38288=>"111000010",
  38289=>"101111000",
  38290=>"011100011",
  38291=>"011011011",
  38292=>"011000010",
  38293=>"001100000",
  38294=>"111010101",
  38295=>"101100011",
  38296=>"111111000",
  38297=>"011111111",
  38298=>"111111001",
  38299=>"111100111",
  38300=>"101101111",
  38301=>"011111111",
  38302=>"011010101",
  38303=>"111101101",
  38304=>"011011101",
  38305=>"100010101",
  38306=>"010110111",
  38307=>"001010111",
  38308=>"111001000",
  38309=>"101101000",
  38310=>"010110101",
  38311=>"101011100",
  38312=>"000100011",
  38313=>"101001001",
  38314=>"111101010",
  38315=>"000011110",
  38316=>"011111101",
  38317=>"011010101",
  38318=>"001100111",
  38319=>"100100100",
  38320=>"100011010",
  38321=>"100111010",
  38322=>"001000101",
  38323=>"111010011",
  38324=>"011001010",
  38325=>"101010011",
  38326=>"001101101",
  38327=>"111111100",
  38328=>"000000000",
  38329=>"000011001",
  38330=>"000000000",
  38331=>"011000000",
  38332=>"111000010",
  38333=>"100101100",
  38334=>"101110110",
  38335=>"111110111",
  38336=>"011011101",
  38337=>"110100011",
  38338=>"000110010",
  38339=>"111011001",
  38340=>"000000111",
  38341=>"011110000",
  38342=>"111101111",
  38343=>"111001000",
  38344=>"010001101",
  38345=>"100101110",
  38346=>"011010111",
  38347=>"111011011",
  38348=>"011100100",
  38349=>"100110101",
  38350=>"011011100",
  38351=>"100101100",
  38352=>"001101101",
  38353=>"011011011",
  38354=>"110010001",
  38355=>"000100010",
  38356=>"011000100",
  38357=>"000000100",
  38358=>"111011000",
  38359=>"111011011",
  38360=>"111001011",
  38361=>"100111001",
  38362=>"010001011",
  38363=>"101010001",
  38364=>"010001001",
  38365=>"001010011",
  38366=>"011001111",
  38367=>"011010111",
  38368=>"000001000",
  38369=>"010011110",
  38370=>"110110000",
  38371=>"111010011",
  38372=>"000001101",
  38373=>"001111000",
  38374=>"011000000",
  38375=>"111001000",
  38376=>"110101000",
  38377=>"101010001",
  38378=>"000010100",
  38379=>"111100011",
  38380=>"001000000",
  38381=>"000000000",
  38382=>"000010100",
  38383=>"010101111",
  38384=>"010000000",
  38385=>"000110000",
  38386=>"001100001",
  38387=>"000000001",
  38388=>"101000000",
  38389=>"101111000",
  38390=>"111101001",
  38391=>"111000011",
  38392=>"111010000",
  38393=>"110010100",
  38394=>"101000001",
  38395=>"000101100",
  38396=>"011011111",
  38397=>"101010001",
  38398=>"001000010",
  38399=>"010110111",
  38400=>"011101001",
  38401=>"111001110",
  38402=>"000001001",
  38403=>"100100000",
  38404=>"111000111",
  38405=>"100000010",
  38406=>"001101010",
  38407=>"000111010",
  38408=>"011110010",
  38409=>"101100010",
  38410=>"000101100",
  38411=>"000110000",
  38412=>"000100111",
  38413=>"001001011",
  38414=>"011100001",
  38415=>"111000000",
  38416=>"100000111",
  38417=>"001010011",
  38418=>"010101010",
  38419=>"111010010",
  38420=>"010010100",
  38421=>"001001010",
  38422=>"001101000",
  38423=>"001110110",
  38424=>"000010010",
  38425=>"110101111",
  38426=>"011001010",
  38427=>"110010100",
  38428=>"001111011",
  38429=>"000010101",
  38430=>"111110000",
  38431=>"010101111",
  38432=>"111001011",
  38433=>"000001110",
  38434=>"001011001",
  38435=>"000110000",
  38436=>"000110110",
  38437=>"110010000",
  38438=>"111011100",
  38439=>"011010110",
  38440=>"001001101",
  38441=>"011000110",
  38442=>"111010000",
  38443=>"011010010",
  38444=>"001110001",
  38445=>"101110100",
  38446=>"101010100",
  38447=>"001000101",
  38448=>"011101001",
  38449=>"111110011",
  38450=>"011010001",
  38451=>"010001010",
  38452=>"100011000",
  38453=>"111110010",
  38454=>"100110100",
  38455=>"000010111",
  38456=>"100011101",
  38457=>"100011001",
  38458=>"011101011",
  38459=>"010000010",
  38460=>"000101001",
  38461=>"011111100",
  38462=>"000101110",
  38463=>"111110011",
  38464=>"011011111",
  38465=>"110100001",
  38466=>"100000001",
  38467=>"001111110",
  38468=>"011001101",
  38469=>"011010110",
  38470=>"000011111",
  38471=>"011100001",
  38472=>"010001100",
  38473=>"011000000",
  38474=>"000111010",
  38475=>"101100001",
  38476=>"001100101",
  38477=>"100001000",
  38478=>"010010011",
  38479=>"000110001",
  38480=>"111100111",
  38481=>"011111000",
  38482=>"000000011",
  38483=>"100010000",
  38484=>"100000000",
  38485=>"110000001",
  38486=>"000100010",
  38487=>"101011101",
  38488=>"111111011",
  38489=>"101000100",
  38490=>"011101001",
  38491=>"011101101",
  38492=>"001011100",
  38493=>"100000100",
  38494=>"000010011",
  38495=>"001101111",
  38496=>"111100000",
  38497=>"000001111",
  38498=>"110000101",
  38499=>"000011000",
  38500=>"011000110",
  38501=>"100010010",
  38502=>"010001111",
  38503=>"110100011",
  38504=>"000110100",
  38505=>"101010011",
  38506=>"110100110",
  38507=>"001110111",
  38508=>"000101000",
  38509=>"100001110",
  38510=>"111110101",
  38511=>"100010001",
  38512=>"101011000",
  38513=>"000000001",
  38514=>"010010011",
  38515=>"111110001",
  38516=>"100111001",
  38517=>"100011010",
  38518=>"111001001",
  38519=>"111000001",
  38520=>"000010000",
  38521=>"010001010",
  38522=>"100010100",
  38523=>"010011011",
  38524=>"000101110",
  38525=>"000100010",
  38526=>"010111011",
  38527=>"101111100",
  38528=>"101110101",
  38529=>"011010100",
  38530=>"100000011",
  38531=>"000010011",
  38532=>"000010101",
  38533=>"011000010",
  38534=>"111010000",
  38535=>"111111000",
  38536=>"000101100",
  38537=>"111001111",
  38538=>"001010000",
  38539=>"100100001",
  38540=>"010111110",
  38541=>"010110101",
  38542=>"001010111",
  38543=>"001101110",
  38544=>"101101100",
  38545=>"011111101",
  38546=>"111111011",
  38547=>"101001001",
  38548=>"101001111",
  38549=>"111011000",
  38550=>"110101100",
  38551=>"001101000",
  38552=>"100011011",
  38553=>"101100010",
  38554=>"101010110",
  38555=>"101101100",
  38556=>"000001101",
  38557=>"101011010",
  38558=>"011101001",
  38559=>"010001001",
  38560=>"101001101",
  38561=>"100111001",
  38562=>"011011000",
  38563=>"000101110",
  38564=>"110001001",
  38565=>"100111011",
  38566=>"001000001",
  38567=>"111100000",
  38568=>"011110001",
  38569=>"111101110",
  38570=>"111100010",
  38571=>"111001100",
  38572=>"100101011",
  38573=>"000110111",
  38574=>"010110010",
  38575=>"110000100",
  38576=>"000100000",
  38577=>"001111000",
  38578=>"001100101",
  38579=>"111000111",
  38580=>"101010111",
  38581=>"111100110",
  38582=>"110100000",
  38583=>"100101110",
  38584=>"101001111",
  38585=>"000001110",
  38586=>"000101110",
  38587=>"101110100",
  38588=>"100001001",
  38589=>"000001011",
  38590=>"011001011",
  38591=>"001111111",
  38592=>"000110011",
  38593=>"000110001",
  38594=>"011110111",
  38595=>"101101100",
  38596=>"100000100",
  38597=>"111111101",
  38598=>"110110001",
  38599=>"001001000",
  38600=>"100101011",
  38601=>"001111011",
  38602=>"111110010",
  38603=>"011010010",
  38604=>"001100101",
  38605=>"000010000",
  38606=>"000000010",
  38607=>"011101010",
  38608=>"010010010",
  38609=>"100101010",
  38610=>"000011001",
  38611=>"011101110",
  38612=>"001000110",
  38613=>"000010100",
  38614=>"000010100",
  38615=>"010111001",
  38616=>"011111001",
  38617=>"101110011",
  38618=>"001011101",
  38619=>"011100010",
  38620=>"001001111",
  38621=>"110100110",
  38622=>"000101101",
  38623=>"110011110",
  38624=>"101011000",
  38625=>"101101100",
  38626=>"110010011",
  38627=>"110010010",
  38628=>"101101110",
  38629=>"011101010",
  38630=>"000010101",
  38631=>"101000110",
  38632=>"101000101",
  38633=>"011101101",
  38634=>"010100100",
  38635=>"100100100",
  38636=>"000000011",
  38637=>"011111010",
  38638=>"001000101",
  38639=>"110000011",
  38640=>"111010010",
  38641=>"010011011",
  38642=>"100000010",
  38643=>"100001111",
  38644=>"001001110",
  38645=>"011010011",
  38646=>"110111100",
  38647=>"111110101",
  38648=>"010010001",
  38649=>"101011101",
  38650=>"011011000",
  38651=>"010100010",
  38652=>"000011110",
  38653=>"000010111",
  38654=>"000000100",
  38655=>"001001100",
  38656=>"000011110",
  38657=>"001011001",
  38658=>"101100111",
  38659=>"000011000",
  38660=>"000001110",
  38661=>"110000110",
  38662=>"100010100",
  38663=>"110110011",
  38664=>"001101101",
  38665=>"101000010",
  38666=>"110001100",
  38667=>"101110111",
  38668=>"001101111",
  38669=>"110110110",
  38670=>"000101010",
  38671=>"100101001",
  38672=>"000011000",
  38673=>"000010001",
  38674=>"110011100",
  38675=>"001011000",
  38676=>"010110110",
  38677=>"000100001",
  38678=>"111001101",
  38679=>"001000011",
  38680=>"111111011",
  38681=>"010011010",
  38682=>"000111100",
  38683=>"000111101",
  38684=>"000000001",
  38685=>"111110100",
  38686=>"110100110",
  38687=>"110110101",
  38688=>"010000100",
  38689=>"101011001",
  38690=>"000000010",
  38691=>"011111111",
  38692=>"001101101",
  38693=>"000101011",
  38694=>"111010110",
  38695=>"001100111",
  38696=>"100111110",
  38697=>"001001100",
  38698=>"111111111",
  38699=>"010011001",
  38700=>"101001001",
  38701=>"000110110",
  38702=>"000111010",
  38703=>"001111011",
  38704=>"110000001",
  38705=>"101010001",
  38706=>"101010111",
  38707=>"010010101",
  38708=>"100000001",
  38709=>"000101000",
  38710=>"001000100",
  38711=>"011011110",
  38712=>"100101111",
  38713=>"000000001",
  38714=>"000111010",
  38715=>"001000000",
  38716=>"010011001",
  38717=>"100101100",
  38718=>"111110111",
  38719=>"101100110",
  38720=>"101000100",
  38721=>"010011000",
  38722=>"111100011",
  38723=>"110001011",
  38724=>"000110001",
  38725=>"011110100",
  38726=>"000000100",
  38727=>"110010000",
  38728=>"111000111",
  38729=>"100011101",
  38730=>"110100110",
  38731=>"001111011",
  38732=>"110110011",
  38733=>"101101010",
  38734=>"111110100",
  38735=>"010011110",
  38736=>"100100100",
  38737=>"100110111",
  38738=>"100000001",
  38739=>"010010000",
  38740=>"100011001",
  38741=>"101100101",
  38742=>"100110101",
  38743=>"110010100",
  38744=>"000010001",
  38745=>"001110010",
  38746=>"000000010",
  38747=>"011000101",
  38748=>"010110110",
  38749=>"001010001",
  38750=>"010111101",
  38751=>"010101101",
  38752=>"010000010",
  38753=>"011010010",
  38754=>"001000011",
  38755=>"011000000",
  38756=>"010111011",
  38757=>"000110011",
  38758=>"001000000",
  38759=>"011100110",
  38760=>"010101010",
  38761=>"100010111",
  38762=>"000101101",
  38763=>"011100001",
  38764=>"001001010",
  38765=>"110101100",
  38766=>"110101010",
  38767=>"100000011",
  38768=>"101000011",
  38769=>"100100011",
  38770=>"101111100",
  38771=>"001100000",
  38772=>"011100000",
  38773=>"100000000",
  38774=>"100001111",
  38775=>"100111000",
  38776=>"111100010",
  38777=>"011011000",
  38778=>"110110111",
  38779=>"100011110",
  38780=>"111001111",
  38781=>"111111101",
  38782=>"001001011",
  38783=>"101111101",
  38784=>"111111000",
  38785=>"001110011",
  38786=>"011100001",
  38787=>"001011110",
  38788=>"100001000",
  38789=>"010011110",
  38790=>"101111101",
  38791=>"100100011",
  38792=>"010111111",
  38793=>"010111010",
  38794=>"101010110",
  38795=>"011001011",
  38796=>"000110000",
  38797=>"011010000",
  38798=>"001010111",
  38799=>"100101010",
  38800=>"000000001",
  38801=>"110101100",
  38802=>"100010000",
  38803=>"010110011",
  38804=>"010001000",
  38805=>"011101111",
  38806=>"001111101",
  38807=>"011101101",
  38808=>"011100011",
  38809=>"100011000",
  38810=>"101100110",
  38811=>"001011011",
  38812=>"010011011",
  38813=>"000110010",
  38814=>"100010011",
  38815=>"110001111",
  38816=>"110100100",
  38817=>"110011010",
  38818=>"010011000",
  38819=>"001101011",
  38820=>"000001000",
  38821=>"101101100",
  38822=>"110111101",
  38823=>"000101100",
  38824=>"101110110",
  38825=>"000000101",
  38826=>"010011111",
  38827=>"111100000",
  38828=>"011000110",
  38829=>"110101001",
  38830=>"110100111",
  38831=>"100100010",
  38832=>"010100001",
  38833=>"001111110",
  38834=>"000000011",
  38835=>"000100011",
  38836=>"010110110",
  38837=>"001111101",
  38838=>"011100010",
  38839=>"000000000",
  38840=>"111110000",
  38841=>"000000100",
  38842=>"000110101",
  38843=>"111011101",
  38844=>"010011010",
  38845=>"010111110",
  38846=>"001101101",
  38847=>"101000100",
  38848=>"111111110",
  38849=>"110110111",
  38850=>"011111010",
  38851=>"111100111",
  38852=>"111001000",
  38853=>"000100011",
  38854=>"001110011",
  38855=>"100110001",
  38856=>"000010111",
  38857=>"100010000",
  38858=>"111110000",
  38859=>"010000100",
  38860=>"011101010",
  38861=>"101011001",
  38862=>"101110110",
  38863=>"011010010",
  38864=>"110000011",
  38865=>"100111001",
  38866=>"100110011",
  38867=>"010110101",
  38868=>"000100011",
  38869=>"111001111",
  38870=>"110100100",
  38871=>"100000100",
  38872=>"100000011",
  38873=>"000110111",
  38874=>"010010000",
  38875=>"010011000",
  38876=>"111101110",
  38877=>"111110110",
  38878=>"001010100",
  38879=>"111100110",
  38880=>"010010101",
  38881=>"011000000",
  38882=>"100111111",
  38883=>"001010101",
  38884=>"111101001",
  38885=>"110100100",
  38886=>"110010110",
  38887=>"000101110",
  38888=>"101000101",
  38889=>"100011110",
  38890=>"110011011",
  38891=>"011000111",
  38892=>"001110001",
  38893=>"101000010",
  38894=>"010001000",
  38895=>"000010010",
  38896=>"010111010",
  38897=>"001111111",
  38898=>"111101111",
  38899=>"000000101",
  38900=>"010101000",
  38901=>"001011000",
  38902=>"001010001",
  38903=>"110001010",
  38904=>"001011010",
  38905=>"001010111",
  38906=>"001111111",
  38907=>"111111000",
  38908=>"100100100",
  38909=>"111110100",
  38910=>"000010110",
  38911=>"100010011",
  38912=>"111100111",
  38913=>"110010010",
  38914=>"111100100",
  38915=>"100001111",
  38916=>"001000111",
  38917=>"111001011",
  38918=>"010001001",
  38919=>"100111010",
  38920=>"100101101",
  38921=>"001010001",
  38922=>"100001100",
  38923=>"110100011",
  38924=>"101110010",
  38925=>"010101101",
  38926=>"001011111",
  38927=>"100000000",
  38928=>"111110001",
  38929=>"100101110",
  38930=>"101010101",
  38931=>"010100100",
  38932=>"101100010",
  38933=>"000000001",
  38934=>"110011111",
  38935=>"010011001",
  38936=>"111000010",
  38937=>"111101111",
  38938=>"010010000",
  38939=>"001010011",
  38940=>"001110001",
  38941=>"101001010",
  38942=>"001001001",
  38943=>"101011011",
  38944=>"010011001",
  38945=>"000110110",
  38946=>"000000110",
  38947=>"110110111",
  38948=>"011100000",
  38949=>"001110101",
  38950=>"011111000",
  38951=>"000111110",
  38952=>"011111010",
  38953=>"101101010",
  38954=>"101000000",
  38955=>"011100000",
  38956=>"011100111",
  38957=>"111011011",
  38958=>"101111001",
  38959=>"001110110",
  38960=>"111010110",
  38961=>"000000011",
  38962=>"001010001",
  38963=>"111111010",
  38964=>"101110111",
  38965=>"010110110",
  38966=>"100111000",
  38967=>"001001000",
  38968=>"000101000",
  38969=>"110101100",
  38970=>"001101111",
  38971=>"010100101",
  38972=>"110001010",
  38973=>"010110001",
  38974=>"100100111",
  38975=>"000111011",
  38976=>"101011100",
  38977=>"010100011",
  38978=>"001101000",
  38979=>"010101110",
  38980=>"000000100",
  38981=>"000100101",
  38982=>"000101000",
  38983=>"101100011",
  38984=>"111110011",
  38985=>"101000101",
  38986=>"000110111",
  38987=>"000110110",
  38988=>"111100111",
  38989=>"101111010",
  38990=>"100000100",
  38991=>"001011001",
  38992=>"010111011",
  38993=>"011001110",
  38994=>"011011010",
  38995=>"111001111",
  38996=>"100001110",
  38997=>"101100011",
  38998=>"000110101",
  38999=>"001001011",
  39000=>"011100011",
  39001=>"001011001",
  39002=>"011001110",
  39003=>"011000010",
  39004=>"010100010",
  39005=>"000100000",
  39006=>"100111100",
  39007=>"100001100",
  39008=>"000001010",
  39009=>"100011011",
  39010=>"001000000",
  39011=>"000101100",
  39012=>"010000010",
  39013=>"101100010",
  39014=>"100010100",
  39015=>"001111000",
  39016=>"101100111",
  39017=>"101001000",
  39018=>"001110011",
  39019=>"111101111",
  39020=>"101101010",
  39021=>"011111110",
  39022=>"111010001",
  39023=>"000110010",
  39024=>"001001100",
  39025=>"001010100",
  39026=>"001101011",
  39027=>"100110110",
  39028=>"000010000",
  39029=>"100101101",
  39030=>"010111101",
  39031=>"010101011",
  39032=>"101101010",
  39033=>"010111010",
  39034=>"100010100",
  39035=>"101011111",
  39036=>"110111011",
  39037=>"010011100",
  39038=>"110111010",
  39039=>"111011110",
  39040=>"111011000",
  39041=>"100010001",
  39042=>"001001000",
  39043=>"111001010",
  39044=>"101001010",
  39045=>"111100001",
  39046=>"111010010",
  39047=>"000100001",
  39048=>"000110100",
  39049=>"001100011",
  39050=>"011100000",
  39051=>"100011111",
  39052=>"101111001",
  39053=>"100111010",
  39054=>"100111001",
  39055=>"110100100",
  39056=>"110101111",
  39057=>"111011010",
  39058=>"011110000",
  39059=>"110110000",
  39060=>"000101001",
  39061=>"010010111",
  39062=>"010010111",
  39063=>"000010100",
  39064=>"111000110",
  39065=>"100000111",
  39066=>"010000111",
  39067=>"000110100",
  39068=>"001100011",
  39069=>"000010101",
  39070=>"100101101",
  39071=>"011010010",
  39072=>"011000111",
  39073=>"000011110",
  39074=>"001110010",
  39075=>"111001101",
  39076=>"010001001",
  39077=>"010111010",
  39078=>"111101100",
  39079=>"010010000",
  39080=>"001100111",
  39081=>"000010000",
  39082=>"010001000",
  39083=>"111101110",
  39084=>"110110001",
  39085=>"010110100",
  39086=>"011101001",
  39087=>"010011001",
  39088=>"110101101",
  39089=>"100001001",
  39090=>"001011100",
  39091=>"011001001",
  39092=>"101101111",
  39093=>"010000111",
  39094=>"100010100",
  39095=>"110000000",
  39096=>"000111010",
  39097=>"001001111",
  39098=>"100100011",
  39099=>"100000001",
  39100=>"001010101",
  39101=>"110110101",
  39102=>"011001010",
  39103=>"101110011",
  39104=>"100100101",
  39105=>"111110010",
  39106=>"000110000",
  39107=>"011010000",
  39108=>"001011111",
  39109=>"000000010",
  39110=>"001100000",
  39111=>"100010111",
  39112=>"100010011",
  39113=>"111101100",
  39114=>"010000100",
  39115=>"001110011",
  39116=>"111101100",
  39117=>"010011101",
  39118=>"010011110",
  39119=>"010001110",
  39120=>"000011101",
  39121=>"100101101",
  39122=>"010100001",
  39123=>"001010000",
  39124=>"011000110",
  39125=>"001011011",
  39126=>"100101000",
  39127=>"111101011",
  39128=>"111000000",
  39129=>"111101000",
  39130=>"111001101",
  39131=>"000000110",
  39132=>"010011000",
  39133=>"011000001",
  39134=>"101100000",
  39135=>"000100010",
  39136=>"100000110",
  39137=>"011111001",
  39138=>"000100100",
  39139=>"001000100",
  39140=>"110011101",
  39141=>"001011001",
  39142=>"101010110",
  39143=>"110001110",
  39144=>"100011111",
  39145=>"001010011",
  39146=>"011111110",
  39147=>"011100101",
  39148=>"111010111",
  39149=>"001000101",
  39150=>"001110010",
  39151=>"111101000",
  39152=>"000000011",
  39153=>"100010001",
  39154=>"101110111",
  39155=>"011010111",
  39156=>"101010101",
  39157=>"011100100",
  39158=>"011111110",
  39159=>"100000010",
  39160=>"111110111",
  39161=>"101000010",
  39162=>"110111101",
  39163=>"010001110",
  39164=>"001111100",
  39165=>"000001000",
  39166=>"000101010",
  39167=>"001111101",
  39168=>"111110100",
  39169=>"000111001",
  39170=>"011001110",
  39171=>"111011010",
  39172=>"001101001",
  39173=>"101101001",
  39174=>"001110000",
  39175=>"100011000",
  39176=>"000111111",
  39177=>"000010100",
  39178=>"100101000",
  39179=>"000111101",
  39180=>"010101111",
  39181=>"000011011",
  39182=>"001000111",
  39183=>"100110101",
  39184=>"001101001",
  39185=>"111110111",
  39186=>"000001000",
  39187=>"111001111",
  39188=>"101110100",
  39189=>"111001001",
  39190=>"010000111",
  39191=>"001101010",
  39192=>"101100100",
  39193=>"001110011",
  39194=>"000110000",
  39195=>"110101001",
  39196=>"101010101",
  39197=>"010111110",
  39198=>"010101010",
  39199=>"101100101",
  39200=>"100111010",
  39201=>"111111011",
  39202=>"110011011",
  39203=>"000101111",
  39204=>"100011110",
  39205=>"010110010",
  39206=>"011110111",
  39207=>"111001100",
  39208=>"000101111",
  39209=>"010110010",
  39210=>"011010101",
  39211=>"011111100",
  39212=>"111011101",
  39213=>"100010100",
  39214=>"011111110",
  39215=>"011100110",
  39216=>"000001101",
  39217=>"101100100",
  39218=>"011100111",
  39219=>"110001001",
  39220=>"010110011",
  39221=>"001101011",
  39222=>"101000101",
  39223=>"111111111",
  39224=>"010100011",
  39225=>"001100000",
  39226=>"111011010",
  39227=>"011110101",
  39228=>"011010100",
  39229=>"010110011",
  39230=>"000000110",
  39231=>"010101000",
  39232=>"101100011",
  39233=>"000101011",
  39234=>"111110111",
  39235=>"100010111",
  39236=>"111110011",
  39237=>"110101001",
  39238=>"001111001",
  39239=>"110011001",
  39240=>"010110100",
  39241=>"101111011",
  39242=>"011101010",
  39243=>"011010001",
  39244=>"001100110",
  39245=>"011010011",
  39246=>"001000000",
  39247=>"011000001",
  39248=>"110110010",
  39249=>"101100011",
  39250=>"111100111",
  39251=>"011101110",
  39252=>"000010001",
  39253=>"001110011",
  39254=>"000110000",
  39255=>"000011010",
  39256=>"011000000",
  39257=>"000000000",
  39258=>"110010101",
  39259=>"000100110",
  39260=>"010001110",
  39261=>"001000000",
  39262=>"000111010",
  39263=>"010110101",
  39264=>"110101101",
  39265=>"101011111",
  39266=>"100101001",
  39267=>"001111111",
  39268=>"100101100",
  39269=>"111000111",
  39270=>"011111101",
  39271=>"001111111",
  39272=>"000110001",
  39273=>"000001010",
  39274=>"101101000",
  39275=>"000111101",
  39276=>"101111111",
  39277=>"110111100",
  39278=>"001000011",
  39279=>"111000001",
  39280=>"101111111",
  39281=>"100001001",
  39282=>"001000101",
  39283=>"000000110",
  39284=>"110010101",
  39285=>"010011110",
  39286=>"010011111",
  39287=>"111111110",
  39288=>"010011011",
  39289=>"011000100",
  39290=>"000100011",
  39291=>"111010010",
  39292=>"001111000",
  39293=>"100011101",
  39294=>"110110010",
  39295=>"110110110",
  39296=>"110110110",
  39297=>"000000101",
  39298=>"000000010",
  39299=>"101111000",
  39300=>"100101010",
  39301=>"110001101",
  39302=>"100111010",
  39303=>"111000100",
  39304=>"110100011",
  39305=>"000110000",
  39306=>"111010101",
  39307=>"010100101",
  39308=>"110100100",
  39309=>"011111010",
  39310=>"011100001",
  39311=>"001110111",
  39312=>"010111010",
  39313=>"010101100",
  39314=>"000100100",
  39315=>"001110100",
  39316=>"110100100",
  39317=>"110011010",
  39318=>"110011110",
  39319=>"011100101",
  39320=>"101001101",
  39321=>"001100000",
  39322=>"001000001",
  39323=>"110111101",
  39324=>"011000110",
  39325=>"101000111",
  39326=>"111001110",
  39327=>"011111011",
  39328=>"010100000",
  39329=>"111111001",
  39330=>"101101011",
  39331=>"100011000",
  39332=>"100001001",
  39333=>"101001111",
  39334=>"101110110",
  39335=>"101100000",
  39336=>"100011100",
  39337=>"110010000",
  39338=>"010010100",
  39339=>"111111010",
  39340=>"101001011",
  39341=>"101111011",
  39342=>"111010111",
  39343=>"110010010",
  39344=>"100010101",
  39345=>"011100001",
  39346=>"101010111",
  39347=>"101111101",
  39348=>"000011100",
  39349=>"111111010",
  39350=>"001001111",
  39351=>"110110111",
  39352=>"100100011",
  39353=>"011100000",
  39354=>"000011011",
  39355=>"010001100",
  39356=>"011001110",
  39357=>"011010000",
  39358=>"110101110",
  39359=>"101001011",
  39360=>"001000100",
  39361=>"110011101",
  39362=>"000111010",
  39363=>"101001010",
  39364=>"011011011",
  39365=>"001001000",
  39366=>"000000110",
  39367=>"111011100",
  39368=>"111111011",
  39369=>"100001101",
  39370=>"010010010",
  39371=>"110101100",
  39372=>"000000010",
  39373=>"001000001",
  39374=>"110001001",
  39375=>"010001000",
  39376=>"101111000",
  39377=>"000001100",
  39378=>"011011101",
  39379=>"011101010",
  39380=>"001001101",
  39381=>"010101010",
  39382=>"100011001",
  39383=>"111011000",
  39384=>"011001000",
  39385=>"111010011",
  39386=>"011010000",
  39387=>"010010111",
  39388=>"110111010",
  39389=>"000010000",
  39390=>"001000111",
  39391=>"010100010",
  39392=>"000101100",
  39393=>"011101010",
  39394=>"001000101",
  39395=>"010111100",
  39396=>"101001101",
  39397=>"100111011",
  39398=>"110011110",
  39399=>"011100101",
  39400=>"011101100",
  39401=>"000101001",
  39402=>"000110010",
  39403=>"001001110",
  39404=>"000010011",
  39405=>"010111110",
  39406=>"000111011",
  39407=>"001010000",
  39408=>"010001001",
  39409=>"001101000",
  39410=>"101001011",
  39411=>"101101100",
  39412=>"110100010",
  39413=>"100101000",
  39414=>"101010010",
  39415=>"111011000",
  39416=>"110100101",
  39417=>"011001001",
  39418=>"000110100",
  39419=>"100111100",
  39420=>"111110000",
  39421=>"011100001",
  39422=>"111000000",
  39423=>"101001011",
  39424=>"110000100",
  39425=>"100100101",
  39426=>"010010010",
  39427=>"110110110",
  39428=>"100101001",
  39429=>"100000100",
  39430=>"110100111",
  39431=>"100001000",
  39432=>"000011011",
  39433=>"000011110",
  39434=>"010111011",
  39435=>"001010110",
  39436=>"000001011",
  39437=>"010100101",
  39438=>"111101011",
  39439=>"001010100",
  39440=>"100010110",
  39441=>"100100011",
  39442=>"100001010",
  39443=>"000101110",
  39444=>"000000011",
  39445=>"111011111",
  39446=>"011101010",
  39447=>"110011000",
  39448=>"101001010",
  39449=>"110100010",
  39450=>"010011110",
  39451=>"011010000",
  39452=>"000011100",
  39453=>"111001101",
  39454=>"001111000",
  39455=>"010110000",
  39456=>"011011111",
  39457=>"101001010",
  39458=>"001110110",
  39459=>"000101011",
  39460=>"100101011",
  39461=>"001110001",
  39462=>"100101100",
  39463=>"111001100",
  39464=>"010010011",
  39465=>"001110011",
  39466=>"110001010",
  39467=>"111110101",
  39468=>"100000000",
  39469=>"100001000",
  39470=>"010001101",
  39471=>"101101011",
  39472=>"100010000",
  39473=>"011111000",
  39474=>"101001010",
  39475=>"100100110",
  39476=>"010100100",
  39477=>"000101011",
  39478=>"011101100",
  39479=>"110100011",
  39480=>"100110100",
  39481=>"001100101",
  39482=>"001000101",
  39483=>"010001010",
  39484=>"010111110",
  39485=>"011011000",
  39486=>"101110010",
  39487=>"101011011",
  39488=>"001011001",
  39489=>"101000011",
  39490=>"101111110",
  39491=>"000011001",
  39492=>"001001010",
  39493=>"001011111",
  39494=>"011000001",
  39495=>"110000101",
  39496=>"110110110",
  39497=>"110001001",
  39498=>"010001000",
  39499=>"011100010",
  39500=>"110001010",
  39501=>"100100101",
  39502=>"110010111",
  39503=>"010010110",
  39504=>"011001001",
  39505=>"010111111",
  39506=>"000010101",
  39507=>"100010001",
  39508=>"101111101",
  39509=>"000011110",
  39510=>"000001011",
  39511=>"101101010",
  39512=>"011101111",
  39513=>"111110011",
  39514=>"011101111",
  39515=>"011010101",
  39516=>"111101000",
  39517=>"101000101",
  39518=>"110011001",
  39519=>"010000100",
  39520=>"001011000",
  39521=>"000000000",
  39522=>"000010001",
  39523=>"011110010",
  39524=>"100010111",
  39525=>"100000000",
  39526=>"010010001",
  39527=>"001101111",
  39528=>"000000001",
  39529=>"111010011",
  39530=>"001000101",
  39531=>"100000000",
  39532=>"101010111",
  39533=>"101111110",
  39534=>"100000101",
  39535=>"111001000",
  39536=>"001011010",
  39537=>"001001111",
  39538=>"000000111",
  39539=>"011111001",
  39540=>"101001011",
  39541=>"111111110",
  39542=>"100000010",
  39543=>"001101111",
  39544=>"010010001",
  39545=>"110010011",
  39546=>"101001100",
  39547=>"011111011",
  39548=>"001001000",
  39549=>"000100111",
  39550=>"101110100",
  39551=>"110111101",
  39552=>"110010111",
  39553=>"010100001",
  39554=>"111111111",
  39555=>"011100000",
  39556=>"100001010",
  39557=>"110100000",
  39558=>"010001010",
  39559=>"101011001",
  39560=>"010110000",
  39561=>"001111111",
  39562=>"110101001",
  39563=>"011101010",
  39564=>"000011001",
  39565=>"101110011",
  39566=>"001100110",
  39567=>"110001000",
  39568=>"101101011",
  39569=>"000100000",
  39570=>"110010111",
  39571=>"101010100",
  39572=>"010001101",
  39573=>"010110101",
  39574=>"010110110",
  39575=>"101010101",
  39576=>"001000110",
  39577=>"110000101",
  39578=>"111111101",
  39579=>"001110111",
  39580=>"111000111",
  39581=>"001100000",
  39582=>"010111111",
  39583=>"111001111",
  39584=>"110001001",
  39585=>"011101000",
  39586=>"010011000",
  39587=>"111110001",
  39588=>"101011001",
  39589=>"101111001",
  39590=>"011010101",
  39591=>"000000000",
  39592=>"001111111",
  39593=>"111101101",
  39594=>"001001011",
  39595=>"101011101",
  39596=>"110010000",
  39597=>"110101101",
  39598=>"111010010",
  39599=>"111000111",
  39600=>"011111010",
  39601=>"100000011",
  39602=>"101110100",
  39603=>"111110100",
  39604=>"000100110",
  39605=>"100110011",
  39606=>"000000011",
  39607=>"101010111",
  39608=>"000000000",
  39609=>"001010100",
  39610=>"100011000",
  39611=>"001100010",
  39612=>"100111000",
  39613=>"011101101",
  39614=>"000111100",
  39615=>"110000000",
  39616=>"010111011",
  39617=>"001100001",
  39618=>"111100101",
  39619=>"011100110",
  39620=>"011001000",
  39621=>"101010111",
  39622=>"011000110",
  39623=>"010000000",
  39624=>"010100010",
  39625=>"010100000",
  39626=>"000000010",
  39627=>"101101000",
  39628=>"000111000",
  39629=>"100110111",
  39630=>"110111100",
  39631=>"000111110",
  39632=>"101111010",
  39633=>"000001110",
  39634=>"011001001",
  39635=>"101011110",
  39636=>"001110010",
  39637=>"100010010",
  39638=>"000011100",
  39639=>"110101000",
  39640=>"101100001",
  39641=>"010000100",
  39642=>"000110011",
  39643=>"011000000",
  39644=>"001000111",
  39645=>"010110110",
  39646=>"100000011",
  39647=>"011100010",
  39648=>"100010110",
  39649=>"011000010",
  39650=>"110001111",
  39651=>"100011111",
  39652=>"001000111",
  39653=>"001110110",
  39654=>"110011001",
  39655=>"000000100",
  39656=>"010000110",
  39657=>"111000101",
  39658=>"010000100",
  39659=>"100100100",
  39660=>"100101001",
  39661=>"010011011",
  39662=>"000000111",
  39663=>"001101110",
  39664=>"101010010",
  39665=>"011000110",
  39666=>"001111101",
  39667=>"111100000",
  39668=>"001101110",
  39669=>"001111011",
  39670=>"001011110",
  39671=>"011010010",
  39672=>"000011001",
  39673=>"000000000",
  39674=>"100110100",
  39675=>"110000100",
  39676=>"110111100",
  39677=>"111000000",
  39678=>"010001011",
  39679=>"000011010",
  39680=>"010011110",
  39681=>"000011110",
  39682=>"000001000",
  39683=>"001001100",
  39684=>"100100101",
  39685=>"100111000",
  39686=>"001011001",
  39687=>"100000001",
  39688=>"110111010",
  39689=>"111010100",
  39690=>"110001100",
  39691=>"110100111",
  39692=>"011111011",
  39693=>"111110100",
  39694=>"111010011",
  39695=>"110010101",
  39696=>"010101011",
  39697=>"001111111",
  39698=>"010101001",
  39699=>"000101111",
  39700=>"011100101",
  39701=>"000100010",
  39702=>"011101110",
  39703=>"111111011",
  39704=>"100010110",
  39705=>"010100100",
  39706=>"110111000",
  39707=>"101000111",
  39708=>"100010010",
  39709=>"100110111",
  39710=>"111110111",
  39711=>"111001100",
  39712=>"110000000",
  39713=>"111011010",
  39714=>"010000110",
  39715=>"111011111",
  39716=>"000000010",
  39717=>"001111001",
  39718=>"011011001",
  39719=>"010101001",
  39720=>"111111110",
  39721=>"100100111",
  39722=>"000010100",
  39723=>"010000110",
  39724=>"111100101",
  39725=>"111111111",
  39726=>"101001111",
  39727=>"011000111",
  39728=>"101001001",
  39729=>"000100101",
  39730=>"001000100",
  39731=>"000101100",
  39732=>"111011000",
  39733=>"111001101",
  39734=>"000100101",
  39735=>"110011010",
  39736=>"101110010",
  39737=>"011011100",
  39738=>"100010111",
  39739=>"001001110",
  39740=>"000100001",
  39741=>"111000010",
  39742=>"100101011",
  39743=>"101001101",
  39744=>"101100001",
  39745=>"111011001",
  39746=>"001110101",
  39747=>"011111111",
  39748=>"010001100",
  39749=>"010010110",
  39750=>"101101000",
  39751=>"101100100",
  39752=>"111001001",
  39753=>"100001111",
  39754=>"001001000",
  39755=>"101011011",
  39756=>"000110110",
  39757=>"011110101",
  39758=>"001100111",
  39759=>"001101010",
  39760=>"000101100",
  39761=>"111100100",
  39762=>"111111011",
  39763=>"011100010",
  39764=>"111000001",
  39765=>"011110100",
  39766=>"000011110",
  39767=>"010111101",
  39768=>"100000011",
  39769=>"000111110",
  39770=>"110110101",
  39771=>"011010100",
  39772=>"100111010",
  39773=>"100000011",
  39774=>"111000000",
  39775=>"000010010",
  39776=>"011000100",
  39777=>"110001011",
  39778=>"110100110",
  39779=>"011111001",
  39780=>"010110101",
  39781=>"000000111",
  39782=>"010011001",
  39783=>"010000111",
  39784=>"101110111",
  39785=>"010111001",
  39786=>"010110110",
  39787=>"001101111",
  39788=>"011110111",
  39789=>"100101001",
  39790=>"000001101",
  39791=>"110011100",
  39792=>"101100110",
  39793=>"111010101",
  39794=>"000000100",
  39795=>"011110000",
  39796=>"001001011",
  39797=>"001110010",
  39798=>"111110011",
  39799=>"010001001",
  39800=>"000100100",
  39801=>"010100001",
  39802=>"111000101",
  39803=>"000001101",
  39804=>"001001000",
  39805=>"011000110",
  39806=>"011001011",
  39807=>"000110100",
  39808=>"000110011",
  39809=>"000010101",
  39810=>"110111100",
  39811=>"010100011",
  39812=>"001100010",
  39813=>"110001110",
  39814=>"001001111",
  39815=>"111110011",
  39816=>"000110101",
  39817=>"110001101",
  39818=>"000000010",
  39819=>"000110100",
  39820=>"000010100",
  39821=>"111101010",
  39822=>"110100111",
  39823=>"010110100",
  39824=>"000100011",
  39825=>"000011111",
  39826=>"100010100",
  39827=>"010011101",
  39828=>"011010110",
  39829=>"001111000",
  39830=>"111100001",
  39831=>"001010011",
  39832=>"101110101",
  39833=>"000001001",
  39834=>"010001100",
  39835=>"000010101",
  39836=>"100110101",
  39837=>"000011111",
  39838=>"110010000",
  39839=>"110111111",
  39840=>"101100110",
  39841=>"110111001",
  39842=>"111111011",
  39843=>"000101110",
  39844=>"101100000",
  39845=>"110111110",
  39846=>"100100011",
  39847=>"001010110",
  39848=>"011111011",
  39849=>"111000101",
  39850=>"000111110",
  39851=>"110011111",
  39852=>"000110001",
  39853=>"111010011",
  39854=>"100100000",
  39855=>"101101001",
  39856=>"011101001",
  39857=>"000111010",
  39858=>"010011010",
  39859=>"010010100",
  39860=>"111101011",
  39861=>"100000000",
  39862=>"010001000",
  39863=>"010101001",
  39864=>"111111010",
  39865=>"101011101",
  39866=>"011111100",
  39867=>"111100001",
  39868=>"101111100",
  39869=>"110011000",
  39870=>"111100100",
  39871=>"010111100",
  39872=>"100011001",
  39873=>"110001000",
  39874=>"110110110",
  39875=>"001001100",
  39876=>"001001010",
  39877=>"000110110",
  39878=>"011101000",
  39879=>"100011010",
  39880=>"100100010",
  39881=>"011111001",
  39882=>"010010011",
  39883=>"011111100",
  39884=>"011000110",
  39885=>"100001010",
  39886=>"000110011",
  39887=>"010010110",
  39888=>"010010101",
  39889=>"101111101",
  39890=>"011110111",
  39891=>"010001001",
  39892=>"111110001",
  39893=>"100000100",
  39894=>"001101001",
  39895=>"011101101",
  39896=>"000000000",
  39897=>"100110100",
  39898=>"011010001",
  39899=>"101001100",
  39900=>"111000111",
  39901=>"000011010",
  39902=>"111011000",
  39903=>"001000011",
  39904=>"000001011",
  39905=>"100100110",
  39906=>"111101100",
  39907=>"001011111",
  39908=>"100010010",
  39909=>"100011110",
  39910=>"110100011",
  39911=>"001111111",
  39912=>"000101101",
  39913=>"101111011",
  39914=>"010001111",
  39915=>"101010110",
  39916=>"101101001",
  39917=>"000011111",
  39918=>"111000001",
  39919=>"111100110",
  39920=>"000000000",
  39921=>"111100010",
  39922=>"000001001",
  39923=>"000010110",
  39924=>"001001010",
  39925=>"100010111",
  39926=>"011110101",
  39927=>"011101111",
  39928=>"111100110",
  39929=>"101010101",
  39930=>"100101111",
  39931=>"110111000",
  39932=>"111000101",
  39933=>"101101000",
  39934=>"111110001",
  39935=>"101010011",
  39936=>"010101111",
  39937=>"110111111",
  39938=>"110110010",
  39939=>"111101100",
  39940=>"011001000",
  39941=>"011000001",
  39942=>"001000011",
  39943=>"111001010",
  39944=>"100010111",
  39945=>"001000010",
  39946=>"100000001",
  39947=>"011010010",
  39948=>"010100101",
  39949=>"111001011",
  39950=>"010000001",
  39951=>"010010010",
  39952=>"001000101",
  39953=>"100000110",
  39954=>"111000100",
  39955=>"100010110",
  39956=>"010100011",
  39957=>"000100110",
  39958=>"011011011",
  39959=>"111100101",
  39960=>"000111000",
  39961=>"000101000",
  39962=>"011101101",
  39963=>"001100001",
  39964=>"000001111",
  39965=>"000010111",
  39966=>"010000001",
  39967=>"000011001",
  39968=>"001101010",
  39969=>"001100111",
  39970=>"111111111",
  39971=>"000000000",
  39972=>"100101001",
  39973=>"000101010",
  39974=>"000000011",
  39975=>"001100011",
  39976=>"111110001",
  39977=>"100111100",
  39978=>"000001001",
  39979=>"011011001",
  39980=>"011110011",
  39981=>"111001100",
  39982=>"010001101",
  39983=>"000110100",
  39984=>"010111110",
  39985=>"101010001",
  39986=>"011101110",
  39987=>"111110101",
  39988=>"001010011",
  39989=>"001101101",
  39990=>"001010101",
  39991=>"001100101",
  39992=>"001000001",
  39993=>"011111001",
  39994=>"000110111",
  39995=>"101011000",
  39996=>"010110011",
  39997=>"001011000",
  39998=>"100001110",
  39999=>"111100000",
  40000=>"011001011",
  40001=>"111000100",
  40002=>"001111010",
  40003=>"100110111",
  40004=>"110011101",
  40005=>"010000111",
  40006=>"100111111",
  40007=>"101101100",
  40008=>"100100101",
  40009=>"100000110",
  40010=>"111100011",
  40011=>"011010010",
  40012=>"001000010",
  40013=>"100000111",
  40014=>"001100101",
  40015=>"110100000",
  40016=>"100101100",
  40017=>"001101101",
  40018=>"110010100",
  40019=>"010111100",
  40020=>"101101001",
  40021=>"011011110",
  40022=>"111011110",
  40023=>"001101000",
  40024=>"011101100",
  40025=>"000111111",
  40026=>"000011100",
  40027=>"101101001",
  40028=>"111000011",
  40029=>"001001001",
  40030=>"001011010",
  40031=>"010111111",
  40032=>"101000011",
  40033=>"011111000",
  40034=>"001001100",
  40035=>"010000100",
  40036=>"101010001",
  40037=>"111010101",
  40038=>"011100100",
  40039=>"000010000",
  40040=>"111011111",
  40041=>"101011101",
  40042=>"110110100",
  40043=>"001010011",
  40044=>"000101101",
  40045=>"000111101",
  40046=>"011011001",
  40047=>"101001110",
  40048=>"000001101",
  40049=>"000000111",
  40050=>"111110111",
  40051=>"100110000",
  40052=>"010101001",
  40053=>"101111101",
  40054=>"000011010",
  40055=>"010110010",
  40056=>"111101011",
  40057=>"101011110",
  40058=>"001101000",
  40059=>"010110000",
  40060=>"110101110",
  40061=>"010100101",
  40062=>"001011010",
  40063=>"111100000",
  40064=>"110111100",
  40065=>"110001001",
  40066=>"010001100",
  40067=>"000011010",
  40068=>"001001110",
  40069=>"101101111",
  40070=>"000010110",
  40071=>"001100010",
  40072=>"010010000",
  40073=>"110000110",
  40074=>"000011011",
  40075=>"010000111",
  40076=>"110001010",
  40077=>"101100110",
  40078=>"001101111",
  40079=>"100011100",
  40080=>"111100111",
  40081=>"011011110",
  40082=>"000110100",
  40083=>"101110110",
  40084=>"010011111",
  40085=>"101001011",
  40086=>"110111111",
  40087=>"110111011",
  40088=>"010110100",
  40089=>"100010111",
  40090=>"011100100",
  40091=>"101001001",
  40092=>"011101011",
  40093=>"011010100",
  40094=>"011011010",
  40095=>"101100001",
  40096=>"100111010",
  40097=>"111011110",
  40098=>"100010101",
  40099=>"011101001",
  40100=>"010111010",
  40101=>"010010000",
  40102=>"011110111",
  40103=>"001001000",
  40104=>"110010110",
  40105=>"010010010",
  40106=>"101011010",
  40107=>"000010101",
  40108=>"111110101",
  40109=>"000010101",
  40110=>"000100011",
  40111=>"010101101",
  40112=>"101001101",
  40113=>"111100001",
  40114=>"001110111",
  40115=>"101011001",
  40116=>"110010111",
  40117=>"010000111",
  40118=>"000111101",
  40119=>"001011101",
  40120=>"010000000",
  40121=>"100101111",
  40122=>"111001001",
  40123=>"001101010",
  40124=>"110100011",
  40125=>"010000110",
  40126=>"001001000",
  40127=>"011000111",
  40128=>"011010011",
  40129=>"001111000",
  40130=>"111110000",
  40131=>"110010011",
  40132=>"100010100",
  40133=>"010101011",
  40134=>"011111100",
  40135=>"100010110",
  40136=>"010000110",
  40137=>"110000011",
  40138=>"011010001",
  40139=>"111100010",
  40140=>"000100000",
  40141=>"000100101",
  40142=>"100001010",
  40143=>"100011010",
  40144=>"000101001",
  40145=>"001010011",
  40146=>"011001100",
  40147=>"110111010",
  40148=>"011111111",
  40149=>"000101000",
  40150=>"101001000",
  40151=>"000101001",
  40152=>"011001011",
  40153=>"001111011",
  40154=>"101000010",
  40155=>"011111001",
  40156=>"001011010",
  40157=>"001000000",
  40158=>"010101011",
  40159=>"100101000",
  40160=>"100000011",
  40161=>"011001111",
  40162=>"101111010",
  40163=>"010000001",
  40164=>"100101111",
  40165=>"011011111",
  40166=>"110111110",
  40167=>"000111001",
  40168=>"000010110",
  40169=>"111000011",
  40170=>"011101110",
  40171=>"111000001",
  40172=>"110100000",
  40173=>"110011100",
  40174=>"001001001",
  40175=>"010011110",
  40176=>"100111110",
  40177=>"111101110",
  40178=>"101100111",
  40179=>"001101110",
  40180=>"111010110",
  40181=>"010100010",
  40182=>"110100111",
  40183=>"111000010",
  40184=>"101010111",
  40185=>"101010001",
  40186=>"100010101",
  40187=>"010001011",
  40188=>"101001001",
  40189=>"110001110",
  40190=>"001110100",
  40191=>"000011101",
  40192=>"111100110",
  40193=>"011110101",
  40194=>"001010011",
  40195=>"100011100",
  40196=>"111111010",
  40197=>"000101110",
  40198=>"011111011",
  40199=>"110101110",
  40200=>"100100001",
  40201=>"110010110",
  40202=>"101010110",
  40203=>"001101100",
  40204=>"000000100",
  40205=>"000010010",
  40206=>"101111111",
  40207=>"001110001",
  40208=>"111110010",
  40209=>"011000001",
  40210=>"110100110",
  40211=>"000010111",
  40212=>"010011101",
  40213=>"101110000",
  40214=>"010101100",
  40215=>"101000000",
  40216=>"000100100",
  40217=>"100110000",
  40218=>"100110001",
  40219=>"110111110",
  40220=>"000010110",
  40221=>"111101001",
  40222=>"101000010",
  40223=>"011010001",
  40224=>"101010010",
  40225=>"011110110",
  40226=>"000101111",
  40227=>"110010101",
  40228=>"001110000",
  40229=>"101101110",
  40230=>"101010000",
  40231=>"100101000",
  40232=>"110101100",
  40233=>"010000010",
  40234=>"111001110",
  40235=>"010110101",
  40236=>"011011010",
  40237=>"000101001",
  40238=>"011111010",
  40239=>"001100101",
  40240=>"000011011",
  40241=>"101101010",
  40242=>"111101001",
  40243=>"110101001",
  40244=>"100110110",
  40245=>"010011000",
  40246=>"110100101",
  40247=>"101001000",
  40248=>"011000001",
  40249=>"001000111",
  40250=>"111100001",
  40251=>"101101010",
  40252=>"000011101",
  40253=>"100100110",
  40254=>"011111100",
  40255=>"011010100",
  40256=>"000110000",
  40257=>"001111001",
  40258=>"011000100",
  40259=>"000000100",
  40260=>"001010000",
  40261=>"011101111",
  40262=>"100000011",
  40263=>"100011110",
  40264=>"000100110",
  40265=>"101100101",
  40266=>"010101000",
  40267=>"001000000",
  40268=>"110010101",
  40269=>"010101010",
  40270=>"101110111",
  40271=>"101010010",
  40272=>"110010111",
  40273=>"010001100",
  40274=>"101111011",
  40275=>"011110000",
  40276=>"001011010",
  40277=>"010010000",
  40278=>"010111111",
  40279=>"011100100",
  40280=>"011011001",
  40281=>"101000000",
  40282=>"001100011",
  40283=>"100101101",
  40284=>"011010111",
  40285=>"000100101",
  40286=>"000101001",
  40287=>"010100110",
  40288=>"100110100",
  40289=>"110101110",
  40290=>"110010111",
  40291=>"111000000",
  40292=>"011111000",
  40293=>"001111111",
  40294=>"000011010",
  40295=>"010100011",
  40296=>"100100110",
  40297=>"000111001",
  40298=>"101101011",
  40299=>"001011010",
  40300=>"111111111",
  40301=>"100101001",
  40302=>"110111101",
  40303=>"011000100",
  40304=>"100110111",
  40305=>"010100000",
  40306=>"111100110",
  40307=>"111101001",
  40308=>"110000011",
  40309=>"100000010",
  40310=>"001110011",
  40311=>"101011011",
  40312=>"001110010",
  40313=>"000110100",
  40314=>"001010111",
  40315=>"101001101",
  40316=>"000111110",
  40317=>"100011011",
  40318=>"010111111",
  40319=>"010111100",
  40320=>"100100110",
  40321=>"111011001",
  40322=>"111010011",
  40323=>"111000001",
  40324=>"100101110",
  40325=>"110000010",
  40326=>"001110001",
  40327=>"101101101",
  40328=>"010000011",
  40329=>"110101111",
  40330=>"101000110",
  40331=>"100000001",
  40332=>"101011001",
  40333=>"010111110",
  40334=>"111111000",
  40335=>"010101111",
  40336=>"001101000",
  40337=>"011000100",
  40338=>"100111011",
  40339=>"100000001",
  40340=>"000111010",
  40341=>"001101111",
  40342=>"000011111",
  40343=>"000101110",
  40344=>"111000110",
  40345=>"001001001",
  40346=>"010011011",
  40347=>"111110111",
  40348=>"000111001",
  40349=>"111010110",
  40350=>"011110001",
  40351=>"110010000",
  40352=>"100101000",
  40353=>"110000011",
  40354=>"100011010",
  40355=>"100001101",
  40356=>"010100100",
  40357=>"111000101",
  40358=>"011101010",
  40359=>"100111100",
  40360=>"010001010",
  40361=>"000010000",
  40362=>"110100101",
  40363=>"100101000",
  40364=>"011010110",
  40365=>"101010101",
  40366=>"101111101",
  40367=>"100111110",
  40368=>"111101110",
  40369=>"101111011",
  40370=>"101111110",
  40371=>"000001101",
  40372=>"110110101",
  40373=>"110101100",
  40374=>"010100111",
  40375=>"111100101",
  40376=>"010101100",
  40377=>"000100101",
  40378=>"010101010",
  40379=>"100110100",
  40380=>"101101010",
  40381=>"110000100",
  40382=>"000100101",
  40383=>"101010110",
  40384=>"110100010",
  40385=>"010001110",
  40386=>"110110100",
  40387=>"110111000",
  40388=>"100101110",
  40389=>"110101011",
  40390=>"001011111",
  40391=>"101101000",
  40392=>"001001011",
  40393=>"001000010",
  40394=>"100010111",
  40395=>"110000101",
  40396=>"011001001",
  40397=>"001001011",
  40398=>"101100100",
  40399=>"101110110",
  40400=>"010101000",
  40401=>"011010100",
  40402=>"111001110",
  40403=>"000010110",
  40404=>"111100110",
  40405=>"110011111",
  40406=>"100100010",
  40407=>"001001001",
  40408=>"010001000",
  40409=>"101100100",
  40410=>"010001010",
  40411=>"110001111",
  40412=>"101110011",
  40413=>"100010001",
  40414=>"111000101",
  40415=>"000111101",
  40416=>"010001101",
  40417=>"010111111",
  40418=>"110010110",
  40419=>"110010010",
  40420=>"010111100",
  40421=>"011100110",
  40422=>"010010110",
  40423=>"110001000",
  40424=>"000010001",
  40425=>"000000000",
  40426=>"110100011",
  40427=>"000110011",
  40428=>"011111011",
  40429=>"100110001",
  40430=>"101101100",
  40431=>"001101000",
  40432=>"011001100",
  40433=>"111001101",
  40434=>"110010001",
  40435=>"111100100",
  40436=>"110101110",
  40437=>"110100000",
  40438=>"111011011",
  40439=>"101111011",
  40440=>"110100010",
  40441=>"100111001",
  40442=>"100001001",
  40443=>"011000110",
  40444=>"110101010",
  40445=>"110001101",
  40446=>"100011111",
  40447=>"110010000",
  40448=>"111011100",
  40449=>"000010011",
  40450=>"100001111",
  40451=>"000000000",
  40452=>"010001101",
  40453=>"111000001",
  40454=>"101001111",
  40455=>"100011110",
  40456=>"011100011",
  40457=>"110010101",
  40458=>"010010011",
  40459=>"011010111",
  40460=>"011001011",
  40461=>"001101101",
  40462=>"101001000",
  40463=>"110111000",
  40464=>"111011101",
  40465=>"101010110",
  40466=>"000011001",
  40467=>"011010011",
  40468=>"111000101",
  40469=>"101011010",
  40470=>"010110100",
  40471=>"101001000",
  40472=>"001001100",
  40473=>"011001011",
  40474=>"010001001",
  40475=>"111010110",
  40476=>"000010000",
  40477=>"010011001",
  40478=>"101000100",
  40479=>"010001110",
  40480=>"111101100",
  40481=>"000011101",
  40482=>"001001101",
  40483=>"010100101",
  40484=>"111000101",
  40485=>"001101100",
  40486=>"010011100",
  40487=>"110010101",
  40488=>"111110101",
  40489=>"101110100",
  40490=>"110110110",
  40491=>"110000101",
  40492=>"010001001",
  40493=>"100111011",
  40494=>"100000101",
  40495=>"101101010",
  40496=>"101111101",
  40497=>"110111010",
  40498=>"101001100",
  40499=>"100000111",
  40500=>"111000110",
  40501=>"111000001",
  40502=>"001001000",
  40503=>"101000110",
  40504=>"001001010",
  40505=>"111110110",
  40506=>"001011010",
  40507=>"110111100",
  40508=>"100100001",
  40509=>"101110000",
  40510=>"100101011",
  40511=>"111100100",
  40512=>"011000100",
  40513=>"100000001",
  40514=>"101010111",
  40515=>"010011111",
  40516=>"011011010",
  40517=>"100010100",
  40518=>"111011001",
  40519=>"011111000",
  40520=>"000011011",
  40521=>"100100101",
  40522=>"011100101",
  40523=>"001010101",
  40524=>"001000100",
  40525=>"111100111",
  40526=>"011010101",
  40527=>"111100011",
  40528=>"001010000",
  40529=>"000110111",
  40530=>"011101000",
  40531=>"101010001",
  40532=>"111000111",
  40533=>"100100001",
  40534=>"001001001",
  40535=>"011001111",
  40536=>"101100001",
  40537=>"010101011",
  40538=>"010000001",
  40539=>"100101110",
  40540=>"111101001",
  40541=>"110100100",
  40542=>"101011101",
  40543=>"011110011",
  40544=>"011111101",
  40545=>"110011100",
  40546=>"000110000",
  40547=>"101001000",
  40548=>"100100100",
  40549=>"110111110",
  40550=>"001101111",
  40551=>"011111001",
  40552=>"001110101",
  40553=>"000101011",
  40554=>"000110001",
  40555=>"100010001",
  40556=>"100000001",
  40557=>"001001011",
  40558=>"011010010",
  40559=>"110101100",
  40560=>"100101001",
  40561=>"011101100",
  40562=>"110110001",
  40563=>"110011001",
  40564=>"110110110",
  40565=>"100100001",
  40566=>"111101011",
  40567=>"100101011",
  40568=>"011000100",
  40569=>"101100110",
  40570=>"011111110",
  40571=>"111101101",
  40572=>"001010100",
  40573=>"010011001",
  40574=>"110100000",
  40575=>"111101001",
  40576=>"000011001",
  40577=>"110010101",
  40578=>"001000000",
  40579=>"101000101",
  40580=>"111001011",
  40581=>"110100000",
  40582=>"100011111",
  40583=>"100100000",
  40584=>"111110100",
  40585=>"010001101",
  40586=>"001000110",
  40587=>"111101100",
  40588=>"011001011",
  40589=>"001001001",
  40590=>"101010100",
  40591=>"101100111",
  40592=>"100000010",
  40593=>"101110110",
  40594=>"110000001",
  40595=>"110000111",
  40596=>"100010010",
  40597=>"011011111",
  40598=>"001110001",
  40599=>"111011101",
  40600=>"100000111",
  40601=>"101011111",
  40602=>"011001011",
  40603=>"001100000",
  40604=>"101110001",
  40605=>"110100010",
  40606=>"010011111",
  40607=>"001010010",
  40608=>"110110000",
  40609=>"010101101",
  40610=>"001001011",
  40611=>"000010000",
  40612=>"000100101",
  40613=>"100110011",
  40614=>"110100000",
  40615=>"111101110",
  40616=>"111101111",
  40617=>"000100000",
  40618=>"101011111",
  40619=>"001100010",
  40620=>"001000100",
  40621=>"110001001",
  40622=>"100011111",
  40623=>"101110111",
  40624=>"000001000",
  40625=>"010100001",
  40626=>"001011110",
  40627=>"010010001",
  40628=>"000111110",
  40629=>"001001101",
  40630=>"000111111",
  40631=>"101010010",
  40632=>"001100000",
  40633=>"011100001",
  40634=>"000100001",
  40635=>"110001101",
  40636=>"110010000",
  40637=>"111001111",
  40638=>"011001000",
  40639=>"101100110",
  40640=>"111001101",
  40641=>"011010111",
  40642=>"100001111",
  40643=>"001100101",
  40644=>"001000110",
  40645=>"010110110",
  40646=>"111010110",
  40647=>"001001000",
  40648=>"111111111",
  40649=>"000010001",
  40650=>"110001101",
  40651=>"001001101",
  40652=>"100100010",
  40653=>"001001101",
  40654=>"010001111",
  40655=>"100000001",
  40656=>"101001011",
  40657=>"101111111",
  40658=>"001010100",
  40659=>"100001000",
  40660=>"110100011",
  40661=>"001101001",
  40662=>"011100010",
  40663=>"111000011",
  40664=>"010111111",
  40665=>"010110110",
  40666=>"110011111",
  40667=>"100110000",
  40668=>"101001001",
  40669=>"110000001",
  40670=>"001011010",
  40671=>"111110111",
  40672=>"001010101",
  40673=>"110101100",
  40674=>"100010111",
  40675=>"010111001",
  40676=>"001011010",
  40677=>"001111001",
  40678=>"010101010",
  40679=>"111001111",
  40680=>"101101001",
  40681=>"101011011",
  40682=>"110010011",
  40683=>"010110001",
  40684=>"001000001",
  40685=>"111111000",
  40686=>"101001101",
  40687=>"000100001",
  40688=>"100100011",
  40689=>"101110101",
  40690=>"001000010",
  40691=>"101101001",
  40692=>"100101111",
  40693=>"100010100",
  40694=>"000101000",
  40695=>"111100010",
  40696=>"010111111",
  40697=>"111010011",
  40698=>"010111110",
  40699=>"110101010",
  40700=>"011011111",
  40701=>"000010100",
  40702=>"011101001",
  40703=>"111000000",
  40704=>"101010111",
  40705=>"000100101",
  40706=>"110001011",
  40707=>"110110111",
  40708=>"100111111",
  40709=>"100101110",
  40710=>"011011000",
  40711=>"101010100",
  40712=>"111010111",
  40713=>"000000010",
  40714=>"110101111",
  40715=>"010010001",
  40716=>"010011101",
  40717=>"010010111",
  40718=>"101000110",
  40719=>"110100110",
  40720=>"101001110",
  40721=>"111011100",
  40722=>"011000101",
  40723=>"110101001",
  40724=>"011100001",
  40725=>"011011000",
  40726=>"110010100",
  40727=>"111011000",
  40728=>"001101111",
  40729=>"010000110",
  40730=>"000011010",
  40731=>"101100110",
  40732=>"100001100",
  40733=>"001000100",
  40734=>"111101101",
  40735=>"000100010",
  40736=>"111011110",
  40737=>"001000000",
  40738=>"000001000",
  40739=>"001101000",
  40740=>"000001110",
  40741=>"100001000",
  40742=>"000000000",
  40743=>"111011110",
  40744=>"001000001",
  40745=>"011010000",
  40746=>"110101010",
  40747=>"000001101",
  40748=>"010111110",
  40749=>"100101000",
  40750=>"001001100",
  40751=>"110110110",
  40752=>"110100101",
  40753=>"000000001",
  40754=>"000011011",
  40755=>"111001000",
  40756=>"001011000",
  40757=>"111111111",
  40758=>"101001100",
  40759=>"110101010",
  40760=>"001100111",
  40761=>"100100101",
  40762=>"101011011",
  40763=>"101011111",
  40764=>"101100100",
  40765=>"000101110",
  40766=>"010111011",
  40767=>"010011101",
  40768=>"100100001",
  40769=>"110010011",
  40770=>"101101100",
  40771=>"111010001",
  40772=>"111101110",
  40773=>"000110110",
  40774=>"001100000",
  40775=>"010100100",
  40776=>"001100111",
  40777=>"100001111",
  40778=>"000011101",
  40779=>"001001001",
  40780=>"011010101",
  40781=>"101001101",
  40782=>"101000111",
  40783=>"010000011",
  40784=>"010100011",
  40785=>"100100011",
  40786=>"101011111",
  40787=>"110000111",
  40788=>"100100110",
  40789=>"101100000",
  40790=>"011001010",
  40791=>"110010010",
  40792=>"100100110",
  40793=>"011010010",
  40794=>"010001000",
  40795=>"111001001",
  40796=>"100011010",
  40797=>"100101100",
  40798=>"011000101",
  40799=>"001010111",
  40800=>"000101111",
  40801=>"110011100",
  40802=>"001101110",
  40803=>"100011111",
  40804=>"011111110",
  40805=>"110110001",
  40806=>"111001011",
  40807=>"111010100",
  40808=>"101011010",
  40809=>"100100000",
  40810=>"000111000",
  40811=>"111001011",
  40812=>"110111010",
  40813=>"101001011",
  40814=>"101000101",
  40815=>"100010110",
  40816=>"001101001",
  40817=>"111010111",
  40818=>"001110100",
  40819=>"011010011",
  40820=>"111111101",
  40821=>"100101101",
  40822=>"001101100",
  40823=>"110000001",
  40824=>"111010000",
  40825=>"010101111",
  40826=>"100001010",
  40827=>"111001001",
  40828=>"001111001",
  40829=>"101111000",
  40830=>"000010001",
  40831=>"110111001",
  40832=>"100101010",
  40833=>"010011111",
  40834=>"010000011",
  40835=>"100101011",
  40836=>"100000000",
  40837=>"101010011",
  40838=>"111100100",
  40839=>"000100100",
  40840=>"011011100",
  40841=>"011001000",
  40842=>"011101110",
  40843=>"110111101",
  40844=>"111100101",
  40845=>"001111011",
  40846=>"100110010",
  40847=>"100100100",
  40848=>"101101110",
  40849=>"000010110",
  40850=>"111111000",
  40851=>"110110101",
  40852=>"111111011",
  40853=>"010110000",
  40854=>"010000001",
  40855=>"011000100",
  40856=>"000101001",
  40857=>"100001000",
  40858=>"010000111",
  40859=>"101010011",
  40860=>"101001100",
  40861=>"111001000",
  40862=>"011110110",
  40863=>"000100010",
  40864=>"110011010",
  40865=>"100011001",
  40866=>"101101110",
  40867=>"111001101",
  40868=>"100101100",
  40869=>"101100001",
  40870=>"011010010",
  40871=>"110111101",
  40872=>"101011101",
  40873=>"111110100",
  40874=>"000101110",
  40875=>"010100100",
  40876=>"101001100",
  40877=>"010110101",
  40878=>"000011100",
  40879=>"001011000",
  40880=>"111001110",
  40881=>"001011010",
  40882=>"011011101",
  40883=>"001001000",
  40884=>"111100101",
  40885=>"000011010",
  40886=>"111111111",
  40887=>"110101100",
  40888=>"100011101",
  40889=>"000001111",
  40890=>"010011011",
  40891=>"000011100",
  40892=>"111000111",
  40893=>"110101101",
  40894=>"010001001",
  40895=>"001101110",
  40896=>"101001101",
  40897=>"101110110",
  40898=>"001010000",
  40899=>"011010101",
  40900=>"100100010",
  40901=>"011100011",
  40902=>"111111100",
  40903=>"110010100",
  40904=>"000001100",
  40905=>"001111101",
  40906=>"010110100",
  40907=>"100000101",
  40908=>"011100011",
  40909=>"110001101",
  40910=>"000100100",
  40911=>"010100111",
  40912=>"001100111",
  40913=>"100110110",
  40914=>"001100101",
  40915=>"001101101",
  40916=>"010111110",
  40917=>"101010101",
  40918=>"010001101",
  40919=>"111101100",
  40920=>"001011101",
  40921=>"100100011",
  40922=>"111111001",
  40923=>"001011011",
  40924=>"101001100",
  40925=>"000111111",
  40926=>"011111100",
  40927=>"100101111",
  40928=>"001101011",
  40929=>"010111011",
  40930=>"101001011",
  40931=>"100011010",
  40932=>"011110100",
  40933=>"100011010",
  40934=>"111111010",
  40935=>"100001011",
  40936=>"111111100",
  40937=>"001001010",
  40938=>"110110100",
  40939=>"000111111",
  40940=>"001010010",
  40941=>"100100101",
  40942=>"000001000",
  40943=>"010010001",
  40944=>"001111111",
  40945=>"010010001",
  40946=>"001100110",
  40947=>"001101101",
  40948=>"010100001",
  40949=>"101010000",
  40950=>"110010101",
  40951=>"010000101",
  40952=>"101111101",
  40953=>"110101001",
  40954=>"001111100",
  40955=>"010001110",
  40956=>"101011111",
  40957=>"110100000",
  40958=>"010000101",
  40959=>"101011001",
  40960=>"111101011",
  40961=>"000110010",
  40962=>"001101111",
  40963=>"110000000",
  40964=>"011000001",
  40965=>"000111001",
  40966=>"001110001",
  40967=>"011110111",
  40968=>"111101110",
  40969=>"010010110",
  40970=>"000000101",
  40971=>"101001111",
  40972=>"101110111",
  40973=>"110010101",
  40974=>"111110010",
  40975=>"010000111",
  40976=>"111010010",
  40977=>"000000111",
  40978=>"101010011",
  40979=>"110000001",
  40980=>"000110011",
  40981=>"110011001",
  40982=>"011000011",
  40983=>"010001001",
  40984=>"010000111",
  40985=>"011011101",
  40986=>"100110111",
  40987=>"000111011",
  40988=>"100011011",
  40989=>"001000111",
  40990=>"001001001",
  40991=>"100010111",
  40992=>"010100110",
  40993=>"100100011",
  40994=>"011100001",
  40995=>"111111110",
  40996=>"001000100",
  40997=>"011111110",
  40998=>"010011001",
  40999=>"111110111",
  41000=>"001001001",
  41001=>"100100001",
  41002=>"101101100",
  41003=>"110100001",
  41004=>"101000010",
  41005=>"111010000",
  41006=>"010110101",
  41007=>"111110110",
  41008=>"100010111",
  41009=>"000100010",
  41010=>"101000001",
  41011=>"010100100",
  41012=>"011111000",
  41013=>"110001000",
  41014=>"100010111",
  41015=>"011110111",
  41016=>"100101011",
  41017=>"100111000",
  41018=>"110001111",
  41019=>"000000101",
  41020=>"000000111",
  41021=>"000110010",
  41022=>"000101111",
  41023=>"100110100",
  41024=>"110101110",
  41025=>"111000010",
  41026=>"011011001",
  41027=>"111110100",
  41028=>"001111111",
  41029=>"101101100",
  41030=>"111001010",
  41031=>"011100011",
  41032=>"000010011",
  41033=>"100001111",
  41034=>"101110110",
  41035=>"001111111",
  41036=>"010011011",
  41037=>"110100100",
  41038=>"111010101",
  41039=>"101011110",
  41040=>"010001101",
  41041=>"111111111",
  41042=>"010011100",
  41043=>"011111100",
  41044=>"110110001",
  41045=>"100100110",
  41046=>"100011100",
  41047=>"001000111",
  41048=>"100001000",
  41049=>"000101000",
  41050=>"111011100",
  41051=>"010000100",
  41052=>"001000100",
  41053=>"100100001",
  41054=>"011001010",
  41055=>"101101110",
  41056=>"010001111",
  41057=>"101100110",
  41058=>"000110011",
  41059=>"001000010",
  41060=>"011001000",
  41061=>"011101111",
  41062=>"010001100",
  41063=>"000101010",
  41064=>"010001000",
  41065=>"001011011",
  41066=>"010000010",
  41067=>"000001010",
  41068=>"001110011",
  41069=>"100000101",
  41070=>"100001110",
  41071=>"010100000",
  41072=>"101001010",
  41073=>"001101011",
  41074=>"100110110",
  41075=>"001111001",
  41076=>"000011010",
  41077=>"110110110",
  41078=>"111001111",
  41079=>"010000110",
  41080=>"111100000",
  41081=>"111111011",
  41082=>"110011010",
  41083=>"111100001",
  41084=>"101111110",
  41085=>"110000001",
  41086=>"011011101",
  41087=>"111010110",
  41088=>"001111111",
  41089=>"111101100",
  41090=>"000010110",
  41091=>"001000011",
  41092=>"111011101",
  41093=>"101101000",
  41094=>"111111110",
  41095=>"101111111",
  41096=>"010100001",
  41097=>"010100001",
  41098=>"111101110",
  41099=>"010011010",
  41100=>"110110011",
  41101=>"011010101",
  41102=>"101110010",
  41103=>"011010100",
  41104=>"001110011",
  41105=>"010101010",
  41106=>"101101101",
  41107=>"100101101",
  41108=>"000011111",
  41109=>"011001111",
  41110=>"000011011",
  41111=>"111011110",
  41112=>"000001010",
  41113=>"111101101",
  41114=>"011010110",
  41115=>"111100001",
  41116=>"010001011",
  41117=>"000110110",
  41118=>"010011001",
  41119=>"010101011",
  41120=>"011010010",
  41121=>"100111010",
  41122=>"111111111",
  41123=>"110000011",
  41124=>"100101000",
  41125=>"100001011",
  41126=>"110100111",
  41127=>"001010111",
  41128=>"011110101",
  41129=>"011010101",
  41130=>"111111111",
  41131=>"101110110",
  41132=>"100011000",
  41133=>"101000000",
  41134=>"010001100",
  41135=>"110000110",
  41136=>"101011010",
  41137=>"010101000",
  41138=>"111110101",
  41139=>"110000110",
  41140=>"010100000",
  41141=>"001100010",
  41142=>"000000001",
  41143=>"000000000",
  41144=>"100001001",
  41145=>"101011110",
  41146=>"011000110",
  41147=>"111010111",
  41148=>"010011110",
  41149=>"100010110",
  41150=>"011101000",
  41151=>"010101000",
  41152=>"000000100",
  41153=>"101100111",
  41154=>"001111001",
  41155=>"010011001",
  41156=>"110100101",
  41157=>"111011010",
  41158=>"110111011",
  41159=>"101110100",
  41160=>"011110010",
  41161=>"011010110",
  41162=>"111010100",
  41163=>"111000101",
  41164=>"001111010",
  41165=>"101000101",
  41166=>"011011101",
  41167=>"001000111",
  41168=>"101100100",
  41169=>"101100100",
  41170=>"000010011",
  41171=>"111101000",
  41172=>"010101001",
  41173=>"110101110",
  41174=>"011100011",
  41175=>"011000001",
  41176=>"100110001",
  41177=>"000110001",
  41178=>"000010101",
  41179=>"001000110",
  41180=>"101001010",
  41181=>"111000100",
  41182=>"001010110",
  41183=>"000000110",
  41184=>"001100011",
  41185=>"100110001",
  41186=>"001001000",
  41187=>"000101000",
  41188=>"010001011",
  41189=>"011110100",
  41190=>"111111011",
  41191=>"101011111",
  41192=>"111010110",
  41193=>"000111011",
  41194=>"011101110",
  41195=>"000000100",
  41196=>"000001101",
  41197=>"010011110",
  41198=>"111100111",
  41199=>"001000011",
  41200=>"001110000",
  41201=>"010101000",
  41202=>"000101111",
  41203=>"011111110",
  41204=>"010000100",
  41205=>"001111110",
  41206=>"101001101",
  41207=>"101011100",
  41208=>"101101010",
  41209=>"111101110",
  41210=>"110001001",
  41211=>"100000101",
  41212=>"111000101",
  41213=>"110101000",
  41214=>"110001100",
  41215=>"111101010",
  41216=>"110000101",
  41217=>"101101110",
  41218=>"111011100",
  41219=>"001000001",
  41220=>"110000011",
  41221=>"110010010",
  41222=>"100001111",
  41223=>"100001100",
  41224=>"000100011",
  41225=>"110111011",
  41226=>"110111101",
  41227=>"110001110",
  41228=>"101001110",
  41229=>"111011010",
  41230=>"111111111",
  41231=>"001011000",
  41232=>"101011111",
  41233=>"101000111",
  41234=>"111001110",
  41235=>"000101100",
  41236=>"000011101",
  41237=>"111100011",
  41238=>"100000111",
  41239=>"101110000",
  41240=>"000101110",
  41241=>"011010010",
  41242=>"110001001",
  41243=>"001011111",
  41244=>"000110111",
  41245=>"101010101",
  41246=>"100010111",
  41247=>"000000100",
  41248=>"100110001",
  41249=>"000001110",
  41250=>"110111010",
  41251=>"111101011",
  41252=>"001010011",
  41253=>"110110011",
  41254=>"000101001",
  41255=>"001101101",
  41256=>"011111010",
  41257=>"011000010",
  41258=>"100100000",
  41259=>"010011100",
  41260=>"110101001",
  41261=>"101101010",
  41262=>"000001011",
  41263=>"100111011",
  41264=>"000010101",
  41265=>"000110010",
  41266=>"001100100",
  41267=>"000011010",
  41268=>"011100110",
  41269=>"110110010",
  41270=>"001010000",
  41271=>"100001000",
  41272=>"111101110",
  41273=>"011000010",
  41274=>"110111010",
  41275=>"000000000",
  41276=>"101110101",
  41277=>"100011111",
  41278=>"101101010",
  41279=>"001111100",
  41280=>"001101101",
  41281=>"101110110",
  41282=>"100110001",
  41283=>"010011101",
  41284=>"100001010",
  41285=>"010101111",
  41286=>"000101011",
  41287=>"101000110",
  41288=>"011100110",
  41289=>"100110010",
  41290=>"011110100",
  41291=>"101111101",
  41292=>"101000010",
  41293=>"011111011",
  41294=>"000000010",
  41295=>"011110110",
  41296=>"010000110",
  41297=>"101000010",
  41298=>"100111110",
  41299=>"001101100",
  41300=>"000010100",
  41301=>"100001000",
  41302=>"100010101",
  41303=>"101001001",
  41304=>"001100000",
  41305=>"000000001",
  41306=>"110001101",
  41307=>"110011010",
  41308=>"101000100",
  41309=>"011101010",
  41310=>"110010100",
  41311=>"001100010",
  41312=>"011110011",
  41313=>"010000111",
  41314=>"100111100",
  41315=>"001101010",
  41316=>"001101001",
  41317=>"100110111",
  41318=>"110100111",
  41319=>"000000001",
  41320=>"110010000",
  41321=>"100100100",
  41322=>"011111010",
  41323=>"001001110",
  41324=>"000101110",
  41325=>"011000111",
  41326=>"011111001",
  41327=>"110101111",
  41328=>"001111111",
  41329=>"111010101",
  41330=>"100010110",
  41331=>"001001101",
  41332=>"101000101",
  41333=>"101110111",
  41334=>"101001000",
  41335=>"100011101",
  41336=>"110110111",
  41337=>"111111010",
  41338=>"111010010",
  41339=>"010011001",
  41340=>"010001110",
  41341=>"011001110",
  41342=>"101000011",
  41343=>"111001001",
  41344=>"110001100",
  41345=>"101101000",
  41346=>"011101101",
  41347=>"000000000",
  41348=>"001011110",
  41349=>"101001000",
  41350=>"110110100",
  41351=>"101111110",
  41352=>"101001000",
  41353=>"111000100",
  41354=>"100001011",
  41355=>"001100000",
  41356=>"001110001",
  41357=>"010000101",
  41358=>"100100001",
  41359=>"000111111",
  41360=>"011010000",
  41361=>"101010001",
  41362=>"111011000",
  41363=>"001111010",
  41364=>"000010010",
  41365=>"001000011",
  41366=>"101111100",
  41367=>"010010111",
  41368=>"011000101",
  41369=>"001000111",
  41370=>"000110001",
  41371=>"110100000",
  41372=>"001001001",
  41373=>"011000110",
  41374=>"100100011",
  41375=>"110010110",
  41376=>"101101000",
  41377=>"111100000",
  41378=>"011101000",
  41379=>"101000110",
  41380=>"000011100",
  41381=>"100010100",
  41382=>"101110111",
  41383=>"111011000",
  41384=>"110111110",
  41385=>"111011001",
  41386=>"010010110",
  41387=>"000110011",
  41388=>"000010010",
  41389=>"111101011",
  41390=>"010101100",
  41391=>"111111110",
  41392=>"000100110",
  41393=>"101100101",
  41394=>"111111110",
  41395=>"000000001",
  41396=>"010110001",
  41397=>"111101110",
  41398=>"111010000",
  41399=>"111010011",
  41400=>"010011100",
  41401=>"000110100",
  41402=>"011111010",
  41403=>"111100100",
  41404=>"100001000",
  41405=>"111010010",
  41406=>"011101011",
  41407=>"100010110",
  41408=>"011101111",
  41409=>"100110011",
  41410=>"101100100",
  41411=>"111010101",
  41412=>"110101001",
  41413=>"111101100",
  41414=>"011010000",
  41415=>"111100001",
  41416=>"101100011",
  41417=>"111111001",
  41418=>"001101000",
  41419=>"100100110",
  41420=>"000110100",
  41421=>"100000011",
  41422=>"111111000",
  41423=>"110010000",
  41424=>"101100011",
  41425=>"110001110",
  41426=>"010111111",
  41427=>"000111011",
  41428=>"000011010",
  41429=>"011001110",
  41430=>"110110110",
  41431=>"000000011",
  41432=>"101010100",
  41433=>"100101111",
  41434=>"001111110",
  41435=>"111110101",
  41436=>"111001001",
  41437=>"101001111",
  41438=>"111111101",
  41439=>"111010001",
  41440=>"101110101",
  41441=>"000101010",
  41442=>"111001110",
  41443=>"100110110",
  41444=>"100001101",
  41445=>"111111111",
  41446=>"001101111",
  41447=>"101111100",
  41448=>"110000001",
  41449=>"110101000",
  41450=>"000101011",
  41451=>"011010101",
  41452=>"010100101",
  41453=>"001010011",
  41454=>"000100000",
  41455=>"000000001",
  41456=>"111000001",
  41457=>"110000101",
  41458=>"000011010",
  41459=>"001001101",
  41460=>"000111010",
  41461=>"111011000",
  41462=>"000110110",
  41463=>"010001010",
  41464=>"001111010",
  41465=>"000011011",
  41466=>"101111101",
  41467=>"010001111",
  41468=>"000000001",
  41469=>"010000101",
  41470=>"010100111",
  41471=>"001111110",
  41472=>"100110010",
  41473=>"011010101",
  41474=>"100010111",
  41475=>"111111001",
  41476=>"111100000",
  41477=>"110111010",
  41478=>"011101010",
  41479=>"010010110",
  41480=>"011001110",
  41481=>"010111001",
  41482=>"011010110",
  41483=>"010111001",
  41484=>"101000011",
  41485=>"001100010",
  41486=>"010010110",
  41487=>"010110011",
  41488=>"101000001",
  41489=>"110011101",
  41490=>"100100000",
  41491=>"100010001",
  41492=>"001110000",
  41493=>"011100010",
  41494=>"100111101",
  41495=>"011110110",
  41496=>"110101111",
  41497=>"101111011",
  41498=>"111010111",
  41499=>"001011101",
  41500=>"000011010",
  41501=>"000010000",
  41502=>"111101010",
  41503=>"101111011",
  41504=>"010100010",
  41505=>"101110011",
  41506=>"000100010",
  41507=>"111110111",
  41508=>"000010011",
  41509=>"001111001",
  41510=>"011110010",
  41511=>"110100100",
  41512=>"000100011",
  41513=>"011000101",
  41514=>"101011111",
  41515=>"110011001",
  41516=>"010111101",
  41517=>"111110011",
  41518=>"101010001",
  41519=>"000101000",
  41520=>"011100111",
  41521=>"101111101",
  41522=>"101001101",
  41523=>"010010110",
  41524=>"001001101",
  41525=>"100001000",
  41526=>"010101101",
  41527=>"010001101",
  41528=>"000011000",
  41529=>"101000000",
  41530=>"010001100",
  41531=>"000000010",
  41532=>"110000111",
  41533=>"100101110",
  41534=>"101101010",
  41535=>"011010100",
  41536=>"011000001",
  41537=>"011010011",
  41538=>"110100001",
  41539=>"100101000",
  41540=>"000100110",
  41541=>"111010000",
  41542=>"101101110",
  41543=>"111111110",
  41544=>"100100110",
  41545=>"100010000",
  41546=>"001110110",
  41547=>"101010011",
  41548=>"100111110",
  41549=>"011111001",
  41550=>"101101100",
  41551=>"010101010",
  41552=>"111011111",
  41553=>"111000100",
  41554=>"010110111",
  41555=>"101110100",
  41556=>"011111010",
  41557=>"000100000",
  41558=>"001001011",
  41559=>"001110010",
  41560=>"000001100",
  41561=>"011001111",
  41562=>"101000000",
  41563=>"000111000",
  41564=>"001101110",
  41565=>"001101000",
  41566=>"101100000",
  41567=>"011100101",
  41568=>"011000010",
  41569=>"001010001",
  41570=>"000101001",
  41571=>"111010110",
  41572=>"010010001",
  41573=>"100010111",
  41574=>"101101100",
  41575=>"111011000",
  41576=>"100100011",
  41577=>"100110000",
  41578=>"111111100",
  41579=>"011000000",
  41580=>"000000110",
  41581=>"010000000",
  41582=>"110110001",
  41583=>"100111011",
  41584=>"100110101",
  41585=>"000101011",
  41586=>"101010111",
  41587=>"110001110",
  41588=>"011100010",
  41589=>"010100101",
  41590=>"111010010",
  41591=>"011010010",
  41592=>"010110111",
  41593=>"101101010",
  41594=>"000001011",
  41595=>"010110001",
  41596=>"010110110",
  41597=>"010010001",
  41598=>"000111111",
  41599=>"110110011",
  41600=>"100000011",
  41601=>"110010010",
  41602=>"101100100",
  41603=>"100101011",
  41604=>"010000000",
  41605=>"101100100",
  41606=>"001100111",
  41607=>"000100010",
  41608=>"101101010",
  41609=>"100010101",
  41610=>"101011110",
  41611=>"111001101",
  41612=>"011000111",
  41613=>"000101000",
  41614=>"111000101",
  41615=>"001011100",
  41616=>"001011011",
  41617=>"010010000",
  41618=>"111100111",
  41619=>"001011111",
  41620=>"101101110",
  41621=>"000110000",
  41622=>"101100111",
  41623=>"000100101",
  41624=>"010000110",
  41625=>"100001111",
  41626=>"111000001",
  41627=>"010100011",
  41628=>"010111011",
  41629=>"100100000",
  41630=>"010101000",
  41631=>"001100001",
  41632=>"110100011",
  41633=>"001011100",
  41634=>"101110100",
  41635=>"001110011",
  41636=>"101011101",
  41637=>"110011110",
  41638=>"100001001",
  41639=>"000011110",
  41640=>"011010010",
  41641=>"001000000",
  41642=>"111100000",
  41643=>"111011111",
  41644=>"000011000",
  41645=>"001000010",
  41646=>"010000111",
  41647=>"000101010",
  41648=>"001111011",
  41649=>"110000111",
  41650=>"100111100",
  41651=>"100110011",
  41652=>"100100001",
  41653=>"000010111",
  41654=>"001010000",
  41655=>"011011101",
  41656=>"010100100",
  41657=>"001100111",
  41658=>"000010101",
  41659=>"100101101",
  41660=>"010001000",
  41661=>"010110000",
  41662=>"001100001",
  41663=>"101111111",
  41664=>"011101111",
  41665=>"000100100",
  41666=>"101001110",
  41667=>"010110110",
  41668=>"000111111",
  41669=>"000000000",
  41670=>"010001111",
  41671=>"000111011",
  41672=>"100101001",
  41673=>"111011001",
  41674=>"101100101",
  41675=>"100000111",
  41676=>"000001000",
  41677=>"100001010",
  41678=>"010001101",
  41679=>"110101101",
  41680=>"100001111",
  41681=>"011100101",
  41682=>"001101011",
  41683=>"110111111",
  41684=>"010000110",
  41685=>"010111010",
  41686=>"101111110",
  41687=>"001000011",
  41688=>"110110101",
  41689=>"011001011",
  41690=>"010000000",
  41691=>"001101001",
  41692=>"001001101",
  41693=>"111000110",
  41694=>"101100111",
  41695=>"111111111",
  41696=>"001111001",
  41697=>"101001000",
  41698=>"110000101",
  41699=>"010111001",
  41700=>"011011111",
  41701=>"101101111",
  41702=>"101111100",
  41703=>"111010100",
  41704=>"010100111",
  41705=>"000000010",
  41706=>"010000000",
  41707=>"000111100",
  41708=>"000101001",
  41709=>"101100011",
  41710=>"010101100",
  41711=>"111001011",
  41712=>"100111110",
  41713=>"011101110",
  41714=>"010111011",
  41715=>"011111001",
  41716=>"010011010",
  41717=>"000011000",
  41718=>"000011101",
  41719=>"101001100",
  41720=>"110110010",
  41721=>"101000000",
  41722=>"000100111",
  41723=>"010100100",
  41724=>"000000000",
  41725=>"010101001",
  41726=>"111100000",
  41727=>"010010000",
  41728=>"011111010",
  41729=>"011100001",
  41730=>"101100010",
  41731=>"011000110",
  41732=>"101100000",
  41733=>"011000111",
  41734=>"100010011",
  41735=>"111111100",
  41736=>"000100000",
  41737=>"110010001",
  41738=>"101110001",
  41739=>"000001101",
  41740=>"101110010",
  41741=>"000000010",
  41742=>"011000101",
  41743=>"101010011",
  41744=>"111000110",
  41745=>"011101001",
  41746=>"000000110",
  41747=>"111111110",
  41748=>"111110111",
  41749=>"000011100",
  41750=>"001001011",
  41751=>"110101001",
  41752=>"101001101",
  41753=>"100100100",
  41754=>"000001001",
  41755=>"001000100",
  41756=>"100111111",
  41757=>"100011011",
  41758=>"100001111",
  41759=>"001000011",
  41760=>"001001001",
  41761=>"111100101",
  41762=>"110001111",
  41763=>"100101001",
  41764=>"110011011",
  41765=>"101111100",
  41766=>"010110111",
  41767=>"111011100",
  41768=>"011011011",
  41769=>"101011011",
  41770=>"111000010",
  41771=>"101111011",
  41772=>"010001001",
  41773=>"110100100",
  41774=>"101101001",
  41775=>"011010011",
  41776=>"000000111",
  41777=>"111001000",
  41778=>"011000000",
  41779=>"010000010",
  41780=>"100101110",
  41781=>"101000101",
  41782=>"010010010",
  41783=>"100101100",
  41784=>"110100011",
  41785=>"011010000",
  41786=>"110011011",
  41787=>"001011000",
  41788=>"111000100",
  41789=>"011001110",
  41790=>"011000101",
  41791=>"110100000",
  41792=>"001101000",
  41793=>"011111011",
  41794=>"011000101",
  41795=>"100000100",
  41796=>"110111101",
  41797=>"011110101",
  41798=>"011101010",
  41799=>"101110100",
  41800=>"100001111",
  41801=>"001001011",
  41802=>"100000100",
  41803=>"000010100",
  41804=>"101001110",
  41805=>"110101100",
  41806=>"001101101",
  41807=>"111110110",
  41808=>"100101111",
  41809=>"100010110",
  41810=>"101101110",
  41811=>"010000011",
  41812=>"111110100",
  41813=>"010000111",
  41814=>"000110011",
  41815=>"101111010",
  41816=>"111100111",
  41817=>"111100110",
  41818=>"110010000",
  41819=>"111100001",
  41820=>"101010001",
  41821=>"010010000",
  41822=>"001100101",
  41823=>"101101000",
  41824=>"111101011",
  41825=>"101010100",
  41826=>"010111111",
  41827=>"010101000",
  41828=>"101001100",
  41829=>"111010010",
  41830=>"110100111",
  41831=>"001110010",
  41832=>"011110111",
  41833=>"111010101",
  41834=>"110101101",
  41835=>"111000011",
  41836=>"100100101",
  41837=>"001111001",
  41838=>"000100100",
  41839=>"110101111",
  41840=>"010110111",
  41841=>"000010010",
  41842=>"101110110",
  41843=>"111111000",
  41844=>"000101100",
  41845=>"010000101",
  41846=>"110001110",
  41847=>"101100001",
  41848=>"000111110",
  41849=>"111110011",
  41850=>"111001101",
  41851=>"111110101",
  41852=>"111110101",
  41853=>"001111101",
  41854=>"111000111",
  41855=>"001101011",
  41856=>"000010110",
  41857=>"000011110",
  41858=>"001000000",
  41859=>"110101100",
  41860=>"001011111",
  41861=>"010110010",
  41862=>"101010110",
  41863=>"011000101",
  41864=>"111011101",
  41865=>"011010111",
  41866=>"001101010",
  41867=>"110000010",
  41868=>"111011000",
  41869=>"000001010",
  41870=>"000011000",
  41871=>"001100100",
  41872=>"101111001",
  41873=>"101010010",
  41874=>"101100100",
  41875=>"101001100",
  41876=>"010001010",
  41877=>"100100010",
  41878=>"000001000",
  41879=>"101010111",
  41880=>"000111100",
  41881=>"111110111",
  41882=>"111011110",
  41883=>"110011100",
  41884=>"001110100",
  41885=>"000001000",
  41886=>"100110000",
  41887=>"101000101",
  41888=>"000001110",
  41889=>"101011011",
  41890=>"111111010",
  41891=>"111010101",
  41892=>"011101000",
  41893=>"110100111",
  41894=>"100011111",
  41895=>"101110001",
  41896=>"001101111",
  41897=>"001111010",
  41898=>"010110101",
  41899=>"100010011",
  41900=>"110111000",
  41901=>"010110111",
  41902=>"010110000",
  41903=>"011001100",
  41904=>"011101010",
  41905=>"111011000",
  41906=>"001101100",
  41907=>"011000111",
  41908=>"101110011",
  41909=>"100010000",
  41910=>"100111010",
  41911=>"111100011",
  41912=>"101101100",
  41913=>"101001000",
  41914=>"010010000",
  41915=>"110001001",
  41916=>"111010000",
  41917=>"101110011",
  41918=>"001011000",
  41919=>"000000000",
  41920=>"110101010",
  41921=>"000000010",
  41922=>"100111001",
  41923=>"011010001",
  41924=>"000110011",
  41925=>"000011110",
  41926=>"111010001",
  41927=>"100001100",
  41928=>"000000100",
  41929=>"011101011",
  41930=>"011000000",
  41931=>"010101000",
  41932=>"111110111",
  41933=>"000111101",
  41934=>"011111001",
  41935=>"100111111",
  41936=>"101110110",
  41937=>"010110101",
  41938=>"000011001",
  41939=>"010001110",
  41940=>"001011100",
  41941=>"010000000",
  41942=>"001111000",
  41943=>"010000001",
  41944=>"100001001",
  41945=>"110101001",
  41946=>"000110111",
  41947=>"001000000",
  41948=>"001101010",
  41949=>"000001000",
  41950=>"110000010",
  41951=>"110111111",
  41952=>"101101011",
  41953=>"110010001",
  41954=>"110011110",
  41955=>"110111000",
  41956=>"001001101",
  41957=>"010101100",
  41958=>"110100011",
  41959=>"101000110",
  41960=>"010010110",
  41961=>"111001100",
  41962=>"100000001",
  41963=>"010110010",
  41964=>"011100111",
  41965=>"010010000",
  41966=>"100011010",
  41967=>"000100001",
  41968=>"011100100",
  41969=>"111101110",
  41970=>"100010111",
  41971=>"101000000",
  41972=>"001001110",
  41973=>"010000000",
  41974=>"111000111",
  41975=>"101111010",
  41976=>"010001110",
  41977=>"100000000",
  41978=>"000101000",
  41979=>"010111111",
  41980=>"101111000",
  41981=>"000101000",
  41982=>"100010001",
  41983=>"100110010",
  41984=>"011011010",
  41985=>"110011010",
  41986=>"101011111",
  41987=>"000010111",
  41988=>"110110010",
  41989=>"100010100",
  41990=>"010100010",
  41991=>"110011100",
  41992=>"001111100",
  41993=>"010001001",
  41994=>"000010011",
  41995=>"111010100",
  41996=>"110011100",
  41997=>"010101111",
  41998=>"110111010",
  41999=>"111111110",
  42000=>"111000000",
  42001=>"001101110",
  42002=>"000111001",
  42003=>"110000110",
  42004=>"101001010",
  42005=>"101111001",
  42006=>"110100011",
  42007=>"111101011",
  42008=>"011011001",
  42009=>"110110101",
  42010=>"100111011",
  42011=>"111101001",
  42012=>"001100010",
  42013=>"001101010",
  42014=>"100100000",
  42015=>"000001000",
  42016=>"011101111",
  42017=>"011010111",
  42018=>"000001100",
  42019=>"101111101",
  42020=>"110010011",
  42021=>"111011100",
  42022=>"101111110",
  42023=>"000001000",
  42024=>"011001111",
  42025=>"110001000",
  42026=>"000010101",
  42027=>"010000100",
  42028=>"111111000",
  42029=>"101001011",
  42030=>"101010100",
  42031=>"111001100",
  42032=>"000101010",
  42033=>"000111101",
  42034=>"111000001",
  42035=>"100101011",
  42036=>"101001001",
  42037=>"100001010",
  42038=>"110111101",
  42039=>"001001101",
  42040=>"110101101",
  42041=>"101000010",
  42042=>"110011010",
  42043=>"101111100",
  42044=>"000001111",
  42045=>"001010010",
  42046=>"010011011",
  42047=>"101100001",
  42048=>"101100111",
  42049=>"000001000",
  42050=>"010101001",
  42051=>"000000011",
  42052=>"000001101",
  42053=>"000010111",
  42054=>"101001110",
  42055=>"101010010",
  42056=>"111110001",
  42057=>"100001010",
  42058=>"111100111",
  42059=>"101000000",
  42060=>"000001100",
  42061=>"001000001",
  42062=>"000001111",
  42063=>"111010110",
  42064=>"001110101",
  42065=>"111011111",
  42066=>"110101000",
  42067=>"100010100",
  42068=>"000001010",
  42069=>"110010000",
  42070=>"000000000",
  42071=>"101001100",
  42072=>"000100011",
  42073=>"101110010",
  42074=>"100101100",
  42075=>"011001110",
  42076=>"111111000",
  42077=>"000000000",
  42078=>"111101101",
  42079=>"000000111",
  42080=>"000110100",
  42081=>"010110000",
  42082=>"110100001",
  42083=>"100010100",
  42084=>"100100010",
  42085=>"101001110",
  42086=>"000100000",
  42087=>"111111011",
  42088=>"011000011",
  42089=>"011001001",
  42090=>"101111011",
  42091=>"010010010",
  42092=>"100011101",
  42093=>"011011100",
  42094=>"101001001",
  42095=>"000011111",
  42096=>"110110111",
  42097=>"110000010",
  42098=>"111010110",
  42099=>"000011100",
  42100=>"100111100",
  42101=>"101110100",
  42102=>"111000000",
  42103=>"011111101",
  42104=>"110001100",
  42105=>"110110100",
  42106=>"000010100",
  42107=>"000111000",
  42108=>"100010010",
  42109=>"111101100",
  42110=>"001000100",
  42111=>"100100001",
  42112=>"110100011",
  42113=>"010110100",
  42114=>"010011100",
  42115=>"110001101",
  42116=>"100000011",
  42117=>"110010111",
  42118=>"000001110",
  42119=>"100101010",
  42120=>"011000000",
  42121=>"001010000",
  42122=>"000101101",
  42123=>"111110100",
  42124=>"011101000",
  42125=>"011011000",
  42126=>"100101011",
  42127=>"111111100",
  42128=>"010100000",
  42129=>"111110100",
  42130=>"011100101",
  42131=>"010100100",
  42132=>"001010101",
  42133=>"010011100",
  42134=>"011101101",
  42135=>"100000100",
  42136=>"010110011",
  42137=>"010010110",
  42138=>"001010011",
  42139=>"000011100",
  42140=>"010011010",
  42141=>"010000111",
  42142=>"101000111",
  42143=>"110010011",
  42144=>"100000011",
  42145=>"010000010",
  42146=>"001001100",
  42147=>"101010100",
  42148=>"000011001",
  42149=>"101001011",
  42150=>"111100110",
  42151=>"100011111",
  42152=>"101110011",
  42153=>"001100100",
  42154=>"101100100",
  42155=>"110010000",
  42156=>"000010101",
  42157=>"000111011",
  42158=>"100101110",
  42159=>"110010010",
  42160=>"011011101",
  42161=>"000101010",
  42162=>"101001110",
  42163=>"011000100",
  42164=>"110110110",
  42165=>"011100110",
  42166=>"000000010",
  42167=>"010011101",
  42168=>"101100101",
  42169=>"010001000",
  42170=>"110011011",
  42171=>"010000111",
  42172=>"101111001",
  42173=>"101010000",
  42174=>"011111110",
  42175=>"011111001",
  42176=>"111110110",
  42177=>"000000000",
  42178=>"100111100",
  42179=>"010110111",
  42180=>"101111000",
  42181=>"011111100",
  42182=>"010010111",
  42183=>"110010000",
  42184=>"001111000",
  42185=>"100001011",
  42186=>"011101011",
  42187=>"001000000",
  42188=>"100101001",
  42189=>"011110010",
  42190=>"010100110",
  42191=>"010011111",
  42192=>"010100000",
  42193=>"111011011",
  42194=>"100000000",
  42195=>"101001101",
  42196=>"111010011",
  42197=>"110110001",
  42198=>"110011001",
  42199=>"111111100",
  42200=>"001011111",
  42201=>"111101101",
  42202=>"000100100",
  42203=>"110110100",
  42204=>"011100011",
  42205=>"011000011",
  42206=>"011000000",
  42207=>"100100001",
  42208=>"111111011",
  42209=>"110100011",
  42210=>"101000110",
  42211=>"111011011",
  42212=>"110100010",
  42213=>"110010100",
  42214=>"000011000",
  42215=>"100110111",
  42216=>"000111100",
  42217=>"101101010",
  42218=>"011111101",
  42219=>"000110011",
  42220=>"110100000",
  42221=>"010110001",
  42222=>"101000010",
  42223=>"101111001",
  42224=>"111010001",
  42225=>"111001010",
  42226=>"000100100",
  42227=>"000111101",
  42228=>"110111001",
  42229=>"001000011",
  42230=>"010001001",
  42231=>"011110100",
  42232=>"110011011",
  42233=>"001000100",
  42234=>"111010011",
  42235=>"001010100",
  42236=>"110010111",
  42237=>"010011111",
  42238=>"010111101",
  42239=>"000001000",
  42240=>"101001100",
  42241=>"111011101",
  42242=>"000010000",
  42243=>"111001010",
  42244=>"101100101",
  42245=>"100001001",
  42246=>"011100111",
  42247=>"010010100",
  42248=>"111101101",
  42249=>"100010001",
  42250=>"111100000",
  42251=>"011111111",
  42252=>"001011100",
  42253=>"111100111",
  42254=>"110001000",
  42255=>"010001010",
  42256=>"101100000",
  42257=>"100000000",
  42258=>"010100011",
  42259=>"110001101",
  42260=>"101000111",
  42261=>"110010100",
  42262=>"101110111",
  42263=>"001010000",
  42264=>"111111110",
  42265=>"001001101",
  42266=>"011000010",
  42267=>"100011100",
  42268=>"001111011",
  42269=>"011010011",
  42270=>"100110100",
  42271=>"000101000",
  42272=>"110110000",
  42273=>"101010100",
  42274=>"101010111",
  42275=>"010111010",
  42276=>"001011001",
  42277=>"011001101",
  42278=>"000011010",
  42279=>"000100000",
  42280=>"110011100",
  42281=>"101010010",
  42282=>"101110100",
  42283=>"101000000",
  42284=>"000000011",
  42285=>"001010010",
  42286=>"011101011",
  42287=>"010111101",
  42288=>"000111111",
  42289=>"100001110",
  42290=>"001010100",
  42291=>"110010001",
  42292=>"111011010",
  42293=>"001001101",
  42294=>"010011010",
  42295=>"110100111",
  42296=>"100100101",
  42297=>"101000101",
  42298=>"000011110",
  42299=>"011001111",
  42300=>"000001011",
  42301=>"110100110",
  42302=>"010111011",
  42303=>"001000100",
  42304=>"011111011",
  42305=>"000011001",
  42306=>"011100100",
  42307=>"110110000",
  42308=>"011100000",
  42309=>"011111111",
  42310=>"101100100",
  42311=>"111111011",
  42312=>"110101101",
  42313=>"110001011",
  42314=>"111100010",
  42315=>"101011111",
  42316=>"000101011",
  42317=>"111000101",
  42318=>"001001110",
  42319=>"100010101",
  42320=>"000000001",
  42321=>"011010100",
  42322=>"001010001",
  42323=>"010100000",
  42324=>"110011111",
  42325=>"000010111",
  42326=>"010010010",
  42327=>"001010000",
  42328=>"010001000",
  42329=>"110101110",
  42330=>"001000010",
  42331=>"000010000",
  42332=>"011000001",
  42333=>"010010101",
  42334=>"011011100",
  42335=>"101100111",
  42336=>"101001000",
  42337=>"100111010",
  42338=>"111111100",
  42339=>"011101001",
  42340=>"000101110",
  42341=>"011110010",
  42342=>"010101011",
  42343=>"011011010",
  42344=>"011011010",
  42345=>"000000000",
  42346=>"000001000",
  42347=>"000001100",
  42348=>"110000001",
  42349=>"101000111",
  42350=>"000110011",
  42351=>"100001000",
  42352=>"010010111",
  42353=>"011101010",
  42354=>"111110110",
  42355=>"111100101",
  42356=>"000000110",
  42357=>"000011000",
  42358=>"010001110",
  42359=>"110101001",
  42360=>"111100111",
  42361=>"111010000",
  42362=>"001001011",
  42363=>"111101010",
  42364=>"111001001",
  42365=>"010000110",
  42366=>"011101111",
  42367=>"011000001",
  42368=>"000111100",
  42369=>"111110111",
  42370=>"011010100",
  42371=>"011110111",
  42372=>"111101101",
  42373=>"011100000",
  42374=>"101100100",
  42375=>"111010111",
  42376=>"111111011",
  42377=>"100111011",
  42378=>"111111000",
  42379=>"101001011",
  42380=>"111101001",
  42381=>"001010110",
  42382=>"010111010",
  42383=>"001101001",
  42384=>"001011001",
  42385=>"000010101",
  42386=>"111011110",
  42387=>"000100110",
  42388=>"111001110",
  42389=>"111010010",
  42390=>"010111111",
  42391=>"011001010",
  42392=>"101011101",
  42393=>"000100111",
  42394=>"011010101",
  42395=>"110011010",
  42396=>"011101001",
  42397=>"011000101",
  42398=>"010001010",
  42399=>"101100111",
  42400=>"111111011",
  42401=>"010011010",
  42402=>"100110100",
  42403=>"000110000",
  42404=>"011000101",
  42405=>"001011011",
  42406=>"001100100",
  42407=>"111001001",
  42408=>"111110000",
  42409=>"010000011",
  42410=>"111010000",
  42411=>"000100111",
  42412=>"000101111",
  42413=>"101101110",
  42414=>"111000110",
  42415=>"110110100",
  42416=>"110010001",
  42417=>"000000110",
  42418=>"100001011",
  42419=>"011101110",
  42420=>"110101110",
  42421=>"101001001",
  42422=>"011111101",
  42423=>"010010111",
  42424=>"010011111",
  42425=>"001000000",
  42426=>"010010100",
  42427=>"010110101",
  42428=>"001111110",
  42429=>"010010010",
  42430=>"010111001",
  42431=>"000110001",
  42432=>"001001100",
  42433=>"000001000",
  42434=>"101101101",
  42435=>"011111000",
  42436=>"000100100",
  42437=>"001111100",
  42438=>"010111000",
  42439=>"001111110",
  42440=>"111111100",
  42441=>"110100111",
  42442=>"111000111",
  42443=>"110111010",
  42444=>"111000010",
  42445=>"110101010",
  42446=>"001000010",
  42447=>"001110011",
  42448=>"101010100",
  42449=>"001100110",
  42450=>"010100110",
  42451=>"001100000",
  42452=>"100111111",
  42453=>"000010010",
  42454=>"000011001",
  42455=>"110100100",
  42456=>"011010010",
  42457=>"111101010",
  42458=>"111111001",
  42459=>"010101010",
  42460=>"111101001",
  42461=>"010111110",
  42462=>"001011111",
  42463=>"110000101",
  42464=>"111011000",
  42465=>"011110000",
  42466=>"000000101",
  42467=>"010101100",
  42468=>"101110000",
  42469=>"100101010",
  42470=>"011010010",
  42471=>"000000010",
  42472=>"000101010",
  42473=>"000010100",
  42474=>"111011001",
  42475=>"101010010",
  42476=>"100000101",
  42477=>"000000000",
  42478=>"110011111",
  42479=>"101101010",
  42480=>"011011010",
  42481=>"111011111",
  42482=>"000001010",
  42483=>"000100010",
  42484=>"001011000",
  42485=>"101010010",
  42486=>"010100111",
  42487=>"010010000",
  42488=>"000001100",
  42489=>"011000000",
  42490=>"001100100",
  42491=>"110110010",
  42492=>"111011111",
  42493=>"000000000",
  42494=>"011111110",
  42495=>"010101111",
  42496=>"111111000",
  42497=>"100010100",
  42498=>"001101110",
  42499=>"010001111",
  42500=>"110000000",
  42501=>"000111101",
  42502=>"001000111",
  42503=>"011010111",
  42504=>"001110000",
  42505=>"000101000",
  42506=>"111001111",
  42507=>"100110110",
  42508=>"101101010",
  42509=>"000100110",
  42510=>"100000110",
  42511=>"001000000",
  42512=>"000001100",
  42513=>"001110111",
  42514=>"000011010",
  42515=>"000101010",
  42516=>"100110101",
  42517=>"101001110",
  42518=>"111000100",
  42519=>"001011010",
  42520=>"111101111",
  42521=>"000000011",
  42522=>"010000001",
  42523=>"001000111",
  42524=>"111101000",
  42525=>"001011100",
  42526=>"101101011",
  42527=>"101111101",
  42528=>"010101001",
  42529=>"100010100",
  42530=>"001010111",
  42531=>"000101011",
  42532=>"010110010",
  42533=>"000111101",
  42534=>"010010110",
  42535=>"100100011",
  42536=>"011100000",
  42537=>"111000110",
  42538=>"000100101",
  42539=>"000100100",
  42540=>"001100010",
  42541=>"110011100",
  42542=>"000000001",
  42543=>"100000010",
  42544=>"100101010",
  42545=>"100001011",
  42546=>"101101110",
  42547=>"011100100",
  42548=>"001110110",
  42549=>"001111111",
  42550=>"100100010",
  42551=>"110010100",
  42552=>"110011011",
  42553=>"010110011",
  42554=>"111110110",
  42555=>"000110011",
  42556=>"110001001",
  42557=>"111110001",
  42558=>"111101011",
  42559=>"010010101",
  42560=>"111000010",
  42561=>"000010110",
  42562=>"110010011",
  42563=>"111000010",
  42564=>"000010000",
  42565=>"111100000",
  42566=>"010001110",
  42567=>"011100000",
  42568=>"110010011",
  42569=>"010001100",
  42570=>"100111101",
  42571=>"100110011",
  42572=>"000110100",
  42573=>"101011100",
  42574=>"000001001",
  42575=>"101000101",
  42576=>"001011101",
  42577=>"000100000",
  42578=>"010101011",
  42579=>"110010010",
  42580=>"000111111",
  42581=>"001000111",
  42582=>"010000001",
  42583=>"110111100",
  42584=>"000000000",
  42585=>"100000010",
  42586=>"111010101",
  42587=>"110000000",
  42588=>"101011000",
  42589=>"011101001",
  42590=>"100001010",
  42591=>"000001100",
  42592=>"111110000",
  42593=>"101101110",
  42594=>"011110000",
  42595=>"111010000",
  42596=>"011100100",
  42597=>"010010011",
  42598=>"001101111",
  42599=>"000011111",
  42600=>"100000100",
  42601=>"111111111",
  42602=>"111110010",
  42603=>"011101000",
  42604=>"000101001",
  42605=>"111100011",
  42606=>"010101010",
  42607=>"101110101",
  42608=>"111110111",
  42609=>"010100010",
  42610=>"001010011",
  42611=>"000000110",
  42612=>"011011011",
  42613=>"111111101",
  42614=>"111111111",
  42615=>"000000000",
  42616=>"111010000",
  42617=>"110101111",
  42618=>"011111000",
  42619=>"001010000",
  42620=>"111110111",
  42621=>"100000011",
  42622=>"000000010",
  42623=>"010000001",
  42624=>"001010100",
  42625=>"101101111",
  42626=>"010111101",
  42627=>"001111101",
  42628=>"101000010",
  42629=>"111101001",
  42630=>"001010000",
  42631=>"111101111",
  42632=>"000010000",
  42633=>"100110101",
  42634=>"001011110",
  42635=>"110010001",
  42636=>"110111111",
  42637=>"101100001",
  42638=>"011100111",
  42639=>"110010000",
  42640=>"011110000",
  42641=>"010010000",
  42642=>"001011100",
  42643=>"101001010",
  42644=>"001000100",
  42645=>"101011001",
  42646=>"000100100",
  42647=>"110000111",
  42648=>"011010001",
  42649=>"000110010",
  42650=>"011101011",
  42651=>"111111100",
  42652=>"110010111",
  42653=>"111000111",
  42654=>"101110001",
  42655=>"100011100",
  42656=>"111110110",
  42657=>"011111000",
  42658=>"000111110",
  42659=>"010100101",
  42660=>"000100001",
  42661=>"111001110",
  42662=>"001011110",
  42663=>"000010111",
  42664=>"001000000",
  42665=>"111110100",
  42666=>"001010110",
  42667=>"111011111",
  42668=>"001111001",
  42669=>"101100111",
  42670=>"000100100",
  42671=>"101100101",
  42672=>"010100101",
  42673=>"000100010",
  42674=>"110101100",
  42675=>"110001110",
  42676=>"111111011",
  42677=>"101111100",
  42678=>"110111011",
  42679=>"101001111",
  42680=>"000000001",
  42681=>"000001001",
  42682=>"011011010",
  42683=>"100010000",
  42684=>"011010101",
  42685=>"000100011",
  42686=>"111101101",
  42687=>"110101001",
  42688=>"111010011",
  42689=>"110100001",
  42690=>"100100010",
  42691=>"110111111",
  42692=>"100001010",
  42693=>"110110000",
  42694=>"010010001",
  42695=>"000011001",
  42696=>"111110101",
  42697=>"000100100",
  42698=>"110000100",
  42699=>"010011100",
  42700=>"101101010",
  42701=>"000100011",
  42702=>"010001101",
  42703=>"010110111",
  42704=>"010111101",
  42705=>"011010010",
  42706=>"000010000",
  42707=>"011011100",
  42708=>"000011010",
  42709=>"011011000",
  42710=>"101110000",
  42711=>"010011110",
  42712=>"011010011",
  42713=>"001001110",
  42714=>"000011110",
  42715=>"001111100",
  42716=>"000000100",
  42717=>"110111010",
  42718=>"111100011",
  42719=>"101010010",
  42720=>"001100111",
  42721=>"001001001",
  42722=>"010011111",
  42723=>"110011111",
  42724=>"001001011",
  42725=>"110101001",
  42726=>"000001101",
  42727=>"000000111",
  42728=>"011000010",
  42729=>"011111101",
  42730=>"100000001",
  42731=>"000001000",
  42732=>"001011001",
  42733=>"000011000",
  42734=>"110100100",
  42735=>"010110110",
  42736=>"011010101",
  42737=>"100100110",
  42738=>"000110110",
  42739=>"101110010",
  42740=>"100111110",
  42741=>"011000110",
  42742=>"101100010",
  42743=>"100001111",
  42744=>"010011001",
  42745=>"111111010",
  42746=>"101110001",
  42747=>"100010000",
  42748=>"011001110",
  42749=>"101100110",
  42750=>"000111001",
  42751=>"000111001",
  42752=>"000111110",
  42753=>"110110010",
  42754=>"111110100",
  42755=>"000001110",
  42756=>"111110110",
  42757=>"001001100",
  42758=>"000011111",
  42759=>"011100101",
  42760=>"111000001",
  42761=>"101011010",
  42762=>"010011100",
  42763=>"010010110",
  42764=>"111001000",
  42765=>"100001100",
  42766=>"100111110",
  42767=>"010001000",
  42768=>"111011010",
  42769=>"111000011",
  42770=>"011100100",
  42771=>"100010101",
  42772=>"101000111",
  42773=>"100100000",
  42774=>"011011011",
  42775=>"001000001",
  42776=>"101000110",
  42777=>"101000110",
  42778=>"101010101",
  42779=>"100111010",
  42780=>"000111010",
  42781=>"111101110",
  42782=>"000101111",
  42783=>"011100011",
  42784=>"111000001",
  42785=>"010111100",
  42786=>"101011011",
  42787=>"111000111",
  42788=>"101101011",
  42789=>"010001011",
  42790=>"101111011",
  42791=>"011001100",
  42792=>"001000011",
  42793=>"110111000",
  42794=>"010110111",
  42795=>"000010000",
  42796=>"010001101",
  42797=>"001110110",
  42798=>"011010010",
  42799=>"010001100",
  42800=>"111010011",
  42801=>"111010010",
  42802=>"111000000",
  42803=>"101101001",
  42804=>"010001110",
  42805=>"000010001",
  42806=>"111110000",
  42807=>"001110010",
  42808=>"010110010",
  42809=>"110001010",
  42810=>"100001101",
  42811=>"011111111",
  42812=>"010001000",
  42813=>"000000110",
  42814=>"111011101",
  42815=>"000000100",
  42816=>"111111010",
  42817=>"110000010",
  42818=>"010100101",
  42819=>"111010100",
  42820=>"111011111",
  42821=>"101100001",
  42822=>"101001100",
  42823=>"101010001",
  42824=>"111101100",
  42825=>"110100100",
  42826=>"100111010",
  42827=>"000001110",
  42828=>"111100010",
  42829=>"011011111",
  42830=>"011101101",
  42831=>"101000111",
  42832=>"011000110",
  42833=>"101110111",
  42834=>"000000010",
  42835=>"100100110",
  42836=>"111010111",
  42837=>"010110001",
  42838=>"110111011",
  42839=>"011111010",
  42840=>"000110010",
  42841=>"111011001",
  42842=>"011011111",
  42843=>"011000101",
  42844=>"000100001",
  42845=>"110011000",
  42846=>"010100110",
  42847=>"011001000",
  42848=>"111001001",
  42849=>"011101001",
  42850=>"101000000",
  42851=>"011010111",
  42852=>"101011011",
  42853=>"100110010",
  42854=>"010011101",
  42855=>"101110111",
  42856=>"100100110",
  42857=>"111100000",
  42858=>"001101111",
  42859=>"111001000",
  42860=>"101011111",
  42861=>"000110010",
  42862=>"100010001",
  42863=>"110100100",
  42864=>"100010101",
  42865=>"010101110",
  42866=>"110001100",
  42867=>"011010000",
  42868=>"111110100",
  42869=>"011111111",
  42870=>"001001011",
  42871=>"010010001",
  42872=>"010100001",
  42873=>"001101110",
  42874=>"111001000",
  42875=>"000010101",
  42876=>"011010110",
  42877=>"110100000",
  42878=>"111101010",
  42879=>"001100100",
  42880=>"100011001",
  42881=>"110101001",
  42882=>"001110011",
  42883=>"000100100",
  42884=>"110001100",
  42885=>"110111001",
  42886=>"100001000",
  42887=>"100100011",
  42888=>"001010000",
  42889=>"000010100",
  42890=>"011000011",
  42891=>"110111101",
  42892=>"000111100",
  42893=>"010110101",
  42894=>"110111101",
  42895=>"011100011",
  42896=>"111011110",
  42897=>"000000000",
  42898=>"011001101",
  42899=>"100101001",
  42900=>"010110110",
  42901=>"100010111",
  42902=>"000101010",
  42903=>"100010001",
  42904=>"101111111",
  42905=>"101100001",
  42906=>"000001111",
  42907=>"101101110",
  42908=>"011100111",
  42909=>"111100110",
  42910=>"101101010",
  42911=>"101000100",
  42912=>"000100110",
  42913=>"011111001",
  42914=>"001110111",
  42915=>"110000111",
  42916=>"111100001",
  42917=>"111101011",
  42918=>"111011011",
  42919=>"000100001",
  42920=>"110000000",
  42921=>"011011011",
  42922=>"100001001",
  42923=>"001001010",
  42924=>"000101111",
  42925=>"110011110",
  42926=>"000011011",
  42927=>"001111101",
  42928=>"110000101",
  42929=>"101111111",
  42930=>"000000011",
  42931=>"001001100",
  42932=>"011111110",
  42933=>"110101000",
  42934=>"001100110",
  42935=>"111111111",
  42936=>"001110010",
  42937=>"111110111",
  42938=>"011101101",
  42939=>"010101111",
  42940=>"000011111",
  42941=>"011000010",
  42942=>"001100000",
  42943=>"100110110",
  42944=>"100111010",
  42945=>"111010010",
  42946=>"111111000",
  42947=>"000110001",
  42948=>"010000011",
  42949=>"000101000",
  42950=>"101111011",
  42951=>"000000110",
  42952=>"010010111",
  42953=>"000100000",
  42954=>"011100010",
  42955=>"110101111",
  42956=>"110011101",
  42957=>"111101101",
  42958=>"010101100",
  42959=>"101011000",
  42960=>"000111110",
  42961=>"111011000",
  42962=>"100110000",
  42963=>"111110010",
  42964=>"100011111",
  42965=>"101110110",
  42966=>"000000100",
  42967=>"111001000",
  42968=>"100000000",
  42969=>"110110001",
  42970=>"100001001",
  42971=>"110010001",
  42972=>"111011001",
  42973=>"010110111",
  42974=>"010111100",
  42975=>"010100101",
  42976=>"100011111",
  42977=>"000000001",
  42978=>"000101101",
  42979=>"000111111",
  42980=>"111011111",
  42981=>"000010001",
  42982=>"011010111",
  42983=>"101001111",
  42984=>"111001101",
  42985=>"100100111",
  42986=>"000010000",
  42987=>"111010011",
  42988=>"000000110",
  42989=>"100110100",
  42990=>"000110000",
  42991=>"111110110",
  42992=>"010110000",
  42993=>"010101111",
  42994=>"001000010",
  42995=>"000111100",
  42996=>"000010010",
  42997=>"110100110",
  42998=>"000000011",
  42999=>"000000010",
  43000=>"010111100",
  43001=>"001101011",
  43002=>"111110001",
  43003=>"000111010",
  43004=>"111010010",
  43005=>"101001000",
  43006=>"101011011",
  43007=>"110000001",
  43008=>"111100111",
  43009=>"110011110",
  43010=>"011010111",
  43011=>"100101110",
  43012=>"110001110",
  43013=>"101000000",
  43014=>"101000110",
  43015=>"001101100",
  43016=>"101001100",
  43017=>"011100100",
  43018=>"110101111",
  43019=>"011100000",
  43020=>"000111101",
  43021=>"110010001",
  43022=>"100001001",
  43023=>"010100111",
  43024=>"000101000",
  43025=>"000101010",
  43026=>"110111101",
  43027=>"011100100",
  43028=>"111100101",
  43029=>"000000010",
  43030=>"010010001",
  43031=>"001111010",
  43032=>"111001100",
  43033=>"111100001",
  43034=>"101011100",
  43035=>"100000001",
  43036=>"110101111",
  43037=>"010001100",
  43038=>"000101101",
  43039=>"000001001",
  43040=>"001001001",
  43041=>"110111011",
  43042=>"001110011",
  43043=>"111100000",
  43044=>"110110100",
  43045=>"000111111",
  43046=>"010100110",
  43047=>"111101010",
  43048=>"100101000",
  43049=>"011100010",
  43050=>"101000101",
  43051=>"110101011",
  43052=>"110000100",
  43053=>"010001001",
  43054=>"110101111",
  43055=>"010010010",
  43056=>"111100000",
  43057=>"110100110",
  43058=>"001001010",
  43059=>"100010110",
  43060=>"111110011",
  43061=>"010011010",
  43062=>"101011011",
  43063=>"000100100",
  43064=>"101000110",
  43065=>"010110010",
  43066=>"000010111",
  43067=>"001010110",
  43068=>"001001010",
  43069=>"100110110",
  43070=>"100000100",
  43071=>"001011010",
  43072=>"010101100",
  43073=>"011001100",
  43074=>"100101110",
  43075=>"011101010",
  43076=>"100110100",
  43077=>"010011111",
  43078=>"100110101",
  43079=>"111100100",
  43080=>"110000111",
  43081=>"111101110",
  43082=>"001010001",
  43083=>"101000101",
  43084=>"010000101",
  43085=>"100101111",
  43086=>"010101001",
  43087=>"110001010",
  43088=>"111101100",
  43089=>"100001110",
  43090=>"001011001",
  43091=>"001100011",
  43092=>"011011000",
  43093=>"111100110",
  43094=>"100110100",
  43095=>"100001010",
  43096=>"010011000",
  43097=>"001101101",
  43098=>"010010001",
  43099=>"011010001",
  43100=>"011010011",
  43101=>"001100011",
  43102=>"100101010",
  43103=>"111011111",
  43104=>"000010011",
  43105=>"000011011",
  43106=>"111000110",
  43107=>"111111101",
  43108=>"010110000",
  43109=>"100101010",
  43110=>"111110100",
  43111=>"110101001",
  43112=>"111000001",
  43113=>"110001110",
  43114=>"010010100",
  43115=>"100100000",
  43116=>"101000000",
  43117=>"101011000",
  43118=>"101101010",
  43119=>"100011101",
  43120=>"100000000",
  43121=>"110101001",
  43122=>"010001100",
  43123=>"001001000",
  43124=>"101100010",
  43125=>"101010101",
  43126=>"110000100",
  43127=>"001110000",
  43128=>"010100010",
  43129=>"110010110",
  43130=>"111101111",
  43131=>"110100111",
  43132=>"010001011",
  43133=>"111010110",
  43134=>"111111111",
  43135=>"101010111",
  43136=>"011000110",
  43137=>"011100110",
  43138=>"111101010",
  43139=>"000111110",
  43140=>"010001010",
  43141=>"111011100",
  43142=>"111010110",
  43143=>"110110110",
  43144=>"100101110",
  43145=>"111010010",
  43146=>"111100011",
  43147=>"011111100",
  43148=>"001100011",
  43149=>"011000000",
  43150=>"000010101",
  43151=>"001010001",
  43152=>"100010001",
  43153=>"001011110",
  43154=>"111000011",
  43155=>"100011100",
  43156=>"101001010",
  43157=>"000101100",
  43158=>"110100011",
  43159=>"101110110",
  43160=>"110010010",
  43161=>"010001001",
  43162=>"111001111",
  43163=>"110101111",
  43164=>"010111100",
  43165=>"111000110",
  43166=>"000111111",
  43167=>"110011001",
  43168=>"000101011",
  43169=>"010001110",
  43170=>"010001010",
  43171=>"001011000",
  43172=>"000001110",
  43173=>"001111010",
  43174=>"001000101",
  43175=>"111111110",
  43176=>"111111100",
  43177=>"011010010",
  43178=>"011001100",
  43179=>"100111010",
  43180=>"000111100",
  43181=>"100010011",
  43182=>"011101100",
  43183=>"010000110",
  43184=>"100111001",
  43185=>"000111000",
  43186=>"101011101",
  43187=>"100011011",
  43188=>"111011100",
  43189=>"101100111",
  43190=>"100110111",
  43191=>"000001111",
  43192=>"001110001",
  43193=>"010010000",
  43194=>"110100011",
  43195=>"100101000",
  43196=>"111001110",
  43197=>"100001011",
  43198=>"110110101",
  43199=>"011000010",
  43200=>"110110010",
  43201=>"100111011",
  43202=>"001011110",
  43203=>"010101100",
  43204=>"000000000",
  43205=>"101010010",
  43206=>"001010101",
  43207=>"010110101",
  43208=>"101011110",
  43209=>"001100011",
  43210=>"000000110",
  43211=>"100101010",
  43212=>"010110001",
  43213=>"100100000",
  43214=>"000000111",
  43215=>"000001101",
  43216=>"011111110",
  43217=>"011110001",
  43218=>"010101010",
  43219=>"100001110",
  43220=>"011110111",
  43221=>"110011111",
  43222=>"010011101",
  43223=>"101111100",
  43224=>"110110100",
  43225=>"110100000",
  43226=>"111011010",
  43227=>"101000000",
  43228=>"110110100",
  43229=>"000100001",
  43230=>"111001111",
  43231=>"000001001",
  43232=>"001110000",
  43233=>"001101000",
  43234=>"110110100",
  43235=>"100011000",
  43236=>"111001010",
  43237=>"100100111",
  43238=>"111000100",
  43239=>"001001010",
  43240=>"011010000",
  43241=>"111011000",
  43242=>"010111110",
  43243=>"011011000",
  43244=>"001010000",
  43245=>"010001101",
  43246=>"110100101",
  43247=>"110011000",
  43248=>"111110101",
  43249=>"101000001",
  43250=>"001000000",
  43251=>"101011000",
  43252=>"101011000",
  43253=>"101000000",
  43254=>"111011111",
  43255=>"001110111",
  43256=>"010110111",
  43257=>"111110011",
  43258=>"001111110",
  43259=>"100010101",
  43260=>"110000001",
  43261=>"001100001",
  43262=>"001111100",
  43263=>"011111000",
  43264=>"001010110",
  43265=>"000101000",
  43266=>"001101010",
  43267=>"000000010",
  43268=>"111111010",
  43269=>"101001100",
  43270=>"001000001",
  43271=>"100100110",
  43272=>"001110001",
  43273=>"000011000",
  43274=>"000100010",
  43275=>"100101100",
  43276=>"110110000",
  43277=>"110001101",
  43278=>"101010000",
  43279=>"111110011",
  43280=>"110101000",
  43281=>"100010010",
  43282=>"001110011",
  43283=>"111010000",
  43284=>"100111101",
  43285=>"011011111",
  43286=>"110100001",
  43287=>"011110010",
  43288=>"111111011",
  43289=>"100000110",
  43290=>"001100111",
  43291=>"011110101",
  43292=>"111100110",
  43293=>"110011111",
  43294=>"011011101",
  43295=>"001000111",
  43296=>"011000100",
  43297=>"011011100",
  43298=>"101001111",
  43299=>"011110001",
  43300=>"000111010",
  43301=>"000000000",
  43302=>"010100010",
  43303=>"101111000",
  43304=>"111010000",
  43305=>"100100000",
  43306=>"110010111",
  43307=>"011110010",
  43308=>"000000111",
  43309=>"110100111",
  43310=>"011100101",
  43311=>"011011000",
  43312=>"101111101",
  43313=>"100100000",
  43314=>"000100111",
  43315=>"000110010",
  43316=>"000110011",
  43317=>"000110111",
  43318=>"010001010",
  43319=>"100110000",
  43320=>"111101111",
  43321=>"010011011",
  43322=>"100011010",
  43323=>"001010100",
  43324=>"100110011",
  43325=>"101100001",
  43326=>"111001100",
  43327=>"000110011",
  43328=>"001001110",
  43329=>"111100111",
  43330=>"110011001",
  43331=>"111110010",
  43332=>"011011110",
  43333=>"001000100",
  43334=>"111100010",
  43335=>"011101000",
  43336=>"101111111",
  43337=>"101000000",
  43338=>"001001110",
  43339=>"001101100",
  43340=>"010111011",
  43341=>"110010111",
  43342=>"101110010",
  43343=>"010010001",
  43344=>"111010111",
  43345=>"111100000",
  43346=>"011010100",
  43347=>"010010101",
  43348=>"010011000",
  43349=>"110110101",
  43350=>"100101001",
  43351=>"101101100",
  43352=>"011010100",
  43353=>"101111111",
  43354=>"000010100",
  43355=>"111100111",
  43356=>"000100110",
  43357=>"100111111",
  43358=>"111101011",
  43359=>"010011001",
  43360=>"100011000",
  43361=>"110000110",
  43362=>"010101001",
  43363=>"111110111",
  43364=>"100011001",
  43365=>"111110101",
  43366=>"010110111",
  43367=>"111110110",
  43368=>"100011110",
  43369=>"000111111",
  43370=>"100100000",
  43371=>"110110000",
  43372=>"111010011",
  43373=>"101100111",
  43374=>"100010011",
  43375=>"111011100",
  43376=>"000111111",
  43377=>"100101100",
  43378=>"110010111",
  43379=>"111111010",
  43380=>"001000010",
  43381=>"010110010",
  43382=>"001000100",
  43383=>"001110000",
  43384=>"010110011",
  43385=>"010000000",
  43386=>"100110100",
  43387=>"110010000",
  43388=>"001011101",
  43389=>"100100001",
  43390=>"011100000",
  43391=>"011001101",
  43392=>"011000000",
  43393=>"011000011",
  43394=>"110101001",
  43395=>"000110010",
  43396=>"000111111",
  43397=>"001011011",
  43398=>"010000011",
  43399=>"011010001",
  43400=>"001001111",
  43401=>"110100100",
  43402=>"010011100",
  43403=>"101101000",
  43404=>"001101011",
  43405=>"001100111",
  43406=>"100101110",
  43407=>"101000101",
  43408=>"110001011",
  43409=>"110001100",
  43410=>"110100101",
  43411=>"000110000",
  43412=>"010110111",
  43413=>"000111111",
  43414=>"000110000",
  43415=>"011010001",
  43416=>"100110111",
  43417=>"100100101",
  43418=>"000101011",
  43419=>"101010001",
  43420=>"100011111",
  43421=>"011110110",
  43422=>"100010110",
  43423=>"001101010",
  43424=>"110101011",
  43425=>"111111010",
  43426=>"010010100",
  43427=>"111001111",
  43428=>"001111011",
  43429=>"111110111",
  43430=>"001010000",
  43431=>"111111010",
  43432=>"101100000",
  43433=>"111111001",
  43434=>"101110010",
  43435=>"000000001",
  43436=>"110011111",
  43437=>"011001011",
  43438=>"001101111",
  43439=>"000111101",
  43440=>"110000011",
  43441=>"000010001",
  43442=>"001011101",
  43443=>"001011000",
  43444=>"101010111",
  43445=>"000110101",
  43446=>"010011110",
  43447=>"100111101",
  43448=>"111011011",
  43449=>"101111110",
  43450=>"010110100",
  43451=>"010001110",
  43452=>"000110101",
  43453=>"001111100",
  43454=>"100101000",
  43455=>"110000010",
  43456=>"000011001",
  43457=>"100110011",
  43458=>"111111101",
  43459=>"011000110",
  43460=>"101101111",
  43461=>"011111100",
  43462=>"000000101",
  43463=>"000000111",
  43464=>"110011100",
  43465=>"001100011",
  43466=>"110111111",
  43467=>"000111000",
  43468=>"000111100",
  43469=>"101100100",
  43470=>"001110100",
  43471=>"000010101",
  43472=>"111110001",
  43473=>"001101101",
  43474=>"111001111",
  43475=>"010100101",
  43476=>"010110111",
  43477=>"001111011",
  43478=>"001000101",
  43479=>"100100010",
  43480=>"000011011",
  43481=>"100111000",
  43482=>"111011000",
  43483=>"010010001",
  43484=>"100011111",
  43485=>"101011101",
  43486=>"100111000",
  43487=>"101011101",
  43488=>"100011001",
  43489=>"101110111",
  43490=>"011001111",
  43491=>"101110000",
  43492=>"000100010",
  43493=>"000010010",
  43494=>"110111111",
  43495=>"101100000",
  43496=>"010101101",
  43497=>"100100100",
  43498=>"111110101",
  43499=>"100011100",
  43500=>"000111000",
  43501=>"100101111",
  43502=>"101000111",
  43503=>"100100000",
  43504=>"111100000",
  43505=>"100000011",
  43506=>"001010010",
  43507=>"011010111",
  43508=>"110000010",
  43509=>"010101101",
  43510=>"110010001",
  43511=>"000011010",
  43512=>"010100000",
  43513=>"001110000",
  43514=>"001111101",
  43515=>"100010001",
  43516=>"011011111",
  43517=>"010011011",
  43518=>"011100001",
  43519=>"111000110",
  43520=>"111111101",
  43521=>"110111000",
  43522=>"000110111",
  43523=>"000000000",
  43524=>"100010001",
  43525=>"111001111",
  43526=>"110011000",
  43527=>"100101011",
  43528=>"011100111",
  43529=>"000101111",
  43530=>"001110110",
  43531=>"111110110",
  43532=>"100100101",
  43533=>"111100011",
  43534=>"000001011",
  43535=>"101001010",
  43536=>"111110001",
  43537=>"101010011",
  43538=>"101011000",
  43539=>"100000111",
  43540=>"000010100",
  43541=>"011111100",
  43542=>"011100111",
  43543=>"001110011",
  43544=>"011000000",
  43545=>"011110110",
  43546=>"111100101",
  43547=>"010000110",
  43548=>"100001111",
  43549=>"100010011",
  43550=>"010110010",
  43551=>"010101100",
  43552=>"100001001",
  43553=>"000100001",
  43554=>"001000111",
  43555=>"001101011",
  43556=>"010111011",
  43557=>"111010000",
  43558=>"101000000",
  43559=>"101110000",
  43560=>"111100100",
  43561=>"100011110",
  43562=>"010011010",
  43563=>"001011010",
  43564=>"110101000",
  43565=>"100100011",
  43566=>"111011001",
  43567=>"011000110",
  43568=>"111110001",
  43569=>"010011111",
  43570=>"110111001",
  43571=>"001111110",
  43572=>"010100000",
  43573=>"100110001",
  43574=>"100111000",
  43575=>"000001001",
  43576=>"000100011",
  43577=>"010010000",
  43578=>"010001100",
  43579=>"000011011",
  43580=>"011001011",
  43581=>"100101010",
  43582=>"000011110",
  43583=>"000011010",
  43584=>"101111111",
  43585=>"101001011",
  43586=>"001011101",
  43587=>"101001110",
  43588=>"110110111",
  43589=>"100101110",
  43590=>"100010101",
  43591=>"000110101",
  43592=>"000100001",
  43593=>"111101001",
  43594=>"001000010",
  43595=>"010100010",
  43596=>"111000001",
  43597=>"000110110",
  43598=>"110011111",
  43599=>"111001011",
  43600=>"010001001",
  43601=>"011110110",
  43602=>"001011000",
  43603=>"001100001",
  43604=>"010100010",
  43605=>"111111101",
  43606=>"011110000",
  43607=>"111000101",
  43608=>"011001010",
  43609=>"010101111",
  43610=>"100011111",
  43611=>"111010001",
  43612=>"001100110",
  43613=>"110100100",
  43614=>"100001001",
  43615=>"111011101",
  43616=>"101000011",
  43617=>"100000010",
  43618=>"101100000",
  43619=>"100101001",
  43620=>"110011010",
  43621=>"000110000",
  43622=>"111001000",
  43623=>"000110011",
  43624=>"010000001",
  43625=>"010111110",
  43626=>"100111100",
  43627=>"110110001",
  43628=>"101011111",
  43629=>"000111110",
  43630=>"001100100",
  43631=>"010101010",
  43632=>"000111011",
  43633=>"110111110",
  43634=>"011010101",
  43635=>"011100111",
  43636=>"111010010",
  43637=>"001000011",
  43638=>"010110000",
  43639=>"101011100",
  43640=>"001010010",
  43641=>"010001100",
  43642=>"111100110",
  43643=>"010011000",
  43644=>"001111100",
  43645=>"110100101",
  43646=>"110100100",
  43647=>"110011011",
  43648=>"011001110",
  43649=>"111100000",
  43650=>"101000111",
  43651=>"101011000",
  43652=>"010010000",
  43653=>"010100010",
  43654=>"011100011",
  43655=>"100001001",
  43656=>"010110010",
  43657=>"100001100",
  43658=>"111111100",
  43659=>"101000110",
  43660=>"110001011",
  43661=>"000101100",
  43662=>"111101111",
  43663=>"101000001",
  43664=>"101110111",
  43665=>"100101101",
  43666=>"110101011",
  43667=>"111100101",
  43668=>"011100000",
  43669=>"110101100",
  43670=>"011011000",
  43671=>"000100111",
  43672=>"101000010",
  43673=>"111110101",
  43674=>"000000101",
  43675=>"010111011",
  43676=>"000111101",
  43677=>"100110001",
  43678=>"000100011",
  43679=>"101001101",
  43680=>"110110101",
  43681=>"001111110",
  43682=>"111111010",
  43683=>"111011000",
  43684=>"011001110",
  43685=>"010111110",
  43686=>"100011010",
  43687=>"100110010",
  43688=>"010110001",
  43689=>"100000000",
  43690=>"010000011",
  43691=>"000100001",
  43692=>"000001101",
  43693=>"010101110",
  43694=>"110000001",
  43695=>"101001001",
  43696=>"010100110",
  43697=>"011110011",
  43698=>"101001000",
  43699=>"010010110",
  43700=>"101111000",
  43701=>"110000011",
  43702=>"010001101",
  43703=>"110001010",
  43704=>"110011110",
  43705=>"011111001",
  43706=>"111010100",
  43707=>"100000011",
  43708=>"100100010",
  43709=>"000010000",
  43710=>"101000011",
  43711=>"010010101",
  43712=>"100101001",
  43713=>"110100111",
  43714=>"010001000",
  43715=>"100111110",
  43716=>"110011110",
  43717=>"100110100",
  43718=>"111001011",
  43719=>"000010101",
  43720=>"001011001",
  43721=>"001000100",
  43722=>"100000110",
  43723=>"011011101",
  43724=>"100101001",
  43725=>"100011110",
  43726=>"100011010",
  43727=>"111110100",
  43728=>"110100110",
  43729=>"101100001",
  43730=>"111101100",
  43731=>"110001100",
  43732=>"100010111",
  43733=>"010001100",
  43734=>"000110001",
  43735=>"000100101",
  43736=>"000110111",
  43737=>"111000100",
  43738=>"110100111",
  43739=>"100101110",
  43740=>"001101110",
  43741=>"100110110",
  43742=>"011001000",
  43743=>"100001011",
  43744=>"100100010",
  43745=>"001011010",
  43746=>"100010000",
  43747=>"000111011",
  43748=>"011000001",
  43749=>"101001011",
  43750=>"101010111",
  43751=>"011111101",
  43752=>"101100111",
  43753=>"110010011",
  43754=>"000001000",
  43755=>"010111010",
  43756=>"001001000",
  43757=>"110010111",
  43758=>"011111101",
  43759=>"110000010",
  43760=>"111001010",
  43761=>"100010001",
  43762=>"111010011",
  43763=>"110110100",
  43764=>"011100011",
  43765=>"011100101",
  43766=>"111011110",
  43767=>"110001111",
  43768=>"000110111",
  43769=>"100111000",
  43770=>"111101111",
  43771=>"011010011",
  43772=>"110000100",
  43773=>"000111000",
  43774=>"000111111",
  43775=>"100111111",
  43776=>"000000100",
  43777=>"100011010",
  43778=>"100000010",
  43779=>"001001010",
  43780=>"110001100",
  43781=>"111001010",
  43782=>"100101001",
  43783=>"011110110",
  43784=>"001001000",
  43785=>"010000111",
  43786=>"000010101",
  43787=>"111001001",
  43788=>"111000011",
  43789=>"111111101",
  43790=>"110011111",
  43791=>"101101101",
  43792=>"110000100",
  43793=>"100100010",
  43794=>"111001101",
  43795=>"110011101",
  43796=>"110000011",
  43797=>"000101011",
  43798=>"010001011",
  43799=>"100010111",
  43800=>"101101000",
  43801=>"110001100",
  43802=>"001101001",
  43803=>"101111010",
  43804=>"001101010",
  43805=>"000111111",
  43806=>"000000111",
  43807=>"100011010",
  43808=>"110100011",
  43809=>"101101110",
  43810=>"111111111",
  43811=>"100000000",
  43812=>"000000110",
  43813=>"001000011",
  43814=>"110001100",
  43815=>"110000001",
  43816=>"100000110",
  43817=>"010111000",
  43818=>"110110000",
  43819=>"111011110",
  43820=>"101000000",
  43821=>"111100000",
  43822=>"000101000",
  43823=>"011001110",
  43824=>"010111010",
  43825=>"000101111",
  43826=>"000111010",
  43827=>"111101011",
  43828=>"111000000",
  43829=>"111100001",
  43830=>"100011111",
  43831=>"111010011",
  43832=>"001001010",
  43833=>"000100000",
  43834=>"101111100",
  43835=>"000111101",
  43836=>"001011111",
  43837=>"101101101",
  43838=>"000101000",
  43839=>"010001100",
  43840=>"001101000",
  43841=>"111001011",
  43842=>"001011101",
  43843=>"000100010",
  43844=>"000010000",
  43845=>"100100111",
  43846=>"011001001",
  43847=>"101000010",
  43848=>"100001010",
  43849=>"010000000",
  43850=>"110101000",
  43851=>"010010110",
  43852=>"110100110",
  43853=>"110001100",
  43854=>"100110101",
  43855=>"010000101",
  43856=>"101111101",
  43857=>"000011110",
  43858=>"100000101",
  43859=>"011111111",
  43860=>"110000111",
  43861=>"000111000",
  43862=>"111010011",
  43863=>"010010011",
  43864=>"010001000",
  43865=>"001101001",
  43866=>"010001100",
  43867=>"001110011",
  43868=>"101000011",
  43869=>"110001110",
  43870=>"000001000",
  43871=>"110110101",
  43872=>"000010100",
  43873=>"111100011",
  43874=>"100001010",
  43875=>"001001110",
  43876=>"111001010",
  43877=>"111001001",
  43878=>"010111101",
  43879=>"011110010",
  43880=>"001011110",
  43881=>"101000101",
  43882=>"010111001",
  43883=>"001101010",
  43884=>"110000101",
  43885=>"110101111",
  43886=>"000010001",
  43887=>"110011011",
  43888=>"000100010",
  43889=>"000101000",
  43890=>"001101010",
  43891=>"110101101",
  43892=>"001000100",
  43893=>"000111100",
  43894=>"111011000",
  43895=>"000101111",
  43896=>"100110000",
  43897=>"000010011",
  43898=>"000000100",
  43899=>"010010000",
  43900=>"110100010",
  43901=>"000000010",
  43902=>"001111110",
  43903=>"011111101",
  43904=>"011101101",
  43905=>"110011010",
  43906=>"101001100",
  43907=>"101000111",
  43908=>"111000110",
  43909=>"011111110",
  43910=>"000011100",
  43911=>"100010011",
  43912=>"101110101",
  43913=>"010011101",
  43914=>"011100111",
  43915=>"111010110",
  43916=>"110111000",
  43917=>"110101011",
  43918=>"001011011",
  43919=>"000101111",
  43920=>"011010000",
  43921=>"010101111",
  43922=>"000000101",
  43923=>"000010101",
  43924=>"011100100",
  43925=>"010000101",
  43926=>"010001111",
  43927=>"100110000",
  43928=>"111010000",
  43929=>"001000011",
  43930=>"110000100",
  43931=>"111010110",
  43932=>"100010101",
  43933=>"011110111",
  43934=>"001001000",
  43935=>"100101100",
  43936=>"011011100",
  43937=>"000110100",
  43938=>"010100100",
  43939=>"001110010",
  43940=>"001000101",
  43941=>"110100101",
  43942=>"011101010",
  43943=>"011110111",
  43944=>"001101010",
  43945=>"000010100",
  43946=>"000111011",
  43947=>"111010110",
  43948=>"001100110",
  43949=>"100011010",
  43950=>"100110010",
  43951=>"110100101",
  43952=>"001001101",
  43953=>"111011001",
  43954=>"100111110",
  43955=>"000111100",
  43956=>"001010010",
  43957=>"101011111",
  43958=>"010011000",
  43959=>"010000110",
  43960=>"001010011",
  43961=>"000101100",
  43962=>"010010101",
  43963=>"100100110",
  43964=>"111100111",
  43965=>"001101101",
  43966=>"001101001",
  43967=>"111111110",
  43968=>"001000010",
  43969=>"111100000",
  43970=>"000111101",
  43971=>"111101000",
  43972=>"111011011",
  43973=>"011010111",
  43974=>"101010100",
  43975=>"111000110",
  43976=>"010111001",
  43977=>"111001000",
  43978=>"101100111",
  43979=>"100010100",
  43980=>"010000110",
  43981=>"011000100",
  43982=>"010010110",
  43983=>"010100011",
  43984=>"010100101",
  43985=>"100000011",
  43986=>"100110001",
  43987=>"110100010",
  43988=>"111110110",
  43989=>"100110010",
  43990=>"100011101",
  43991=>"111100010",
  43992=>"111011101",
  43993=>"111001101",
  43994=>"001011011",
  43995=>"101111010",
  43996=>"100011101",
  43997=>"010100100",
  43998=>"000100110",
  43999=>"001000110",
  44000=>"000000000",
  44001=>"111100110",
  44002=>"011011000",
  44003=>"111011111",
  44004=>"101000101",
  44005=>"001010000",
  44006=>"000011001",
  44007=>"001101000",
  44008=>"100100000",
  44009=>"111110010",
  44010=>"000101011",
  44011=>"001101110",
  44012=>"011101100",
  44013=>"100000101",
  44014=>"010110101",
  44015=>"010000101",
  44016=>"111010111",
  44017=>"101001100",
  44018=>"001101001",
  44019=>"001101110",
  44020=>"101100011",
  44021=>"111011111",
  44022=>"010010010",
  44023=>"101001111",
  44024=>"010110110",
  44025=>"011101011",
  44026=>"110111011",
  44027=>"011001110",
  44028=>"111111111",
  44029=>"100010110",
  44030=>"001001111",
  44031=>"001001011",
  44032=>"100010010",
  44033=>"001000101",
  44034=>"100001000",
  44035=>"111001111",
  44036=>"110010011",
  44037=>"010100010",
  44038=>"001000001",
  44039=>"001101001",
  44040=>"001000001",
  44041=>"001110100",
  44042=>"011011011",
  44043=>"101110000",
  44044=>"001010010",
  44045=>"011010101",
  44046=>"011100111",
  44047=>"101000101",
  44048=>"001000110",
  44049=>"101110010",
  44050=>"100110001",
  44051=>"110000011",
  44052=>"001011011",
  44053=>"101011001",
  44054=>"111101100",
  44055=>"011001111",
  44056=>"100011111",
  44057=>"101010010",
  44058=>"100111101",
  44059=>"001001100",
  44060=>"000110100",
  44061=>"000011010",
  44062=>"001011111",
  44063=>"110111011",
  44064=>"110001101",
  44065=>"000111010",
  44066=>"111111110",
  44067=>"001110010",
  44068=>"001110001",
  44069=>"101110101",
  44070=>"101111111",
  44071=>"011101011",
  44072=>"100011110",
  44073=>"101101100",
  44074=>"110010100",
  44075=>"110000110",
  44076=>"001111110",
  44077=>"100110100",
  44078=>"001111101",
  44079=>"101010011",
  44080=>"000010100",
  44081=>"111101011",
  44082=>"111100001",
  44083=>"111101111",
  44084=>"001011100",
  44085=>"010110000",
  44086=>"101100011",
  44087=>"001011101",
  44088=>"000000000",
  44089=>"110110100",
  44090=>"010001000",
  44091=>"101000110",
  44092=>"010000011",
  44093=>"100000000",
  44094=>"100110011",
  44095=>"100101001",
  44096=>"010000001",
  44097=>"010011001",
  44098=>"100000000",
  44099=>"000101110",
  44100=>"011001101",
  44101=>"001000000",
  44102=>"101001000",
  44103=>"110101001",
  44104=>"010101001",
  44105=>"001100000",
  44106=>"010100000",
  44107=>"110110100",
  44108=>"000111011",
  44109=>"100111110",
  44110=>"111011100",
  44111=>"000000101",
  44112=>"101001010",
  44113=>"000001011",
  44114=>"010101011",
  44115=>"010010110",
  44116=>"110001010",
  44117=>"110110011",
  44118=>"110001000",
  44119=>"001101101",
  44120=>"010110110",
  44121=>"011101001",
  44122=>"001000010",
  44123=>"011000101",
  44124=>"000111011",
  44125=>"110111101",
  44126=>"001010101",
  44127=>"110111101",
  44128=>"010111100",
  44129=>"100111001",
  44130=>"011011001",
  44131=>"110011111",
  44132=>"001000111",
  44133=>"011001011",
  44134=>"111110110",
  44135=>"011000111",
  44136=>"110001000",
  44137=>"001101110",
  44138=>"000001001",
  44139=>"010110100",
  44140=>"111011010",
  44141=>"111111101",
  44142=>"100010101",
  44143=>"101011110",
  44144=>"111000001",
  44145=>"100000111",
  44146=>"100100110",
  44147=>"110001110",
  44148=>"101100100",
  44149=>"011010010",
  44150=>"101110110",
  44151=>"101000000",
  44152=>"101101001",
  44153=>"110111100",
  44154=>"000001000",
  44155=>"010111011",
  44156=>"110100101",
  44157=>"010000000",
  44158=>"110111001",
  44159=>"110010110",
  44160=>"100000110",
  44161=>"001110101",
  44162=>"110011110",
  44163=>"010111001",
  44164=>"101000111",
  44165=>"010000111",
  44166=>"000000100",
  44167=>"010100101",
  44168=>"101110011",
  44169=>"001111000",
  44170=>"011010110",
  44171=>"001101011",
  44172=>"111100001",
  44173=>"111110010",
  44174=>"111110000",
  44175=>"111011101",
  44176=>"001111010",
  44177=>"110011110",
  44178=>"101010101",
  44179=>"101001011",
  44180=>"010010001",
  44181=>"000101010",
  44182=>"001011000",
  44183=>"010111000",
  44184=>"011001010",
  44185=>"111001001",
  44186=>"000010000",
  44187=>"100110000",
  44188=>"011110001",
  44189=>"000001100",
  44190=>"101010010",
  44191=>"101010000",
  44192=>"110010110",
  44193=>"110111110",
  44194=>"011111001",
  44195=>"001000011",
  44196=>"111101000",
  44197=>"111101111",
  44198=>"101010100",
  44199=>"110001101",
  44200=>"100000110",
  44201=>"111000000",
  44202=>"000011000",
  44203=>"000001001",
  44204=>"001110001",
  44205=>"001100000",
  44206=>"111001100",
  44207=>"110001000",
  44208=>"110000010",
  44209=>"010010100",
  44210=>"111101010",
  44211=>"100001011",
  44212=>"011000010",
  44213=>"000100100",
  44214=>"110110010",
  44215=>"101001011",
  44216=>"100111010",
  44217=>"011100101",
  44218=>"011000011",
  44219=>"100111111",
  44220=>"101110001",
  44221=>"000001101",
  44222=>"111100011",
  44223=>"011011110",
  44224=>"011001001",
  44225=>"110110100",
  44226=>"110110100",
  44227=>"010100100",
  44228=>"011011111",
  44229=>"000001111",
  44230=>"001011111",
  44231=>"010110001",
  44232=>"110111111",
  44233=>"111010000",
  44234=>"100101001",
  44235=>"011100001",
  44236=>"101111101",
  44237=>"101001000",
  44238=>"001101000",
  44239=>"101111111",
  44240=>"001110101",
  44241=>"101111000",
  44242=>"010110001",
  44243=>"110100111",
  44244=>"110110110",
  44245=>"011100011",
  44246=>"011111101",
  44247=>"111100101",
  44248=>"011100010",
  44249=>"011001100",
  44250=>"111010111",
  44251=>"010000110",
  44252=>"111001001",
  44253=>"101111101",
  44254=>"011000111",
  44255=>"101100100",
  44256=>"111001001",
  44257=>"000100111",
  44258=>"000100001",
  44259=>"000111010",
  44260=>"100000000",
  44261=>"010010010",
  44262=>"011001010",
  44263=>"110010110",
  44264=>"111100110",
  44265=>"010111000",
  44266=>"000001111",
  44267=>"110010111",
  44268=>"000010001",
  44269=>"000000101",
  44270=>"010000011",
  44271=>"001100011",
  44272=>"101110101",
  44273=>"111100001",
  44274=>"000000001",
  44275=>"000101000",
  44276=>"000011001",
  44277=>"110100100",
  44278=>"101000100",
  44279=>"101111101",
  44280=>"100011001",
  44281=>"000011101",
  44282=>"100010100",
  44283=>"101010110",
  44284=>"111111101",
  44285=>"011111010",
  44286=>"110000110",
  44287=>"111000110",
  44288=>"010000111",
  44289=>"110110110",
  44290=>"100001111",
  44291=>"001111111",
  44292=>"001000101",
  44293=>"100101001",
  44294=>"110110001",
  44295=>"101101001",
  44296=>"100000100",
  44297=>"111000110",
  44298=>"110110001",
  44299=>"010010101",
  44300=>"110001110",
  44301=>"001101100",
  44302=>"001010011",
  44303=>"001111010",
  44304=>"010001010",
  44305=>"110001101",
  44306=>"010111101",
  44307=>"101101001",
  44308=>"100100000",
  44309=>"010110110",
  44310=>"101011011",
  44311=>"110010111",
  44312=>"111111010",
  44313=>"010101010",
  44314=>"000100011",
  44315=>"101011011",
  44316=>"010011010",
  44317=>"100000111",
  44318=>"000011110",
  44319=>"000111011",
  44320=>"101111101",
  44321=>"111111110",
  44322=>"100110000",
  44323=>"100101001",
  44324=>"000101010",
  44325=>"111000101",
  44326=>"100100111",
  44327=>"101100110",
  44328=>"001110000",
  44329=>"101101101",
  44330=>"111001010",
  44331=>"110100011",
  44332=>"101010001",
  44333=>"111101010",
  44334=>"000001000",
  44335=>"000000010",
  44336=>"110010010",
  44337=>"001000111",
  44338=>"101110100",
  44339=>"010010101",
  44340=>"101001010",
  44341=>"001000010",
  44342=>"010100101",
  44343=>"100111010",
  44344=>"010011001",
  44345=>"011111001",
  44346=>"011010001",
  44347=>"111011011",
  44348=>"110101010",
  44349=>"110000001",
  44350=>"011011010",
  44351=>"111110110",
  44352=>"011111011",
  44353=>"100111111",
  44354=>"110111001",
  44355=>"110010000",
  44356=>"100001101",
  44357=>"010110111",
  44358=>"100001110",
  44359=>"111010100",
  44360=>"010000111",
  44361=>"011101001",
  44362=>"101010001",
  44363=>"010101100",
  44364=>"000101000",
  44365=>"101000110",
  44366=>"110100100",
  44367=>"101110111",
  44368=>"111000011",
  44369=>"000000111",
  44370=>"100001111",
  44371=>"110011011",
  44372=>"010100011",
  44373=>"000101101",
  44374=>"101000010",
  44375=>"011101101",
  44376=>"000110111",
  44377=>"111010101",
  44378=>"010111001",
  44379=>"001000010",
  44380=>"010100100",
  44381=>"101000011",
  44382=>"001011010",
  44383=>"101100110",
  44384=>"001101010",
  44385=>"000100011",
  44386=>"010101011",
  44387=>"111010011",
  44388=>"111001010",
  44389=>"000001010",
  44390=>"100101001",
  44391=>"111110110",
  44392=>"000111001",
  44393=>"000001001",
  44394=>"010011110",
  44395=>"000010100",
  44396=>"011000000",
  44397=>"011001110",
  44398=>"101000011",
  44399=>"100011110",
  44400=>"101011100",
  44401=>"001110000",
  44402=>"110111110",
  44403=>"100000000",
  44404=>"011101000",
  44405=>"010100101",
  44406=>"111100110",
  44407=>"010010001",
  44408=>"111110001",
  44409=>"101111010",
  44410=>"011001111",
  44411=>"110101000",
  44412=>"011010110",
  44413=>"001111111",
  44414=>"010011000",
  44415=>"000101000",
  44416=>"110111000",
  44417=>"010101010",
  44418=>"100101010",
  44419=>"000010000",
  44420=>"001001001",
  44421=>"100000101",
  44422=>"100001011",
  44423=>"101101100",
  44424=>"000101001",
  44425=>"101010101",
  44426=>"100010010",
  44427=>"000001101",
  44428=>"010001011",
  44429=>"111011010",
  44430=>"000111100",
  44431=>"101110101",
  44432=>"110000011",
  44433=>"011100001",
  44434=>"010000111",
  44435=>"010111010",
  44436=>"001010100",
  44437=>"011110100",
  44438=>"010011010",
  44439=>"010010101",
  44440=>"101000001",
  44441=>"001101001",
  44442=>"110111011",
  44443=>"001010010",
  44444=>"111101001",
  44445=>"100001100",
  44446=>"000000011",
  44447=>"001111000",
  44448=>"101001001",
  44449=>"011111110",
  44450=>"110100010",
  44451=>"010001110",
  44452=>"001000101",
  44453=>"111011011",
  44454=>"101100011",
  44455=>"001000011",
  44456=>"111111011",
  44457=>"110000011",
  44458=>"000000110",
  44459=>"000111100",
  44460=>"010010001",
  44461=>"101111000",
  44462=>"101001000",
  44463=>"110101101",
  44464=>"000101010",
  44465=>"010010001",
  44466=>"001000101",
  44467=>"010000010",
  44468=>"110000111",
  44469=>"010110001",
  44470=>"110011111",
  44471=>"101001000",
  44472=>"011001010",
  44473=>"001011000",
  44474=>"110000000",
  44475=>"111111111",
  44476=>"000110010",
  44477=>"000110110",
  44478=>"010001111",
  44479=>"111111000",
  44480=>"000100110",
  44481=>"111111101",
  44482=>"001100101",
  44483=>"010000011",
  44484=>"000000101",
  44485=>"110010110",
  44486=>"101100011",
  44487=>"111111001",
  44488=>"011000000",
  44489=>"000101110",
  44490=>"000011110",
  44491=>"110111011",
  44492=>"100100000",
  44493=>"100000000",
  44494=>"001110101",
  44495=>"111101110",
  44496=>"111111010",
  44497=>"001011001",
  44498=>"010001111",
  44499=>"111011110",
  44500=>"000111000",
  44501=>"001110011",
  44502=>"101100011",
  44503=>"000101010",
  44504=>"101001001",
  44505=>"100010101",
  44506=>"000110010",
  44507=>"111010111",
  44508=>"111001111",
  44509=>"000011111",
  44510=>"111110101",
  44511=>"110010100",
  44512=>"111101100",
  44513=>"011011101",
  44514=>"101101100",
  44515=>"100011001",
  44516=>"101100110",
  44517=>"100011001",
  44518=>"100000100",
  44519=>"110000101",
  44520=>"000010000",
  44521=>"101001101",
  44522=>"110011000",
  44523=>"100111001",
  44524=>"001101011",
  44525=>"000011110",
  44526=>"010110000",
  44527=>"110011111",
  44528=>"101101110",
  44529=>"011000100",
  44530=>"001000110",
  44531=>"001000000",
  44532=>"000110110",
  44533=>"000110010",
  44534=>"111111110",
  44535=>"111001000",
  44536=>"010101010",
  44537=>"000011101",
  44538=>"011010010",
  44539=>"100011010",
  44540=>"101001111",
  44541=>"001111010",
  44542=>"010000110",
  44543=>"010111000",
  44544=>"011110111",
  44545=>"011100111",
  44546=>"000010100",
  44547=>"010001100",
  44548=>"010100101",
  44549=>"110101111",
  44550=>"100001100",
  44551=>"000000000",
  44552=>"010100101",
  44553=>"010010011",
  44554=>"101010010",
  44555=>"000110001",
  44556=>"100110111",
  44557=>"010111111",
  44558=>"010101010",
  44559=>"001001011",
  44560=>"000000111",
  44561=>"001010101",
  44562=>"111011000",
  44563=>"011111010",
  44564=>"000010110",
  44565=>"010001111",
  44566=>"111110001",
  44567=>"001111011",
  44568=>"110000101",
  44569=>"000010011",
  44570=>"100101001",
  44571=>"001111001",
  44572=>"110000110",
  44573=>"101101010",
  44574=>"001111111",
  44575=>"001101110",
  44576=>"000000011",
  44577=>"001111011",
  44578=>"010001111",
  44579=>"000110000",
  44580=>"110011000",
  44581=>"100011111",
  44582=>"011110110",
  44583=>"100001000",
  44584=>"011001100",
  44585=>"001111010",
  44586=>"011010111",
  44587=>"011110001",
  44588=>"110111000",
  44589=>"101110010",
  44590=>"101000100",
  44591=>"000000110",
  44592=>"000010001",
  44593=>"111100101",
  44594=>"000111000",
  44595=>"010000101",
  44596=>"110101000",
  44597=>"111111111",
  44598=>"101111111",
  44599=>"011110001",
  44600=>"101001111",
  44601=>"011000101",
  44602=>"101101000",
  44603=>"000101001",
  44604=>"101001011",
  44605=>"010000010",
  44606=>"101110001",
  44607=>"001001100",
  44608=>"010001010",
  44609=>"111010001",
  44610=>"011101100",
  44611=>"100000010",
  44612=>"000011000",
  44613=>"001111111",
  44614=>"001101000",
  44615=>"010101100",
  44616=>"111011111",
  44617=>"000101111",
  44618=>"100000010",
  44619=>"100010111",
  44620=>"111001100",
  44621=>"010010010",
  44622=>"000100000",
  44623=>"000010110",
  44624=>"100110111",
  44625=>"111001001",
  44626=>"100110010",
  44627=>"001111110",
  44628=>"001101000",
  44629=>"010001000",
  44630=>"111110001",
  44631=>"101001100",
  44632=>"101001000",
  44633=>"010001010",
  44634=>"011110111",
  44635=>"111011111",
  44636=>"101100100",
  44637=>"110011111",
  44638=>"001101110",
  44639=>"101100110",
  44640=>"011100110",
  44641=>"111000000",
  44642=>"100011001",
  44643=>"001111000",
  44644=>"101100110",
  44645=>"111110100",
  44646=>"101111000",
  44647=>"001011111",
  44648=>"011000000",
  44649=>"100011000",
  44650=>"000101111",
  44651=>"000000001",
  44652=>"011111011",
  44653=>"010110011",
  44654=>"111100110",
  44655=>"011100000",
  44656=>"010111011",
  44657=>"111111111",
  44658=>"110011100",
  44659=>"010111010",
  44660=>"010101101",
  44661=>"101010000",
  44662=>"011000100",
  44663=>"010111100",
  44664=>"000000110",
  44665=>"000100011",
  44666=>"100001010",
  44667=>"111110101",
  44668=>"111011110",
  44669=>"101101100",
  44670=>"010111000",
  44671=>"011011101",
  44672=>"011110110",
  44673=>"101111000",
  44674=>"011010010",
  44675=>"101000111",
  44676=>"010001010",
  44677=>"111001100",
  44678=>"000001100",
  44679=>"100111111",
  44680=>"011110111",
  44681=>"011101000",
  44682=>"011011100",
  44683=>"001101101",
  44684=>"000100100",
  44685=>"101101010",
  44686=>"011001010",
  44687=>"010010111",
  44688=>"001110010",
  44689=>"111011101",
  44690=>"101101011",
  44691=>"110010000",
  44692=>"101100111",
  44693=>"111110011",
  44694=>"010100110",
  44695=>"101111000",
  44696=>"101010000",
  44697=>"001110001",
  44698=>"000110001",
  44699=>"010000011",
  44700=>"001100000",
  44701=>"111000101",
  44702=>"101100111",
  44703=>"011101110",
  44704=>"001010000",
  44705=>"010111101",
  44706=>"001110101",
  44707=>"000001011",
  44708=>"011101001",
  44709=>"010010110",
  44710=>"001100011",
  44711=>"011100101",
  44712=>"000010110",
  44713=>"011011110",
  44714=>"000000010",
  44715=>"011100100",
  44716=>"010011101",
  44717=>"100101101",
  44718=>"101000101",
  44719=>"011010000",
  44720=>"101001101",
  44721=>"010010011",
  44722=>"111110110",
  44723=>"010010101",
  44724=>"101011100",
  44725=>"000110111",
  44726=>"101001011",
  44727=>"111000010",
  44728=>"100001000",
  44729=>"011010011",
  44730=>"101010000",
  44731=>"000100101",
  44732=>"000110111",
  44733=>"111011100",
  44734=>"000001111",
  44735=>"111000010",
  44736=>"000000011",
  44737=>"101111111",
  44738=>"111010010",
  44739=>"000011111",
  44740=>"010010001",
  44741=>"100110101",
  44742=>"001011101",
  44743=>"010110010",
  44744=>"001001110",
  44745=>"110011011",
  44746=>"000110001",
  44747=>"011110000",
  44748=>"111011100",
  44749=>"110011100",
  44750=>"100010010",
  44751=>"000010010",
  44752=>"010001010",
  44753=>"001011101",
  44754=>"100011100",
  44755=>"100110010",
  44756=>"001011111",
  44757=>"101011010",
  44758=>"101000001",
  44759=>"011110011",
  44760=>"001000011",
  44761=>"011111000",
  44762=>"101111001",
  44763=>"110010011",
  44764=>"000010101",
  44765=>"011011100",
  44766=>"100001111",
  44767=>"100011110",
  44768=>"111011100",
  44769=>"001010000",
  44770=>"011010000",
  44771=>"101000110",
  44772=>"100110010",
  44773=>"000110000",
  44774=>"101101101",
  44775=>"011011000",
  44776=>"110101010",
  44777=>"101111111",
  44778=>"011011100",
  44779=>"000100000",
  44780=>"100101101",
  44781=>"010010011",
  44782=>"100011011",
  44783=>"100011010",
  44784=>"100100100",
  44785=>"101100110",
  44786=>"110000101",
  44787=>"011001111",
  44788=>"010011101",
  44789=>"001100111",
  44790=>"000101010",
  44791=>"010010011",
  44792=>"010001111",
  44793=>"010111111",
  44794=>"101110010",
  44795=>"000101100",
  44796=>"101100000",
  44797=>"111100000",
  44798=>"100000010",
  44799=>"011000000",
  44800=>"000110110",
  44801=>"100011110",
  44802=>"101001000",
  44803=>"000001111",
  44804=>"000100000",
  44805=>"011010000",
  44806=>"111011110",
  44807=>"011010100",
  44808=>"111011101",
  44809=>"101001101",
  44810=>"011100101",
  44811=>"111010100",
  44812=>"111000100",
  44813=>"011001011",
  44814=>"100101101",
  44815=>"101010011",
  44816=>"011101010",
  44817=>"101110010",
  44818=>"001010001",
  44819=>"001001001",
  44820=>"011001001",
  44821=>"010100110",
  44822=>"110100000",
  44823=>"111100001",
  44824=>"101010001",
  44825=>"010010111",
  44826=>"110000011",
  44827=>"011110001",
  44828=>"110000111",
  44829=>"000100011",
  44830=>"111000010",
  44831=>"000000111",
  44832=>"111010111",
  44833=>"110000010",
  44834=>"110001111",
  44835=>"111000001",
  44836=>"010110001",
  44837=>"001101101",
  44838=>"000000110",
  44839=>"000111011",
  44840=>"110001000",
  44841=>"100111100",
  44842=>"100001001",
  44843=>"010100011",
  44844=>"000010110",
  44845=>"100101101",
  44846=>"101000111",
  44847=>"000001011",
  44848=>"100111001",
  44849=>"101000011",
  44850=>"111111010",
  44851=>"101010101",
  44852=>"001000010",
  44853=>"001000100",
  44854=>"000110011",
  44855=>"100001000",
  44856=>"010001101",
  44857=>"011000000",
  44858=>"101010001",
  44859=>"001110110",
  44860=>"111001001",
  44861=>"111100110",
  44862=>"010000110",
  44863=>"010001110",
  44864=>"111110100",
  44865=>"001011111",
  44866=>"001000011",
  44867=>"011000100",
  44868=>"100001000",
  44869=>"001000001",
  44870=>"111100111",
  44871=>"001001110",
  44872=>"101000010",
  44873=>"011011100",
  44874=>"100001111",
  44875=>"110011011",
  44876=>"011101100",
  44877=>"010101010",
  44878=>"011111111",
  44879=>"100011101",
  44880=>"010001110",
  44881=>"011000000",
  44882=>"001101110",
  44883=>"111100111",
  44884=>"110000111",
  44885=>"000000001",
  44886=>"001100010",
  44887=>"000001110",
  44888=>"111100111",
  44889=>"101001100",
  44890=>"001111100",
  44891=>"011101101",
  44892=>"110010100",
  44893=>"101100111",
  44894=>"001110111",
  44895=>"000111010",
  44896=>"101001110",
  44897=>"101110000",
  44898=>"001001000",
  44899=>"001110011",
  44900=>"010000100",
  44901=>"111001100",
  44902=>"111111100",
  44903=>"000111110",
  44904=>"000000000",
  44905=>"011000100",
  44906=>"110111001",
  44907=>"110001111",
  44908=>"110001001",
  44909=>"000000000",
  44910=>"011011011",
  44911=>"010100000",
  44912=>"001010101",
  44913=>"010000000",
  44914=>"111001101",
  44915=>"000101000",
  44916=>"101011001",
  44917=>"111110100",
  44918=>"110000110",
  44919=>"000111011",
  44920=>"000001110",
  44921=>"000010100",
  44922=>"111101010",
  44923=>"000010010",
  44924=>"000010100",
  44925=>"000010010",
  44926=>"101010110",
  44927=>"001100110",
  44928=>"101101110",
  44929=>"010010001",
  44930=>"001001101",
  44931=>"110000101",
  44932=>"100100101",
  44933=>"010100001",
  44934=>"000011110",
  44935=>"100000110",
  44936=>"010011011",
  44937=>"110000000",
  44938=>"100111011",
  44939=>"111000001",
  44940=>"110110110",
  44941=>"111111001",
  44942=>"111111001",
  44943=>"000001100",
  44944=>"000100001",
  44945=>"000001111",
  44946=>"011101111",
  44947=>"100011001",
  44948=>"110001101",
  44949=>"011001111",
  44950=>"110111010",
  44951=>"111100111",
  44952=>"011001101",
  44953=>"010000001",
  44954=>"001011010",
  44955=>"100011101",
  44956=>"001111010",
  44957=>"101001011",
  44958=>"100010000",
  44959=>"100001010",
  44960=>"101001110",
  44961=>"010110111",
  44962=>"011100110",
  44963=>"101101001",
  44964=>"010001000",
  44965=>"001000011",
  44966=>"001111001",
  44967=>"001011000",
  44968=>"010110110",
  44969=>"100001000",
  44970=>"101000010",
  44971=>"010000111",
  44972=>"101011010",
  44973=>"011111110",
  44974=>"101101011",
  44975=>"000001001",
  44976=>"010011100",
  44977=>"111111100",
  44978=>"001010100",
  44979=>"000100101",
  44980=>"110010011",
  44981=>"001010100",
  44982=>"100000001",
  44983=>"111111010",
  44984=>"001100110",
  44985=>"111011111",
  44986=>"101011100",
  44987=>"100111111",
  44988=>"001101000",
  44989=>"001111101",
  44990=>"101111111",
  44991=>"011011000",
  44992=>"010111110",
  44993=>"111111010",
  44994=>"101000100",
  44995=>"110000100",
  44996=>"010110000",
  44997=>"111001110",
  44998=>"010010000",
  44999=>"101111110",
  45000=>"000000100",
  45001=>"111000001",
  45002=>"111001101",
  45003=>"010101101",
  45004=>"001101101",
  45005=>"001100001",
  45006=>"000001100",
  45007=>"110110011",
  45008=>"110110000",
  45009=>"111000001",
  45010=>"010010101",
  45011=>"001101010",
  45012=>"001111001",
  45013=>"001111100",
  45014=>"110101011",
  45015=>"101001110",
  45016=>"010011001",
  45017=>"111011011",
  45018=>"011111111",
  45019=>"011111110",
  45020=>"000010000",
  45021=>"111111011",
  45022=>"101101011",
  45023=>"001011111",
  45024=>"001010001",
  45025=>"110000000",
  45026=>"110010000",
  45027=>"110010000",
  45028=>"000100001",
  45029=>"000101111",
  45030=>"001001001",
  45031=>"101010000",
  45032=>"111000100",
  45033=>"101100110",
  45034=>"101010001",
  45035=>"000010000",
  45036=>"110100101",
  45037=>"110100110",
  45038=>"111011100",
  45039=>"111110110",
  45040=>"000111010",
  45041=>"011100010",
  45042=>"111011111",
  45043=>"110111110",
  45044=>"101011111",
  45045=>"111111111",
  45046=>"000111011",
  45047=>"111011011",
  45048=>"010100101",
  45049=>"110001000",
  45050=>"001101100",
  45051=>"011011001",
  45052=>"000010010",
  45053=>"100001001",
  45054=>"100011111",
  45055=>"100010000",
  45056=>"000000010",
  45057=>"101111001",
  45058=>"111011001",
  45059=>"111000000",
  45060=>"000100000",
  45061=>"000100111",
  45062=>"100011000",
  45063=>"100001000",
  45064=>"010110111",
  45065=>"010110000",
  45066=>"011101101",
  45067=>"100111011",
  45068=>"101001101",
  45069=>"000101010",
  45070=>"011000100",
  45071=>"101011101",
  45072=>"110100010",
  45073=>"000000100",
  45074=>"010001110",
  45075=>"011000001",
  45076=>"111010010",
  45077=>"010110101",
  45078=>"010110000",
  45079=>"101001000",
  45080=>"010111011",
  45081=>"001001010",
  45082=>"000011100",
  45083=>"110111101",
  45084=>"111001000",
  45085=>"100010110",
  45086=>"111110000",
  45087=>"111101011",
  45088=>"001000100",
  45089=>"000010101",
  45090=>"010100100",
  45091=>"010010011",
  45092=>"101001011",
  45093=>"010110011",
  45094=>"001011111",
  45095=>"010000100",
  45096=>"101100000",
  45097=>"111101110",
  45098=>"110000001",
  45099=>"011101111",
  45100=>"000000000",
  45101=>"001111110",
  45102=>"100011101",
  45103=>"101001010",
  45104=>"011011100",
  45105=>"011011101",
  45106=>"100101011",
  45107=>"011111111",
  45108=>"101010000",
  45109=>"100111101",
  45110=>"011000111",
  45111=>"010011100",
  45112=>"001001000",
  45113=>"010001111",
  45114=>"010110001",
  45115=>"111010101",
  45116=>"001000010",
  45117=>"000101000",
  45118=>"101011011",
  45119=>"010100011",
  45120=>"110011010",
  45121=>"100000010",
  45122=>"110001100",
  45123=>"111001100",
  45124=>"110110101",
  45125=>"001011011",
  45126=>"110101110",
  45127=>"111000110",
  45128=>"010100110",
  45129=>"000111011",
  45130=>"111010101",
  45131=>"001000101",
  45132=>"001110101",
  45133=>"010110010",
  45134=>"010111011",
  45135=>"001110110",
  45136=>"001010001",
  45137=>"001010100",
  45138=>"000111101",
  45139=>"010011110",
  45140=>"000010100",
  45141=>"010001000",
  45142=>"011001000",
  45143=>"110000110",
  45144=>"011111000",
  45145=>"100010010",
  45146=>"101000010",
  45147=>"000011101",
  45148=>"111011111",
  45149=>"000000011",
  45150=>"000001111",
  45151=>"100000111",
  45152=>"111011001",
  45153=>"001111000",
  45154=>"010000001",
  45155=>"000000100",
  45156=>"110001000",
  45157=>"100011011",
  45158=>"000011010",
  45159=>"010101010",
  45160=>"110110011",
  45161=>"001010101",
  45162=>"111000111",
  45163=>"000011010",
  45164=>"110010000",
  45165=>"001000100",
  45166=>"010100110",
  45167=>"101001111",
  45168=>"010001001",
  45169=>"001101111",
  45170=>"111101101",
  45171=>"001000010",
  45172=>"111011001",
  45173=>"110000001",
  45174=>"010010000",
  45175=>"100011011",
  45176=>"111111000",
  45177=>"010011011",
  45178=>"001100111",
  45179=>"011011000",
  45180=>"110001011",
  45181=>"011100100",
  45182=>"110110011",
  45183=>"000100000",
  45184=>"011111111",
  45185=>"111101010",
  45186=>"000110001",
  45187=>"011101101",
  45188=>"010001000",
  45189=>"000100110",
  45190=>"111011001",
  45191=>"111000001",
  45192=>"011111101",
  45193=>"011010101",
  45194=>"000011100",
  45195=>"011111110",
  45196=>"011011001",
  45197=>"011100101",
  45198=>"111010110",
  45199=>"001011111",
  45200=>"010000000",
  45201=>"001000001",
  45202=>"110110101",
  45203=>"111100010",
  45204=>"000000001",
  45205=>"110011011",
  45206=>"110101000",
  45207=>"100000000",
  45208=>"010001011",
  45209=>"011010111",
  45210=>"001100110",
  45211=>"101111000",
  45212=>"110010100",
  45213=>"010101011",
  45214=>"111001011",
  45215=>"111110010",
  45216=>"111100101",
  45217=>"010001111",
  45218=>"111111000",
  45219=>"001010101",
  45220=>"001111100",
  45221=>"001011111",
  45222=>"010011000",
  45223=>"110001111",
  45224=>"100101001",
  45225=>"001001010",
  45226=>"101011011",
  45227=>"010100010",
  45228=>"001101100",
  45229=>"010000101",
  45230=>"001100100",
  45231=>"110011001",
  45232=>"110001011",
  45233=>"110010111",
  45234=>"001000111",
  45235=>"010010000",
  45236=>"011000000",
  45237=>"110111000",
  45238=>"111101011",
  45239=>"111101101",
  45240=>"001100101",
  45241=>"001001000",
  45242=>"001110100",
  45243=>"000001110",
  45244=>"100101000",
  45245=>"010010110",
  45246=>"000011111",
  45247=>"100001000",
  45248=>"011010100",
  45249=>"101000011",
  45250=>"111000000",
  45251=>"111101000",
  45252=>"011111010",
  45253=>"101101011",
  45254=>"111110010",
  45255=>"111000110",
  45256=>"100111101",
  45257=>"010001001",
  45258=>"010011011",
  45259=>"011111111",
  45260=>"000101100",
  45261=>"010011010",
  45262=>"100101010",
  45263=>"001101111",
  45264=>"110101000",
  45265=>"111001000",
  45266=>"010001000",
  45267=>"111111110",
  45268=>"011000010",
  45269=>"000000010",
  45270=>"110111101",
  45271=>"000111100",
  45272=>"100111101",
  45273=>"010000001",
  45274=>"010100101",
  45275=>"011100011",
  45276=>"111011101",
  45277=>"011111111",
  45278=>"000101000",
  45279=>"101101111",
  45280=>"100111111",
  45281=>"010010000",
  45282=>"011100110",
  45283=>"101000110",
  45284=>"111000110",
  45285=>"100010000",
  45286=>"000000000",
  45287=>"100110100",
  45288=>"000111110",
  45289=>"010111000",
  45290=>"001000100",
  45291=>"111101110",
  45292=>"010010001",
  45293=>"001010010",
  45294=>"000100010",
  45295=>"001000101",
  45296=>"111010001",
  45297=>"101010111",
  45298=>"100000011",
  45299=>"100001000",
  45300=>"010001001",
  45301=>"100010000",
  45302=>"111000000",
  45303=>"010011110",
  45304=>"101011110",
  45305=>"011100110",
  45306=>"100010010",
  45307=>"010000110",
  45308=>"111011000",
  45309=>"100001110",
  45310=>"111000001",
  45311=>"000011100",
  45312=>"101111100",
  45313=>"011111111",
  45314=>"100001011",
  45315=>"100010110",
  45316=>"110000111",
  45317=>"000001000",
  45318=>"011011011",
  45319=>"011111011",
  45320=>"101000000",
  45321=>"001011110",
  45322=>"100111001",
  45323=>"100100010",
  45324=>"001110111",
  45325=>"010010000",
  45326=>"010011011",
  45327=>"000001100",
  45328=>"110110001",
  45329=>"100100011",
  45330=>"101101000",
  45331=>"100000110",
  45332=>"100100011",
  45333=>"001010110",
  45334=>"001000110",
  45335=>"101001001",
  45336=>"101101001",
  45337=>"000101110",
  45338=>"101100101",
  45339=>"010000101",
  45340=>"010000010",
  45341=>"000000001",
  45342=>"010001110",
  45343=>"001101101",
  45344=>"010110101",
  45345=>"001011101",
  45346=>"111110010",
  45347=>"101011000",
  45348=>"000001110",
  45349=>"000010101",
  45350=>"000000001",
  45351=>"100110011",
  45352=>"110110100",
  45353=>"001000100",
  45354=>"111100111",
  45355=>"101110101",
  45356=>"001100000",
  45357=>"011000001",
  45358=>"101101000",
  45359=>"000010001",
  45360=>"001001000",
  45361=>"111110000",
  45362=>"011001101",
  45363=>"100011000",
  45364=>"010110001",
  45365=>"010011001",
  45366=>"011010100",
  45367=>"010010101",
  45368=>"010100101",
  45369=>"111011111",
  45370=>"111110001",
  45371=>"000010011",
  45372=>"100001000",
  45373=>"010000100",
  45374=>"010001001",
  45375=>"110111001",
  45376=>"100101010",
  45377=>"110010100",
  45378=>"011110011",
  45379=>"001000101",
  45380=>"001010000",
  45381=>"010100101",
  45382=>"000010001",
  45383=>"011001101",
  45384=>"111111011",
  45385=>"001001010",
  45386=>"110000010",
  45387=>"000111110",
  45388=>"000110100",
  45389=>"001101011",
  45390=>"000101111",
  45391=>"111011010",
  45392=>"100111100",
  45393=>"010100010",
  45394=>"010000001",
  45395=>"111010001",
  45396=>"000000100",
  45397=>"000100000",
  45398=>"010011111",
  45399=>"100111101",
  45400=>"100011100",
  45401=>"100010010",
  45402=>"010110100",
  45403=>"000000001",
  45404=>"000010100",
  45405=>"010011000",
  45406=>"101110010",
  45407=>"001011001",
  45408=>"110011001",
  45409=>"000101001",
  45410=>"100111010",
  45411=>"001000100",
  45412=>"010111000",
  45413=>"110000011",
  45414=>"101010010",
  45415=>"011000111",
  45416=>"001010000",
  45417=>"110100101",
  45418=>"101001111",
  45419=>"101011001",
  45420=>"110011110",
  45421=>"000000101",
  45422=>"101001111",
  45423=>"100000011",
  45424=>"110001000",
  45425=>"111101010",
  45426=>"010110010",
  45427=>"000001001",
  45428=>"001011110",
  45429=>"011110111",
  45430=>"011101000",
  45431=>"100010000",
  45432=>"100111011",
  45433=>"011010011",
  45434=>"011010110",
  45435=>"010111101",
  45436=>"000010000",
  45437=>"001011010",
  45438=>"110010011",
  45439=>"111000110",
  45440=>"110101010",
  45441=>"111000000",
  45442=>"001110110",
  45443=>"000010101",
  45444=>"111011100",
  45445=>"000000001",
  45446=>"101100110",
  45447=>"111111011",
  45448=>"011010011",
  45449=>"010000001",
  45450=>"001111000",
  45451=>"111101001",
  45452=>"101010001",
  45453=>"111001010",
  45454=>"111101111",
  45455=>"000111110",
  45456=>"001010001",
  45457=>"101101111",
  45458=>"111011011",
  45459=>"101011010",
  45460=>"100111011",
  45461=>"011010101",
  45462=>"001000111",
  45463=>"111111111",
  45464=>"001010110",
  45465=>"111101010",
  45466=>"011000011",
  45467=>"000011110",
  45468=>"110100011",
  45469=>"101011001",
  45470=>"110101001",
  45471=>"011111011",
  45472=>"000101110",
  45473=>"001101011",
  45474=>"111101110",
  45475=>"110000000",
  45476=>"010110100",
  45477=>"000101101",
  45478=>"010110010",
  45479=>"011110011",
  45480=>"000011110",
  45481=>"001111000",
  45482=>"110101001",
  45483=>"100001111",
  45484=>"000001001",
  45485=>"000011010",
  45486=>"100100010",
  45487=>"100010101",
  45488=>"101011111",
  45489=>"000000010",
  45490=>"110010010",
  45491=>"010001110",
  45492=>"110100010",
  45493=>"100111111",
  45494=>"101110110",
  45495=>"001001000",
  45496=>"101000000",
  45497=>"001111001",
  45498=>"100101110",
  45499=>"100100100",
  45500=>"001110111",
  45501=>"100010011",
  45502=>"000001011",
  45503=>"100111011",
  45504=>"110101100",
  45505=>"000001011",
  45506=>"000101101",
  45507=>"110111101",
  45508=>"100111100",
  45509=>"000000101",
  45510=>"000010000",
  45511=>"101011111",
  45512=>"010101111",
  45513=>"100110110",
  45514=>"111110110",
  45515=>"001101011",
  45516=>"100100101",
  45517=>"111011000",
  45518=>"010000001",
  45519=>"000000010",
  45520=>"001001110",
  45521=>"001011000",
  45522=>"000101110",
  45523=>"111000111",
  45524=>"011101000",
  45525=>"001011111",
  45526=>"101101010",
  45527=>"101010000",
  45528=>"100010000",
  45529=>"111101110",
  45530=>"101000101",
  45531=>"010001101",
  45532=>"111111100",
  45533=>"110100011",
  45534=>"100101011",
  45535=>"100101110",
  45536=>"101110101",
  45537=>"110111100",
  45538=>"001000001",
  45539=>"010100110",
  45540=>"100000111",
  45541=>"010010000",
  45542=>"001001011",
  45543=>"101101011",
  45544=>"101010000",
  45545=>"100010011",
  45546=>"111001011",
  45547=>"111101111",
  45548=>"111011110",
  45549=>"110011100",
  45550=>"101001001",
  45551=>"111001100",
  45552=>"111111001",
  45553=>"111100010",
  45554=>"011011100",
  45555=>"010000000",
  45556=>"000110110",
  45557=>"000101111",
  45558=>"011101010",
  45559=>"110100010",
  45560=>"010110111",
  45561=>"111001110",
  45562=>"010000010",
  45563=>"010001101",
  45564=>"011101011",
  45565=>"000010001",
  45566=>"000100101",
  45567=>"111110111",
  45568=>"100000101",
  45569=>"000111000",
  45570=>"001101111",
  45571=>"000100011",
  45572=>"111111110",
  45573=>"111111011",
  45574=>"001111010",
  45575=>"000000010",
  45576=>"010011011",
  45577=>"100010110",
  45578=>"101010101",
  45579=>"100001011",
  45580=>"100101111",
  45581=>"111100100",
  45582=>"010110010",
  45583=>"110110101",
  45584=>"100011101",
  45585=>"010011001",
  45586=>"101010100",
  45587=>"100011110",
  45588=>"011110100",
  45589=>"110000110",
  45590=>"011001110",
  45591=>"010111101",
  45592=>"001000110",
  45593=>"001111000",
  45594=>"110001010",
  45595=>"011011101",
  45596=>"110101001",
  45597=>"101001001",
  45598=>"010100000",
  45599=>"000110001",
  45600=>"101100010",
  45601=>"101111101",
  45602=>"011000101",
  45603=>"100110011",
  45604=>"000111000",
  45605=>"000101100",
  45606=>"110111100",
  45607=>"001100001",
  45608=>"101111000",
  45609=>"010010001",
  45610=>"001000111",
  45611=>"111010010",
  45612=>"011011000",
  45613=>"011001100",
  45614=>"010100011",
  45615=>"110010010",
  45616=>"100010010",
  45617=>"101010001",
  45618=>"000001111",
  45619=>"110010111",
  45620=>"110111110",
  45621=>"000110011",
  45622=>"100000101",
  45623=>"111110111",
  45624=>"101101000",
  45625=>"000000001",
  45626=>"010110001",
  45627=>"010100111",
  45628=>"010100001",
  45629=>"001001101",
  45630=>"101000101",
  45631=>"000100100",
  45632=>"010111001",
  45633=>"000111101",
  45634=>"000110010",
  45635=>"111011011",
  45636=>"000000001",
  45637=>"011000110",
  45638=>"100111001",
  45639=>"010110010",
  45640=>"010001011",
  45641=>"100010010",
  45642=>"001000101",
  45643=>"100110100",
  45644=>"101000110",
  45645=>"000010010",
  45646=>"011111010",
  45647=>"000101110",
  45648=>"011000010",
  45649=>"111111011",
  45650=>"111000000",
  45651=>"010110100",
  45652=>"000001111",
  45653=>"101000111",
  45654=>"011000100",
  45655=>"010101001",
  45656=>"100101011",
  45657=>"100000011",
  45658=>"111101110",
  45659=>"000001100",
  45660=>"111000100",
  45661=>"111100000",
  45662=>"000011101",
  45663=>"100110100",
  45664=>"101000001",
  45665=>"111100101",
  45666=>"101111011",
  45667=>"100010100",
  45668=>"011101101",
  45669=>"000000001",
  45670=>"000101100",
  45671=>"001000011",
  45672=>"101101100",
  45673=>"111110000",
  45674=>"111011110",
  45675=>"100010000",
  45676=>"000001011",
  45677=>"100111010",
  45678=>"000110111",
  45679=>"100101111",
  45680=>"101111001",
  45681=>"010001100",
  45682=>"111110001",
  45683=>"101111110",
  45684=>"011100010",
  45685=>"110001011",
  45686=>"000111110",
  45687=>"000011110",
  45688=>"000101101",
  45689=>"101001101",
  45690=>"111110101",
  45691=>"011101111",
  45692=>"000010010",
  45693=>"010100110",
  45694=>"000010000",
  45695=>"011010011",
  45696=>"000101000",
  45697=>"011100111",
  45698=>"100011110",
  45699=>"001000001",
  45700=>"101110111",
  45701=>"101100101",
  45702=>"101001100",
  45703=>"000101111",
  45704=>"001100000",
  45705=>"100000001",
  45706=>"101111011",
  45707=>"100101100",
  45708=>"100000100",
  45709=>"001100101",
  45710=>"000111111",
  45711=>"111110001",
  45712=>"100011110",
  45713=>"010111010",
  45714=>"111100111",
  45715=>"001100100",
  45716=>"100101000",
  45717=>"000111000",
  45718=>"100100010",
  45719=>"110100101",
  45720=>"111010001",
  45721=>"010000001",
  45722=>"100000001",
  45723=>"001110110",
  45724=>"000110000",
  45725=>"100001100",
  45726=>"110010000",
  45727=>"001100001",
  45728=>"001010110",
  45729=>"111100001",
  45730=>"010100110",
  45731=>"010111101",
  45732=>"000110000",
  45733=>"010001000",
  45734=>"111110110",
  45735=>"000110000",
  45736=>"110111010",
  45737=>"001010111",
  45738=>"101000010",
  45739=>"001011000",
  45740=>"001001100",
  45741=>"000110100",
  45742=>"000111000",
  45743=>"111001111",
  45744=>"000100100",
  45745=>"100001010",
  45746=>"101010000",
  45747=>"010001111",
  45748=>"100101010",
  45749=>"111011101",
  45750=>"101011110",
  45751=>"000111010",
  45752=>"111101110",
  45753=>"000001100",
  45754=>"111001101",
  45755=>"110010101",
  45756=>"010001111",
  45757=>"110000000",
  45758=>"001000110",
  45759=>"011010101",
  45760=>"000010000",
  45761=>"111000010",
  45762=>"000110000",
  45763=>"000010000",
  45764=>"111110111",
  45765=>"000000100",
  45766=>"111110110",
  45767=>"000001010",
  45768=>"111011111",
  45769=>"100011100",
  45770=>"100101011",
  45771=>"001100001",
  45772=>"110100110",
  45773=>"000100001",
  45774=>"100011101",
  45775=>"000100001",
  45776=>"111111110",
  45777=>"100010100",
  45778=>"010110111",
  45779=>"110101100",
  45780=>"000000100",
  45781=>"000000100",
  45782=>"110011110",
  45783=>"101011101",
  45784=>"000000100",
  45785=>"011111110",
  45786=>"100000101",
  45787=>"111101011",
  45788=>"100001100",
  45789=>"011000110",
  45790=>"111110100",
  45791=>"001100101",
  45792=>"100110111",
  45793=>"010001100",
  45794=>"000010010",
  45795=>"101100111",
  45796=>"111010001",
  45797=>"110110101",
  45798=>"010100010",
  45799=>"001110110",
  45800=>"101110110",
  45801=>"111111111",
  45802=>"010100000",
  45803=>"000110001",
  45804=>"111110010",
  45805=>"001101101",
  45806=>"100111001",
  45807=>"011001111",
  45808=>"010000100",
  45809=>"101001011",
  45810=>"100010010",
  45811=>"110111000",
  45812=>"111011111",
  45813=>"100011110",
  45814=>"110110111",
  45815=>"111011010",
  45816=>"100110000",
  45817=>"100001001",
  45818=>"000000001",
  45819=>"010001101",
  45820=>"101000011",
  45821=>"011001001",
  45822=>"110110001",
  45823=>"110010001",
  45824=>"000000011",
  45825=>"000011011",
  45826=>"110101111",
  45827=>"001010101",
  45828=>"001101100",
  45829=>"000011001",
  45830=>"001010111",
  45831=>"110010001",
  45832=>"110001010",
  45833=>"101110110",
  45834=>"000001010",
  45835=>"100111101",
  45836=>"011011001",
  45837=>"100011101",
  45838=>"111011000",
  45839=>"011001110",
  45840=>"101010011",
  45841=>"101110000",
  45842=>"010110010",
  45843=>"010100111",
  45844=>"000000010",
  45845=>"100101010",
  45846=>"000101100",
  45847=>"110100111",
  45848=>"110000100",
  45849=>"000101000",
  45850=>"000000110",
  45851=>"100011010",
  45852=>"101011010",
  45853=>"111011100",
  45854=>"001000010",
  45855=>"101110111",
  45856=>"011001101",
  45857=>"101110110",
  45858=>"000110110",
  45859=>"110100000",
  45860=>"001111001",
  45861=>"100100110",
  45862=>"001111000",
  45863=>"111011001",
  45864=>"010000000",
  45865=>"100100110",
  45866=>"000100110",
  45867=>"001100111",
  45868=>"111111000",
  45869=>"010011011",
  45870=>"111111011",
  45871=>"000100011",
  45872=>"010111101",
  45873=>"001101011",
  45874=>"100101000",
  45875=>"011001010",
  45876=>"010101111",
  45877=>"110011000",
  45878=>"010000000",
  45879=>"011111101",
  45880=>"010100001",
  45881=>"100101010",
  45882=>"011111001",
  45883=>"111011110",
  45884=>"000000100",
  45885=>"001111000",
  45886=>"000111011",
  45887=>"010000111",
  45888=>"001100110",
  45889=>"000100110",
  45890=>"100100011",
  45891=>"001011000",
  45892=>"111101010",
  45893=>"010100001",
  45894=>"010010001",
  45895=>"010001001",
  45896=>"101110110",
  45897=>"000001110",
  45898=>"001011000",
  45899=>"110101001",
  45900=>"101111000",
  45901=>"011110011",
  45902=>"010010101",
  45903=>"110100000",
  45904=>"110010011",
  45905=>"111011110",
  45906=>"111000101",
  45907=>"000001101",
  45908=>"010010000",
  45909=>"110010000",
  45910=>"000000101",
  45911=>"011110000",
  45912=>"000100011",
  45913=>"110101111",
  45914=>"011101100",
  45915=>"100011000",
  45916=>"111101101",
  45917=>"110000110",
  45918=>"000001001",
  45919=>"000000101",
  45920=>"111001001",
  45921=>"001100010",
  45922=>"111000101",
  45923=>"000010001",
  45924=>"100110010",
  45925=>"000100100",
  45926=>"000101111",
  45927=>"001100111",
  45928=>"111001100",
  45929=>"011100011",
  45930=>"111110010",
  45931=>"000011000",
  45932=>"011001011",
  45933=>"001011100",
  45934=>"001000000",
  45935=>"100111001",
  45936=>"001111011",
  45937=>"011111111",
  45938=>"000000111",
  45939=>"000000010",
  45940=>"111111010",
  45941=>"100001111",
  45942=>"111101111",
  45943=>"010001000",
  45944=>"110011001",
  45945=>"110010100",
  45946=>"010101000",
  45947=>"010000110",
  45948=>"000001000",
  45949=>"111100110",
  45950=>"101100111",
  45951=>"100111010",
  45952=>"100010110",
  45953=>"010000000",
  45954=>"111000101",
  45955=>"111011011",
  45956=>"100001000",
  45957=>"010000011",
  45958=>"110101000",
  45959=>"000100000",
  45960=>"100011001",
  45961=>"001000110",
  45962=>"100001100",
  45963=>"100001000",
  45964=>"101110010",
  45965=>"111111100",
  45966=>"100101001",
  45967=>"011110011",
  45968=>"001010011",
  45969=>"000011100",
  45970=>"011111000",
  45971=>"000010001",
  45972=>"110110000",
  45973=>"001011000",
  45974=>"000000011",
  45975=>"000011010",
  45976=>"101100111",
  45977=>"111100111",
  45978=>"011111110",
  45979=>"101111100",
  45980=>"110000101",
  45981=>"111010110",
  45982=>"010100101",
  45983=>"110010001",
  45984=>"111001111",
  45985=>"110100110",
  45986=>"110110011",
  45987=>"011110111",
  45988=>"111000110",
  45989=>"110111000",
  45990=>"010011010",
  45991=>"111111100",
  45992=>"110101101",
  45993=>"101110010",
  45994=>"011011000",
  45995=>"010011010",
  45996=>"010010011",
  45997=>"001111011",
  45998=>"101101010",
  45999=>"111011000",
  46000=>"001010001",
  46001=>"011111100",
  46002=>"101001000",
  46003=>"100011101",
  46004=>"110100010",
  46005=>"001101000",
  46006=>"110011111",
  46007=>"000000010",
  46008=>"111100011",
  46009=>"100111111",
  46010=>"100111101",
  46011=>"110100101",
  46012=>"111001010",
  46013=>"011001010",
  46014=>"001100111",
  46015=>"010100010",
  46016=>"110111000",
  46017=>"000111000",
  46018=>"100001110",
  46019=>"111010010",
  46020=>"000101010",
  46021=>"000100111",
  46022=>"000100001",
  46023=>"001101010",
  46024=>"101100010",
  46025=>"101000000",
  46026=>"110101001",
  46027=>"011011010",
  46028=>"110101011",
  46029=>"100100110",
  46030=>"101000011",
  46031=>"001011101",
  46032=>"110100111",
  46033=>"100100010",
  46034=>"111011001",
  46035=>"111100001",
  46036=>"100000110",
  46037=>"010000000",
  46038=>"010111000",
  46039=>"111111011",
  46040=>"111110110",
  46041=>"101101100",
  46042=>"101000101",
  46043=>"001100001",
  46044=>"011111100",
  46045=>"000101001",
  46046=>"011001101",
  46047=>"000110110",
  46048=>"101111001",
  46049=>"011001000",
  46050=>"000101001",
  46051=>"010000101",
  46052=>"010000010",
  46053=>"001001110",
  46054=>"011011110",
  46055=>"101011001",
  46056=>"001001100",
  46057=>"101100101",
  46058=>"001010010",
  46059=>"111111011",
  46060=>"011001000",
  46061=>"011101001",
  46062=>"100000011",
  46063=>"001100111",
  46064=>"010000010",
  46065=>"000010011",
  46066=>"101100111",
  46067=>"111101011",
  46068=>"011010111",
  46069=>"101100011",
  46070=>"000011110",
  46071=>"111101111",
  46072=>"000001011",
  46073=>"110001001",
  46074=>"000010000",
  46075=>"111100010",
  46076=>"000011110",
  46077=>"001101001",
  46078=>"001011011",
  46079=>"001111100",
  46080=>"100110110",
  46081=>"110101111",
  46082=>"111011001",
  46083=>"101001001",
  46084=>"000010110",
  46085=>"111100110",
  46086=>"100001001",
  46087=>"110111100",
  46088=>"000011000",
  46089=>"111110100",
  46090=>"000000010",
  46091=>"111011010",
  46092=>"000000000",
  46093=>"011101111",
  46094=>"111110001",
  46095=>"100001000",
  46096=>"011011101",
  46097=>"000010100",
  46098=>"110111110",
  46099=>"100001111",
  46100=>"100111110",
  46101=>"011110010",
  46102=>"101001010",
  46103=>"011101000",
  46104=>"111011100",
  46105=>"100100110",
  46106=>"110000010",
  46107=>"011010011",
  46108=>"110010101",
  46109=>"010011100",
  46110=>"001101110",
  46111=>"110111110",
  46112=>"000011000",
  46113=>"110100110",
  46114=>"011110100",
  46115=>"011110101",
  46116=>"111001010",
  46117=>"001011010",
  46118=>"100100011",
  46119=>"100100101",
  46120=>"011011100",
  46121=>"001110000",
  46122=>"010011001",
  46123=>"111011100",
  46124=>"000110111",
  46125=>"110000011",
  46126=>"001100000",
  46127=>"111001011",
  46128=>"000000100",
  46129=>"110000010",
  46130=>"001101011",
  46131=>"111001110",
  46132=>"101001010",
  46133=>"111010011",
  46134=>"001001101",
  46135=>"001111010",
  46136=>"001101110",
  46137=>"011100100",
  46138=>"101010110",
  46139=>"100010111",
  46140=>"110011010",
  46141=>"000110100",
  46142=>"101001100",
  46143=>"001011101",
  46144=>"100101010",
  46145=>"110111111",
  46146=>"101111001",
  46147=>"011000001",
  46148=>"100111000",
  46149=>"101010011",
  46150=>"111111111",
  46151=>"110011111",
  46152=>"100010000",
  46153=>"001010110",
  46154=>"110111000",
  46155=>"001101111",
  46156=>"110101101",
  46157=>"110010101",
  46158=>"111111100",
  46159=>"100101101",
  46160=>"000000011",
  46161=>"110000100",
  46162=>"101110110",
  46163=>"111101100",
  46164=>"111100001",
  46165=>"101001101",
  46166=>"000010000",
  46167=>"001010100",
  46168=>"000101100",
  46169=>"000000110",
  46170=>"110011101",
  46171=>"010010010",
  46172=>"001101011",
  46173=>"000111011",
  46174=>"111001111",
  46175=>"110111001",
  46176=>"100100110",
  46177=>"010101111",
  46178=>"110000001",
  46179=>"000010000",
  46180=>"110100101",
  46181=>"111110000",
  46182=>"100110000",
  46183=>"011011111",
  46184=>"101100100",
  46185=>"101100011",
  46186=>"010101001",
  46187=>"110101100",
  46188=>"010101001",
  46189=>"111111101",
  46190=>"101001010",
  46191=>"000110100",
  46192=>"011100000",
  46193=>"011001011",
  46194=>"001011110",
  46195=>"100010001",
  46196=>"001100010",
  46197=>"011100011",
  46198=>"000111110",
  46199=>"001011100",
  46200=>"011111111",
  46201=>"100000110",
  46202=>"100011010",
  46203=>"110100110",
  46204=>"000110101",
  46205=>"100001101",
  46206=>"110010111",
  46207=>"011011111",
  46208=>"101011000",
  46209=>"000100011",
  46210=>"100000111",
  46211=>"111110110",
  46212=>"100101010",
  46213=>"001100011",
  46214=>"001010111",
  46215=>"000110101",
  46216=>"111101001",
  46217=>"101001010",
  46218=>"111110001",
  46219=>"010101011",
  46220=>"101111001",
  46221=>"100101101",
  46222=>"100110110",
  46223=>"010111110",
  46224=>"000101100",
  46225=>"010101000",
  46226=>"111011011",
  46227=>"100100000",
  46228=>"100110101",
  46229=>"011001001",
  46230=>"000110111",
  46231=>"011110010",
  46232=>"101001100",
  46233=>"000000111",
  46234=>"111000010",
  46235=>"000111110",
  46236=>"100100110",
  46237=>"011010111",
  46238=>"100110110",
  46239=>"101011011",
  46240=>"010100001",
  46241=>"101100011",
  46242=>"001110010",
  46243=>"101110011",
  46244=>"100110011",
  46245=>"011100110",
  46246=>"111110101",
  46247=>"111000001",
  46248=>"111011110",
  46249=>"101001001",
  46250=>"110111110",
  46251=>"101110110",
  46252=>"011110110",
  46253=>"011011101",
  46254=>"011110001",
  46255=>"110010100",
  46256=>"010001100",
  46257=>"111101010",
  46258=>"000111011",
  46259=>"010110001",
  46260=>"110100000",
  46261=>"110110110",
  46262=>"010001011",
  46263=>"110011001",
  46264=>"001110110",
  46265=>"011111110",
  46266=>"011001101",
  46267=>"011010101",
  46268=>"101000010",
  46269=>"001001010",
  46270=>"111100001",
  46271=>"110010011",
  46272=>"010111101",
  46273=>"100100010",
  46274=>"010100100",
  46275=>"011001011",
  46276=>"001010110",
  46277=>"100011101",
  46278=>"111110100",
  46279=>"110101111",
  46280=>"001000000",
  46281=>"110111010",
  46282=>"101001111",
  46283=>"100011000",
  46284=>"110100001",
  46285=>"000101000",
  46286=>"010011101",
  46287=>"001110110",
  46288=>"110101010",
  46289=>"011001100",
  46290=>"110001011",
  46291=>"100100000",
  46292=>"000000110",
  46293=>"100100001",
  46294=>"110010111",
  46295=>"010111011",
  46296=>"010111101",
  46297=>"000000001",
  46298=>"111110111",
  46299=>"111011000",
  46300=>"000101011",
  46301=>"010010001",
  46302=>"110011011",
  46303=>"000001100",
  46304=>"100001111",
  46305=>"100110100",
  46306=>"110011010",
  46307=>"000101110",
  46308=>"010011010",
  46309=>"000110011",
  46310=>"110110100",
  46311=>"000110010",
  46312=>"111011101",
  46313=>"101111011",
  46314=>"000110001",
  46315=>"011111010",
  46316=>"111111100",
  46317=>"100110000",
  46318=>"001010101",
  46319=>"101100011",
  46320=>"110011110",
  46321=>"010000111",
  46322=>"000100101",
  46323=>"101100101",
  46324=>"011001100",
  46325=>"111110010",
  46326=>"110100110",
  46327=>"100100100",
  46328=>"110100110",
  46329=>"100010000",
  46330=>"101010010",
  46331=>"100110000",
  46332=>"010110100",
  46333=>"000100000",
  46334=>"000111010",
  46335=>"010100010",
  46336=>"110110001",
  46337=>"010100111",
  46338=>"000100010",
  46339=>"011100101",
  46340=>"000111101",
  46341=>"101010011",
  46342=>"010001011",
  46343=>"111010111",
  46344=>"000011001",
  46345=>"000110110",
  46346=>"011000010",
  46347=>"001000001",
  46348=>"011110010",
  46349=>"010100011",
  46350=>"101010011",
  46351=>"000001101",
  46352=>"001001011",
  46353=>"111001010",
  46354=>"110101100",
  46355=>"100101110",
  46356=>"010101100",
  46357=>"011000001",
  46358=>"011010000",
  46359=>"010000010",
  46360=>"000001010",
  46361=>"100000100",
  46362=>"101001101",
  46363=>"100011100",
  46364=>"111000011",
  46365=>"111101111",
  46366=>"101001111",
  46367=>"000111010",
  46368=>"101000000",
  46369=>"100001010",
  46370=>"001110000",
  46371=>"111000101",
  46372=>"011110100",
  46373=>"101111111",
  46374=>"110100110",
  46375=>"000110001",
  46376=>"100110100",
  46377=>"101010111",
  46378=>"100100011",
  46379=>"011000111",
  46380=>"011101110",
  46381=>"101001000",
  46382=>"110111101",
  46383=>"111110100",
  46384=>"110111101",
  46385=>"110110001",
  46386=>"101001111",
  46387=>"001001101",
  46388=>"111111110",
  46389=>"010111111",
  46390=>"111110000",
  46391=>"000110111",
  46392=>"000110101",
  46393=>"011011101",
  46394=>"111111101",
  46395=>"100110111",
  46396=>"010000110",
  46397=>"100110111",
  46398=>"100010100",
  46399=>"111100001",
  46400=>"100101000",
  46401=>"100010111",
  46402=>"001101111",
  46403=>"110000101",
  46404=>"110100011",
  46405=>"011011100",
  46406=>"011001110",
  46407=>"010000110",
  46408=>"101000101",
  46409=>"100010011",
  46410=>"011010010",
  46411=>"000010001",
  46412=>"101000100",
  46413=>"101000010",
  46414=>"010100110",
  46415=>"100000010",
  46416=>"111111000",
  46417=>"100011000",
  46418=>"111110110",
  46419=>"001111001",
  46420=>"011010011",
  46421=>"001000011",
  46422=>"111100011",
  46423=>"110100101",
  46424=>"111100000",
  46425=>"100110101",
  46426=>"010010000",
  46427=>"001000010",
  46428=>"001101000",
  46429=>"010110011",
  46430=>"000010001",
  46431=>"100110001",
  46432=>"100010110",
  46433=>"100101001",
  46434=>"011010000",
  46435=>"100000000",
  46436=>"101001110",
  46437=>"101110101",
  46438=>"000011101",
  46439=>"110010010",
  46440=>"000000000",
  46441=>"000000011",
  46442=>"101101101",
  46443=>"000010111",
  46444=>"111011101",
  46445=>"100011001",
  46446=>"111101100",
  46447=>"110010000",
  46448=>"000000010",
  46449=>"000110101",
  46450=>"010000011",
  46451=>"011110001",
  46452=>"101011011",
  46453=>"000000011",
  46454=>"000000100",
  46455=>"100001100",
  46456=>"010011100",
  46457=>"110110010",
  46458=>"110101001",
  46459=>"000110110",
  46460=>"001011000",
  46461=>"010111011",
  46462=>"010111000",
  46463=>"111110101",
  46464=>"001001011",
  46465=>"000000100",
  46466=>"000111000",
  46467=>"010001101",
  46468=>"001011010",
  46469=>"110010010",
  46470=>"001011111",
  46471=>"111111110",
  46472=>"000000100",
  46473=>"010010101",
  46474=>"000110101",
  46475=>"011101110",
  46476=>"100110010",
  46477=>"010011101",
  46478=>"101010001",
  46479=>"010011110",
  46480=>"011101000",
  46481=>"101110100",
  46482=>"011110100",
  46483=>"000001010",
  46484=>"111111110",
  46485=>"001110101",
  46486=>"100110110",
  46487=>"100110010",
  46488=>"001110101",
  46489=>"110110111",
  46490=>"100010110",
  46491=>"010110010",
  46492=>"101111000",
  46493=>"100001101",
  46494=>"011111100",
  46495=>"011001101",
  46496=>"110101111",
  46497=>"110110111",
  46498=>"101000110",
  46499=>"101010001",
  46500=>"101101101",
  46501=>"100000000",
  46502=>"001010101",
  46503=>"001100110",
  46504=>"101011000",
  46505=>"101100100",
  46506=>"110101100",
  46507=>"101011101",
  46508=>"110101101",
  46509=>"011001100",
  46510=>"110100001",
  46511=>"011000001",
  46512=>"001100100",
  46513=>"110110100",
  46514=>"011110111",
  46515=>"000000101",
  46516=>"100111011",
  46517=>"010111011",
  46518=>"000011110",
  46519=>"010110000",
  46520=>"110001011",
  46521=>"011110110",
  46522=>"000110011",
  46523=>"111011001",
  46524=>"011101110",
  46525=>"111000010",
  46526=>"000110110",
  46527=>"000100010",
  46528=>"000000101",
  46529=>"001001000",
  46530=>"110101101",
  46531=>"111111011",
  46532=>"111100011",
  46533=>"110011100",
  46534=>"000011010",
  46535=>"111110101",
  46536=>"000110101",
  46537=>"111100101",
  46538=>"011111101",
  46539=>"001001010",
  46540=>"111101111",
  46541=>"110101010",
  46542=>"000111011",
  46543=>"001110111",
  46544=>"101010101",
  46545=>"000110000",
  46546=>"000000110",
  46547=>"001001111",
  46548=>"001000110",
  46549=>"000100100",
  46550=>"100000101",
  46551=>"100000110",
  46552=>"011111100",
  46553=>"100000001",
  46554=>"110100010",
  46555=>"011010101",
  46556=>"110010010",
  46557=>"100100111",
  46558=>"111100100",
  46559=>"001001001",
  46560=>"001100010",
  46561=>"110000100",
  46562=>"110100111",
  46563=>"101110111",
  46564=>"110100100",
  46565=>"111000001",
  46566=>"011110111",
  46567=>"101100000",
  46568=>"001111100",
  46569=>"100110001",
  46570=>"010111111",
  46571=>"001111011",
  46572=>"101010000",
  46573=>"111101111",
  46574=>"101000010",
  46575=>"001101101",
  46576=>"010101001",
  46577=>"010100111",
  46578=>"110010110",
  46579=>"100100110",
  46580=>"110111100",
  46581=>"011111110",
  46582=>"101100000",
  46583=>"010111100",
  46584=>"100001000",
  46585=>"011011011",
  46586=>"111101111",
  46587=>"110100011",
  46588=>"010101000",
  46589=>"010100111",
  46590=>"111110001",
  46591=>"110000010",
  46592=>"001101101",
  46593=>"001111100",
  46594=>"011101111",
  46595=>"100110110",
  46596=>"001011101",
  46597=>"001000100",
  46598=>"111101000",
  46599=>"011100100",
  46600=>"100000001",
  46601=>"000011000",
  46602=>"110000000",
  46603=>"011111010",
  46604=>"110111111",
  46605=>"100001101",
  46606=>"111011000",
  46607=>"111100000",
  46608=>"100110101",
  46609=>"011000000",
  46610=>"100011000",
  46611=>"110100110",
  46612=>"010100100",
  46613=>"000101100",
  46614=>"111100001",
  46615=>"001100000",
  46616=>"001000110",
  46617=>"101110001",
  46618=>"100100011",
  46619=>"001101111",
  46620=>"100011011",
  46621=>"101100110",
  46622=>"000110010",
  46623=>"101000010",
  46624=>"010110000",
  46625=>"101101110",
  46626=>"010110101",
  46627=>"100100011",
  46628=>"110110001",
  46629=>"101000011",
  46630=>"100010111",
  46631=>"110110101",
  46632=>"100101001",
  46633=>"111101111",
  46634=>"100000101",
  46635=>"111111010",
  46636=>"010000001",
  46637=>"010101001",
  46638=>"010010111",
  46639=>"110100111",
  46640=>"101000011",
  46641=>"011101001",
  46642=>"000010100",
  46643=>"000110010",
  46644=>"000100100",
  46645=>"000011101",
  46646=>"010100111",
  46647=>"100001101",
  46648=>"110001110",
  46649=>"100110110",
  46650=>"010011010",
  46651=>"011010011",
  46652=>"000001000",
  46653=>"010001101",
  46654=>"010000100",
  46655=>"101101110",
  46656=>"100110110",
  46657=>"100010111",
  46658=>"110010101",
  46659=>"100000010",
  46660=>"011100001",
  46661=>"010000011",
  46662=>"000101001",
  46663=>"110100100",
  46664=>"001111010",
  46665=>"100100100",
  46666=>"101110011",
  46667=>"110100000",
  46668=>"111111100",
  46669=>"100110100",
  46670=>"000110111",
  46671=>"111100001",
  46672=>"011101000",
  46673=>"011010010",
  46674=>"100110101",
  46675=>"111100011",
  46676=>"001101111",
  46677=>"010110110",
  46678=>"010110100",
  46679=>"001111110",
  46680=>"000111110",
  46681=>"010011110",
  46682=>"111111111",
  46683=>"100100101",
  46684=>"000100100",
  46685=>"011100001",
  46686=>"011101111",
  46687=>"000110100",
  46688=>"000000000",
  46689=>"000000010",
  46690=>"111110100",
  46691=>"101010101",
  46692=>"101011000",
  46693=>"000101000",
  46694=>"110010001",
  46695=>"011100001",
  46696=>"000011001",
  46697=>"011111001",
  46698=>"101001001",
  46699=>"000010110",
  46700=>"110010001",
  46701=>"011010001",
  46702=>"000001100",
  46703=>"010011011",
  46704=>"101111000",
  46705=>"101011100",
  46706=>"011101001",
  46707=>"111100010",
  46708=>"000110010",
  46709=>"011110010",
  46710=>"011010000",
  46711=>"000110100",
  46712=>"110111000",
  46713=>"110011000",
  46714=>"001110101",
  46715=>"001000101",
  46716=>"110011001",
  46717=>"100000001",
  46718=>"101111100",
  46719=>"101101111",
  46720=>"110111110",
  46721=>"100011010",
  46722=>"110110100",
  46723=>"011000000",
  46724=>"000101011",
  46725=>"001110111",
  46726=>"000010011",
  46727=>"111111011",
  46728=>"110111001",
  46729=>"110100110",
  46730=>"110001001",
  46731=>"100001111",
  46732=>"111011011",
  46733=>"111011001",
  46734=>"111100100",
  46735=>"100111101",
  46736=>"010110001",
  46737=>"100110100",
  46738=>"100110011",
  46739=>"110011100",
  46740=>"100000010",
  46741=>"000011011",
  46742=>"111000010",
  46743=>"100101111",
  46744=>"001011000",
  46745=>"100111011",
  46746=>"001010111",
  46747=>"101001101",
  46748=>"111100100",
  46749=>"101111111",
  46750=>"011100111",
  46751=>"110000100",
  46752=>"001100110",
  46753=>"100010011",
  46754=>"110000100",
  46755=>"001000100",
  46756=>"101100100",
  46757=>"011101111",
  46758=>"100110111",
  46759=>"011011000",
  46760=>"001001011",
  46761=>"010000011",
  46762=>"111100111",
  46763=>"010010100",
  46764=>"010001000",
  46765=>"010000110",
  46766=>"101101000",
  46767=>"000101001",
  46768=>"011101101",
  46769=>"110011110",
  46770=>"110000001",
  46771=>"000101110",
  46772=>"000000100",
  46773=>"111101010",
  46774=>"100001101",
  46775=>"111101111",
  46776=>"001001000",
  46777=>"000001001",
  46778=>"111111100",
  46779=>"101000001",
  46780=>"011100000",
  46781=>"010010000",
  46782=>"100110111",
  46783=>"100110110",
  46784=>"100000100",
  46785=>"011111010",
  46786=>"100001110",
  46787=>"001010011",
  46788=>"010100000",
  46789=>"101110100",
  46790=>"110000010",
  46791=>"100100010",
  46792=>"111110100",
  46793=>"110010110",
  46794=>"111111001",
  46795=>"001011100",
  46796=>"110100011",
  46797=>"011101000",
  46798=>"100011010",
  46799=>"000100100",
  46800=>"010111110",
  46801=>"110001111",
  46802=>"011000111",
  46803=>"100010010",
  46804=>"100101110",
  46805=>"011001011",
  46806=>"011011110",
  46807=>"101110110",
  46808=>"001110001",
  46809=>"000011011",
  46810=>"101100100",
  46811=>"111011101",
  46812=>"000100101",
  46813=>"111101111",
  46814=>"000100000",
  46815=>"110101111",
  46816=>"111100001",
  46817=>"000010000",
  46818=>"000100111",
  46819=>"110011000",
  46820=>"010101101",
  46821=>"011000111",
  46822=>"110001000",
  46823=>"000001100",
  46824=>"100010111",
  46825=>"101000101",
  46826=>"001000001",
  46827=>"010101110",
  46828=>"001000011",
  46829=>"100000110",
  46830=>"011010001",
  46831=>"110111100",
  46832=>"110010010",
  46833=>"110010111",
  46834=>"011011101",
  46835=>"110011000",
  46836=>"010100111",
  46837=>"011000001",
  46838=>"000111100",
  46839=>"000110010",
  46840=>"000111001",
  46841=>"010110100",
  46842=>"100001010",
  46843=>"111000011",
  46844=>"110001100",
  46845=>"101011101",
  46846=>"011001011",
  46847=>"010110101",
  46848=>"110010110",
  46849=>"000000001",
  46850=>"010010100",
  46851=>"001000101",
  46852=>"011100101",
  46853=>"010001101",
  46854=>"001010101",
  46855=>"010000010",
  46856=>"001111011",
  46857=>"100110000",
  46858=>"011100000",
  46859=>"001100100",
  46860=>"001000111",
  46861=>"011001001",
  46862=>"000110101",
  46863=>"110100101",
  46864=>"101100111",
  46865=>"100110110",
  46866=>"110110100",
  46867=>"111011001",
  46868=>"101110100",
  46869=>"111111100",
  46870=>"000010110",
  46871=>"101011001",
  46872=>"000011000",
  46873=>"000001100",
  46874=>"100010001",
  46875=>"001111101",
  46876=>"110110010",
  46877=>"011001100",
  46878=>"110110010",
  46879=>"010111011",
  46880=>"010111000",
  46881=>"111010100",
  46882=>"111101001",
  46883=>"000110000",
  46884=>"000000111",
  46885=>"110011000",
  46886=>"111011000",
  46887=>"000111110",
  46888=>"001000001",
  46889=>"101100110",
  46890=>"100110000",
  46891=>"100101101",
  46892=>"010111111",
  46893=>"000001110",
  46894=>"100111110",
  46895=>"110010010",
  46896=>"001000010",
  46897=>"100100010",
  46898=>"110101001",
  46899=>"001101110",
  46900=>"111100111",
  46901=>"111100010",
  46902=>"100011111",
  46903=>"001100111",
  46904=>"011111011",
  46905=>"111101000",
  46906=>"001001101",
  46907=>"111011110",
  46908=>"011000001",
  46909=>"111010100",
  46910=>"110101101",
  46911=>"000010001",
  46912=>"001101101",
  46913=>"111110111",
  46914=>"101111000",
  46915=>"101010111",
  46916=>"100110110",
  46917=>"111010001",
  46918=>"111110110",
  46919=>"110001100",
  46920=>"010000000",
  46921=>"011100110",
  46922=>"001001111",
  46923=>"100111110",
  46924=>"111010010",
  46925=>"010011000",
  46926=>"001110101",
  46927=>"110101111",
  46928=>"101111111",
  46929=>"111111010",
  46930=>"100100000",
  46931=>"010001101",
  46932=>"000000001",
  46933=>"101010111",
  46934=>"011000001",
  46935=>"010010001",
  46936=>"111100000",
  46937=>"001011011",
  46938=>"101101111",
  46939=>"101110001",
  46940=>"001010010",
  46941=>"001110101",
  46942=>"100010000",
  46943=>"100010100",
  46944=>"010010011",
  46945=>"110000101",
  46946=>"110100000",
  46947=>"000101110",
  46948=>"110101100",
  46949=>"110110000",
  46950=>"111111111",
  46951=>"000001010",
  46952=>"111110111",
  46953=>"110000010",
  46954=>"010101101",
  46955=>"110110011",
  46956=>"110110010",
  46957=>"001000011",
  46958=>"101000110",
  46959=>"001001100",
  46960=>"100010011",
  46961=>"000011101",
  46962=>"000011010",
  46963=>"100100000",
  46964=>"110100001",
  46965=>"001111110",
  46966=>"010111110",
  46967=>"111110100",
  46968=>"110110011",
  46969=>"100101010",
  46970=>"111000101",
  46971=>"101000100",
  46972=>"100100000",
  46973=>"100001001",
  46974=>"111010100",
  46975=>"110011000",
  46976=>"000011001",
  46977=>"000000011",
  46978=>"100001000",
  46979=>"100010100",
  46980=>"110001110",
  46981=>"011001011",
  46982=>"010110110",
  46983=>"110100000",
  46984=>"010010101",
  46985=>"110010101",
  46986=>"011110110",
  46987=>"101101100",
  46988=>"000001011",
  46989=>"010011011",
  46990=>"000000011",
  46991=>"101110001",
  46992=>"110110111",
  46993=>"111010111",
  46994=>"111010000",
  46995=>"110111000",
  46996=>"011010100",
  46997=>"011010101",
  46998=>"010001100",
  46999=>"000010010",
  47000=>"000110110",
  47001=>"100100110",
  47002=>"010001000",
  47003=>"011010111",
  47004=>"000101010",
  47005=>"011101000",
  47006=>"101010000",
  47007=>"101000110",
  47008=>"101000000",
  47009=>"101010111",
  47010=>"110000111",
  47011=>"111001110",
  47012=>"010110010",
  47013=>"110110111",
  47014=>"000110111",
  47015=>"000010110",
  47016=>"000011110",
  47017=>"010110011",
  47018=>"001000110",
  47019=>"011011100",
  47020=>"110000111",
  47021=>"110000001",
  47022=>"001100111",
  47023=>"110010110",
  47024=>"001011000",
  47025=>"101111001",
  47026=>"011110111",
  47027=>"100010000",
  47028=>"111111011",
  47029=>"011101001",
  47030=>"100000100",
  47031=>"001000101",
  47032=>"101000001",
  47033=>"010110110",
  47034=>"010111111",
  47035=>"011010100",
  47036=>"010010011",
  47037=>"111110000",
  47038=>"101011010",
  47039=>"100101110",
  47040=>"110101011",
  47041=>"111100110",
  47042=>"000100011",
  47043=>"100011101",
  47044=>"101000101",
  47045=>"111000100",
  47046=>"000110000",
  47047=>"100111010",
  47048=>"111110001",
  47049=>"010111011",
  47050=>"011100101",
  47051=>"101100011",
  47052=>"011110000",
  47053=>"101110101",
  47054=>"100111110",
  47055=>"101011110",
  47056=>"011011101",
  47057=>"111110000",
  47058=>"111000001",
  47059=>"000001001",
  47060=>"000110101",
  47061=>"111100101",
  47062=>"110110100",
  47063=>"001001101",
  47064=>"111100100",
  47065=>"010111010",
  47066=>"001100001",
  47067=>"011011101",
  47068=>"010111111",
  47069=>"100011101",
  47070=>"111111010",
  47071=>"111110011",
  47072=>"000011111",
  47073=>"110010000",
  47074=>"101001111",
  47075=>"100110110",
  47076=>"110111100",
  47077=>"101110110",
  47078=>"001101110",
  47079=>"110010101",
  47080=>"011001110",
  47081=>"000001010",
  47082=>"111000110",
  47083=>"001110010",
  47084=>"111011000",
  47085=>"001000011",
  47086=>"101001111",
  47087=>"011110010",
  47088=>"000011000",
  47089=>"100000100",
  47090=>"100000101",
  47091=>"011110101",
  47092=>"100011000",
  47093=>"000110000",
  47094=>"110000000",
  47095=>"000001000",
  47096=>"011000011",
  47097=>"100101011",
  47098=>"111101000",
  47099=>"111001001",
  47100=>"110010001",
  47101=>"000000100",
  47102=>"000100010",
  47103=>"110100000",
  47104=>"000001100",
  47105=>"110101010",
  47106=>"101001110",
  47107=>"010001010",
  47108=>"011011111",
  47109=>"011111010",
  47110=>"011011110",
  47111=>"001000101",
  47112=>"010010100",
  47113=>"111011100",
  47114=>"101111001",
  47115=>"000011111",
  47116=>"111000100",
  47117=>"000011011",
  47118=>"101100101",
  47119=>"010011010",
  47120=>"111101101",
  47121=>"010011010",
  47122=>"010100001",
  47123=>"001111001",
  47124=>"000010100",
  47125=>"001000101",
  47126=>"110101111",
  47127=>"010000000",
  47128=>"110011000",
  47129=>"000010110",
  47130=>"001001111",
  47131=>"001000100",
  47132=>"001010101",
  47133=>"011011010",
  47134=>"001100100",
  47135=>"001110100",
  47136=>"000000101",
  47137=>"010111111",
  47138=>"100111110",
  47139=>"111101000",
  47140=>"111000111",
  47141=>"001111010",
  47142=>"100000100",
  47143=>"100110000",
  47144=>"010001010",
  47145=>"010011110",
  47146=>"100101011",
  47147=>"101011011",
  47148=>"001011100",
  47149=>"110101001",
  47150=>"011101110",
  47151=>"101000100",
  47152=>"100110111",
  47153=>"010010001",
  47154=>"101011011",
  47155=>"011110011",
  47156=>"001010101",
  47157=>"101011100",
  47158=>"001100111",
  47159=>"110111111",
  47160=>"001001011",
  47161=>"110100100",
  47162=>"110110011",
  47163=>"000111100",
  47164=>"100101110",
  47165=>"110001001",
  47166=>"111011110",
  47167=>"000101111",
  47168=>"011110111",
  47169=>"001000010",
  47170=>"111100010",
  47171=>"000101110",
  47172=>"110101110",
  47173=>"011010100",
  47174=>"110001000",
  47175=>"111010010",
  47176=>"001001111",
  47177=>"010110110",
  47178=>"100110111",
  47179=>"000001010",
  47180=>"010111100",
  47181=>"100010110",
  47182=>"100100011",
  47183=>"011000010",
  47184=>"011111111",
  47185=>"010010001",
  47186=>"111111001",
  47187=>"101110100",
  47188=>"011000000",
  47189=>"110111001",
  47190=>"101100001",
  47191=>"011001100",
  47192=>"011010001",
  47193=>"000101111",
  47194=>"111100111",
  47195=>"001001001",
  47196=>"010010010",
  47197=>"010011000",
  47198=>"110000111",
  47199=>"011000010",
  47200=>"100001000",
  47201=>"011100101",
  47202=>"001010001",
  47203=>"100000011",
  47204=>"100111101",
  47205=>"000001111",
  47206=>"000010000",
  47207=>"110001100",
  47208=>"010000001",
  47209=>"110001110",
  47210=>"101010101",
  47211=>"001011111",
  47212=>"001001000",
  47213=>"101011100",
  47214=>"011111100",
  47215=>"000010011",
  47216=>"100000000",
  47217=>"100011011",
  47218=>"100010111",
  47219=>"111111100",
  47220=>"010011011",
  47221=>"110111101",
  47222=>"101101000",
  47223=>"011010110",
  47224=>"100100111",
  47225=>"001000101",
  47226=>"001010010",
  47227=>"110101111",
  47228=>"110001010",
  47229=>"100011000",
  47230=>"000001110",
  47231=>"110100111",
  47232=>"101110100",
  47233=>"000011011",
  47234=>"000101111",
  47235=>"011001001",
  47236=>"101101111",
  47237=>"101000100",
  47238=>"100001011",
  47239=>"101011100",
  47240=>"101110000",
  47241=>"001111001",
  47242=>"001001000",
  47243=>"001001001",
  47244=>"011100001",
  47245=>"001000111",
  47246=>"000101000",
  47247=>"110101011",
  47248=>"001000010",
  47249=>"001111000",
  47250=>"001000001",
  47251=>"110100101",
  47252=>"000111100",
  47253=>"101100011",
  47254=>"011010110",
  47255=>"001010011",
  47256=>"010101010",
  47257=>"011011100",
  47258=>"001000001",
  47259=>"011010001",
  47260=>"000110010",
  47261=>"110010001",
  47262=>"010011001",
  47263=>"100011100",
  47264=>"110110000",
  47265=>"101110100",
  47266=>"100010000",
  47267=>"101000010",
  47268=>"100111000",
  47269=>"001111111",
  47270=>"111100000",
  47271=>"100000000",
  47272=>"001110111",
  47273=>"110100111",
  47274=>"010000100",
  47275=>"100111000",
  47276=>"011000000",
  47277=>"110101000",
  47278=>"111111100",
  47279=>"110110110",
  47280=>"000100010",
  47281=>"110100100",
  47282=>"001011001",
  47283=>"101000000",
  47284=>"100000101",
  47285=>"110110011",
  47286=>"001001001",
  47287=>"011110010",
  47288=>"010000011",
  47289=>"111010010",
  47290=>"110000010",
  47291=>"010001101",
  47292=>"111100011",
  47293=>"110100010",
  47294=>"010011100",
  47295=>"111010001",
  47296=>"010101010",
  47297=>"010110100",
  47298=>"100000010",
  47299=>"100000000",
  47300=>"001011101",
  47301=>"001000101",
  47302=>"010010101",
  47303=>"101110101",
  47304=>"101101110",
  47305=>"100010011",
  47306=>"111100001",
  47307=>"011001100",
  47308=>"101111110",
  47309=>"100001000",
  47310=>"000010110",
  47311=>"110010100",
  47312=>"111000010",
  47313=>"011000111",
  47314=>"001100001",
  47315=>"110001110",
  47316=>"010000000",
  47317=>"001010100",
  47318=>"011011010",
  47319=>"011011011",
  47320=>"010100001",
  47321=>"101000101",
  47322=>"011110100",
  47323=>"001111011",
  47324=>"000011110",
  47325=>"011000100",
  47326=>"010011011",
  47327=>"110101010",
  47328=>"010010001",
  47329=>"101001111",
  47330=>"111111111",
  47331=>"010110000",
  47332=>"110010011",
  47333=>"110101011",
  47334=>"100011001",
  47335=>"010000001",
  47336=>"101001101",
  47337=>"100100100",
  47338=>"100010110",
  47339=>"100101000",
  47340=>"110000100",
  47341=>"000010100",
  47342=>"100000000",
  47343=>"011010001",
  47344=>"111001011",
  47345=>"100000001",
  47346=>"010101000",
  47347=>"011111001",
  47348=>"011101100",
  47349=>"011001011",
  47350=>"010110000",
  47351=>"100100011",
  47352=>"010111011",
  47353=>"101100000",
  47354=>"000000000",
  47355=>"010010001",
  47356=>"001100101",
  47357=>"100011100",
  47358=>"110011111",
  47359=>"101100101",
  47360=>"111011111",
  47361=>"001100010",
  47362=>"000100111",
  47363=>"100011000",
  47364=>"110001000",
  47365=>"100100001",
  47366=>"010011100",
  47367=>"101000111",
  47368=>"001100100",
  47369=>"001110001",
  47370=>"011111011",
  47371=>"000000100",
  47372=>"100001100",
  47373=>"000110111",
  47374=>"110100001",
  47375=>"001111000",
  47376=>"110110110",
  47377=>"111111111",
  47378=>"011100111",
  47379=>"100001111",
  47380=>"101001100",
  47381=>"110110110",
  47382=>"010000101",
  47383=>"101101001",
  47384=>"110001101",
  47385=>"111000101",
  47386=>"011011101",
  47387=>"011010011",
  47388=>"000001100",
  47389=>"010000101",
  47390=>"100001110",
  47391=>"000010010",
  47392=>"000000000",
  47393=>"101001000",
  47394=>"000100101",
  47395=>"000000100",
  47396=>"011110100",
  47397=>"000101001",
  47398=>"011010100",
  47399=>"111001111",
  47400=>"001011100",
  47401=>"011100100",
  47402=>"000110100",
  47403=>"110001000",
  47404=>"000101101",
  47405=>"000010100",
  47406=>"100010110",
  47407=>"011111100",
  47408=>"000001110",
  47409=>"001001110",
  47410=>"101001101",
  47411=>"011001110",
  47412=>"110111001",
  47413=>"111011110",
  47414=>"110110101",
  47415=>"101000000",
  47416=>"100100001",
  47417=>"001010110",
  47418=>"100100001",
  47419=>"000101011",
  47420=>"100111111",
  47421=>"110100001",
  47422=>"101011010",
  47423=>"001000011",
  47424=>"101000010",
  47425=>"110000100",
  47426=>"101100100",
  47427=>"000000110",
  47428=>"001110100",
  47429=>"101000100",
  47430=>"010001000",
  47431=>"001101011",
  47432=>"000100101",
  47433=>"101001011",
  47434=>"011010111",
  47435=>"111101100",
  47436=>"011111010",
  47437=>"000101101",
  47438=>"100001111",
  47439=>"101101011",
  47440=>"001101000",
  47441=>"011111111",
  47442=>"111101100",
  47443=>"010001111",
  47444=>"000101001",
  47445=>"100110010",
  47446=>"001010001",
  47447=>"111101100",
  47448=>"100010110",
  47449=>"000100000",
  47450=>"111011100",
  47451=>"100100011",
  47452=>"111111101",
  47453=>"010100011",
  47454=>"011001011",
  47455=>"011000101",
  47456=>"100111111",
  47457=>"001001100",
  47458=>"001001000",
  47459=>"010001001",
  47460=>"000000000",
  47461=>"000011000",
  47462=>"110110111",
  47463=>"010110101",
  47464=>"100101001",
  47465=>"100001101",
  47466=>"001010001",
  47467=>"000000111",
  47468=>"011111011",
  47469=>"111010100",
  47470=>"000011000",
  47471=>"010101000",
  47472=>"100110000",
  47473=>"100001101",
  47474=>"111110001",
  47475=>"011100000",
  47476=>"010010011",
  47477=>"010101011",
  47478=>"000101110",
  47479=>"101000010",
  47480=>"100101011",
  47481=>"101101100",
  47482=>"100100001",
  47483=>"110110100",
  47484=>"110011000",
  47485=>"001011110",
  47486=>"100000010",
  47487=>"110001100",
  47488=>"000101010",
  47489=>"000000100",
  47490=>"110000001",
  47491=>"000111000",
  47492=>"110001111",
  47493=>"100000111",
  47494=>"100010000",
  47495=>"011100100",
  47496=>"001010000",
  47497=>"010110011",
  47498=>"110111011",
  47499=>"001101111",
  47500=>"110000001",
  47501=>"000011110",
  47502=>"010000010",
  47503=>"000100001",
  47504=>"011001111",
  47505=>"000100111",
  47506=>"111110010",
  47507=>"001100010",
  47508=>"001110010",
  47509=>"111101110",
  47510=>"100100111",
  47511=>"101001111",
  47512=>"000000010",
  47513=>"001011110",
  47514=>"100100000",
  47515=>"000110011",
  47516=>"011011010",
  47517=>"000001011",
  47518=>"110101110",
  47519=>"010010001",
  47520=>"000101011",
  47521=>"101110011",
  47522=>"110000001",
  47523=>"010000000",
  47524=>"000100000",
  47525=>"101001001",
  47526=>"111001001",
  47527=>"111010000",
  47528=>"010111010",
  47529=>"111010100",
  47530=>"010010001",
  47531=>"010000011",
  47532=>"110011111",
  47533=>"011001100",
  47534=>"100110100",
  47535=>"000100001",
  47536=>"001000001",
  47537=>"100101010",
  47538=>"111001011",
  47539=>"000010110",
  47540=>"110010001",
  47541=>"101001101",
  47542=>"101110101",
  47543=>"000110111",
  47544=>"011110101",
  47545=>"001110100",
  47546=>"100001100",
  47547=>"100110000",
  47548=>"100000101",
  47549=>"000011100",
  47550=>"011010001",
  47551=>"010010111",
  47552=>"110110000",
  47553=>"000001111",
  47554=>"010101010",
  47555=>"000001101",
  47556=>"101101100",
  47557=>"100000010",
  47558=>"011100100",
  47559=>"001110110",
  47560=>"010100101",
  47561=>"100010001",
  47562=>"010100110",
  47563=>"111101011",
  47564=>"010101000",
  47565=>"000010010",
  47566=>"000001110",
  47567=>"011100001",
  47568=>"110001101",
  47569=>"000010100",
  47570=>"100100101",
  47571=>"001001001",
  47572=>"000111101",
  47573=>"010010111",
  47574=>"001101101",
  47575=>"010011010",
  47576=>"100000101",
  47577=>"100101001",
  47578=>"010010100",
  47579=>"001010000",
  47580=>"101011001",
  47581=>"111111011",
  47582=>"101101011",
  47583=>"000110011",
  47584=>"100101011",
  47585=>"000111001",
  47586=>"110100101",
  47587=>"101101101",
  47588=>"111011000",
  47589=>"011100011",
  47590=>"110100011",
  47591=>"011100110",
  47592=>"011110111",
  47593=>"010100101",
  47594=>"000000001",
  47595=>"111000011",
  47596=>"000000000",
  47597=>"001011101",
  47598=>"011101111",
  47599=>"011100000",
  47600=>"011100000",
  47601=>"101101100",
  47602=>"110011010",
  47603=>"111100001",
  47604=>"001010100",
  47605=>"100001011",
  47606=>"010000111",
  47607=>"001100111",
  47608=>"100000001",
  47609=>"001011011",
  47610=>"111110011",
  47611=>"110111111",
  47612=>"000001000",
  47613=>"101110110",
  47614=>"110101100",
  47615=>"110000011",
  47616=>"110010100",
  47617=>"011101100",
  47618=>"100010001",
  47619=>"100000001",
  47620=>"100111100",
  47621=>"010101100",
  47622=>"111100101",
  47623=>"011000000",
  47624=>"111000111",
  47625=>"000101010",
  47626=>"010110111",
  47627=>"011011101",
  47628=>"010111110",
  47629=>"110101011",
  47630=>"010010110",
  47631=>"110111011",
  47632=>"010100110",
  47633=>"000001000",
  47634=>"100100111",
  47635=>"011100000",
  47636=>"000010010",
  47637=>"000111101",
  47638=>"111101011",
  47639=>"110101000",
  47640=>"011101110",
  47641=>"011010100",
  47642=>"100010010",
  47643=>"111001111",
  47644=>"100000101",
  47645=>"000010100",
  47646=>"111001101",
  47647=>"011000100",
  47648=>"101110110",
  47649=>"001000001",
  47650=>"000111100",
  47651=>"001000010",
  47652=>"111010111",
  47653=>"001100100",
  47654=>"011111001",
  47655=>"110100111",
  47656=>"011101100",
  47657=>"000010111",
  47658=>"100010101",
  47659=>"101101001",
  47660=>"011010001",
  47661=>"011001010",
  47662=>"101000011",
  47663=>"101000100",
  47664=>"100110001",
  47665=>"010101000",
  47666=>"001000100",
  47667=>"000000001",
  47668=>"111011001",
  47669=>"011010001",
  47670=>"011100110",
  47671=>"000110101",
  47672=>"010011011",
  47673=>"111011101",
  47674=>"001111001",
  47675=>"001010010",
  47676=>"011101001",
  47677=>"001000101",
  47678=>"000110110",
  47679=>"010011001",
  47680=>"101000001",
  47681=>"010001010",
  47682=>"110111101",
  47683=>"100100100",
  47684=>"111001001",
  47685=>"111000110",
  47686=>"000101000",
  47687=>"011001001",
  47688=>"000101000",
  47689=>"111100000",
  47690=>"000110011",
  47691=>"110100010",
  47692=>"001010011",
  47693=>"000100010",
  47694=>"000000010",
  47695=>"000101111",
  47696=>"010000000",
  47697=>"100110010",
  47698=>"000111010",
  47699=>"111011110",
  47700=>"010111100",
  47701=>"100010101",
  47702=>"011100011",
  47703=>"010100100",
  47704=>"100110001",
  47705=>"100001100",
  47706=>"101110001",
  47707=>"001010111",
  47708=>"010100001",
  47709=>"101110000",
  47710=>"000101011",
  47711=>"111111111",
  47712=>"011101001",
  47713=>"110111100",
  47714=>"011100010",
  47715=>"101000001",
  47716=>"010011011",
  47717=>"101001001",
  47718=>"110001110",
  47719=>"111011011",
  47720=>"000110000",
  47721=>"011000001",
  47722=>"100110111",
  47723=>"001100011",
  47724=>"000111110",
  47725=>"101110110",
  47726=>"101110111",
  47727=>"110101000",
  47728=>"110010000",
  47729=>"001000010",
  47730=>"111101001",
  47731=>"001111100",
  47732=>"001000010",
  47733=>"101110000",
  47734=>"011110100",
  47735=>"000100111",
  47736=>"111101100",
  47737=>"111001001",
  47738=>"110000111",
  47739=>"111100011",
  47740=>"000100110",
  47741=>"001010001",
  47742=>"110110010",
  47743=>"101110101",
  47744=>"010100100",
  47745=>"111101111",
  47746=>"000110111",
  47747=>"001111001",
  47748=>"001110011",
  47749=>"100000000",
  47750=>"010001101",
  47751=>"101011001",
  47752=>"010010111",
  47753=>"011001100",
  47754=>"000111001",
  47755=>"111110011",
  47756=>"000110101",
  47757=>"001000100",
  47758=>"110001101",
  47759=>"001110001",
  47760=>"010000011",
  47761=>"000100110",
  47762=>"101110001",
  47763=>"011001011",
  47764=>"000001010",
  47765=>"011101111",
  47766=>"111011010",
  47767=>"101110001",
  47768=>"000011100",
  47769=>"101011111",
  47770=>"010011000",
  47771=>"100001000",
  47772=>"001011010",
  47773=>"011101100",
  47774=>"000101001",
  47775=>"110111100",
  47776=>"100011101",
  47777=>"000111010",
  47778=>"100100000",
  47779=>"110111001",
  47780=>"111100101",
  47781=>"100001101",
  47782=>"100101001",
  47783=>"000100010",
  47784=>"110111100",
  47785=>"110101100",
  47786=>"000010011",
  47787=>"110101010",
  47788=>"011011100",
  47789=>"111110010",
  47790=>"111010101",
  47791=>"111001001",
  47792=>"001001000",
  47793=>"000100111",
  47794=>"001000101",
  47795=>"110011001",
  47796=>"101010110",
  47797=>"100100011",
  47798=>"110001010",
  47799=>"110101010",
  47800=>"101000000",
  47801=>"001000111",
  47802=>"011001011",
  47803=>"100001001",
  47804=>"001110101",
  47805=>"110011010",
  47806=>"000000011",
  47807=>"111110110",
  47808=>"000101100",
  47809=>"000000011",
  47810=>"111010011",
  47811=>"000000100",
  47812=>"111100101",
  47813=>"010010110",
  47814=>"101110000",
  47815=>"000010000",
  47816=>"001100001",
  47817=>"111000101",
  47818=>"001111001",
  47819=>"101100101",
  47820=>"000000100",
  47821=>"000110100",
  47822=>"010000000",
  47823=>"010011010",
  47824=>"110110101",
  47825=>"101000000",
  47826=>"011110010",
  47827=>"000011101",
  47828=>"000100101",
  47829=>"000111011",
  47830=>"111101011",
  47831=>"000110010",
  47832=>"000001111",
  47833=>"111001101",
  47834=>"111011100",
  47835=>"111011101",
  47836=>"000000011",
  47837=>"111101011",
  47838=>"100000110",
  47839=>"101101010",
  47840=>"001001000",
  47841=>"001000001",
  47842=>"100011101",
  47843=>"111110101",
  47844=>"001011011",
  47845=>"101100111",
  47846=>"000011011",
  47847=>"101011101",
  47848=>"000001001",
  47849=>"110010100",
  47850=>"011100001",
  47851=>"111000100",
  47852=>"011110110",
  47853=>"000011101",
  47854=>"011101101",
  47855=>"010101010",
  47856=>"111111000",
  47857=>"101101110",
  47858=>"011001001",
  47859=>"011100000",
  47860=>"000000011",
  47861=>"001010110",
  47862=>"001100001",
  47863=>"101100100",
  47864=>"000011100",
  47865=>"110001100",
  47866=>"110000011",
  47867=>"011000000",
  47868=>"100010101",
  47869=>"111110110",
  47870=>"010011100",
  47871=>"010111110",
  47872=>"010100010",
  47873=>"111111110",
  47874=>"111100001",
  47875=>"101100001",
  47876=>"011110000",
  47877=>"100001110",
  47878=>"101111110",
  47879=>"011101001",
  47880=>"000000000",
  47881=>"000111001",
  47882=>"100100110",
  47883=>"000001010",
  47884=>"100000110",
  47885=>"110010011",
  47886=>"001111010",
  47887=>"000010101",
  47888=>"101011100",
  47889=>"100111010",
  47890=>"101001001",
  47891=>"010010110",
  47892=>"100001001",
  47893=>"100100101",
  47894=>"011011001",
  47895=>"101110001",
  47896=>"100001110",
  47897=>"000100100",
  47898=>"100000010",
  47899=>"010101011",
  47900=>"011010010",
  47901=>"001000110",
  47902=>"101011000",
  47903=>"100001010",
  47904=>"111000100",
  47905=>"110011101",
  47906=>"110100111",
  47907=>"100110110",
  47908=>"010101010",
  47909=>"100000000",
  47910=>"110000100",
  47911=>"111000101",
  47912=>"000001111",
  47913=>"101111100",
  47914=>"010010101",
  47915=>"011000110",
  47916=>"001001011",
  47917=>"111011000",
  47918=>"101000010",
  47919=>"000111000",
  47920=>"000100100",
  47921=>"110010101",
  47922=>"011001011",
  47923=>"001001100",
  47924=>"100110110",
  47925=>"011101001",
  47926=>"001111100",
  47927=>"110101010",
  47928=>"111110010",
  47929=>"000101000",
  47930=>"111010101",
  47931=>"011110100",
  47932=>"101011010",
  47933=>"000100000",
  47934=>"011111000",
  47935=>"001100101",
  47936=>"010111101",
  47937=>"111110110",
  47938=>"001110001",
  47939=>"111000010",
  47940=>"111011001",
  47941=>"010101011",
  47942=>"000110110",
  47943=>"000100010",
  47944=>"010100110",
  47945=>"011000001",
  47946=>"011100110",
  47947=>"001001111",
  47948=>"110110111",
  47949=>"001101101",
  47950=>"111111100",
  47951=>"010011111",
  47952=>"111010011",
  47953=>"101100000",
  47954=>"100001011",
  47955=>"000011000",
  47956=>"001101010",
  47957=>"001101101",
  47958=>"110000000",
  47959=>"001000010",
  47960=>"000010000",
  47961=>"011110110",
  47962=>"000001010",
  47963=>"000000111",
  47964=>"110101010",
  47965=>"110111101",
  47966=>"110111011",
  47967=>"000001001",
  47968=>"001110110",
  47969=>"001000111",
  47970=>"011100111",
  47971=>"010001011",
  47972=>"110100101",
  47973=>"111111101",
  47974=>"100011101",
  47975=>"101011011",
  47976=>"101010100",
  47977=>"001001101",
  47978=>"001110000",
  47979=>"111101011",
  47980=>"100011000",
  47981=>"110010011",
  47982=>"000001011",
  47983=>"001110010",
  47984=>"010111101",
  47985=>"101101111",
  47986=>"101001100",
  47987=>"110011001",
  47988=>"011010000",
  47989=>"010001101",
  47990=>"000100000",
  47991=>"000000011",
  47992=>"000110000",
  47993=>"100111100",
  47994=>"010001111",
  47995=>"100101001",
  47996=>"000001110",
  47997=>"111110001",
  47998=>"010100101",
  47999=>"111101011",
  48000=>"001100110",
  48001=>"101000111",
  48002=>"010001011",
  48003=>"000001101",
  48004=>"011111000",
  48005=>"110100101",
  48006=>"111110100",
  48007=>"100000001",
  48008=>"111101110",
  48009=>"010101101",
  48010=>"011010101",
  48011=>"110011011",
  48012=>"011011100",
  48013=>"100110011",
  48014=>"000011000",
  48015=>"010011100",
  48016=>"101111100",
  48017=>"010100110",
  48018=>"001000000",
  48019=>"011101010",
  48020=>"011110110",
  48021=>"011100011",
  48022=>"000000111",
  48023=>"101000100",
  48024=>"000001000",
  48025=>"111000100",
  48026=>"000011110",
  48027=>"000010001",
  48028=>"100101100",
  48029=>"100001010",
  48030=>"001000101",
  48031=>"011000000",
  48032=>"101010000",
  48033=>"010011000",
  48034=>"000000000",
  48035=>"101111101",
  48036=>"101011111",
  48037=>"101110010",
  48038=>"010101000",
  48039=>"100010001",
  48040=>"101011000",
  48041=>"100101001",
  48042=>"000100000",
  48043=>"011010001",
  48044=>"010101111",
  48045=>"011100000",
  48046=>"111000011",
  48047=>"011001111",
  48048=>"010000101",
  48049=>"100001101",
  48050=>"001111111",
  48051=>"001110011",
  48052=>"111110010",
  48053=>"000010101",
  48054=>"101111000",
  48055=>"111000011",
  48056=>"001010001",
  48057=>"100110001",
  48058=>"101001000",
  48059=>"110111000",
  48060=>"011101000",
  48061=>"000101110",
  48062=>"111110100",
  48063=>"100011110",
  48064=>"110111010",
  48065=>"011011100",
  48066=>"001011101",
  48067=>"100110001",
  48068=>"001011010",
  48069=>"110001101",
  48070=>"101011010",
  48071=>"101100011",
  48072=>"001001101",
  48073=>"011000110",
  48074=>"100010111",
  48075=>"010111101",
  48076=>"010100101",
  48077=>"000110110",
  48078=>"111010110",
  48079=>"000101010",
  48080=>"000110111",
  48081=>"001101011",
  48082=>"100100001",
  48083=>"000011011",
  48084=>"000011010",
  48085=>"010110111",
  48086=>"110001101",
  48087=>"010001011",
  48088=>"110000011",
  48089=>"010000101",
  48090=>"101111011",
  48091=>"111111111",
  48092=>"000010110",
  48093=>"101011010",
  48094=>"110110001",
  48095=>"001101000",
  48096=>"000001010",
  48097=>"110011111",
  48098=>"001000011",
  48099=>"010100010",
  48100=>"111000010",
  48101=>"001110100",
  48102=>"010100010",
  48103=>"101010000",
  48104=>"000000000",
  48105=>"001000000",
  48106=>"001111010",
  48107=>"110011010",
  48108=>"010111011",
  48109=>"001011001",
  48110=>"001001100",
  48111=>"101110000",
  48112=>"010100101",
  48113=>"111000011",
  48114=>"111100100",
  48115=>"011010011",
  48116=>"000010000",
  48117=>"001100111",
  48118=>"010010111",
  48119=>"010001011",
  48120=>"010101101",
  48121=>"011000001",
  48122=>"000010001",
  48123=>"110100100",
  48124=>"010000100",
  48125=>"011100011",
  48126=>"110010001",
  48127=>"011011100",
  48128=>"101001100",
  48129=>"110010101",
  48130=>"011110110",
  48131=>"000000000",
  48132=>"111010001",
  48133=>"000001110",
  48134=>"001010000",
  48135=>"101000100",
  48136=>"011011001",
  48137=>"100101110",
  48138=>"110011101",
  48139=>"100001101",
  48140=>"010100111",
  48141=>"000000101",
  48142=>"010010001",
  48143=>"010111100",
  48144=>"001110101",
  48145=>"101101001",
  48146=>"011011110",
  48147=>"001100001",
  48148=>"100000000",
  48149=>"001011010",
  48150=>"110010000",
  48151=>"010111101",
  48152=>"111000011",
  48153=>"000010110",
  48154=>"011010010",
  48155=>"010111101",
  48156=>"110001101",
  48157=>"010010110",
  48158=>"101001000",
  48159=>"010011010",
  48160=>"011111000",
  48161=>"000000011",
  48162=>"001001100",
  48163=>"110000110",
  48164=>"010101011",
  48165=>"000000010",
  48166=>"101001001",
  48167=>"111001000",
  48168=>"001110010",
  48169=>"010010110",
  48170=>"101101000",
  48171=>"000011010",
  48172=>"110100001",
  48173=>"001111111",
  48174=>"001000111",
  48175=>"010000110",
  48176=>"101000100",
  48177=>"111011001",
  48178=>"101100011",
  48179=>"010001110",
  48180=>"010011111",
  48181=>"000010110",
  48182=>"010000100",
  48183=>"110111101",
  48184=>"001000000",
  48185=>"001100110",
  48186=>"100000110",
  48187=>"010000010",
  48188=>"111110000",
  48189=>"000101011",
  48190=>"001100011",
  48191=>"100111010",
  48192=>"100010000",
  48193=>"001110111",
  48194=>"001111100",
  48195=>"010000001",
  48196=>"011110010",
  48197=>"001001111",
  48198=>"010101101",
  48199=>"110110111",
  48200=>"110101110",
  48201=>"101001011",
  48202=>"001100000",
  48203=>"011011110",
  48204=>"011001111",
  48205=>"100101101",
  48206=>"100010010",
  48207=>"000111001",
  48208=>"001101111",
  48209=>"000000000",
  48210=>"110101110",
  48211=>"000011111",
  48212=>"101111101",
  48213=>"100010000",
  48214=>"111000111",
  48215=>"000101011",
  48216=>"001101001",
  48217=>"100100110",
  48218=>"111000110",
  48219=>"011011111",
  48220=>"100111100",
  48221=>"110001101",
  48222=>"010010000",
  48223=>"000001011",
  48224=>"011001000",
  48225=>"000010100",
  48226=>"000001101",
  48227=>"111110101",
  48228=>"110111010",
  48229=>"000110001",
  48230=>"100011010",
  48231=>"101110110",
  48232=>"000111100",
  48233=>"001000111",
  48234=>"010001111",
  48235=>"000011100",
  48236=>"001101010",
  48237=>"001000100",
  48238=>"101100011",
  48239=>"000010001",
  48240=>"011000111",
  48241=>"001001001",
  48242=>"001000011",
  48243=>"110011010",
  48244=>"000010000",
  48245=>"001001100",
  48246=>"111111101",
  48247=>"101110011",
  48248=>"101010110",
  48249=>"111010000",
  48250=>"111111101",
  48251=>"011000011",
  48252=>"001001000",
  48253=>"101001110",
  48254=>"010110000",
  48255=>"000001010",
  48256=>"101000011",
  48257=>"000000100",
  48258=>"110010101",
  48259=>"011001110",
  48260=>"101100100",
  48261=>"001000100",
  48262=>"010011100",
  48263=>"011011000",
  48264=>"101001110",
  48265=>"001111011",
  48266=>"101001011",
  48267=>"101010100",
  48268=>"100101011",
  48269=>"000101000",
  48270=>"001100000",
  48271=>"010000001",
  48272=>"011101101",
  48273=>"110110100",
  48274=>"111001010",
  48275=>"110011110",
  48276=>"100011111",
  48277=>"101001000",
  48278=>"101101110",
  48279=>"001100111",
  48280=>"101001101",
  48281=>"111100001",
  48282=>"111011001",
  48283=>"000010101",
  48284=>"010111101",
  48285=>"111101000",
  48286=>"111011111",
  48287=>"011110010",
  48288=>"110111101",
  48289=>"100001110",
  48290=>"001110010",
  48291=>"111111000",
  48292=>"000011001",
  48293=>"011100011",
  48294=>"001011010",
  48295=>"011011001",
  48296=>"010111101",
  48297=>"111000010",
  48298=>"101000100",
  48299=>"111100100",
  48300=>"111011001",
  48301=>"010011010",
  48302=>"111011101",
  48303=>"001010000",
  48304=>"110110001",
  48305=>"111001100",
  48306=>"001001011",
  48307=>"001010100",
  48308=>"001100100",
  48309=>"000001010",
  48310=>"001101101",
  48311=>"000100000",
  48312=>"011101011",
  48313=>"101111100",
  48314=>"100110100",
  48315=>"010100000",
  48316=>"000001101",
  48317=>"000001010",
  48318=>"111111100",
  48319=>"110000001",
  48320=>"011011100",
  48321=>"001110111",
  48322=>"000100100",
  48323=>"010111111",
  48324=>"101110110",
  48325=>"101110000",
  48326=>"001001011",
  48327=>"001011011",
  48328=>"000100101",
  48329=>"100011010",
  48330=>"000101011",
  48331=>"110101011",
  48332=>"001010100",
  48333=>"010010101",
  48334=>"110001011",
  48335=>"110101101",
  48336=>"111110101",
  48337=>"110101101",
  48338=>"001001101",
  48339=>"010010010",
  48340=>"000000110",
  48341=>"001010001",
  48342=>"100110011",
  48343=>"010001111",
  48344=>"101000110",
  48345=>"010011110",
  48346=>"111000000",
  48347=>"100110001",
  48348=>"111110010",
  48349=>"100111111",
  48350=>"111101111",
  48351=>"100110010",
  48352=>"110000000",
  48353=>"111110001",
  48354=>"101011000",
  48355=>"001000000",
  48356=>"010010000",
  48357=>"111000110",
  48358=>"011111100",
  48359=>"011110001",
  48360=>"001000101",
  48361=>"010100011",
  48362=>"011001110",
  48363=>"011000101",
  48364=>"000111001",
  48365=>"001000011",
  48366=>"101111111",
  48367=>"110000000",
  48368=>"010100101",
  48369=>"010110000",
  48370=>"111111110",
  48371=>"101110011",
  48372=>"000001001",
  48373=>"101011000",
  48374=>"110111100",
  48375=>"100110100",
  48376=>"111011011",
  48377=>"110001000",
  48378=>"010011101",
  48379=>"011001110",
  48380=>"001000001",
  48381=>"111111000",
  48382=>"011111101",
  48383=>"010000001",
  48384=>"100010010",
  48385=>"100000100",
  48386=>"100110100",
  48387=>"110100000",
  48388=>"011011110",
  48389=>"000001100",
  48390=>"100011111",
  48391=>"100000111",
  48392=>"101101010",
  48393=>"000001001",
  48394=>"111111001",
  48395=>"100011111",
  48396=>"000000010",
  48397=>"111011111",
  48398=>"011000100",
  48399=>"110100011",
  48400=>"010101011",
  48401=>"010100110",
  48402=>"101010000",
  48403=>"000111000",
  48404=>"100100100",
  48405=>"000110000",
  48406=>"100010101",
  48407=>"000100111",
  48408=>"111011001",
  48409=>"111000111",
  48410=>"100010101",
  48411=>"101110000",
  48412=>"111100001",
  48413=>"111001101",
  48414=>"111110000",
  48415=>"110101001",
  48416=>"000100111",
  48417=>"001111000",
  48418=>"111101100",
  48419=>"100001101",
  48420=>"111011011",
  48421=>"110001000",
  48422=>"110011000",
  48423=>"010001111",
  48424=>"010111000",
  48425=>"110010111",
  48426=>"101101101",
  48427=>"000010010",
  48428=>"010010111",
  48429=>"100100111",
  48430=>"000111000",
  48431=>"111100011",
  48432=>"101100010",
  48433=>"101000000",
  48434=>"110010110",
  48435=>"000011111",
  48436=>"111000010",
  48437=>"001111010",
  48438=>"011111111",
  48439=>"010000001",
  48440=>"000110000",
  48441=>"111101110",
  48442=>"000011000",
  48443=>"000101111",
  48444=>"110100100",
  48445=>"111100010",
  48446=>"110110010",
  48447=>"000100001",
  48448=>"010011000",
  48449=>"101100101",
  48450=>"000111100",
  48451=>"000110101",
  48452=>"110100011",
  48453=>"011010111",
  48454=>"111110110",
  48455=>"100011010",
  48456=>"000101111",
  48457=>"011100001",
  48458=>"010000100",
  48459=>"110110001",
  48460=>"011010111",
  48461=>"100110111",
  48462=>"001000000",
  48463=>"100101101",
  48464=>"100110010",
  48465=>"011111101",
  48466=>"011000000",
  48467=>"011111101",
  48468=>"100101000",
  48469=>"001100110",
  48470=>"101000000",
  48471=>"001011000",
  48472=>"001101000",
  48473=>"111011101",
  48474=>"111110011",
  48475=>"001101101",
  48476=>"110101111",
  48477=>"111000010",
  48478=>"001000101",
  48479=>"100011010",
  48480=>"011110110",
  48481=>"110110101",
  48482=>"110000000",
  48483=>"000011000",
  48484=>"011111111",
  48485=>"001100111",
  48486=>"011000011",
  48487=>"110000101",
  48488=>"010101011",
  48489=>"110100000",
  48490=>"000001110",
  48491=>"001111001",
  48492=>"100100110",
  48493=>"111000011",
  48494=>"000000010",
  48495=>"110010101",
  48496=>"010111100",
  48497=>"101110100",
  48498=>"001110100",
  48499=>"010100100",
  48500=>"111011101",
  48501=>"001110000",
  48502=>"000010000",
  48503=>"101110010",
  48504=>"010100000",
  48505=>"101101110",
  48506=>"001101011",
  48507=>"101101001",
  48508=>"100011110",
  48509=>"111111001",
  48510=>"111110101",
  48511=>"011101011",
  48512=>"010010101",
  48513=>"100001010",
  48514=>"100010101",
  48515=>"010011110",
  48516=>"111101110",
  48517=>"001110011",
  48518=>"010100101",
  48519=>"101000011",
  48520=>"111110100",
  48521=>"011010001",
  48522=>"000000001",
  48523=>"011000100",
  48524=>"011000000",
  48525=>"110001001",
  48526=>"111011111",
  48527=>"010010100",
  48528=>"001000100",
  48529=>"010001111",
  48530=>"000000010",
  48531=>"010111001",
  48532=>"100111100",
  48533=>"000010101",
  48534=>"001011101",
  48535=>"110100110",
  48536=>"110111011",
  48537=>"011101000",
  48538=>"011001010",
  48539=>"111111000",
  48540=>"110011011",
  48541=>"001101011",
  48542=>"011010000",
  48543=>"110000110",
  48544=>"010011001",
  48545=>"110011111",
  48546=>"001110100",
  48547=>"110001001",
  48548=>"110001111",
  48549=>"001111111",
  48550=>"011111101",
  48551=>"111101110",
  48552=>"101000101",
  48553=>"100000010",
  48554=>"100011101",
  48555=>"100010100",
  48556=>"000110011",
  48557=>"010111101",
  48558=>"100110010",
  48559=>"110101010",
  48560=>"001001101",
  48561=>"010011000",
  48562=>"101001111",
  48563=>"100011001",
  48564=>"000110001",
  48565=>"110111001",
  48566=>"111011001",
  48567=>"101100010",
  48568=>"010111100",
  48569=>"101011111",
  48570=>"001010000",
  48571=>"001101101",
  48572=>"101001001",
  48573=>"101111110",
  48574=>"110101110",
  48575=>"000110010",
  48576=>"011010111",
  48577=>"100001101",
  48578=>"011001101",
  48579=>"111000011",
  48580=>"110011110",
  48581=>"000000111",
  48582=>"101001111",
  48583=>"000011000",
  48584=>"100110001",
  48585=>"101110001",
  48586=>"111111111",
  48587=>"110010000",
  48588=>"010010001",
  48589=>"111011100",
  48590=>"101111101",
  48591=>"000010001",
  48592=>"000010001",
  48593=>"100000010",
  48594=>"111111110",
  48595=>"100111111",
  48596=>"111110110",
  48597=>"010111001",
  48598=>"110001010",
  48599=>"110111001",
  48600=>"001010110",
  48601=>"010101000",
  48602=>"010011000",
  48603=>"000011110",
  48604=>"101100100",
  48605=>"111011001",
  48606=>"101110010",
  48607=>"101001100",
  48608=>"111011010",
  48609=>"010111011",
  48610=>"011010110",
  48611=>"110000110",
  48612=>"101101011",
  48613=>"000110011",
  48614=>"111100000",
  48615=>"000010010",
  48616=>"010111110",
  48617=>"100101010",
  48618=>"010100101",
  48619=>"000100000",
  48620=>"100001111",
  48621=>"111111101",
  48622=>"010011101",
  48623=>"101000010",
  48624=>"101100010",
  48625=>"011001111",
  48626=>"101000001",
  48627=>"001000110",
  48628=>"100000000",
  48629=>"101010010",
  48630=>"111000000",
  48631=>"100110110",
  48632=>"010110101",
  48633=>"100110000",
  48634=>"001111101",
  48635=>"001101100",
  48636=>"101010110",
  48637=>"001110011",
  48638=>"010111000",
  48639=>"000010000",
  48640=>"000011100",
  48641=>"100111111",
  48642=>"110100010",
  48643=>"110001010",
  48644=>"001100101",
  48645=>"100010000",
  48646=>"011001001",
  48647=>"110001110",
  48648=>"010110100",
  48649=>"101110101",
  48650=>"000000100",
  48651=>"001000100",
  48652=>"010010010",
  48653=>"110011111",
  48654=>"101010100",
  48655=>"001001110",
  48656=>"010111111",
  48657=>"000100100",
  48658=>"101000010",
  48659=>"110000011",
  48660=>"010001101",
  48661=>"110010001",
  48662=>"000100011",
  48663=>"010110010",
  48664=>"100100110",
  48665=>"110101010",
  48666=>"011001011",
  48667=>"010111001",
  48668=>"101110111",
  48669=>"110000000",
  48670=>"101011111",
  48671=>"110100010",
  48672=>"011110100",
  48673=>"001000010",
  48674=>"011101110",
  48675=>"000100101",
  48676=>"001100000",
  48677=>"011010011",
  48678=>"111011000",
  48679=>"000000010",
  48680=>"001000010",
  48681=>"100101101",
  48682=>"001011101",
  48683=>"001110001",
  48684=>"011101101",
  48685=>"010000110",
  48686=>"011111001",
  48687=>"010001110",
  48688=>"111100100",
  48689=>"000011001",
  48690=>"110110100",
  48691=>"110101011",
  48692=>"001101111",
  48693=>"111010001",
  48694=>"000011000",
  48695=>"000010101",
  48696=>"011111010",
  48697=>"011001011",
  48698=>"001100111",
  48699=>"001111000",
  48700=>"101011111",
  48701=>"100100011",
  48702=>"111011000",
  48703=>"011010011",
  48704=>"100100011",
  48705=>"101110000",
  48706=>"001110110",
  48707=>"001010111",
  48708=>"011011001",
  48709=>"011000001",
  48710=>"111101101",
  48711=>"010100100",
  48712=>"001111001",
  48713=>"101111111",
  48714=>"010001111",
  48715=>"010010100",
  48716=>"000110110",
  48717=>"101111101",
  48718=>"011010011",
  48719=>"000110110",
  48720=>"011110100",
  48721=>"010000110",
  48722=>"101111100",
  48723=>"100011110",
  48724=>"000110010",
  48725=>"001001000",
  48726=>"011001011",
  48727=>"010001010",
  48728=>"110111001",
  48729=>"001101000",
  48730=>"010110000",
  48731=>"001111101",
  48732=>"001010000",
  48733=>"100001010",
  48734=>"000101010",
  48735=>"000101000",
  48736=>"001110001",
  48737=>"100001111",
  48738=>"001001111",
  48739=>"000110100",
  48740=>"100100000",
  48741=>"001000110",
  48742=>"100111110",
  48743=>"000000110",
  48744=>"000110011",
  48745=>"101110100",
  48746=>"011010001",
  48747=>"000101010",
  48748=>"001011001",
  48749=>"101110000",
  48750=>"101111010",
  48751=>"110100010",
  48752=>"011101010",
  48753=>"000000000",
  48754=>"011101100",
  48755=>"001001100",
  48756=>"010010100",
  48757=>"100000100",
  48758=>"010101000",
  48759=>"001110100",
  48760=>"010011010",
  48761=>"011100001",
  48762=>"010100010",
  48763=>"111100010",
  48764=>"110000110",
  48765=>"001110100",
  48766=>"010110001",
  48767=>"110010010",
  48768=>"010101010",
  48769=>"011111100",
  48770=>"011101100",
  48771=>"110001011",
  48772=>"101100100",
  48773=>"011100110",
  48774=>"001100110",
  48775=>"010000100",
  48776=>"000110000",
  48777=>"001010101",
  48778=>"010110001",
  48779=>"100110101",
  48780=>"100101110",
  48781=>"110000110",
  48782=>"110010001",
  48783=>"101100111",
  48784=>"111100010",
  48785=>"011011010",
  48786=>"110100110",
  48787=>"110001110",
  48788=>"110001000",
  48789=>"110111111",
  48790=>"101001111",
  48791=>"010111111",
  48792=>"110111001",
  48793=>"110011011",
  48794=>"101010101",
  48795=>"000011010",
  48796=>"100000110",
  48797=>"010111010",
  48798=>"111001000",
  48799=>"001000111",
  48800=>"110010101",
  48801=>"010100010",
  48802=>"001001010",
  48803=>"100010100",
  48804=>"000000001",
  48805=>"010111001",
  48806=>"000100100",
  48807=>"111101000",
  48808=>"111000100",
  48809=>"010001011",
  48810=>"110111000",
  48811=>"001110000",
  48812=>"100010100",
  48813=>"010000100",
  48814=>"010111101",
  48815=>"000000101",
  48816=>"010101011",
  48817=>"010011110",
  48818=>"101000000",
  48819=>"101011001",
  48820=>"001011011",
  48821=>"100010000",
  48822=>"111010101",
  48823=>"010000100",
  48824=>"111010100",
  48825=>"100010010",
  48826=>"010000000",
  48827=>"101110101",
  48828=>"101101001",
  48829=>"100110010",
  48830=>"001111111",
  48831=>"011000100",
  48832=>"111011000",
  48833=>"110000100",
  48834=>"100111000",
  48835=>"111010001",
  48836=>"100111110",
  48837=>"000001011",
  48838=>"001011001",
  48839=>"001001011",
  48840=>"000001110",
  48841=>"100110100",
  48842=>"000101010",
  48843=>"011110001",
  48844=>"011111101",
  48845=>"111011111",
  48846=>"111101110",
  48847=>"110100011",
  48848=>"001110010",
  48849=>"110000110",
  48850=>"000100110",
  48851=>"001001100",
  48852=>"111100110",
  48853=>"001010000",
  48854=>"000000001",
  48855=>"101010100",
  48856=>"000011010",
  48857=>"100100010",
  48858=>"011001010",
  48859=>"111101010",
  48860=>"101100001",
  48861=>"010100001",
  48862=>"000110100",
  48863=>"010010011",
  48864=>"111101001",
  48865=>"011110010",
  48866=>"001111100",
  48867=>"101111100",
  48868=>"000111101",
  48869=>"111000111",
  48870=>"111110101",
  48871=>"011110111",
  48872=>"110100010",
  48873=>"000010000",
  48874=>"010100110",
  48875=>"110101000",
  48876=>"001010101",
  48877=>"000000111",
  48878=>"100000000",
  48879=>"111111101",
  48880=>"101101100",
  48881=>"011000101",
  48882=>"101000101",
  48883=>"110001001",
  48884=>"111011100",
  48885=>"001100111",
  48886=>"001111000",
  48887=>"100000000",
  48888=>"001000000",
  48889=>"101000100",
  48890=>"000001100",
  48891=>"010011000",
  48892=>"000010001",
  48893=>"111111000",
  48894=>"000000110",
  48895=>"010110100",
  48896=>"001100010",
  48897=>"001100111",
  48898=>"001010000",
  48899=>"011000100",
  48900=>"010110101",
  48901=>"100100001",
  48902=>"111111010",
  48903=>"000101101",
  48904=>"011110100",
  48905=>"000111111",
  48906=>"101111010",
  48907=>"100000101",
  48908=>"100001001",
  48909=>"010000100",
  48910=>"110111000",
  48911=>"011001011",
  48912=>"111001000",
  48913=>"001010001",
  48914=>"000011011",
  48915=>"101101101",
  48916=>"110110100",
  48917=>"010000001",
  48918=>"111110110",
  48919=>"000100011",
  48920=>"010010100",
  48921=>"001100100",
  48922=>"111110000",
  48923=>"010011001",
  48924=>"101100100",
  48925=>"011010001",
  48926=>"010011000",
  48927=>"011011010",
  48928=>"000000111",
  48929=>"111100101",
  48930=>"110000101",
  48931=>"101101010",
  48932=>"001101100",
  48933=>"000010010",
  48934=>"110100110",
  48935=>"001011111",
  48936=>"010111111",
  48937=>"001010101",
  48938=>"010101011",
  48939=>"000110001",
  48940=>"111100010",
  48941=>"111101111",
  48942=>"111011110",
  48943=>"111110111",
  48944=>"100100001",
  48945=>"010000110",
  48946=>"100000001",
  48947=>"010101100",
  48948=>"000110010",
  48949=>"110101100",
  48950=>"000001000",
  48951=>"010111000",
  48952=>"011101001",
  48953=>"000001011",
  48954=>"110101010",
  48955=>"111101100",
  48956=>"000100001",
  48957=>"010010011",
  48958=>"110101101",
  48959=>"011110111",
  48960=>"010111010",
  48961=>"111000001",
  48962=>"101111100",
  48963=>"010111111",
  48964=>"100110111",
  48965=>"011110111",
  48966=>"001111100",
  48967=>"000010010",
  48968=>"001011011",
  48969=>"001100111",
  48970=>"110000000",
  48971=>"100101100",
  48972=>"101010000",
  48973=>"000010000",
  48974=>"100101110",
  48975=>"110101111",
  48976=>"111000100",
  48977=>"100101001",
  48978=>"000001000",
  48979=>"000100000",
  48980=>"101100001",
  48981=>"101001110",
  48982=>"100010000",
  48983=>"001010110",
  48984=>"010111100",
  48985=>"011110110",
  48986=>"011111101",
  48987=>"100000010",
  48988=>"100000101",
  48989=>"000100100",
  48990=>"010110111",
  48991=>"010010111",
  48992=>"110000110",
  48993=>"100000010",
  48994=>"111100010",
  48995=>"100010000",
  48996=>"100000000",
  48997=>"010110001",
  48998=>"110000101",
  48999=>"101100100",
  49000=>"011001110",
  49001=>"011110100",
  49002=>"010101100",
  49003=>"100000010",
  49004=>"101111101",
  49005=>"001011110",
  49006=>"000101011",
  49007=>"111110101",
  49008=>"101101010",
  49009=>"100110000",
  49010=>"110101001",
  49011=>"101010100",
  49012=>"001000000",
  49013=>"100011000",
  49014=>"010100110",
  49015=>"111001011",
  49016=>"010010011",
  49017=>"100111000",
  49018=>"101101001",
  49019=>"111110101",
  49020=>"000011010",
  49021=>"001011010",
  49022=>"100101010",
  49023=>"110101011",
  49024=>"001101010",
  49025=>"000000100",
  49026=>"010101110",
  49027=>"011001010",
  49028=>"110000000",
  49029=>"100101111",
  49030=>"111000101",
  49031=>"110010010",
  49032=>"001101000",
  49033=>"101110100",
  49034=>"000011010",
  49035=>"000000001",
  49036=>"011010110",
  49037=>"000010111",
  49038=>"101100001",
  49039=>"010111100",
  49040=>"100100011",
  49041=>"111111010",
  49042=>"000000000",
  49043=>"100000000",
  49044=>"100110010",
  49045=>"101000101",
  49046=>"010010110",
  49047=>"011101110",
  49048=>"000100001",
  49049=>"101100111",
  49050=>"001010000",
  49051=>"100000000",
  49052=>"001100110",
  49053=>"010111101",
  49054=>"001100101",
  49055=>"111110000",
  49056=>"100001101",
  49057=>"001100100",
  49058=>"011001001",
  49059=>"010101101",
  49060=>"110000011",
  49061=>"011111001",
  49062=>"111001111",
  49063=>"010011011",
  49064=>"011001110",
  49065=>"010011001",
  49066=>"101101110",
  49067=>"110000010",
  49068=>"111101110",
  49069=>"000001010",
  49070=>"010000111",
  49071=>"101000010",
  49072=>"100010010",
  49073=>"100001110",
  49074=>"000000110",
  49075=>"111111001",
  49076=>"000100010",
  49077=>"011000001",
  49078=>"110100000",
  49079=>"000101101",
  49080=>"000000010",
  49081=>"011000001",
  49082=>"101110001",
  49083=>"101100110",
  49084=>"110000101",
  49085=>"011011111",
  49086=>"100110011",
  49087=>"000101110",
  49088=>"111000100",
  49089=>"101101111",
  49090=>"111110101",
  49091=>"010111000",
  49092=>"100000111",
  49093=>"100100011",
  49094=>"001111000",
  49095=>"011001001",
  49096=>"101000111",
  49097=>"100110010",
  49098=>"110011111",
  49099=>"001101000",
  49100=>"001100110",
  49101=>"001001100",
  49102=>"000111101",
  49103=>"110111111",
  49104=>"100011010",
  49105=>"100001100",
  49106=>"011000110",
  49107=>"000000110",
  49108=>"110100010",
  49109=>"111111011",
  49110=>"111010001",
  49111=>"001110111",
  49112=>"111011001",
  49113=>"101100111",
  49114=>"111111000",
  49115=>"111011110",
  49116=>"010011101",
  49117=>"110000000",
  49118=>"001100101",
  49119=>"011001100",
  49120=>"100001100",
  49121=>"011110010",
  49122=>"110110001",
  49123=>"001000110",
  49124=>"010010001",
  49125=>"111110010",
  49126=>"010110101",
  49127=>"111100000",
  49128=>"001011010",
  49129=>"010100111",
  49130=>"011011110",
  49131=>"001101011",
  49132=>"101110000",
  49133=>"011000000",
  49134=>"111001110",
  49135=>"111100000",
  49136=>"111001111",
  49137=>"011011011",
  49138=>"000001010",
  49139=>"111000111",
  49140=>"100000000",
  49141=>"101000110",
  49142=>"010101110",
  49143=>"001100011",
  49144=>"011001010",
  49145=>"101010010",
  49146=>"101000100",
  49147=>"111000011",
  49148=>"010010010",
  49149=>"100100001",
  49150=>"111010110",
  49151=>"000000010",
  49152=>"111000000",
  49153=>"110110111",
  49154=>"110011100",
  49155=>"000100101",
  49156=>"011101100",
  49157=>"110011111",
  49158=>"010101110",
  49159=>"111001010",
  49160=>"110010001",
  49161=>"101001001",
  49162=>"101011001",
  49163=>"101100111",
  49164=>"111111100",
  49165=>"000001001",
  49166=>"101111010",
  49167=>"100000100",
  49168=>"100000000",
  49169=>"001100100",
  49170=>"111100011",
  49171=>"111101111",
  49172=>"000001000",
  49173=>"010001001",
  49174=>"111000111",
  49175=>"110110001",
  49176=>"010001000",
  49177=>"011100110",
  49178=>"010110110",
  49179=>"011000010",
  49180=>"001100000",
  49181=>"011010111",
  49182=>"100011110",
  49183=>"110010100",
  49184=>"000010000",
  49185=>"111111110",
  49186=>"110001011",
  49187=>"111100011",
  49188=>"011101011",
  49189=>"010101100",
  49190=>"011110110",
  49191=>"010111100",
  49192=>"101100001",
  49193=>"010001001",
  49194=>"011111110",
  49195=>"110110101",
  49196=>"001000111",
  49197=>"101001100",
  49198=>"101110110",
  49199=>"001111100",
  49200=>"000110101",
  49201=>"001111000",
  49202=>"110111111",
  49203=>"011110111",
  49204=>"001101111",
  49205=>"011100110",
  49206=>"001100101",
  49207=>"100100000",
  49208=>"010101101",
  49209=>"111100001",
  49210=>"110000101",
  49211=>"100000000",
  49212=>"010000100",
  49213=>"011100111",
  49214=>"001100000",
  49215=>"010110010",
  49216=>"111011110",
  49217=>"001000000",
  49218=>"111001100",
  49219=>"000000000",
  49220=>"011010010",
  49221=>"011110011",
  49222=>"011100000",
  49223=>"000110100",
  49224=>"001011101",
  49225=>"011110100",
  49226=>"001100000",
  49227=>"010101100",
  49228=>"010110011",
  49229=>"101110111",
  49230=>"110000110",
  49231=>"000000100",
  49232=>"011101101",
  49233=>"101101011",
  49234=>"000110111",
  49235=>"010110111",
  49236=>"001100101",
  49237=>"101111100",
  49238=>"000000010",
  49239=>"101110010",
  49240=>"111100111",
  49241=>"101101110",
  49242=>"100101111",
  49243=>"011101100",
  49244=>"111001010",
  49245=>"101000010",
  49246=>"010111011",
  49247=>"111100010",
  49248=>"010011001",
  49249=>"111010100",
  49250=>"001001100",
  49251=>"000111001",
  49252=>"011100101",
  49253=>"000000100",
  49254=>"100110111",
  49255=>"010000101",
  49256=>"111101101",
  49257=>"001110011",
  49258=>"000010100",
  49259=>"110110000",
  49260=>"101010000",
  49261=>"001011001",
  49262=>"110001001",
  49263=>"110001010",
  49264=>"011001100",
  49265=>"110010111",
  49266=>"100010001",
  49267=>"101111010",
  49268=>"110000110",
  49269=>"100110110",
  49270=>"000101110",
  49271=>"001000111",
  49272=>"100000010",
  49273=>"110110100",
  49274=>"110101100",
  49275=>"000100011",
  49276=>"010001111",
  49277=>"111001001",
  49278=>"010011101",
  49279=>"110010100",
  49280=>"100010000",
  49281=>"011110001",
  49282=>"110011101",
  49283=>"100001110",
  49284=>"110010001",
  49285=>"110111001",
  49286=>"000010110",
  49287=>"001101000",
  49288=>"010110101",
  49289=>"100100111",
  49290=>"001000010",
  49291=>"110000001",
  49292=>"000001011",
  49293=>"000000111",
  49294=>"110010111",
  49295=>"111111111",
  49296=>"001000111",
  49297=>"000100001",
  49298=>"000110010",
  49299=>"010000101",
  49300=>"110100111",
  49301=>"011100001",
  49302=>"011010100",
  49303=>"111011001",
  49304=>"110010010",
  49305=>"010000111",
  49306=>"000101000",
  49307=>"101111000",
  49308=>"000100010",
  49309=>"010011001",
  49310=>"110010000",
  49311=>"110010011",
  49312=>"111100100",
  49313=>"101101011",
  49314=>"000110101",
  49315=>"100100010",
  49316=>"010101100",
  49317=>"001110101",
  49318=>"011010101",
  49319=>"100010011",
  49320=>"000010010",
  49321=>"001001100",
  49322=>"010111011",
  49323=>"101101111",
  49324=>"010111111",
  49325=>"011001101",
  49326=>"010010101",
  49327=>"110101101",
  49328=>"011011001",
  49329=>"110001110",
  49330=>"010010001",
  49331=>"011001100",
  49332=>"001001010",
  49333=>"111000000",
  49334=>"100001010",
  49335=>"100011000",
  49336=>"101101101",
  49337=>"011010001",
  49338=>"010011111",
  49339=>"001110111",
  49340=>"010000101",
  49341=>"000100110",
  49342=>"111001111",
  49343=>"010111001",
  49344=>"000000111",
  49345=>"110000100",
  49346=>"000101101",
  49347=>"111010110",
  49348=>"110010100",
  49349=>"011000001",
  49350=>"110000010",
  49351=>"101110000",
  49352=>"000110111",
  49353=>"111111110",
  49354=>"111100000",
  49355=>"101100010",
  49356=>"110000011",
  49357=>"110010001",
  49358=>"011001100",
  49359=>"000111101",
  49360=>"101100100",
  49361=>"001110010",
  49362=>"010001111",
  49363=>"110101001",
  49364=>"100000110",
  49365=>"110001010",
  49366=>"001000111",
  49367=>"001101001",
  49368=>"111000000",
  49369=>"010101010",
  49370=>"100100100",
  49371=>"100010000",
  49372=>"101000101",
  49373=>"110101101",
  49374=>"010101010",
  49375=>"011001111",
  49376=>"000010010",
  49377=>"000010010",
  49378=>"111010001",
  49379=>"000100000",
  49380=>"000101001",
  49381=>"010111101",
  49382=>"001111000",
  49383=>"110000101",
  49384=>"011001100",
  49385=>"001100101",
  49386=>"000011000",
  49387=>"000101100",
  49388=>"011101100",
  49389=>"110000110",
  49390=>"100110110",
  49391=>"100010111",
  49392=>"100011001",
  49393=>"100011100",
  49394=>"100001111",
  49395=>"010000000",
  49396=>"010110100",
  49397=>"001000001",
  49398=>"000111010",
  49399=>"000010000",
  49400=>"001110111",
  49401=>"111101100",
  49402=>"001011010",
  49403=>"001001000",
  49404=>"010000000",
  49405=>"010000010",
  49406=>"110000011",
  49407=>"011101110",
  49408=>"010100011",
  49409=>"010100111",
  49410=>"111111101",
  49411=>"010101001",
  49412=>"000001000",
  49413=>"110011010",
  49414=>"101111001",
  49415=>"100110101",
  49416=>"001101111",
  49417=>"010011110",
  49418=>"011010110",
  49419=>"100011000",
  49420=>"001001000",
  49421=>"000111101",
  49422=>"110000011",
  49423=>"000001010",
  49424=>"100010000",
  49425=>"010110110",
  49426=>"000010110",
  49427=>"111110111",
  49428=>"000101001",
  49429=>"000101010",
  49430=>"100110001",
  49431=>"101011000",
  49432=>"001111000",
  49433=>"101100111",
  49434=>"100111001",
  49435=>"001010001",
  49436=>"010001001",
  49437=>"111010000",
  49438=>"111011111",
  49439=>"110011001",
  49440=>"001101101",
  49441=>"100011011",
  49442=>"000011011",
  49443=>"100101101",
  49444=>"110010011",
  49445=>"000011011",
  49446=>"010011010",
  49447=>"011101010",
  49448=>"000000110",
  49449=>"011101101",
  49450=>"000000000",
  49451=>"000110111",
  49452=>"010000000",
  49453=>"010101010",
  49454=>"101001010",
  49455=>"010100010",
  49456=>"001000100",
  49457=>"011100001",
  49458=>"000100101",
  49459=>"110010011",
  49460=>"111111100",
  49461=>"010111010",
  49462=>"101110111",
  49463=>"011100100",
  49464=>"000100000",
  49465=>"011010000",
  49466=>"100101101",
  49467=>"100110111",
  49468=>"110001011",
  49469=>"101101110",
  49470=>"011000000",
  49471=>"001001001",
  49472=>"110001001",
  49473=>"001100011",
  49474=>"010000011",
  49475=>"110111001",
  49476=>"100101010",
  49477=>"001001110",
  49478=>"011011000",
  49479=>"011100110",
  49480=>"011000010",
  49481=>"110110111",
  49482=>"000101001",
  49483=>"000110111",
  49484=>"011010001",
  49485=>"001011101",
  49486=>"001110010",
  49487=>"101111010",
  49488=>"001111101",
  49489=>"011000110",
  49490=>"001110001",
  49491=>"110110011",
  49492=>"101001000",
  49493=>"000110101",
  49494=>"100001110",
  49495=>"001001000",
  49496=>"100001010",
  49497=>"011001011",
  49498=>"011001000",
  49499=>"111000110",
  49500=>"011011101",
  49501=>"111111001",
  49502=>"000001100",
  49503=>"011010100",
  49504=>"001000011",
  49505=>"110010001",
  49506=>"010001011",
  49507=>"000100001",
  49508=>"111000111",
  49509=>"100000011",
  49510=>"010001001",
  49511=>"111101000",
  49512=>"101000110",
  49513=>"001011110",
  49514=>"000100110",
  49515=>"001001010",
  49516=>"111110100",
  49517=>"110100010",
  49518=>"010000011",
  49519=>"000000001",
  49520=>"010001001",
  49521=>"111011000",
  49522=>"001110010",
  49523=>"001000010",
  49524=>"101111111",
  49525=>"011000111",
  49526=>"111001100",
  49527=>"001000011",
  49528=>"010011001",
  49529=>"001011011",
  49530=>"011111111",
  49531=>"001010110",
  49532=>"001001011",
  49533=>"110000111",
  49534=>"100011001",
  49535=>"101111100",
  49536=>"001111000",
  49537=>"001010100",
  49538=>"110111010",
  49539=>"000010110",
  49540=>"111101110",
  49541=>"101101011",
  49542=>"000100101",
  49543=>"000011010",
  49544=>"101100001",
  49545=>"000011001",
  49546=>"000001111",
  49547=>"010001001",
  49548=>"110000100",
  49549=>"101111101",
  49550=>"110000010",
  49551=>"001011001",
  49552=>"010100000",
  49553=>"111000000",
  49554=>"000100111",
  49555=>"110111100",
  49556=>"110000111",
  49557=>"000001000",
  49558=>"100010110",
  49559=>"100100000",
  49560=>"101101001",
  49561=>"010000010",
  49562=>"100100000",
  49563=>"001101011",
  49564=>"110100101",
  49565=>"001100000",
  49566=>"000011001",
  49567=>"111110001",
  49568=>"101010010",
  49569=>"111001010",
  49570=>"110100001",
  49571=>"110001011",
  49572=>"010100110",
  49573=>"111001000",
  49574=>"011010000",
  49575=>"010111001",
  49576=>"101101100",
  49577=>"000000101",
  49578=>"110000000",
  49579=>"001100010",
  49580=>"111110000",
  49581=>"001000001",
  49582=>"011110011",
  49583=>"000000101",
  49584=>"010000000",
  49585=>"111111000",
  49586=>"101010110",
  49587=>"110110100",
  49588=>"101001101",
  49589=>"010011000",
  49590=>"010101011",
  49591=>"010110010",
  49592=>"011011001",
  49593=>"001110111",
  49594=>"000010001",
  49595=>"110010000",
  49596=>"101010010",
  49597=>"101001101",
  49598=>"111100011",
  49599=>"111111101",
  49600=>"000001001",
  49601=>"000110111",
  49602=>"000110111",
  49603=>"000111011",
  49604=>"011101011",
  49605=>"011101101",
  49606=>"011111011",
  49607=>"100001010",
  49608=>"100101011",
  49609=>"011111111",
  49610=>"011111011",
  49611=>"011011001",
  49612=>"110110100",
  49613=>"010101000",
  49614=>"100100001",
  49615=>"010111000",
  49616=>"101011011",
  49617=>"001001110",
  49618=>"101000000",
  49619=>"011110110",
  49620=>"111011000",
  49621=>"001011001",
  49622=>"110101000",
  49623=>"100111001",
  49624=>"000010000",
  49625=>"111111101",
  49626=>"110100110",
  49627=>"101010110",
  49628=>"111100000",
  49629=>"101010011",
  49630=>"101110000",
  49631=>"010110011",
  49632=>"010100010",
  49633=>"111000110",
  49634=>"100010110",
  49635=>"111111110",
  49636=>"001110001",
  49637=>"001000101",
  49638=>"010001101",
  49639=>"011001010",
  49640=>"101001011",
  49641=>"001000011",
  49642=>"000001010",
  49643=>"010110001",
  49644=>"110111111",
  49645=>"000000000",
  49646=>"001101111",
  49647=>"101000011",
  49648=>"110111011",
  49649=>"100100111",
  49650=>"100011101",
  49651=>"001100000",
  49652=>"000000010",
  49653=>"100000110",
  49654=>"011010000",
  49655=>"101110100",
  49656=>"100001001",
  49657=>"101011110",
  49658=>"111001110",
  49659=>"001010100",
  49660=>"001000101",
  49661=>"110011101",
  49662=>"110001111",
  49663=>"101010000",
  49664=>"000110100",
  49665=>"110110110",
  49666=>"111010111",
  49667=>"101100000",
  49668=>"100110101",
  49669=>"001010111",
  49670=>"101100100",
  49671=>"111101110",
  49672=>"011011100",
  49673=>"011010101",
  49674=>"110111001",
  49675=>"100000110",
  49676=>"101100100",
  49677=>"000000011",
  49678=>"000001110",
  49679=>"101000011",
  49680=>"110011110",
  49681=>"111100010",
  49682=>"111100110",
  49683=>"101011100",
  49684=>"000000001",
  49685=>"011100011",
  49686=>"010001010",
  49687=>"100001110",
  49688=>"010000110",
  49689=>"010001101",
  49690=>"010011100",
  49691=>"101001101",
  49692=>"100000010",
  49693=>"011011110",
  49694=>"111110011",
  49695=>"111111110",
  49696=>"000110011",
  49697=>"101000010",
  49698=>"000000011",
  49699=>"011000001",
  49700=>"000101111",
  49701=>"011001111",
  49702=>"011000010",
  49703=>"010111010",
  49704=>"001001100",
  49705=>"100110010",
  49706=>"010011111",
  49707=>"000101011",
  49708=>"100001100",
  49709=>"100011001",
  49710=>"001111000",
  49711=>"101100010",
  49712=>"001000100",
  49713=>"111011110",
  49714=>"100011110",
  49715=>"011010001",
  49716=>"111100000",
  49717=>"010000001",
  49718=>"000000011",
  49719=>"111001110",
  49720=>"111100101",
  49721=>"111100010",
  49722=>"010100110",
  49723=>"100110001",
  49724=>"010100100",
  49725=>"100010111",
  49726=>"000001110",
  49727=>"001011010",
  49728=>"110000011",
  49729=>"011110000",
  49730=>"100000000",
  49731=>"111101111",
  49732=>"011001100",
  49733=>"101000010",
  49734=>"001100100",
  49735=>"010001000",
  49736=>"010111110",
  49737=>"101110111",
  49738=>"111001001",
  49739=>"010110100",
  49740=>"101110110",
  49741=>"001101001",
  49742=>"110001111",
  49743=>"100100100",
  49744=>"011010010",
  49745=>"100110100",
  49746=>"101010111",
  49747=>"110110110",
  49748=>"100111000",
  49749=>"100110101",
  49750=>"111010010",
  49751=>"100101000",
  49752=>"110001001",
  49753=>"110010000",
  49754=>"101110111",
  49755=>"110100000",
  49756=>"010001011",
  49757=>"001010001",
  49758=>"001110110",
  49759=>"100111111",
  49760=>"100011001",
  49761=>"010000000",
  49762=>"110101110",
  49763=>"110101010",
  49764=>"100110100",
  49765=>"000001011",
  49766=>"011100101",
  49767=>"001100011",
  49768=>"010011101",
  49769=>"011000011",
  49770=>"001111010",
  49771=>"101010100",
  49772=>"010000110",
  49773=>"111000010",
  49774=>"000010101",
  49775=>"010001100",
  49776=>"011001001",
  49777=>"001001110",
  49778=>"011111101",
  49779=>"100000001",
  49780=>"111110110",
  49781=>"010111000",
  49782=>"001101011",
  49783=>"000111111",
  49784=>"100011011",
  49785=>"010111100",
  49786=>"111011011",
  49787=>"001110001",
  49788=>"001000101",
  49789=>"011000001",
  49790=>"111111001",
  49791=>"111110001",
  49792=>"011110101",
  49793=>"001001110",
  49794=>"101011110",
  49795=>"000001111",
  49796=>"000000110",
  49797=>"000110000",
  49798=>"101000001",
  49799=>"000010011",
  49800=>"011100000",
  49801=>"010000000",
  49802=>"111000101",
  49803=>"111111011",
  49804=>"110101110",
  49805=>"001110101",
  49806=>"110101000",
  49807=>"000101110",
  49808=>"110101010",
  49809=>"001100011",
  49810=>"001001001",
  49811=>"011011101",
  49812=>"110010111",
  49813=>"111011111",
  49814=>"111111000",
  49815=>"110110110",
  49816=>"110000100",
  49817=>"001011100",
  49818=>"011010100",
  49819=>"001011001",
  49820=>"101010011",
  49821=>"100010101",
  49822=>"010000010",
  49823=>"110000010",
  49824=>"011000101",
  49825=>"101101101",
  49826=>"000000111",
  49827=>"001010010",
  49828=>"101101001",
  49829=>"000101010",
  49830=>"111010101",
  49831=>"000001110",
  49832=>"100000101",
  49833=>"001010000",
  49834=>"110001100",
  49835=>"101111000",
  49836=>"110101111",
  49837=>"101000000",
  49838=>"001011010",
  49839=>"010010100",
  49840=>"000001101",
  49841=>"100010011",
  49842=>"110010101",
  49843=>"110001101",
  49844=>"011010010",
  49845=>"001111000",
  49846=>"011011001",
  49847=>"110001001",
  49848=>"111011111",
  49849=>"111011111",
  49850=>"001001011",
  49851=>"010111011",
  49852=>"110001011",
  49853=>"001110010",
  49854=>"000000100",
  49855=>"010100010",
  49856=>"111110111",
  49857=>"101011011",
  49858=>"000110011",
  49859=>"000100101",
  49860=>"010101111",
  49861=>"001011110",
  49862=>"101010001",
  49863=>"001001101",
  49864=>"011010110",
  49865=>"101111110",
  49866=>"001110010",
  49867=>"100100001",
  49868=>"000011011",
  49869=>"100001111",
  49870=>"000000011",
  49871=>"011001101",
  49872=>"000100011",
  49873=>"010001111",
  49874=>"111000010",
  49875=>"011010010",
  49876=>"001101001",
  49877=>"110001000",
  49878=>"011101100",
  49879=>"100100101",
  49880=>"001010000",
  49881=>"110100110",
  49882=>"010000001",
  49883=>"100111111",
  49884=>"101100010",
  49885=>"000001010",
  49886=>"100110110",
  49887=>"111010000",
  49888=>"001101010",
  49889=>"001011000",
  49890=>"000001111",
  49891=>"010001101",
  49892=>"111101010",
  49893=>"000101011",
  49894=>"000000111",
  49895=>"010001100",
  49896=>"000100101",
  49897=>"111001100",
  49898=>"010010010",
  49899=>"011011111",
  49900=>"010001011",
  49901=>"010111011",
  49902=>"000101111",
  49903=>"001001111",
  49904=>"011000000",
  49905=>"100010111",
  49906=>"111011001",
  49907=>"110111110",
  49908=>"110111111",
  49909=>"010000110",
  49910=>"000010011",
  49911=>"001000110",
  49912=>"110001010",
  49913=>"011001101",
  49914=>"111111101",
  49915=>"111100011",
  49916=>"100100110",
  49917=>"011010101",
  49918=>"010100000",
  49919=>"011101000",
  49920=>"000111110",
  49921=>"100100001",
  49922=>"010100011",
  49923=>"000000101",
  49924=>"000101011",
  49925=>"010000110",
  49926=>"100100111",
  49927=>"111101110",
  49928=>"011001110",
  49929=>"101011001",
  49930=>"010110100",
  49931=>"101111100",
  49932=>"111110001",
  49933=>"001111010",
  49934=>"011001011",
  49935=>"011011010",
  49936=>"111000110",
  49937=>"010100011",
  49938=>"111000100",
  49939=>"011001001",
  49940=>"001101111",
  49941=>"000010000",
  49942=>"001111101",
  49943=>"000110101",
  49944=>"011011010",
  49945=>"011000011",
  49946=>"000000111",
  49947=>"111011010",
  49948=>"100001001",
  49949=>"011101101",
  49950=>"101000000",
  49951=>"011111100",
  49952=>"100100000",
  49953=>"100010000",
  49954=>"011000000",
  49955=>"000010001",
  49956=>"001101011",
  49957=>"100100001",
  49958=>"111011001",
  49959=>"101010011",
  49960=>"000001100",
  49961=>"011100100",
  49962=>"111011001",
  49963=>"100010111",
  49964=>"000111011",
  49965=>"000000001",
  49966=>"111010100",
  49967=>"110001111",
  49968=>"000111001",
  49969=>"000110111",
  49970=>"110111001",
  49971=>"111101100",
  49972=>"101001100",
  49973=>"000001010",
  49974=>"111110000",
  49975=>"000110001",
  49976=>"111011011",
  49977=>"110010101",
  49978=>"000000101",
  49979=>"011011111",
  49980=>"001100001",
  49981=>"000000101",
  49982=>"101100101",
  49983=>"011101101",
  49984=>"101110100",
  49985=>"011111001",
  49986=>"100100000",
  49987=>"110001000",
  49988=>"000100001",
  49989=>"010001110",
  49990=>"100110001",
  49991=>"100000111",
  49992=>"101100011",
  49993=>"001111001",
  49994=>"010011001",
  49995=>"101000011",
  49996=>"010000010",
  49997=>"111101100",
  49998=>"001000010",
  49999=>"011101011",
  50000=>"111110000",
  50001=>"000110110",
  50002=>"100101100",
  50003=>"001101010",
  50004=>"001101000",
  50005=>"110000011",
  50006=>"001000000",
  50007=>"010000001",
  50008=>"010111001",
  50009=>"111010011",
  50010=>"110011000",
  50011=>"000010110",
  50012=>"010011011",
  50013=>"000000100",
  50014=>"110100001",
  50015=>"000000000",
  50016=>"010110101",
  50017=>"010001000",
  50018=>"000010000",
  50019=>"100001001",
  50020=>"100000001",
  50021=>"111101111",
  50022=>"100110010",
  50023=>"001011100",
  50024=>"111000000",
  50025=>"100000110",
  50026=>"100011010",
  50027=>"001010111",
  50028=>"110000110",
  50029=>"110001110",
  50030=>"000101000",
  50031=>"110110111",
  50032=>"111000111",
  50033=>"001001111",
  50034=>"000100111",
  50035=>"001100001",
  50036=>"000000011",
  50037=>"001111000",
  50038=>"001100101",
  50039=>"100110011",
  50040=>"100101100",
  50041=>"001010000",
  50042=>"101001010",
  50043=>"001110101",
  50044=>"000000100",
  50045=>"011001001",
  50046=>"111011001",
  50047=>"100111111",
  50048=>"110111001",
  50049=>"100101110",
  50050=>"111001100",
  50051=>"100101101",
  50052=>"000001101",
  50053=>"010100011",
  50054=>"001001110",
  50055=>"110101100",
  50056=>"000010100",
  50057=>"010110101",
  50058=>"010110001",
  50059=>"010000101",
  50060=>"110011100",
  50061=>"001001100",
  50062=>"101001011",
  50063=>"101000110",
  50064=>"111101100",
  50065=>"010001010",
  50066=>"001110001",
  50067=>"111010010",
  50068=>"000011100",
  50069=>"000101110",
  50070=>"110011101",
  50071=>"101000011",
  50072=>"011100010",
  50073=>"111110000",
  50074=>"011010111",
  50075=>"101100011",
  50076=>"010000001",
  50077=>"111011100",
  50078=>"000100110",
  50079=>"100000100",
  50080=>"001000000",
  50081=>"100000000",
  50082=>"110010101",
  50083=>"011001111",
  50084=>"000000101",
  50085=>"010110010",
  50086=>"000110101",
  50087=>"011010000",
  50088=>"100100001",
  50089=>"011010110",
  50090=>"000010000",
  50091=>"011001110",
  50092=>"111000010",
  50093=>"001110110",
  50094=>"000001101",
  50095=>"010010010",
  50096=>"011001010",
  50097=>"010010110",
  50098=>"000100111",
  50099=>"010000111",
  50100=>"011010100",
  50101=>"100001110",
  50102=>"111111011",
  50103=>"011100000",
  50104=>"111110110",
  50105=>"010011000",
  50106=>"100110010",
  50107=>"010010100",
  50108=>"010101000",
  50109=>"111101110",
  50110=>"111101000",
  50111=>"101100100",
  50112=>"000100110",
  50113=>"100100110",
  50114=>"010101011",
  50115=>"001100010",
  50116=>"000100001",
  50117=>"010100011",
  50118=>"111000011",
  50119=>"001110101",
  50120=>"000110000",
  50121=>"110100010",
  50122=>"100011100",
  50123=>"001001001",
  50124=>"000101100",
  50125=>"111001110",
  50126=>"001011000",
  50127=>"010111100",
  50128=>"100101110",
  50129=>"101110100",
  50130=>"110111000",
  50131=>"001011010",
  50132=>"001011011",
  50133=>"001000101",
  50134=>"001101011",
  50135=>"001101011",
  50136=>"010011100",
  50137=>"100001010",
  50138=>"001011110",
  50139=>"111011110",
  50140=>"101111000",
  50141=>"010010011",
  50142=>"011001000",
  50143=>"100010110",
  50144=>"000100111",
  50145=>"010001111",
  50146=>"010110010",
  50147=>"010000111",
  50148=>"010100000",
  50149=>"000000000",
  50150=>"101111001",
  50151=>"100100010",
  50152=>"101101110",
  50153=>"010000001",
  50154=>"100000111",
  50155=>"000101011",
  50156=>"110111000",
  50157=>"000100111",
  50158=>"000111001",
  50159=>"100110101",
  50160=>"100000101",
  50161=>"100000110",
  50162=>"001111000",
  50163=>"001000000",
  50164=>"100011100",
  50165=>"010010111",
  50166=>"100110100",
  50167=>"011100111",
  50168=>"000001011",
  50169=>"011001001",
  50170=>"111000100",
  50171=>"111110101",
  50172=>"110100000",
  50173=>"100011011",
  50174=>"010111111",
  50175=>"001000010",
  50176=>"111111101",
  50177=>"101100111",
  50178=>"100001110",
  50179=>"010101001",
  50180=>"001111011",
  50181=>"111001101",
  50182=>"000110100",
  50183=>"101001000",
  50184=>"010011101",
  50185=>"110000101",
  50186=>"100001110",
  50187=>"011110101",
  50188=>"000011100",
  50189=>"100101001",
  50190=>"100010110",
  50191=>"110000110",
  50192=>"100100011",
  50193=>"011100010",
  50194=>"001001100",
  50195=>"001011110",
  50196=>"101001001",
  50197=>"000111000",
  50198=>"010010110",
  50199=>"101100101",
  50200=>"111010000",
  50201=>"001001000",
  50202=>"110100100",
  50203=>"011110010",
  50204=>"001001000",
  50205=>"011110111",
  50206=>"001010000",
  50207=>"000010001",
  50208=>"000000000",
  50209=>"000100110",
  50210=>"110001010",
  50211=>"111000001",
  50212=>"010110101",
  50213=>"100000100",
  50214=>"000011111",
  50215=>"100101001",
  50216=>"000011101",
  50217=>"010111101",
  50218=>"100011110",
  50219=>"000010001",
  50220=>"110101111",
  50221=>"111011101",
  50222=>"001011111",
  50223=>"101111111",
  50224=>"100101101",
  50225=>"110110011",
  50226=>"001001011",
  50227=>"010001101",
  50228=>"110000011",
  50229=>"000100011",
  50230=>"000100011",
  50231=>"011000000",
  50232=>"110000110",
  50233=>"001100000",
  50234=>"010111010",
  50235=>"001101000",
  50236=>"000100110",
  50237=>"011010000",
  50238=>"010000001",
  50239=>"000010010",
  50240=>"110000100",
  50241=>"011010101",
  50242=>"011100111",
  50243=>"001001111",
  50244=>"110111111",
  50245=>"101100001",
  50246=>"011011000",
  50247=>"111010010",
  50248=>"001101010",
  50249=>"100010011",
  50250=>"110100111",
  50251=>"001101010",
  50252=>"000110101",
  50253=>"110101000",
  50254=>"001111000",
  50255=>"010100110",
  50256=>"011111111",
  50257=>"110111110",
  50258=>"100110010",
  50259=>"100000001",
  50260=>"111110010",
  50261=>"101100010",
  50262=>"000011110",
  50263=>"100100101",
  50264=>"001011010",
  50265=>"011011000",
  50266=>"110001010",
  50267=>"110111001",
  50268=>"010001011",
  50269=>"001101110",
  50270=>"101011111",
  50271=>"011010001",
  50272=>"000100101",
  50273=>"111111001",
  50274=>"000110110",
  50275=>"000100001",
  50276=>"001101011",
  50277=>"101111101",
  50278=>"011001010",
  50279=>"110011010",
  50280=>"000101110",
  50281=>"010010110",
  50282=>"100001111",
  50283=>"001111101",
  50284=>"010100111",
  50285=>"001000000",
  50286=>"010000011",
  50287=>"100011000",
  50288=>"001000000",
  50289=>"000110000",
  50290=>"101101111",
  50291=>"111110101",
  50292=>"001010111",
  50293=>"011100110",
  50294=>"001111110",
  50295=>"111111011",
  50296=>"010000000",
  50297=>"000001101",
  50298=>"010111001",
  50299=>"011101000",
  50300=>"000100011",
  50301=>"111010101",
  50302=>"110111110",
  50303=>"100100000",
  50304=>"100001011",
  50305=>"100101011",
  50306=>"000010111",
  50307=>"100000111",
  50308=>"100101110",
  50309=>"111011001",
  50310=>"101110100",
  50311=>"100001010",
  50312=>"100010111",
  50313=>"101010011",
  50314=>"000101011",
  50315=>"110111011",
  50316=>"100000010",
  50317=>"011000101",
  50318=>"100000001",
  50319=>"011100110",
  50320=>"000000111",
  50321=>"111011100",
  50322=>"110111000",
  50323=>"001011000",
  50324=>"100000101",
  50325=>"100111000",
  50326=>"101100100",
  50327=>"110111000",
  50328=>"101011011",
  50329=>"001110111",
  50330=>"100101011",
  50331=>"101011101",
  50332=>"001010000",
  50333=>"010100100",
  50334=>"111100011",
  50335=>"001100011",
  50336=>"110001100",
  50337=>"111110111",
  50338=>"110110111",
  50339=>"111110001",
  50340=>"000010010",
  50341=>"011110000",
  50342=>"111001111",
  50343=>"001001011",
  50344=>"101101000",
  50345=>"101010010",
  50346=>"110111010",
  50347=>"010100111",
  50348=>"001100001",
  50349=>"111001110",
  50350=>"011111111",
  50351=>"110000011",
  50352=>"011000111",
  50353=>"000110100",
  50354=>"000100010",
  50355=>"101000011",
  50356=>"110001100",
  50357=>"010100101",
  50358=>"101111100",
  50359=>"010011100",
  50360=>"000101010",
  50361=>"010100101",
  50362=>"011001100",
  50363=>"010100100",
  50364=>"100111010",
  50365=>"111001111",
  50366=>"001111010",
  50367=>"000111011",
  50368=>"010110010",
  50369=>"101100110",
  50370=>"011001001",
  50371=>"011011000",
  50372=>"110010010",
  50373=>"101111001",
  50374=>"110011100",
  50375=>"010111011",
  50376=>"011101010",
  50377=>"101100111",
  50378=>"011101111",
  50379=>"100100010",
  50380=>"110010100",
  50381=>"101001100",
  50382=>"000000011",
  50383=>"100010011",
  50384=>"100100111",
  50385=>"100110100",
  50386=>"110100101",
  50387=>"011110101",
  50388=>"101000000",
  50389=>"110001010",
  50390=>"010000101",
  50391=>"001111100",
  50392=>"101110011",
  50393=>"100100111",
  50394=>"010110110",
  50395=>"100001110",
  50396=>"100010010",
  50397=>"101000001",
  50398=>"001011000",
  50399=>"111111001",
  50400=>"001000101",
  50401=>"010001110",
  50402=>"111111110",
  50403=>"111100100",
  50404=>"101010111",
  50405=>"110010111",
  50406=>"000100100",
  50407=>"010100010",
  50408=>"101011100",
  50409=>"001110011",
  50410=>"001010100",
  50411=>"100000010",
  50412=>"100111101",
  50413=>"110010001",
  50414=>"000111010",
  50415=>"101110011",
  50416=>"000000011",
  50417=>"110011111",
  50418=>"001001001",
  50419=>"011001100",
  50420=>"111111110",
  50421=>"000001001",
  50422=>"001111110",
  50423=>"000000011",
  50424=>"011111001",
  50425=>"100011010",
  50426=>"100011101",
  50427=>"110110100",
  50428=>"000010101",
  50429=>"000001100",
  50430=>"000011100",
  50431=>"101111011",
  50432=>"001000010",
  50433=>"000011100",
  50434=>"111110110",
  50435=>"100010011",
  50436=>"000000111",
  50437=>"000111111",
  50438=>"100010001",
  50439=>"000100111",
  50440=>"000110101",
  50441=>"000011101",
  50442=>"001011000",
  50443=>"110011000",
  50444=>"101101011",
  50445=>"011100101",
  50446=>"111110101",
  50447=>"000101101",
  50448=>"111010000",
  50449=>"101101000",
  50450=>"000011110",
  50451=>"000010101",
  50452=>"010000111",
  50453=>"001000011",
  50454=>"001101011",
  50455=>"010111000",
  50456=>"110000011",
  50457=>"000000101",
  50458=>"001000000",
  50459=>"000010000",
  50460=>"001011100",
  50461=>"111101101",
  50462=>"101100010",
  50463=>"000000001",
  50464=>"010011101",
  50465=>"010011010",
  50466=>"110110000",
  50467=>"000011000",
  50468=>"111101011",
  50469=>"010100110",
  50470=>"001000101",
  50471=>"001001100",
  50472=>"111011101",
  50473=>"101001100",
  50474=>"001111110",
  50475=>"111100110",
  50476=>"000000101",
  50477=>"100001000",
  50478=>"000000110",
  50479=>"010010110",
  50480=>"011111100",
  50481=>"000111110",
  50482=>"100000000",
  50483=>"110011111",
  50484=>"110110101",
  50485=>"100010000",
  50486=>"111101110",
  50487=>"101000001",
  50488=>"000100000",
  50489=>"011110000",
  50490=>"101110110",
  50491=>"100100100",
  50492=>"101111000",
  50493=>"110111110",
  50494=>"110000101",
  50495=>"000010011",
  50496=>"100100000",
  50497=>"110000110",
  50498=>"000000000",
  50499=>"000000011",
  50500=>"010010111",
  50501=>"011110110",
  50502=>"111100010",
  50503=>"000010111",
  50504=>"011010110",
  50505=>"000000001",
  50506=>"001101110",
  50507=>"100000100",
  50508=>"011100010",
  50509=>"101011100",
  50510=>"100010010",
  50511=>"110111101",
  50512=>"101011110",
  50513=>"111011011",
  50514=>"111111111",
  50515=>"101100011",
  50516=>"011100001",
  50517=>"000110010",
  50518=>"001100111",
  50519=>"110101100",
  50520=>"011010111",
  50521=>"010001011",
  50522=>"110110111",
  50523=>"101010101",
  50524=>"110000110",
  50525=>"110101110",
  50526=>"001101000",
  50527=>"010000110",
  50528=>"111101110",
  50529=>"101000001",
  50530=>"101101111",
  50531=>"100001110",
  50532=>"111000100",
  50533=>"010100110",
  50534=>"000001110",
  50535=>"000100111",
  50536=>"110010010",
  50537=>"101001011",
  50538=>"101001010",
  50539=>"010001111",
  50540=>"110111100",
  50541=>"001010110",
  50542=>"100000010",
  50543=>"001111011",
  50544=>"110101100",
  50545=>"000111110",
  50546=>"001000000",
  50547=>"101000101",
  50548=>"001101001",
  50549=>"101101101",
  50550=>"110101111",
  50551=>"010100111",
  50552=>"100110110",
  50553=>"111110110",
  50554=>"000110000",
  50555=>"110010001",
  50556=>"110100011",
  50557=>"101111000",
  50558=>"010100110",
  50559=>"100100101",
  50560=>"100100010",
  50561=>"001110001",
  50562=>"110111100",
  50563=>"100001001",
  50564=>"001111100",
  50565=>"110000111",
  50566=>"110111000",
  50567=>"100001011",
  50568=>"100000111",
  50569=>"111111010",
  50570=>"110101111",
  50571=>"111010001",
  50572=>"011001110",
  50573=>"000011110",
  50574=>"010000000",
  50575=>"010101000",
  50576=>"110000011",
  50577=>"001010110",
  50578=>"111101101",
  50579=>"100100110",
  50580=>"000001111",
  50581=>"100010011",
  50582=>"111100001",
  50583=>"001001101",
  50584=>"011111011",
  50585=>"001000001",
  50586=>"101101100",
  50587=>"010000101",
  50588=>"101110011",
  50589=>"000101000",
  50590=>"001010111",
  50591=>"111101011",
  50592=>"110011001",
  50593=>"010001000",
  50594=>"100101011",
  50595=>"000110100",
  50596=>"111111001",
  50597=>"000100110",
  50598=>"110011100",
  50599=>"010011010",
  50600=>"011001100",
  50601=>"001110101",
  50602=>"010100110",
  50603=>"100000001",
  50604=>"101000111",
  50605=>"001011101",
  50606=>"000100101",
  50607=>"111011011",
  50608=>"010100100",
  50609=>"111000110",
  50610=>"100100110",
  50611=>"011101001",
  50612=>"111101111",
  50613=>"111101010",
  50614=>"101111111",
  50615=>"010001000",
  50616=>"001110010",
  50617=>"000111010",
  50618=>"010101110",
  50619=>"110011110",
  50620=>"000110100",
  50621=>"110001000",
  50622=>"011011111",
  50623=>"010101111",
  50624=>"110001001",
  50625=>"011001001",
  50626=>"101011111",
  50627=>"101001010",
  50628=>"111101101",
  50629=>"010011000",
  50630=>"100010011",
  50631=>"110100000",
  50632=>"000000100",
  50633=>"001101010",
  50634=>"011001000",
  50635=>"111100010",
  50636=>"101110011",
  50637=>"111000101",
  50638=>"010111000",
  50639=>"101011010",
  50640=>"100111111",
  50641=>"011000010",
  50642=>"011010111",
  50643=>"001001011",
  50644=>"111101101",
  50645=>"001100001",
  50646=>"001011111",
  50647=>"111111111",
  50648=>"001000100",
  50649=>"001000001",
  50650=>"011101010",
  50651=>"110011110",
  50652=>"100010011",
  50653=>"010011111",
  50654=>"111000001",
  50655=>"100110101",
  50656=>"000010001",
  50657=>"001010111",
  50658=>"001001111",
  50659=>"110001001",
  50660=>"110010111",
  50661=>"011110000",
  50662=>"101101110",
  50663=>"000011011",
  50664=>"110111011",
  50665=>"000010001",
  50666=>"010010110",
  50667=>"011010010",
  50668=>"101110110",
  50669=>"101011111",
  50670=>"001011000",
  50671=>"110100110",
  50672=>"001000011",
  50673=>"110111001",
  50674=>"001011010",
  50675=>"000100100",
  50676=>"000111011",
  50677=>"111110100",
  50678=>"011100111",
  50679=>"011011001",
  50680=>"010100100",
  50681=>"110101111",
  50682=>"101011000",
  50683=>"101100000",
  50684=>"100100101",
  50685=>"111000011",
  50686=>"011010011",
  50687=>"110100010",
  50688=>"010100000",
  50689=>"111100000",
  50690=>"000001010",
  50691=>"011100000",
  50692=>"011111011",
  50693=>"100011001",
  50694=>"011001110",
  50695=>"100000001",
  50696=>"101101101",
  50697=>"110011011",
  50698=>"000101111",
  50699=>"010110111",
  50700=>"000001011",
  50701=>"110111100",
  50702=>"000011011",
  50703=>"110101111",
  50704=>"101010001",
  50705=>"000011010",
  50706=>"001110001",
  50707=>"101011000",
  50708=>"001000011",
  50709=>"100000100",
  50710=>"001110000",
  50711=>"000111110",
  50712=>"111011110",
  50713=>"010110011",
  50714=>"000000111",
  50715=>"010000010",
  50716=>"100001010",
  50717=>"001001010",
  50718=>"010011101",
  50719=>"100100001",
  50720=>"100110101",
  50721=>"101100101",
  50722=>"011010010",
  50723=>"110001101",
  50724=>"111100000",
  50725=>"101100110",
  50726=>"111111111",
  50727=>"100001001",
  50728=>"010001000",
  50729=>"111101110",
  50730=>"011001011",
  50731=>"010100111",
  50732=>"111100011",
  50733=>"100011100",
  50734=>"001011101",
  50735=>"100011001",
  50736=>"101100000",
  50737=>"101010001",
  50738=>"101000101",
  50739=>"110001010",
  50740=>"100001100",
  50741=>"000000011",
  50742=>"001100000",
  50743=>"010110010",
  50744=>"100010100",
  50745=>"111101111",
  50746=>"010100111",
  50747=>"100011000",
  50748=>"111011000",
  50749=>"011001011",
  50750=>"101001001",
  50751=>"111011100",
  50752=>"111011011",
  50753=>"100011001",
  50754=>"101001000",
  50755=>"000101101",
  50756=>"001001011",
  50757=>"100111001",
  50758=>"100110110",
  50759=>"110011111",
  50760=>"101001101",
  50761=>"110111111",
  50762=>"110001011",
  50763=>"111101111",
  50764=>"010000010",
  50765=>"011100111",
  50766=>"101100111",
  50767=>"110111100",
  50768=>"010010101",
  50769=>"000110010",
  50770=>"010111000",
  50771=>"001000110",
  50772=>"100000111",
  50773=>"011101000",
  50774=>"100100010",
  50775=>"111110111",
  50776=>"010001010",
  50777=>"111111000",
  50778=>"010101110",
  50779=>"110001001",
  50780=>"001101000",
  50781=>"001101101",
  50782=>"101010000",
  50783=>"101110000",
  50784=>"110111010",
  50785=>"111111011",
  50786=>"001100111",
  50787=>"100011111",
  50788=>"001000011",
  50789=>"010101100",
  50790=>"111110011",
  50791=>"010110001",
  50792=>"000010011",
  50793=>"101001101",
  50794=>"001100100",
  50795=>"010001011",
  50796=>"100010011",
  50797=>"010101111",
  50798=>"101110011",
  50799=>"010100100",
  50800=>"010010110",
  50801=>"000000000",
  50802=>"001100000",
  50803=>"001011100",
  50804=>"110101101",
  50805=>"001010111",
  50806=>"011010001",
  50807=>"110011000",
  50808=>"110111000",
  50809=>"000001111",
  50810=>"000110101",
  50811=>"100101011",
  50812=>"101111110",
  50813=>"111011111",
  50814=>"111110011",
  50815=>"011101101",
  50816=>"001011001",
  50817=>"100110011",
  50818=>"110011110",
  50819=>"001011111",
  50820=>"111111001",
  50821=>"000000000",
  50822=>"001010100",
  50823=>"000111011",
  50824=>"001000100",
  50825=>"010110100",
  50826=>"101001001",
  50827=>"110010001",
  50828=>"010000000",
  50829=>"000110111",
  50830=>"101111100",
  50831=>"110100100",
  50832=>"000010010",
  50833=>"000100110",
  50834=>"111100011",
  50835=>"001110110",
  50836=>"001101101",
  50837=>"100101100",
  50838=>"111010101",
  50839=>"011001000",
  50840=>"100010111",
  50841=>"110110110",
  50842=>"110110010",
  50843=>"011100010",
  50844=>"000001110",
  50845=>"101000000",
  50846=>"011001110",
  50847=>"011000010",
  50848=>"100101001",
  50849=>"110101100",
  50850=>"000111010",
  50851=>"010110001",
  50852=>"110110100",
  50853=>"101110111",
  50854=>"101010111",
  50855=>"110110101",
  50856=>"010010001",
  50857=>"101110110",
  50858=>"001010001",
  50859=>"111001100",
  50860=>"001001010",
  50861=>"010011000",
  50862=>"011000011",
  50863=>"101000000",
  50864=>"100011101",
  50865=>"000001011",
  50866=>"010000011",
  50867=>"111000101",
  50868=>"011010100",
  50869=>"001111000",
  50870=>"101001010",
  50871=>"100110100",
  50872=>"100001001",
  50873=>"111111100",
  50874=>"111011101",
  50875=>"101100001",
  50876=>"110010010",
  50877=>"100110101",
  50878=>"000001101",
  50879=>"001010001",
  50880=>"110111011",
  50881=>"011100101",
  50882=>"001000000",
  50883=>"110110111",
  50884=>"110011101",
  50885=>"000100111",
  50886=>"100100011",
  50887=>"010001001",
  50888=>"010000011",
  50889=>"101001111",
  50890=>"001000000",
  50891=>"010000001",
  50892=>"000001111",
  50893=>"011011010",
  50894=>"000010110",
  50895=>"010101100",
  50896=>"001010000",
  50897=>"000000111",
  50898=>"011011101",
  50899=>"000100110",
  50900=>"100101110",
  50901=>"011100010",
  50902=>"111100100",
  50903=>"001011110",
  50904=>"101101100",
  50905=>"011101011",
  50906=>"011111101",
  50907=>"111100110",
  50908=>"101000100",
  50909=>"011000001",
  50910=>"110101000",
  50911=>"110011110",
  50912=>"010101000",
  50913=>"000000111",
  50914=>"101111101",
  50915=>"110001110",
  50916=>"100111010",
  50917=>"101010000",
  50918=>"100010000",
  50919=>"001111010",
  50920=>"110100110",
  50921=>"111010011",
  50922=>"001010000",
  50923=>"010100001",
  50924=>"100100001",
  50925=>"111010010",
  50926=>"000010010",
  50927=>"111001101",
  50928=>"000101000",
  50929=>"100110011",
  50930=>"001111111",
  50931=>"001000000",
  50932=>"010001001",
  50933=>"000000000",
  50934=>"011100000",
  50935=>"110000101",
  50936=>"111011000",
  50937=>"101010110",
  50938=>"101101001",
  50939=>"010001101",
  50940=>"110011110",
  50941=>"011100111",
  50942=>"011101001",
  50943=>"100100101",
  50944=>"000110110",
  50945=>"001011011",
  50946=>"111111010",
  50947=>"111000011",
  50948=>"011110101",
  50949=>"010110110",
  50950=>"011111011",
  50951=>"011000100",
  50952=>"101100010",
  50953=>"000110001",
  50954=>"001000011",
  50955=>"110000000",
  50956=>"100010000",
  50957=>"011011011",
  50958=>"110001010",
  50959=>"110011100",
  50960=>"001010100",
  50961=>"100010100",
  50962=>"110110011",
  50963=>"101101011",
  50964=>"110100110",
  50965=>"000111010",
  50966=>"011101010",
  50967=>"001000011",
  50968=>"000000100",
  50969=>"000001001",
  50970=>"011001001",
  50971=>"110001110",
  50972=>"001111111",
  50973=>"111101010",
  50974=>"010000100",
  50975=>"010011101",
  50976=>"101011001",
  50977=>"110101000",
  50978=>"110000001",
  50979=>"110000000",
  50980=>"011111011",
  50981=>"101011001",
  50982=>"000000010",
  50983=>"101001010",
  50984=>"001001001",
  50985=>"110101000",
  50986=>"011110010",
  50987=>"010110010",
  50988=>"011011110",
  50989=>"010010001",
  50990=>"011011100",
  50991=>"101110011",
  50992=>"010011110",
  50993=>"100111111",
  50994=>"001000010",
  50995=>"000010111",
  50996=>"010101101",
  50997=>"111001011",
  50998=>"111100100",
  50999=>"001010101",
  51000=>"000000010",
  51001=>"001011011",
  51002=>"011111000",
  51003=>"111000000",
  51004=>"001110101",
  51005=>"000000101",
  51006=>"110001011",
  51007=>"101110110",
  51008=>"100010111",
  51009=>"011011010",
  51010=>"110101010",
  51011=>"100110000",
  51012=>"101000001",
  51013=>"101010001",
  51014=>"111001000",
  51015=>"101011101",
  51016=>"001000001",
  51017=>"110000110",
  51018=>"101000100",
  51019=>"100111011",
  51020=>"010011100",
  51021=>"101010100",
  51022=>"000010000",
  51023=>"100110111",
  51024=>"111111011",
  51025=>"011001111",
  51026=>"101101000",
  51027=>"010000110",
  51028=>"010000011",
  51029=>"011100011",
  51030=>"111001001",
  51031=>"101010001",
  51032=>"010011001",
  51033=>"111001110",
  51034=>"100010110",
  51035=>"101101010",
  51036=>"111100111",
  51037=>"100110100",
  51038=>"000010000",
  51039=>"100100101",
  51040=>"010111011",
  51041=>"110100101",
  51042=>"011100101",
  51043=>"011110011",
  51044=>"011111111",
  51045=>"010111000",
  51046=>"100000100",
  51047=>"010010011",
  51048=>"111000101",
  51049=>"100000111",
  51050=>"000110000",
  51051=>"000001111",
  51052=>"001100101",
  51053=>"011100111",
  51054=>"110000001",
  51055=>"000001000",
  51056=>"100100001",
  51057=>"001010010",
  51058=>"110001111",
  51059=>"010000101",
  51060=>"001101001",
  51061=>"110010010",
  51062=>"001010000",
  51063=>"110000011",
  51064=>"000100101",
  51065=>"001011011",
  51066=>"101111101",
  51067=>"010101011",
  51068=>"000010111",
  51069=>"111001001",
  51070=>"110001101",
  51071=>"111110001",
  51072=>"100110001",
  51073=>"001010101",
  51074=>"111100000",
  51075=>"111001111",
  51076=>"101000010",
  51077=>"010010111",
  51078=>"010000111",
  51079=>"001001011",
  51080=>"001101000",
  51081=>"001000011",
  51082=>"011100100",
  51083=>"001010111",
  51084=>"001011110",
  51085=>"000011011",
  51086=>"001000001",
  51087=>"010100110",
  51088=>"000111100",
  51089=>"001001110",
  51090=>"110100111",
  51091=>"011100110",
  51092=>"000010011",
  51093=>"011000101",
  51094=>"101000111",
  51095=>"000011000",
  51096=>"101100011",
  51097=>"101000100",
  51098=>"000101011",
  51099=>"111011100",
  51100=>"110111101",
  51101=>"100010011",
  51102=>"100000011",
  51103=>"000110100",
  51104=>"010101000",
  51105=>"011100101",
  51106=>"100100010",
  51107=>"001010111",
  51108=>"110000111",
  51109=>"111010111",
  51110=>"110010100",
  51111=>"001111011",
  51112=>"001011000",
  51113=>"111101101",
  51114=>"111110111",
  51115=>"000010010",
  51116=>"110011010",
  51117=>"100110100",
  51118=>"101000011",
  51119=>"000000101",
  51120=>"011010100",
  51121=>"011011000",
  51122=>"000100111",
  51123=>"010111100",
  51124=>"011101000",
  51125=>"000010111",
  51126=>"010011010",
  51127=>"000000000",
  51128=>"101000010",
  51129=>"110101101",
  51130=>"100110000",
  51131=>"000101101",
  51132=>"011000001",
  51133=>"011110111",
  51134=>"000000011",
  51135=>"000001010",
  51136=>"001011100",
  51137=>"001011001",
  51138=>"010000101",
  51139=>"100011100",
  51140=>"011010101",
  51141=>"000001100",
  51142=>"100001100",
  51143=>"100010011",
  51144=>"000011011",
  51145=>"011011010",
  51146=>"011110001",
  51147=>"000111010",
  51148=>"101100001",
  51149=>"011010010",
  51150=>"000000100",
  51151=>"000000100",
  51152=>"011111111",
  51153=>"101111111",
  51154=>"010000111",
  51155=>"110011011",
  51156=>"100011110",
  51157=>"001011000",
  51158=>"101110000",
  51159=>"001011111",
  51160=>"000001011",
  51161=>"010000111",
  51162=>"110110111",
  51163=>"011001111",
  51164=>"000100001",
  51165=>"001011000",
  51166=>"010000100",
  51167=>"111001000",
  51168=>"101001111",
  51169=>"110001100",
  51170=>"111101101",
  51171=>"001110011",
  51172=>"010110101",
  51173=>"111011100",
  51174=>"101011001",
  51175=>"000100000",
  51176=>"001011110",
  51177=>"111111100",
  51178=>"001101000",
  51179=>"111001101",
  51180=>"000111011",
  51181=>"001110001",
  51182=>"000101000",
  51183=>"010111100",
  51184=>"101111110",
  51185=>"111010100",
  51186=>"110100011",
  51187=>"111000110",
  51188=>"111010100",
  51189=>"001011111",
  51190=>"001100101",
  51191=>"010011011",
  51192=>"010010000",
  51193=>"110101011",
  51194=>"001001101",
  51195=>"000000000",
  51196=>"110011111",
  51197=>"111100011",
  51198=>"101000110",
  51199=>"000010011",
  51200=>"010000110",
  51201=>"001100101",
  51202=>"000101100",
  51203=>"100111100",
  51204=>"001111011",
  51205=>"100010101",
  51206=>"000101010",
  51207=>"111100000",
  51208=>"101100000",
  51209=>"101110110",
  51210=>"000000000",
  51211=>"111010000",
  51212=>"111100110",
  51213=>"101000110",
  51214=>"100110111",
  51215=>"110111101",
  51216=>"101100100",
  51217=>"110110011",
  51218=>"001111110",
  51219=>"101100000",
  51220=>"011011010",
  51221=>"011000111",
  51222=>"110111000",
  51223=>"010100000",
  51224=>"111101101",
  51225=>"101111110",
  51226=>"011000110",
  51227=>"110101101",
  51228=>"100000010",
  51229=>"001110110",
  51230=>"100001110",
  51231=>"110100111",
  51232=>"100011100",
  51233=>"111010000",
  51234=>"010001110",
  51235=>"001101001",
  51236=>"101101110",
  51237=>"110010010",
  51238=>"011110010",
  51239=>"011110010",
  51240=>"011111110",
  51241=>"000111111",
  51242=>"100000010",
  51243=>"001100111",
  51244=>"100110111",
  51245=>"101011001",
  51246=>"101101111",
  51247=>"100001110",
  51248=>"010111110",
  51249=>"100111011",
  51250=>"100101010",
  51251=>"100101101",
  51252=>"000011001",
  51253=>"011111001",
  51254=>"000011010",
  51255=>"010010111",
  51256=>"000001100",
  51257=>"010000100",
  51258=>"111000100",
  51259=>"011000000",
  51260=>"000000000",
  51261=>"101111001",
  51262=>"010110010",
  51263=>"101000101",
  51264=>"101000110",
  51265=>"011010101",
  51266=>"111101001",
  51267=>"100001001",
  51268=>"101111110",
  51269=>"101111110",
  51270=>"011010010",
  51271=>"101111110",
  51272=>"111101000",
  51273=>"111011110",
  51274=>"000001100",
  51275=>"010101011",
  51276=>"001101010",
  51277=>"100100010",
  51278=>"101111111",
  51279=>"111001011",
  51280=>"111100000",
  51281=>"001010100",
  51282=>"001111011",
  51283=>"110001001",
  51284=>"010100101",
  51285=>"110001100",
  51286=>"000100111",
  51287=>"000111001",
  51288=>"100100100",
  51289=>"010001100",
  51290=>"101011100",
  51291=>"001010000",
  51292=>"000100011",
  51293=>"111101010",
  51294=>"000100110",
  51295=>"011000100",
  51296=>"010100001",
  51297=>"010101100",
  51298=>"001000110",
  51299=>"001101110",
  51300=>"100000100",
  51301=>"100100001",
  51302=>"100110101",
  51303=>"000001100",
  51304=>"111110111",
  51305=>"011110001",
  51306=>"000000010",
  51307=>"101100000",
  51308=>"111011010",
  51309=>"111001001",
  51310=>"011011100",
  51311=>"000000010",
  51312=>"101001111",
  51313=>"010100101",
  51314=>"101111011",
  51315=>"001001000",
  51316=>"111110111",
  51317=>"000110101",
  51318=>"010010101",
  51319=>"001101111",
  51320=>"010011010",
  51321=>"001000110",
  51322=>"000110111",
  51323=>"001110010",
  51324=>"101010111",
  51325=>"001011001",
  51326=>"110000000",
  51327=>"000100001",
  51328=>"101101100",
  51329=>"011011001",
  51330=>"001010000",
  51331=>"110001100",
  51332=>"111000000",
  51333=>"110111100",
  51334=>"001010001",
  51335=>"000110011",
  51336=>"110111011",
  51337=>"110110101",
  51338=>"110100110",
  51339=>"010111110",
  51340=>"110001000",
  51341=>"011000101",
  51342=>"111111000",
  51343=>"001001101",
  51344=>"110001010",
  51345=>"100100000",
  51346=>"001100110",
  51347=>"011010001",
  51348=>"000001010",
  51349=>"100111000",
  51350=>"100000001",
  51351=>"111110001",
  51352=>"010001101",
  51353=>"100110111",
  51354=>"110110100",
  51355=>"110110101",
  51356=>"100111101",
  51357=>"010101010",
  51358=>"001000110",
  51359=>"111011100",
  51360=>"000001100",
  51361=>"001100011",
  51362=>"100010100",
  51363=>"100001011",
  51364=>"100110101",
  51365=>"000011100",
  51366=>"011001110",
  51367=>"010011010",
  51368=>"011001101",
  51369=>"001101100",
  51370=>"111100000",
  51371=>"100110010",
  51372=>"001111011",
  51373=>"010111110",
  51374=>"110110100",
  51375=>"111000110",
  51376=>"111111101",
  51377=>"110101000",
  51378=>"100110000",
  51379=>"110101110",
  51380=>"011001000",
  51381=>"111100111",
  51382=>"000100101",
  51383=>"111000001",
  51384=>"110111001",
  51385=>"011110110",
  51386=>"000100000",
  51387=>"100101101",
  51388=>"001011000",
  51389=>"001100000",
  51390=>"010011100",
  51391=>"111101110",
  51392=>"110000101",
  51393=>"100110001",
  51394=>"001101111",
  51395=>"000011111",
  51396=>"010100000",
  51397=>"010101111",
  51398=>"001001011",
  51399=>"000001000",
  51400=>"011011111",
  51401=>"010010011",
  51402=>"100001100",
  51403=>"101010001",
  51404=>"101110101",
  51405=>"011100010",
  51406=>"100101101",
  51407=>"101001111",
  51408=>"101100101",
  51409=>"101000111",
  51410=>"011000100",
  51411=>"101000011",
  51412=>"111010111",
  51413=>"010001000",
  51414=>"101110100",
  51415=>"110111000",
  51416=>"100001011",
  51417=>"000010000",
  51418=>"000001011",
  51419=>"000110100",
  51420=>"110110101",
  51421=>"100010110",
  51422=>"001010001",
  51423=>"001100110",
  51424=>"100101000",
  51425=>"100001111",
  51426=>"000111101",
  51427=>"111111000",
  51428=>"111011000",
  51429=>"001100101",
  51430=>"011011011",
  51431=>"111110101",
  51432=>"000000111",
  51433=>"110011111",
  51434=>"010100010",
  51435=>"000010010",
  51436=>"100111110",
  51437=>"111000010",
  51438=>"100001011",
  51439=>"001101111",
  51440=>"010010110",
  51441=>"100010111",
  51442=>"011010111",
  51443=>"010100001",
  51444=>"001111101",
  51445=>"010100100",
  51446=>"001101001",
  51447=>"000110010",
  51448=>"000101001",
  51449=>"100100011",
  51450=>"111000011",
  51451=>"000100001",
  51452=>"110100000",
  51453=>"100011001",
  51454=>"011010001",
  51455=>"000000000",
  51456=>"001011001",
  51457=>"001011010",
  51458=>"001010000",
  51459=>"010111001",
  51460=>"010100101",
  51461=>"001111001",
  51462=>"010111010",
  51463=>"101100100",
  51464=>"011000110",
  51465=>"010100110",
  51466=>"110011110",
  51467=>"100000000",
  51468=>"001011111",
  51469=>"111001100",
  51470=>"000001110",
  51471=>"111110000",
  51472=>"011011110",
  51473=>"001011000",
  51474=>"000000000",
  51475=>"111010111",
  51476=>"110110111",
  51477=>"111110011",
  51478=>"100001100",
  51479=>"100110010",
  51480=>"000101110",
  51481=>"000010011",
  51482=>"110100010",
  51483=>"000101101",
  51484=>"110011011",
  51485=>"111000000",
  51486=>"110010000",
  51487=>"100010000",
  51488=>"100000111",
  51489=>"100000001",
  51490=>"111011101",
  51491=>"001000111",
  51492=>"000101001",
  51493=>"010001110",
  51494=>"011000100",
  51495=>"101010000",
  51496=>"011101110",
  51497=>"110011111",
  51498=>"100010011",
  51499=>"100000000",
  51500=>"111010010",
  51501=>"000101110",
  51502=>"100011101",
  51503=>"101111100",
  51504=>"000001000",
  51505=>"110110010",
  51506=>"110100010",
  51507=>"010111000",
  51508=>"110000001",
  51509=>"011000110",
  51510=>"100011001",
  51511=>"010000101",
  51512=>"000111100",
  51513=>"110011000",
  51514=>"011000000",
  51515=>"001100101",
  51516=>"110110111",
  51517=>"000111000",
  51518=>"001110010",
  51519=>"011001100",
  51520=>"100011001",
  51521=>"111100011",
  51522=>"101111001",
  51523=>"110011000",
  51524=>"111101011",
  51525=>"010101111",
  51526=>"001100000",
  51527=>"100000100",
  51528=>"011111011",
  51529=>"001100100",
  51530=>"110101001",
  51531=>"000010010",
  51532=>"000000001",
  51533=>"000000101",
  51534=>"111001011",
  51535=>"000100111",
  51536=>"011100100",
  51537=>"011010100",
  51538=>"100010001",
  51539=>"100000000",
  51540=>"101011101",
  51541=>"001111101",
  51542=>"111100010",
  51543=>"001110010",
  51544=>"101011001",
  51545=>"001110111",
  51546=>"110001000",
  51547=>"101100010",
  51548=>"001001001",
  51549=>"111101011",
  51550=>"111100101",
  51551=>"001111100",
  51552=>"100100010",
  51553=>"111111110",
  51554=>"100101001",
  51555=>"000001101",
  51556=>"111010001",
  51557=>"100000011",
  51558=>"000001011",
  51559=>"100101000",
  51560=>"011011011",
  51561=>"000001111",
  51562=>"011000001",
  51563=>"110111010",
  51564=>"101110000",
  51565=>"011110011",
  51566=>"011011011",
  51567=>"011111111",
  51568=>"111001011",
  51569=>"000000011",
  51570=>"111100000",
  51571=>"001100100",
  51572=>"010101100",
  51573=>"001000111",
  51574=>"101000100",
  51575=>"010111111",
  51576=>"001010010",
  51577=>"010010011",
  51578=>"011110110",
  51579=>"111000010",
  51580=>"110001100",
  51581=>"111111001",
  51582=>"011101110",
  51583=>"011011111",
  51584=>"100111110",
  51585=>"010100111",
  51586=>"110110011",
  51587=>"100110100",
  51588=>"111010010",
  51589=>"100001110",
  51590=>"100000111",
  51591=>"110001101",
  51592=>"100001010",
  51593=>"111001010",
  51594=>"001000000",
  51595=>"001110111",
  51596=>"001000100",
  51597=>"100111100",
  51598=>"011111011",
  51599=>"111110001",
  51600=>"011110110",
  51601=>"111110001",
  51602=>"110101011",
  51603=>"101111101",
  51604=>"001010000",
  51605=>"010110101",
  51606=>"111001011",
  51607=>"010110101",
  51608=>"100110001",
  51609=>"001000000",
  51610=>"010000110",
  51611=>"100101010",
  51612=>"000000100",
  51613=>"000111101",
  51614=>"001000010",
  51615=>"001001010",
  51616=>"100011001",
  51617=>"001001001",
  51618=>"011111001",
  51619=>"000101010",
  51620=>"101011110",
  51621=>"011010010",
  51622=>"010110001",
  51623=>"111000100",
  51624=>"101011101",
  51625=>"000111001",
  51626=>"000101100",
  51627=>"000111100",
  51628=>"000111100",
  51629=>"111000110",
  51630=>"101011111",
  51631=>"111111011",
  51632=>"011111011",
  51633=>"111011111",
  51634=>"000011101",
  51635=>"111010000",
  51636=>"111000101",
  51637=>"100101000",
  51638=>"000101111",
  51639=>"111101111",
  51640=>"000000011",
  51641=>"000001111",
  51642=>"100010000",
  51643=>"101010110",
  51644=>"001100011",
  51645=>"100111101",
  51646=>"000011000",
  51647=>"001000000",
  51648=>"000010000",
  51649=>"100101111",
  51650=>"010000010",
  51651=>"100001010",
  51652=>"001000110",
  51653=>"111011010",
  51654=>"001111110",
  51655=>"000100110",
  51656=>"111100101",
  51657=>"101010101",
  51658=>"101101000",
  51659=>"100111101",
  51660=>"100000000",
  51661=>"000010111",
  51662=>"110010000",
  51663=>"101110100",
  51664=>"001001101",
  51665=>"100100001",
  51666=>"100000100",
  51667=>"000101110",
  51668=>"101100000",
  51669=>"110001110",
  51670=>"000000001",
  51671=>"001011000",
  51672=>"001010101",
  51673=>"100001101",
  51674=>"111100001",
  51675=>"000010101",
  51676=>"110110010",
  51677=>"100000001",
  51678=>"000001010",
  51679=>"111110100",
  51680=>"110001101",
  51681=>"011100011",
  51682=>"111011100",
  51683=>"000101101",
  51684=>"001000000",
  51685=>"000001110",
  51686=>"000011111",
  51687=>"101010101",
  51688=>"100111000",
  51689=>"101000110",
  51690=>"001000000",
  51691=>"110111101",
  51692=>"111001110",
  51693=>"001100000",
  51694=>"111000100",
  51695=>"100011010",
  51696=>"111001100",
  51697=>"010110010",
  51698=>"110110100",
  51699=>"111111111",
  51700=>"001100001",
  51701=>"101101010",
  51702=>"111010101",
  51703=>"111110001",
  51704=>"101100100",
  51705=>"100011010",
  51706=>"101001010",
  51707=>"100111010",
  51708=>"110101100",
  51709=>"111010110",
  51710=>"110110110",
  51711=>"100011001",
  51712=>"100111000",
  51713=>"110000001",
  51714=>"010111111",
  51715=>"000011011",
  51716=>"000010110",
  51717=>"100000100",
  51718=>"110011000",
  51719=>"101101011",
  51720=>"000100000",
  51721=>"100011101",
  51722=>"001010011",
  51723=>"110000100",
  51724=>"001000001",
  51725=>"011010000",
  51726=>"101001000",
  51727=>"100001011",
  51728=>"011101101",
  51729=>"010010010",
  51730=>"101011000",
  51731=>"101000000",
  51732=>"011111000",
  51733=>"000010110",
  51734=>"100110101",
  51735=>"101000000",
  51736=>"100000100",
  51737=>"110100000",
  51738=>"010100000",
  51739=>"110010010",
  51740=>"000100001",
  51741=>"011100110",
  51742=>"000101000",
  51743=>"010001111",
  51744=>"111000110",
  51745=>"111001010",
  51746=>"110000101",
  51747=>"111100100",
  51748=>"001101001",
  51749=>"011001111",
  51750=>"101011010",
  51751=>"001001001",
  51752=>"010111100",
  51753=>"000110100",
  51754=>"001011000",
  51755=>"111110011",
  51756=>"000000100",
  51757=>"100111100",
  51758=>"101000001",
  51759=>"101101110",
  51760=>"011001100",
  51761=>"110001101",
  51762=>"001010011",
  51763=>"001110101",
  51764=>"011101000",
  51765=>"100000011",
  51766=>"100011001",
  51767=>"011100111",
  51768=>"000111010",
  51769=>"111001110",
  51770=>"010000100",
  51771=>"010000010",
  51772=>"010010111",
  51773=>"011000001",
  51774=>"001001000",
  51775=>"111111010",
  51776=>"111000000",
  51777=>"100110011",
  51778=>"001111110",
  51779=>"110100000",
  51780=>"011101010",
  51781=>"111011101",
  51782=>"010100000",
  51783=>"011101110",
  51784=>"010001000",
  51785=>"001111000",
  51786=>"010110110",
  51787=>"100011010",
  51788=>"000111101",
  51789=>"010111111",
  51790=>"101011111",
  51791=>"010111000",
  51792=>"111000110",
  51793=>"011010111",
  51794=>"001111000",
  51795=>"100000111",
  51796=>"010111000",
  51797=>"100110011",
  51798=>"100110011",
  51799=>"011100010",
  51800=>"100001010",
  51801=>"101101110",
  51802=>"000100000",
  51803=>"110010001",
  51804=>"001100110",
  51805=>"000111110",
  51806=>"101110100",
  51807=>"000011101",
  51808=>"110011000",
  51809=>"111110111",
  51810=>"100110111",
  51811=>"001101000",
  51812=>"011111100",
  51813=>"110110100",
  51814=>"101111111",
  51815=>"000100110",
  51816=>"101011001",
  51817=>"111110111",
  51818=>"010111111",
  51819=>"111000011",
  51820=>"101011111",
  51821=>"000011001",
  51822=>"101101111",
  51823=>"101001001",
  51824=>"110101000",
  51825=>"011100010",
  51826=>"111110000",
  51827=>"001100111",
  51828=>"100001000",
  51829=>"110111001",
  51830=>"111111110",
  51831=>"010100011",
  51832=>"111101000",
  51833=>"111001001",
  51834=>"110001010",
  51835=>"001111011",
  51836=>"111100000",
  51837=>"111010010",
  51838=>"011001011",
  51839=>"100011010",
  51840=>"100011000",
  51841=>"110010010",
  51842=>"111001000",
  51843=>"010101110",
  51844=>"001100001",
  51845=>"010000111",
  51846=>"101000111",
  51847=>"100011111",
  51848=>"110010011",
  51849=>"010000011",
  51850=>"011010111",
  51851=>"010110001",
  51852=>"101000111",
  51853=>"111101010",
  51854=>"001000001",
  51855=>"101110011",
  51856=>"100000111",
  51857=>"110010101",
  51858=>"011010000",
  51859=>"010101001",
  51860=>"000111101",
  51861=>"101011010",
  51862=>"010001110",
  51863=>"010100010",
  51864=>"011011100",
  51865=>"000110100",
  51866=>"101101000",
  51867=>"100111111",
  51868=>"111000010",
  51869=>"010111111",
  51870=>"010001000",
  51871=>"011000111",
  51872=>"000010101",
  51873=>"010001010",
  51874=>"110100000",
  51875=>"100010101",
  51876=>"100001111",
  51877=>"110110101",
  51878=>"100000000",
  51879=>"010010000",
  51880=>"011100010",
  51881=>"100001111",
  51882=>"010010111",
  51883=>"001100001",
  51884=>"101100001",
  51885=>"001001010",
  51886=>"000000000",
  51887=>"111100000",
  51888=>"010010011",
  51889=>"100011011",
  51890=>"100011110",
  51891=>"111011011",
  51892=>"101011111",
  51893=>"001001101",
  51894=>"001100001",
  51895=>"011111011",
  51896=>"111111100",
  51897=>"010001111",
  51898=>"100101101",
  51899=>"110010101",
  51900=>"100111011",
  51901=>"111000001",
  51902=>"100011000",
  51903=>"001101101",
  51904=>"011100111",
  51905=>"100111100",
  51906=>"001000000",
  51907=>"011101100",
  51908=>"011111000",
  51909=>"110000001",
  51910=>"000110010",
  51911=>"000000001",
  51912=>"011001000",
  51913=>"110111100",
  51914=>"110000011",
  51915=>"011010001",
  51916=>"010011100",
  51917=>"001110010",
  51918=>"000111101",
  51919=>"001111011",
  51920=>"111001101",
  51921=>"101001101",
  51922=>"011010111",
  51923=>"111110111",
  51924=>"111011100",
  51925=>"000001001",
  51926=>"000010000",
  51927=>"110000001",
  51928=>"110101001",
  51929=>"111001111",
  51930=>"010001110",
  51931=>"110010110",
  51932=>"011011111",
  51933=>"111101000",
  51934=>"100110101",
  51935=>"001100111",
  51936=>"001000110",
  51937=>"001110111",
  51938=>"101001111",
  51939=>"000001111",
  51940=>"001101111",
  51941=>"100110101",
  51942=>"101111110",
  51943=>"100111000",
  51944=>"011100100",
  51945=>"000011100",
  51946=>"111111000",
  51947=>"110110111",
  51948=>"011011101",
  51949=>"111110100",
  51950=>"001000010",
  51951=>"011000110",
  51952=>"100010111",
  51953=>"000000010",
  51954=>"000110110",
  51955=>"011001011",
  51956=>"000011000",
  51957=>"101011101",
  51958=>"110000111",
  51959=>"110101001",
  51960=>"010111010",
  51961=>"001100001",
  51962=>"011101001",
  51963=>"000101010",
  51964=>"001100000",
  51965=>"101010000",
  51966=>"000011100",
  51967=>"101100110",
  51968=>"001110001",
  51969=>"000111000",
  51970=>"010001000",
  51971=>"000100010",
  51972=>"000001001",
  51973=>"111110011",
  51974=>"010010101",
  51975=>"111101001",
  51976=>"001111011",
  51977=>"100110100",
  51978=>"010100101",
  51979=>"011101111",
  51980=>"001100101",
  51981=>"011000101",
  51982=>"010001001",
  51983=>"010011110",
  51984=>"010110111",
  51985=>"001101101",
  51986=>"101100010",
  51987=>"110111010",
  51988=>"011110111",
  51989=>"001100101",
  51990=>"010100101",
  51991=>"001110001",
  51992=>"110011010",
  51993=>"100010111",
  51994=>"001110101",
  51995=>"110111001",
  51996=>"011000111",
  51997=>"010111100",
  51998=>"101001000",
  51999=>"000001111",
  52000=>"101110011",
  52001=>"100000010",
  52002=>"100000000",
  52003=>"001101000",
  52004=>"011000000",
  52005=>"001101110",
  52006=>"011011111",
  52007=>"001010001",
  52008=>"001000101",
  52009=>"111111001",
  52010=>"001011111",
  52011=>"001000011",
  52012=>"011101110",
  52013=>"000000000",
  52014=>"001011011",
  52015=>"010011111",
  52016=>"001010011",
  52017=>"111100111",
  52018=>"000010011",
  52019=>"101110111",
  52020=>"111110111",
  52021=>"100000101",
  52022=>"100111011",
  52023=>"101111111",
  52024=>"110010000",
  52025=>"111011111",
  52026=>"101101110",
  52027=>"001110100",
  52028=>"111100000",
  52029=>"011010110",
  52030=>"101011001",
  52031=>"101110111",
  52032=>"001011000",
  52033=>"101110001",
  52034=>"000011011",
  52035=>"110011010",
  52036=>"110000010",
  52037=>"011011001",
  52038=>"000111111",
  52039=>"010010110",
  52040=>"010010100",
  52041=>"111011100",
  52042=>"010010111",
  52043=>"000101101",
  52044=>"011100101",
  52045=>"011111101",
  52046=>"110100111",
  52047=>"110111000",
  52048=>"100000111",
  52049=>"001001111",
  52050=>"111000110",
  52051=>"000011110",
  52052=>"100111111",
  52053=>"000101111",
  52054=>"101111011",
  52055=>"110011000",
  52056=>"000000101",
  52057=>"110010101",
  52058=>"111011100",
  52059=>"011010100",
  52060=>"001111000",
  52061=>"100010111",
  52062=>"100101010",
  52063=>"101010011",
  52064=>"010100101",
  52065=>"111111111",
  52066=>"000111110",
  52067=>"111110001",
  52068=>"001000111",
  52069=>"110000001",
  52070=>"001000000",
  52071=>"000101111",
  52072=>"100010101",
  52073=>"000100110",
  52074=>"110101000",
  52075=>"111001111",
  52076=>"001100001",
  52077=>"010110010",
  52078=>"110110000",
  52079=>"011000101",
  52080=>"000100000",
  52081=>"001101010",
  52082=>"010110110",
  52083=>"110100011",
  52084=>"000111011",
  52085=>"111100011",
  52086=>"001001101",
  52087=>"100111101",
  52088=>"110000100",
  52089=>"100110111",
  52090=>"011110001",
  52091=>"100011101",
  52092=>"000100010",
  52093=>"000001000",
  52094=>"001110000",
  52095=>"110111111",
  52096=>"000110101",
  52097=>"101000101",
  52098=>"000010011",
  52099=>"001010010",
  52100=>"010100100",
  52101=>"101101111",
  52102=>"110011001",
  52103=>"000001001",
  52104=>"010110000",
  52105=>"100000001",
  52106=>"001010101",
  52107=>"111111111",
  52108=>"101100000",
  52109=>"011000001",
  52110=>"101100111",
  52111=>"100001011",
  52112=>"001011110",
  52113=>"011011010",
  52114=>"000000111",
  52115=>"010111101",
  52116=>"101100100",
  52117=>"000111110",
  52118=>"100011101",
  52119=>"001000100",
  52120=>"010001010",
  52121=>"000001010",
  52122=>"011110110",
  52123=>"110110001",
  52124=>"000100000",
  52125=>"011001010",
  52126=>"011000000",
  52127=>"010100111",
  52128=>"000000010",
  52129=>"010100001",
  52130=>"011111111",
  52131=>"010110001",
  52132=>"001100011",
  52133=>"010101111",
  52134=>"010011111",
  52135=>"001010110",
  52136=>"000100000",
  52137=>"110001011",
  52138=>"001101101",
  52139=>"100000101",
  52140=>"000100100",
  52141=>"100110111",
  52142=>"001100011",
  52143=>"101110100",
  52144=>"111010011",
  52145=>"100000001",
  52146=>"010111101",
  52147=>"011101011",
  52148=>"001011100",
  52149=>"001111110",
  52150=>"011011011",
  52151=>"011001111",
  52152=>"101100110",
  52153=>"111100000",
  52154=>"111111000",
  52155=>"111001000",
  52156=>"111111111",
  52157=>"111110110",
  52158=>"000010000",
  52159=>"111101100",
  52160=>"000101110",
  52161=>"010010000",
  52162=>"110111000",
  52163=>"100000101",
  52164=>"111100110",
  52165=>"001110101",
  52166=>"111111111",
  52167=>"010111011",
  52168=>"000010001",
  52169=>"001011000",
  52170=>"000001100",
  52171=>"110010000",
  52172=>"001110111",
  52173=>"000110011",
  52174=>"110001000",
  52175=>"111011010",
  52176=>"010001100",
  52177=>"100001101",
  52178=>"010111011",
  52179=>"011100000",
  52180=>"101000010",
  52181=>"111100011",
  52182=>"001111011",
  52183=>"110011011",
  52184=>"000100100",
  52185=>"101110101",
  52186=>"000110000",
  52187=>"000100000",
  52188=>"010011010",
  52189=>"010001111",
  52190=>"001010010",
  52191=>"111100011",
  52192=>"110011110",
  52193=>"000000111",
  52194=>"110000011",
  52195=>"010010011",
  52196=>"000001011",
  52197=>"111010100",
  52198=>"001111010",
  52199=>"100011010",
  52200=>"001011101",
  52201=>"110101111",
  52202=>"000111100",
  52203=>"110111101",
  52204=>"010110011",
  52205=>"000111000",
  52206=>"011000110",
  52207=>"000010110",
  52208=>"001100001",
  52209=>"010101001",
  52210=>"001100011",
  52211=>"111101010",
  52212=>"101001111",
  52213=>"010000101",
  52214=>"000001101",
  52215=>"111010010",
  52216=>"110100111",
  52217=>"000000101",
  52218=>"101111100",
  52219=>"101110100",
  52220=>"000100011",
  52221=>"010011111",
  52222=>"010011000",
  52223=>"101000010",
  52224=>"101100000",
  52225=>"101010101",
  52226=>"110011110",
  52227=>"011111001",
  52228=>"111110110",
  52229=>"010001000",
  52230=>"001010000",
  52231=>"001010001",
  52232=>"100110111",
  52233=>"101100001",
  52234=>"101000111",
  52235=>"101000110",
  52236=>"110000100",
  52237=>"011000111",
  52238=>"001100111",
  52239=>"100000111",
  52240=>"111110011",
  52241=>"101110111",
  52242=>"010111110",
  52243=>"011101011",
  52244=>"000110110",
  52245=>"001110001",
  52246=>"101101011",
  52247=>"111101000",
  52248=>"110001000",
  52249=>"110000111",
  52250=>"000100110",
  52251=>"010100110",
  52252=>"011001110",
  52253=>"001010101",
  52254=>"100001011",
  52255=>"111100111",
  52256=>"000000010",
  52257=>"100000000",
  52258=>"110101000",
  52259=>"111000110",
  52260=>"100100100",
  52261=>"111010000",
  52262=>"011000010",
  52263=>"110111001",
  52264=>"000111010",
  52265=>"100010001",
  52266=>"001110010",
  52267=>"111001111",
  52268=>"000101010",
  52269=>"111100100",
  52270=>"001011001",
  52271=>"111000111",
  52272=>"001111111",
  52273=>"101110101",
  52274=>"001011111",
  52275=>"000010000",
  52276=>"000011010",
  52277=>"000101100",
  52278=>"100010101",
  52279=>"000010100",
  52280=>"001100001",
  52281=>"100111100",
  52282=>"000111101",
  52283=>"001010000",
  52284=>"001001011",
  52285=>"010011101",
  52286=>"111110001",
  52287=>"000101010",
  52288=>"011011100",
  52289=>"000000010",
  52290=>"100111001",
  52291=>"101010011",
  52292=>"110011000",
  52293=>"111010101",
  52294=>"100100011",
  52295=>"000001110",
  52296=>"001011100",
  52297=>"001000000",
  52298=>"101100011",
  52299=>"101011011",
  52300=>"101110101",
  52301=>"111000000",
  52302=>"101001011",
  52303=>"110001100",
  52304=>"000100001",
  52305=>"010011000",
  52306=>"000110111",
  52307=>"110010100",
  52308=>"111111000",
  52309=>"011100111",
  52310=>"111000001",
  52311=>"100001001",
  52312=>"111110010",
  52313=>"011100011",
  52314=>"100011111",
  52315=>"011110011",
  52316=>"111000111",
  52317=>"000100010",
  52318=>"100000001",
  52319=>"000011111",
  52320=>"000111001",
  52321=>"111101110",
  52322=>"110000000",
  52323=>"010001011",
  52324=>"011100011",
  52325=>"000011001",
  52326=>"111001101",
  52327=>"001101111",
  52328=>"010101101",
  52329=>"010100110",
  52330=>"111100011",
  52331=>"000110000",
  52332=>"011000101",
  52333=>"000110000",
  52334=>"010011000",
  52335=>"010100001",
  52336=>"010100011",
  52337=>"000011010",
  52338=>"001111011",
  52339=>"110111111",
  52340=>"101101100",
  52341=>"010100110",
  52342=>"110110100",
  52343=>"100100010",
  52344=>"011101001",
  52345=>"110011100",
  52346=>"001011000",
  52347=>"111001111",
  52348=>"101001111",
  52349=>"111111101",
  52350=>"110100111",
  52351=>"000000000",
  52352=>"001100101",
  52353=>"101001100",
  52354=>"111010010",
  52355=>"101001101",
  52356=>"010100111",
  52357=>"001001011",
  52358=>"010101000",
  52359=>"110010001",
  52360=>"100001010",
  52361=>"010000011",
  52362=>"100101010",
  52363=>"001111001",
  52364=>"101011101",
  52365=>"000101110",
  52366=>"100110111",
  52367=>"110110011",
  52368=>"100000111",
  52369=>"010101110",
  52370=>"101111011",
  52371=>"001010001",
  52372=>"010111010",
  52373=>"100000000",
  52374=>"001101010",
  52375=>"100010010",
  52376=>"101110111",
  52377=>"001000111",
  52378=>"100001110",
  52379=>"000110000",
  52380=>"100000000",
  52381=>"000111011",
  52382=>"111001000",
  52383=>"101101101",
  52384=>"001011101",
  52385=>"100100001",
  52386=>"110001101",
  52387=>"110000001",
  52388=>"100101011",
  52389=>"010111111",
  52390=>"010000010",
  52391=>"111000100",
  52392=>"001001000",
  52393=>"100111110",
  52394=>"111000111",
  52395=>"100010010",
  52396=>"111111000",
  52397=>"001001100",
  52398=>"001000001",
  52399=>"001101010",
  52400=>"001000000",
  52401=>"101101000",
  52402=>"100110100",
  52403=>"011101001",
  52404=>"110000001",
  52405=>"000010010",
  52406=>"111111011",
  52407=>"010111010",
  52408=>"000000000",
  52409=>"110001101",
  52410=>"100000111",
  52411=>"111100110",
  52412=>"110111011",
  52413=>"011100011",
  52414=>"010010011",
  52415=>"001011110",
  52416=>"111110010",
  52417=>"010001100",
  52418=>"010101010",
  52419=>"010000111",
  52420=>"101111000",
  52421=>"100100111",
  52422=>"000111110",
  52423=>"101101000",
  52424=>"001011100",
  52425=>"010101010",
  52426=>"101110110",
  52427=>"100000010",
  52428=>"101011001",
  52429=>"110101100",
  52430=>"010000111",
  52431=>"111000111",
  52432=>"010101110",
  52433=>"000101110",
  52434=>"001100000",
  52435=>"111000110",
  52436=>"010000110",
  52437=>"111111111",
  52438=>"010011010",
  52439=>"111101011",
  52440=>"101000110",
  52441=>"111101000",
  52442=>"010001011",
  52443=>"001101101",
  52444=>"011100010",
  52445=>"100101001",
  52446=>"111101011",
  52447=>"000111110",
  52448=>"010101100",
  52449=>"000111001",
  52450=>"000001001",
  52451=>"000000100",
  52452=>"000010001",
  52453=>"001010111",
  52454=>"001001110",
  52455=>"101100010",
  52456=>"100000011",
  52457=>"101011110",
  52458=>"111100001",
  52459=>"110110101",
  52460=>"011011100",
  52461=>"100011110",
  52462=>"011000110",
  52463=>"010110001",
  52464=>"110010010",
  52465=>"011011000",
  52466=>"100000100",
  52467=>"110110111",
  52468=>"001101110",
  52469=>"011100011",
  52470=>"101101111",
  52471=>"010000111",
  52472=>"000101100",
  52473=>"110010011",
  52474=>"111011111",
  52475=>"110100100",
  52476=>"010111111",
  52477=>"010011001",
  52478=>"010100010",
  52479=>"001011111",
  52480=>"111011100",
  52481=>"111010101",
  52482=>"111011011",
  52483=>"010001111",
  52484=>"000110101",
  52485=>"111110001",
  52486=>"001011011",
  52487=>"011101101",
  52488=>"111011000",
  52489=>"100110110",
  52490=>"001011101",
  52491=>"111001010",
  52492=>"000010111",
  52493=>"101000111",
  52494=>"001011110",
  52495=>"010110010",
  52496=>"001000001",
  52497=>"000101101",
  52498=>"111111100",
  52499=>"011011001",
  52500=>"001100001",
  52501=>"010100110",
  52502=>"000000011",
  52503=>"000000001",
  52504=>"000101000",
  52505=>"001100001",
  52506=>"001001000",
  52507=>"100110101",
  52508=>"100110011",
  52509=>"111100000",
  52510=>"011011100",
  52511=>"001110100",
  52512=>"110010001",
  52513=>"110101011",
  52514=>"001111001",
  52515=>"011000110",
  52516=>"100010000",
  52517=>"011100111",
  52518=>"111010100",
  52519=>"100010101",
  52520=>"110000110",
  52521=>"011001000",
  52522=>"101110000",
  52523=>"000011101",
  52524=>"011000001",
  52525=>"010100000",
  52526=>"000000100",
  52527=>"111001011",
  52528=>"100101110",
  52529=>"010101001",
  52530=>"011111100",
  52531=>"001001110",
  52532=>"000011100",
  52533=>"110010011",
  52534=>"111100011",
  52535=>"000001010",
  52536=>"000000000",
  52537=>"010001001",
  52538=>"010110111",
  52539=>"101111110",
  52540=>"010000101",
  52541=>"110101111",
  52542=>"010001110",
  52543=>"010100101",
  52544=>"111000110",
  52545=>"110010111",
  52546=>"101010010",
  52547=>"110110100",
  52548=>"000111111",
  52549=>"111100011",
  52550=>"001111100",
  52551=>"001101000",
  52552=>"000101010",
  52553=>"000000111",
  52554=>"010100010",
  52555=>"001001100",
  52556=>"011101010",
  52557=>"000010010",
  52558=>"010100010",
  52559=>"001010010",
  52560=>"011011110",
  52561=>"101001001",
  52562=>"001101110",
  52563=>"100001011",
  52564=>"111101101",
  52565=>"000111111",
  52566=>"001101101",
  52567=>"011000101",
  52568=>"111110011",
  52569=>"000101111",
  52570=>"100111010",
  52571=>"110101100",
  52572=>"000000100",
  52573=>"010000010",
  52574=>"001011011",
  52575=>"000111100",
  52576=>"000110111",
  52577=>"011011000",
  52578=>"100000011",
  52579=>"000010001",
  52580=>"100010000",
  52581=>"100000001",
  52582=>"111011000",
  52583=>"011100011",
  52584=>"010010001",
  52585=>"000010000",
  52586=>"010111010",
  52587=>"000111111",
  52588=>"111000110",
  52589=>"101111101",
  52590=>"111001010",
  52591=>"001001110",
  52592=>"100000111",
  52593=>"010010011",
  52594=>"000111010",
  52595=>"111000010",
  52596=>"000010101",
  52597=>"111010101",
  52598=>"011111111",
  52599=>"011011000",
  52600=>"111000011",
  52601=>"000011000",
  52602=>"111110000",
  52603=>"000111000",
  52604=>"101110101",
  52605=>"101100110",
  52606=>"100001010",
  52607=>"001100010",
  52608=>"111111111",
  52609=>"101111011",
  52610=>"101010001",
  52611=>"011111101",
  52612=>"001100001",
  52613=>"101110101",
  52614=>"000110011",
  52615=>"111000010",
  52616=>"001001101",
  52617=>"011000111",
  52618=>"101010000",
  52619=>"100001001",
  52620=>"000011111",
  52621=>"001111011",
  52622=>"001110100",
  52623=>"011011011",
  52624=>"010011110",
  52625=>"011000000",
  52626=>"010111001",
  52627=>"001111111",
  52628=>"000010000",
  52629=>"001000100",
  52630=>"100000101",
  52631=>"010110000",
  52632=>"000010100",
  52633=>"000010000",
  52634=>"110001101",
  52635=>"000001111",
  52636=>"010011110",
  52637=>"101110101",
  52638=>"111111100",
  52639=>"111001111",
  52640=>"001010010",
  52641=>"000000000",
  52642=>"000010000",
  52643=>"011000010",
  52644=>"111110110",
  52645=>"010000100",
  52646=>"011011001",
  52647=>"000000010",
  52648=>"010110000",
  52649=>"100001111",
  52650=>"000011000",
  52651=>"101110000",
  52652=>"000000100",
  52653=>"101010111",
  52654=>"000011011",
  52655=>"111010100",
  52656=>"110001100",
  52657=>"010100010",
  52658=>"011011011",
  52659=>"011110101",
  52660=>"010000110",
  52661=>"110101111",
  52662=>"010000110",
  52663=>"110000010",
  52664=>"000100110",
  52665=>"111101101",
  52666=>"000010110",
  52667=>"111010010",
  52668=>"100101101",
  52669=>"010010101",
  52670=>"111010110",
  52671=>"011111111",
  52672=>"000010001",
  52673=>"100111111",
  52674=>"101001111",
  52675=>"010100011",
  52676=>"000000001",
  52677=>"011010011",
  52678=>"011110110",
  52679=>"000001101",
  52680=>"011011001",
  52681=>"011010110",
  52682=>"010010000",
  52683=>"110111111",
  52684=>"111001101",
  52685=>"000001111",
  52686=>"111011010",
  52687=>"101001000",
  52688=>"111100101",
  52689=>"010000010",
  52690=>"011010000",
  52691=>"111010110",
  52692=>"000110101",
  52693=>"000010110",
  52694=>"011111110",
  52695=>"001100000",
  52696=>"101100000",
  52697=>"101001100",
  52698=>"011000010",
  52699=>"100101100",
  52700=>"110001110",
  52701=>"110010101",
  52702=>"000000101",
  52703=>"011111110",
  52704=>"111100000",
  52705=>"111111000",
  52706=>"110011010",
  52707=>"110101100",
  52708=>"111110110",
  52709=>"010010111",
  52710=>"001100000",
  52711=>"101000000",
  52712=>"000010110",
  52713=>"101111110",
  52714=>"010010111",
  52715=>"001110001",
  52716=>"011010110",
  52717=>"101110011",
  52718=>"011001000",
  52719=>"000000010",
  52720=>"101001110",
  52721=>"000010110",
  52722=>"001100001",
  52723=>"111100100",
  52724=>"000100011",
  52725=>"001111110",
  52726=>"110110000",
  52727=>"001000111",
  52728=>"001101101",
  52729=>"110110001",
  52730=>"001101111",
  52731=>"101111001",
  52732=>"100111100",
  52733=>"110001011",
  52734=>"101000101",
  52735=>"001001010",
  52736=>"001100010",
  52737=>"110110001",
  52738=>"100100011",
  52739=>"101001111",
  52740=>"011111000",
  52741=>"010100101",
  52742=>"011011010",
  52743=>"001011101",
  52744=>"011011010",
  52745=>"111000001",
  52746=>"011000011",
  52747=>"000111110",
  52748=>"000100110",
  52749=>"101101101",
  52750=>"110000101",
  52751=>"011000100",
  52752=>"100110010",
  52753=>"010111101",
  52754=>"010000101",
  52755=>"000110111",
  52756=>"100000111",
  52757=>"011111000",
  52758=>"001001011",
  52759=>"100101000",
  52760=>"010101111",
  52761=>"011101110",
  52762=>"101000100",
  52763=>"001000100",
  52764=>"000010001",
  52765=>"000011000",
  52766=>"101111001",
  52767=>"110000011",
  52768=>"110111001",
  52769=>"101011001",
  52770=>"001101110",
  52771=>"011001101",
  52772=>"001101111",
  52773=>"111000011",
  52774=>"110010100",
  52775=>"111011010",
  52776=>"011100110",
  52777=>"110000101",
  52778=>"101001111",
  52779=>"001000101",
  52780=>"110001010",
  52781=>"000001010",
  52782=>"001111010",
  52783=>"010000010",
  52784=>"000010101",
  52785=>"111110111",
  52786=>"101110001",
  52787=>"000110000",
  52788=>"001000000",
  52789=>"010110110",
  52790=>"000111011",
  52791=>"110010101",
  52792=>"001111110",
  52793=>"000100101",
  52794=>"000000111",
  52795=>"000110101",
  52796=>"110001010",
  52797=>"010111000",
  52798=>"011000010",
  52799=>"110110010",
  52800=>"111111010",
  52801=>"100011010",
  52802=>"000011100",
  52803=>"001000100",
  52804=>"000100111",
  52805=>"111101111",
  52806=>"010101000",
  52807=>"100100000",
  52808=>"111010101",
  52809=>"110100110",
  52810=>"101111111",
  52811=>"101001010",
  52812=>"010101011",
  52813=>"011101001",
  52814=>"011111100",
  52815=>"101110000",
  52816=>"000011100",
  52817=>"100110000",
  52818=>"000010101",
  52819=>"111000001",
  52820=>"001100010",
  52821=>"001001001",
  52822=>"111111011",
  52823=>"100110111",
  52824=>"110100110",
  52825=>"000000010",
  52826=>"001100010",
  52827=>"001101001",
  52828=>"001100100",
  52829=>"000001000",
  52830=>"101110110",
  52831=>"100001111",
  52832=>"110001100",
  52833=>"011100000",
  52834=>"110100101",
  52835=>"000000000",
  52836=>"011011001",
  52837=>"110011100",
  52838=>"101011011",
  52839=>"001101111",
  52840=>"000110101",
  52841=>"110101011",
  52842=>"111001000",
  52843=>"010110110",
  52844=>"100101110",
  52845=>"100010101",
  52846=>"011100101",
  52847=>"000011100",
  52848=>"000100100",
  52849=>"100110100",
  52850=>"010001101",
  52851=>"000110101",
  52852=>"001010100",
  52853=>"101001111",
  52854=>"001001000",
  52855=>"011101000",
  52856=>"111010101",
  52857=>"101010010",
  52858=>"001000100",
  52859=>"111000011",
  52860=>"011001011",
  52861=>"100101010",
  52862=>"010100011",
  52863=>"100010010",
  52864=>"001111010",
  52865=>"010101010",
  52866=>"111000111",
  52867=>"110101011",
  52868=>"000000100",
  52869=>"000001001",
  52870=>"010100000",
  52871=>"010101001",
  52872=>"001110000",
  52873=>"000101000",
  52874=>"111101011",
  52875=>"000010010",
  52876=>"001101000",
  52877=>"111000100",
  52878=>"000111100",
  52879=>"010000101",
  52880=>"100001100",
  52881=>"000111001",
  52882=>"101001111",
  52883=>"001010010",
  52884=>"001010001",
  52885=>"100000001",
  52886=>"001100101",
  52887=>"001000001",
  52888=>"010011111",
  52889=>"010000100",
  52890=>"110111100",
  52891=>"101111111",
  52892=>"010101101",
  52893=>"011001101",
  52894=>"111010001",
  52895=>"110000101",
  52896=>"001000001",
  52897=>"000101101",
  52898=>"011101111",
  52899=>"001110100",
  52900=>"101100110",
  52901=>"111111000",
  52902=>"101100111",
  52903=>"101100101",
  52904=>"100011100",
  52905=>"111101110",
  52906=>"110100111",
  52907=>"011111111",
  52908=>"000111000",
  52909=>"000001011",
  52910=>"111000001",
  52911=>"100011100",
  52912=>"000010110",
  52913=>"100100001",
  52914=>"111000110",
  52915=>"001001110",
  52916=>"110010010",
  52917=>"111100111",
  52918=>"100100111",
  52919=>"001110101",
  52920=>"110011100",
  52921=>"010100001",
  52922=>"110010100",
  52923=>"000110101",
  52924=>"111100001",
  52925=>"001110100",
  52926=>"000011101",
  52927=>"101111111",
  52928=>"101110001",
  52929=>"001001011",
  52930=>"010110111",
  52931=>"110111010",
  52932=>"010011100",
  52933=>"110011111",
  52934=>"000111001",
  52935=>"100010111",
  52936=>"110011101",
  52937=>"001000010",
  52938=>"010101111",
  52939=>"001101110",
  52940=>"010000101",
  52941=>"110110001",
  52942=>"000000100",
  52943=>"010110011",
  52944=>"101000001",
  52945=>"010000101",
  52946=>"100011101",
  52947=>"011010001",
  52948=>"110011010",
  52949=>"110100010",
  52950=>"101100100",
  52951=>"000011001",
  52952=>"000000101",
  52953=>"000100011",
  52954=>"101110000",
  52955=>"111100011",
  52956=>"011001011",
  52957=>"111100000",
  52958=>"100000111",
  52959=>"011100001",
  52960=>"100100111",
  52961=>"010000111",
  52962=>"011010101",
  52963=>"101000001",
  52964=>"001100110",
  52965=>"110111011",
  52966=>"110001010",
  52967=>"110100111",
  52968=>"100001011",
  52969=>"000111010",
  52970=>"100100010",
  52971=>"100101000",
  52972=>"100000101",
  52973=>"101100000",
  52974=>"011101000",
  52975=>"000001101",
  52976=>"110110011",
  52977=>"111101010",
  52978=>"000100011",
  52979=>"101111110",
  52980=>"000011001",
  52981=>"101111100",
  52982=>"001011111",
  52983=>"111111100",
  52984=>"100010011",
  52985=>"001010100",
  52986=>"111100010",
  52987=>"000000000",
  52988=>"110111010",
  52989=>"011110011",
  52990=>"101100100",
  52991=>"011111001",
  52992=>"110000010",
  52993=>"101001110",
  52994=>"010101111",
  52995=>"001000101",
  52996=>"011000100",
  52997=>"101111111",
  52998=>"001011100",
  52999=>"001100100",
  53000=>"011100101",
  53001=>"011001111",
  53002=>"101101001",
  53003=>"110101100",
  53004=>"110000111",
  53005=>"111000001",
  53006=>"110101100",
  53007=>"110010111",
  53008=>"110010011",
  53009=>"000001011",
  53010=>"110000101",
  53011=>"001111011",
  53012=>"101111111",
  53013=>"011011011",
  53014=>"001011000",
  53015=>"000000011",
  53016=>"110101100",
  53017=>"100111000",
  53018=>"100010100",
  53019=>"011001011",
  53020=>"100100110",
  53021=>"011011111",
  53022=>"010010000",
  53023=>"111100100",
  53024=>"001111101",
  53025=>"000000000",
  53026=>"010110000",
  53027=>"001110101",
  53028=>"000010100",
  53029=>"000011000",
  53030=>"011111000",
  53031=>"111010001",
  53032=>"101010000",
  53033=>"111000011",
  53034=>"100011101",
  53035=>"110111111",
  53036=>"110110110",
  53037=>"111010110",
  53038=>"000000111",
  53039=>"000001100",
  53040=>"000101100",
  53041=>"100011100",
  53042=>"110101101",
  53043=>"110001000",
  53044=>"111011010",
  53045=>"011011101",
  53046=>"100111010",
  53047=>"111011111",
  53048=>"001100111",
  53049=>"101100111",
  53050=>"111011010",
  53051=>"110100001",
  53052=>"100010100",
  53053=>"101011010",
  53054=>"111011000",
  53055=>"110101110",
  53056=>"000111000",
  53057=>"100011011",
  53058=>"110101110",
  53059=>"000000101",
  53060=>"111111111",
  53061=>"110000111",
  53062=>"000111000",
  53063=>"101110101",
  53064=>"111000111",
  53065=>"100111001",
  53066=>"111001000",
  53067=>"110000011",
  53068=>"101000111",
  53069=>"011011110",
  53070=>"110000111",
  53071=>"000011111",
  53072=>"101010010",
  53073=>"010001111",
  53074=>"111011110",
  53075=>"010011011",
  53076=>"101000010",
  53077=>"101000110",
  53078=>"000111101",
  53079=>"000101100",
  53080=>"001010101",
  53081=>"001011010",
  53082=>"010011111",
  53083=>"010010000",
  53084=>"101101010",
  53085=>"111101001",
  53086=>"111100101",
  53087=>"101010100",
  53088=>"111011010",
  53089=>"111011001",
  53090=>"000010000",
  53091=>"001111101",
  53092=>"000110001",
  53093=>"100110111",
  53094=>"001000011",
  53095=>"101010110",
  53096=>"010010000",
  53097=>"000000011",
  53098=>"010011011",
  53099=>"001001101",
  53100=>"010110000",
  53101=>"100000000",
  53102=>"111011010",
  53103=>"101010010",
  53104=>"100111110",
  53105=>"001000101",
  53106=>"000001010",
  53107=>"100100110",
  53108=>"011111011",
  53109=>"010001110",
  53110=>"110001010",
  53111=>"100111001",
  53112=>"011000101",
  53113=>"010010010",
  53114=>"001000000",
  53115=>"011001111",
  53116=>"000100011",
  53117=>"001100011",
  53118=>"101111110",
  53119=>"011101010",
  53120=>"001000001",
  53121=>"000100001",
  53122=>"010001011",
  53123=>"011000011",
  53124=>"111110110",
  53125=>"110000100",
  53126=>"111111100",
  53127=>"101000001",
  53128=>"100110010",
  53129=>"101110100",
  53130=>"110101110",
  53131=>"010000100",
  53132=>"001101011",
  53133=>"010011001",
  53134=>"000010101",
  53135=>"011110000",
  53136=>"010111000",
  53137=>"110011000",
  53138=>"001000101",
  53139=>"100001001",
  53140=>"000000011",
  53141=>"100001100",
  53142=>"011111010",
  53143=>"110101001",
  53144=>"001101100",
  53145=>"100010101",
  53146=>"100110001",
  53147=>"101100100",
  53148=>"001110101",
  53149=>"101010111",
  53150=>"001110111",
  53151=>"001101011",
  53152=>"100000010",
  53153=>"110010010",
  53154=>"001101100",
  53155=>"001000000",
  53156=>"110011001",
  53157=>"000010011",
  53158=>"101100100",
  53159=>"100011000",
  53160=>"001001111",
  53161=>"101001001",
  53162=>"010011011",
  53163=>"111111111",
  53164=>"110000111",
  53165=>"110000100",
  53166=>"000111010",
  53167=>"100101000",
  53168=>"001111110",
  53169=>"001011011",
  53170=>"000111110",
  53171=>"101110100",
  53172=>"111011000",
  53173=>"110010100",
  53174=>"101110001",
  53175=>"101011100",
  53176=>"100000001",
  53177=>"110100111",
  53178=>"010011110",
  53179=>"010101001",
  53180=>"000001000",
  53181=>"101110110",
  53182=>"011000111",
  53183=>"011001011",
  53184=>"000011111",
  53185=>"010010001",
  53186=>"101001000",
  53187=>"111110100",
  53188=>"101100010",
  53189=>"001011110",
  53190=>"101101100",
  53191=>"100111111",
  53192=>"111001100",
  53193=>"000111011",
  53194=>"100000110",
  53195=>"011011111",
  53196=>"101110110",
  53197=>"110111010",
  53198=>"010001010",
  53199=>"101011011",
  53200=>"001101010",
  53201=>"010010110",
  53202=>"011011101",
  53203=>"111111011",
  53204=>"000111010",
  53205=>"000000001",
  53206=>"101110011",
  53207=>"010100001",
  53208=>"010111000",
  53209=>"000010000",
  53210=>"001001000",
  53211=>"101111000",
  53212=>"110000001",
  53213=>"100110110",
  53214=>"101111110",
  53215=>"001100100",
  53216=>"110010001",
  53217=>"101001101",
  53218=>"010011010",
  53219=>"001111001",
  53220=>"000000000",
  53221=>"011001000",
  53222=>"010101110",
  53223=>"100011000",
  53224=>"000110010",
  53225=>"100011001",
  53226=>"111010010",
  53227=>"010001101",
  53228=>"100001001",
  53229=>"110101000",
  53230=>"010100010",
  53231=>"000111010",
  53232=>"011011010",
  53233=>"011111101",
  53234=>"000001000",
  53235=>"000110001",
  53236=>"010000101",
  53237=>"011100001",
  53238=>"011101111",
  53239=>"101001101",
  53240=>"111101111",
  53241=>"100011100",
  53242=>"100000011",
  53243=>"101001001",
  53244=>"111101111",
  53245=>"111110101",
  53246=>"000101100",
  53247=>"110110101",
  53248=>"111101000",
  53249=>"111011111",
  53250=>"100110011",
  53251=>"000000100",
  53252=>"111011100",
  53253=>"110100100",
  53254=>"100010111",
  53255=>"011101000",
  53256=>"001110101",
  53257=>"001110100",
  53258=>"100001000",
  53259=>"001101010",
  53260=>"111111001",
  53261=>"101000011",
  53262=>"000010010",
  53263=>"100011110",
  53264=>"011110110",
  53265=>"000000110",
  53266=>"111011111",
  53267=>"100010011",
  53268=>"001111111",
  53269=>"001010010",
  53270=>"100000100",
  53271=>"011000111",
  53272=>"110110000",
  53273=>"100100110",
  53274=>"010010110",
  53275=>"111001110",
  53276=>"110001011",
  53277=>"000100000",
  53278=>"001011001",
  53279=>"111011111",
  53280=>"010101001",
  53281=>"000110110",
  53282=>"010111111",
  53283=>"001111010",
  53284=>"110111000",
  53285=>"000000101",
  53286=>"010110101",
  53287=>"100110111",
  53288=>"001111111",
  53289=>"001110000",
  53290=>"101011111",
  53291=>"011001011",
  53292=>"101110001",
  53293=>"010110000",
  53294=>"000001101",
  53295=>"100001010",
  53296=>"011000110",
  53297=>"100000111",
  53298=>"011001011",
  53299=>"011100000",
  53300=>"111111000",
  53301=>"100111000",
  53302=>"101001011",
  53303=>"000011011",
  53304=>"001101110",
  53305=>"001111010",
  53306=>"111110100",
  53307=>"100000110",
  53308=>"010100110",
  53309=>"110110110",
  53310=>"011000000",
  53311=>"000010000",
  53312=>"011000010",
  53313=>"010101100",
  53314=>"111010111",
  53315=>"010000110",
  53316=>"110010111",
  53317=>"001100001",
  53318=>"111110001",
  53319=>"000010010",
  53320=>"111001110",
  53321=>"100110000",
  53322=>"100010111",
  53323=>"001010000",
  53324=>"110110001",
  53325=>"010000110",
  53326=>"000111110",
  53327=>"110010010",
  53328=>"010000100",
  53329=>"101000001",
  53330=>"011111010",
  53331=>"000001110",
  53332=>"101001001",
  53333=>"001000001",
  53334=>"111011000",
  53335=>"000001111",
  53336=>"000001100",
  53337=>"011110011",
  53338=>"101110110",
  53339=>"111000100",
  53340=>"011001000",
  53341=>"001010101",
  53342=>"011011010",
  53343=>"000000101",
  53344=>"001110110",
  53345=>"110011100",
  53346=>"101010100",
  53347=>"001010001",
  53348=>"011001001",
  53349=>"000100100",
  53350=>"000111101",
  53351=>"010110001",
  53352=>"100111110",
  53353=>"010100101",
  53354=>"010011011",
  53355=>"111010111",
  53356=>"001001100",
  53357=>"111001001",
  53358=>"110000001",
  53359=>"111100010",
  53360=>"111001101",
  53361=>"011111011",
  53362=>"100010000",
  53363=>"001111010",
  53364=>"000010000",
  53365=>"010101010",
  53366=>"010000001",
  53367=>"000000111",
  53368=>"100101100",
  53369=>"100110000",
  53370=>"111111111",
  53371=>"100100111",
  53372=>"011101001",
  53373=>"010111101",
  53374=>"101000110",
  53375=>"010110011",
  53376=>"011001010",
  53377=>"010010001",
  53378=>"010111101",
  53379=>"101011011",
  53380=>"110111011",
  53381=>"000010101",
  53382=>"100111000",
  53383=>"010100001",
  53384=>"100011111",
  53385=>"101100110",
  53386=>"111001001",
  53387=>"000000011",
  53388=>"001100110",
  53389=>"111101010",
  53390=>"100111110",
  53391=>"100000010",
  53392=>"010101000",
  53393=>"101100001",
  53394=>"010101101",
  53395=>"011110110",
  53396=>"110100100",
  53397=>"111101001",
  53398=>"011111001",
  53399=>"110000101",
  53400=>"001001111",
  53401=>"101000100",
  53402=>"110000011",
  53403=>"111010110",
  53404=>"010000111",
  53405=>"001101001",
  53406=>"111001000",
  53407=>"000001101",
  53408=>"110111111",
  53409=>"010111001",
  53410=>"000100011",
  53411=>"100101111",
  53412=>"001110110",
  53413=>"100100100",
  53414=>"101100110",
  53415=>"111100110",
  53416=>"011011100",
  53417=>"110111000",
  53418=>"100111100",
  53419=>"001001010",
  53420=>"111000000",
  53421=>"111001100",
  53422=>"101101111",
  53423=>"110010011",
  53424=>"001100001",
  53425=>"111101110",
  53426=>"011101110",
  53427=>"011001011",
  53428=>"110011000",
  53429=>"110110110",
  53430=>"010101000",
  53431=>"101111001",
  53432=>"100100000",
  53433=>"000000011",
  53434=>"001000001",
  53435=>"010110110",
  53436=>"100011110",
  53437=>"101000010",
  53438=>"011001011",
  53439=>"101100001",
  53440=>"011010001",
  53441=>"100010100",
  53442=>"010010001",
  53443=>"010010000",
  53444=>"001111010",
  53445=>"000000011",
  53446=>"111001100",
  53447=>"001011011",
  53448=>"110000000",
  53449=>"111011001",
  53450=>"111101101",
  53451=>"011100011",
  53452=>"010111010",
  53453=>"000010011",
  53454=>"001000010",
  53455=>"001011110",
  53456=>"110010111",
  53457=>"001100110",
  53458=>"010001110",
  53459=>"100100100",
  53460=>"110100110",
  53461=>"110111100",
  53462=>"011000100",
  53463=>"011101101",
  53464=>"101000000",
  53465=>"010010101",
  53466=>"001000110",
  53467=>"110000110",
  53468=>"101000000",
  53469=>"001101011",
  53470=>"101110011",
  53471=>"011011111",
  53472=>"011001101",
  53473=>"010111010",
  53474=>"101110011",
  53475=>"110110000",
  53476=>"101010110",
  53477=>"100010101",
  53478=>"100100100",
  53479=>"000110011",
  53480=>"001001010",
  53481=>"000001111",
  53482=>"011011001",
  53483=>"110001111",
  53484=>"110111011",
  53485=>"111010110",
  53486=>"101011011",
  53487=>"010001000",
  53488=>"100111000",
  53489=>"101110001",
  53490=>"011000101",
  53491=>"110010000",
  53492=>"110010010",
  53493=>"010100111",
  53494=>"001001000",
  53495=>"100100000",
  53496=>"000100100",
  53497=>"111001001",
  53498=>"011110100",
  53499=>"001011000",
  53500=>"111101111",
  53501=>"110110101",
  53502=>"000111011",
  53503=>"000100011",
  53504=>"110110010",
  53505=>"011011001",
  53506=>"010101011",
  53507=>"001000100",
  53508=>"101111110",
  53509=>"010110000",
  53510=>"010000000",
  53511=>"101111111",
  53512=>"000101001",
  53513=>"001010011",
  53514=>"100100000",
  53515=>"101000101",
  53516=>"000000010",
  53517=>"101000111",
  53518=>"011111010",
  53519=>"000001000",
  53520=>"001000010",
  53521=>"010111100",
  53522=>"101110011",
  53523=>"111011011",
  53524=>"010100100",
  53525=>"010000010",
  53526=>"101010010",
  53527=>"010000111",
  53528=>"011010010",
  53529=>"010010001",
  53530=>"111011110",
  53531=>"011111100",
  53532=>"001101111",
  53533=>"111111100",
  53534=>"011010010",
  53535=>"101011001",
  53536=>"100100010",
  53537=>"001001010",
  53538=>"100001001",
  53539=>"010110001",
  53540=>"111010000",
  53541=>"100000100",
  53542=>"111010110",
  53543=>"011100100",
  53544=>"110000010",
  53545=>"101010111",
  53546=>"000100001",
  53547=>"110111010",
  53548=>"111011110",
  53549=>"110100010",
  53550=>"010000001",
  53551=>"000010001",
  53552=>"111011100",
  53553=>"111100100",
  53554=>"101000101",
  53555=>"011111010",
  53556=>"100110100",
  53557=>"100000011",
  53558=>"010010010",
  53559=>"101111011",
  53560=>"000011100",
  53561=>"001101001",
  53562=>"101111111",
  53563=>"101011101",
  53564=>"011011010",
  53565=>"101001101",
  53566=>"110101100",
  53567=>"011100100",
  53568=>"110100111",
  53569=>"011001101",
  53570=>"111101101",
  53571=>"010000011",
  53572=>"011101010",
  53573=>"010100010",
  53574=>"011101011",
  53575=>"000110000",
  53576=>"111011101",
  53577=>"110010100",
  53578=>"000011100",
  53579=>"101000111",
  53580=>"010110001",
  53581=>"011100001",
  53582=>"111111010",
  53583=>"000010010",
  53584=>"100111010",
  53585=>"001001100",
  53586=>"101110011",
  53587=>"001010000",
  53588=>"011111001",
  53589=>"011010001",
  53590=>"111100110",
  53591=>"101011000",
  53592=>"100010010",
  53593=>"001010001",
  53594=>"010100011",
  53595=>"111001111",
  53596=>"000010100",
  53597=>"000111100",
  53598=>"010111010",
  53599=>"010011100",
  53600=>"100111010",
  53601=>"011010001",
  53602=>"111110000",
  53603=>"100001100",
  53604=>"011011101",
  53605=>"011101100",
  53606=>"110010110",
  53607=>"111110100",
  53608=>"100000001",
  53609=>"000000111",
  53610=>"111110101",
  53611=>"011011010",
  53612=>"110111110",
  53613=>"000111110",
  53614=>"111100000",
  53615=>"001001010",
  53616=>"110010000",
  53617=>"001000100",
  53618=>"010011001",
  53619=>"100100101",
  53620=>"111111101",
  53621=>"110010000",
  53622=>"010001111",
  53623=>"100101011",
  53624=>"001001001",
  53625=>"111010000",
  53626=>"110110100",
  53627=>"100111011",
  53628=>"100101001",
  53629=>"001101110",
  53630=>"110011100",
  53631=>"010001011",
  53632=>"001011000",
  53633=>"110111010",
  53634=>"101000001",
  53635=>"000010110",
  53636=>"100110111",
  53637=>"111011111",
  53638=>"100111011",
  53639=>"101110010",
  53640=>"011101000",
  53641=>"000010011",
  53642=>"010101001",
  53643=>"101110000",
  53644=>"111111110",
  53645=>"000101011",
  53646=>"000001111",
  53647=>"110101101",
  53648=>"000100111",
  53649=>"011011011",
  53650=>"101100111",
  53651=>"101001111",
  53652=>"011110001",
  53653=>"001101110",
  53654=>"110111111",
  53655=>"011011010",
  53656=>"001001111",
  53657=>"111101111",
  53658=>"001000010",
  53659=>"101011111",
  53660=>"111000100",
  53661=>"010100101",
  53662=>"110001101",
  53663=>"111101110",
  53664=>"101100011",
  53665=>"101011010",
  53666=>"010110010",
  53667=>"010111100",
  53668=>"001111010",
  53669=>"001010000",
  53670=>"100010011",
  53671=>"011010011",
  53672=>"111010111",
  53673=>"000001011",
  53674=>"000101111",
  53675=>"110100010",
  53676=>"111110101",
  53677=>"000100001",
  53678=>"010000101",
  53679=>"100111101",
  53680=>"010011010",
  53681=>"110100101",
  53682=>"011110010",
  53683=>"000011011",
  53684=>"000000010",
  53685=>"111000010",
  53686=>"101100010",
  53687=>"010111001",
  53688=>"100000100",
  53689=>"010010000",
  53690=>"111001001",
  53691=>"011100000",
  53692=>"101111110",
  53693=>"000011000",
  53694=>"011110111",
  53695=>"000110111",
  53696=>"011010101",
  53697=>"100001001",
  53698=>"111010111",
  53699=>"000000110",
  53700=>"110101000",
  53701=>"011101100",
  53702=>"001101000",
  53703=>"110011000",
  53704=>"011010000",
  53705=>"111001101",
  53706=>"011011001",
  53707=>"010000111",
  53708=>"101000101",
  53709=>"111001010",
  53710=>"001100000",
  53711=>"001011111",
  53712=>"010010000",
  53713=>"100000110",
  53714=>"001000011",
  53715=>"011010110",
  53716=>"110011000",
  53717=>"100100101",
  53718=>"111100111",
  53719=>"110100001",
  53720=>"000000001",
  53721=>"111111010",
  53722=>"111000101",
  53723=>"110011001",
  53724=>"101001001",
  53725=>"111100101",
  53726=>"000111101",
  53727=>"011011001",
  53728=>"011010110",
  53729=>"110010001",
  53730=>"100110100",
  53731=>"101000001",
  53732=>"100011010",
  53733=>"001010101",
  53734=>"110110010",
  53735=>"011011011",
  53736=>"001011101",
  53737=>"000111010",
  53738=>"010000001",
  53739=>"000111011",
  53740=>"111110111",
  53741=>"111100111",
  53742=>"000011000",
  53743=>"111000011",
  53744=>"001011111",
  53745=>"000011101",
  53746=>"000011100",
  53747=>"001010101",
  53748=>"011100011",
  53749=>"000100010",
  53750=>"111110101",
  53751=>"111101000",
  53752=>"101000001",
  53753=>"110000111",
  53754=>"111101111",
  53755=>"000011000",
  53756=>"011100000",
  53757=>"000111101",
  53758=>"111000001",
  53759=>"110111100",
  53760=>"101101101",
  53761=>"010111110",
  53762=>"100110101",
  53763=>"011111010",
  53764=>"000100101",
  53765=>"111010101",
  53766=>"110001101",
  53767=>"110011010",
  53768=>"111010010",
  53769=>"001010001",
  53770=>"011110010",
  53771=>"001010000",
  53772=>"101001101",
  53773=>"001010101",
  53774=>"010111110",
  53775=>"001011001",
  53776=>"111100001",
  53777=>"100110000",
  53778=>"110001010",
  53779=>"111010101",
  53780=>"111101000",
  53781=>"001111101",
  53782=>"111000101",
  53783=>"110011010",
  53784=>"011101111",
  53785=>"101100001",
  53786=>"001011001",
  53787=>"000110100",
  53788=>"000000101",
  53789=>"100010100",
  53790=>"110011000",
  53791=>"100111010",
  53792=>"010000000",
  53793=>"101110100",
  53794=>"011001000",
  53795=>"001011101",
  53796=>"011100010",
  53797=>"110100111",
  53798=>"110010100",
  53799=>"100110100",
  53800=>"110100100",
  53801=>"011111110",
  53802=>"001101001",
  53803=>"111001101",
  53804=>"100101100",
  53805=>"100101101",
  53806=>"101010001",
  53807=>"111101100",
  53808=>"100010001",
  53809=>"110110010",
  53810=>"110100010",
  53811=>"001010011",
  53812=>"001111011",
  53813=>"100111001",
  53814=>"000001111",
  53815=>"011001100",
  53816=>"010100110",
  53817=>"111101100",
  53818=>"001001010",
  53819=>"001001001",
  53820=>"000110000",
  53821=>"100101100",
  53822=>"010111100",
  53823=>"111001111",
  53824=>"000111111",
  53825=>"111011110",
  53826=>"100110000",
  53827=>"110011010",
  53828=>"111000011",
  53829=>"101011001",
  53830=>"011100000",
  53831=>"111010010",
  53832=>"000010010",
  53833=>"110010101",
  53834=>"010101000",
  53835=>"110110111",
  53836=>"001110010",
  53837=>"110100110",
  53838=>"110111110",
  53839=>"110111010",
  53840=>"100110000",
  53841=>"000101110",
  53842=>"001110001",
  53843=>"111001001",
  53844=>"010101000",
  53845=>"101110111",
  53846=>"010000001",
  53847=>"110000100",
  53848=>"001000011",
  53849=>"010100100",
  53850=>"111100110",
  53851=>"100101011",
  53852=>"101000110",
  53853=>"011000011",
  53854=>"000101001",
  53855=>"011101110",
  53856=>"110011001",
  53857=>"001010010",
  53858=>"000000100",
  53859=>"110110110",
  53860=>"001000010",
  53861=>"101000110",
  53862=>"100101011",
  53863=>"110100111",
  53864=>"001000001",
  53865=>"010111101",
  53866=>"101011110",
  53867=>"110000100",
  53868=>"001001101",
  53869=>"001001001",
  53870=>"000000101",
  53871=>"101000010",
  53872=>"010110000",
  53873=>"011111100",
  53874=>"010111111",
  53875=>"101000010",
  53876=>"100000000",
  53877=>"010000011",
  53878=>"011001110",
  53879=>"011111110",
  53880=>"100000010",
  53881=>"100111110",
  53882=>"111111100",
  53883=>"000100001",
  53884=>"110101000",
  53885=>"010011100",
  53886=>"111101101",
  53887=>"001110111",
  53888=>"110101000",
  53889=>"101110001",
  53890=>"000110100",
  53891=>"100000110",
  53892=>"110001010",
  53893=>"111100101",
  53894=>"110010010",
  53895=>"001101110",
  53896=>"010100001",
  53897=>"101011000",
  53898=>"000001000",
  53899=>"011000111",
  53900=>"001111111",
  53901=>"001011100",
  53902=>"111111001",
  53903=>"110100000",
  53904=>"110010110",
  53905=>"100100110",
  53906=>"000100010",
  53907=>"110100111",
  53908=>"000000100",
  53909=>"101100000",
  53910=>"001110101",
  53911=>"001101100",
  53912=>"110010011",
  53913=>"011000111",
  53914=>"010011010",
  53915=>"001001000",
  53916=>"100001010",
  53917=>"001110110",
  53918=>"000001101",
  53919=>"111110110",
  53920=>"111110110",
  53921=>"001100111",
  53922=>"101010011",
  53923=>"001011011",
  53924=>"100100100",
  53925=>"000011010",
  53926=>"111100000",
  53927=>"011110010",
  53928=>"010010010",
  53929=>"100001111",
  53930=>"001100100",
  53931=>"111110000",
  53932=>"001011001",
  53933=>"111000001",
  53934=>"011000001",
  53935=>"110011100",
  53936=>"010110101",
  53937=>"100010000",
  53938=>"111100110",
  53939=>"000100110",
  53940=>"110000001",
  53941=>"000100011",
  53942=>"000100110",
  53943=>"010101100",
  53944=>"010011001",
  53945=>"111101010",
  53946=>"000000111",
  53947=>"000101101",
  53948=>"000001010",
  53949=>"010010000",
  53950=>"011001010",
  53951=>"000111001",
  53952=>"100110101",
  53953=>"100100110",
  53954=>"100100010",
  53955=>"001110010",
  53956=>"100100101",
  53957=>"010111101",
  53958=>"011011011",
  53959=>"111110011",
  53960=>"110111001",
  53961=>"111110101",
  53962=>"110110101",
  53963=>"001011001",
  53964=>"001001000",
  53965=>"110010101",
  53966=>"101000100",
  53967=>"100000010",
  53968=>"111000010",
  53969=>"101111101",
  53970=>"100010000",
  53971=>"110101100",
  53972=>"011001101",
  53973=>"111000000",
  53974=>"101110110",
  53975=>"110000110",
  53976=>"000000011",
  53977=>"000111111",
  53978=>"111000101",
  53979=>"011010110",
  53980=>"010000111",
  53981=>"111111010",
  53982=>"110110111",
  53983=>"001111111",
  53984=>"101110001",
  53985=>"111000000",
  53986=>"000001100",
  53987=>"010010100",
  53988=>"111010010",
  53989=>"101100111",
  53990=>"010100001",
  53991=>"110110010",
  53992=>"010100100",
  53993=>"111101101",
  53994=>"101111011",
  53995=>"000111010",
  53996=>"010100100",
  53997=>"011110111",
  53998=>"011100100",
  53999=>"101100110",
  54000=>"100110001",
  54001=>"000010000",
  54002=>"000000111",
  54003=>"011000101",
  54004=>"101010111",
  54005=>"010001001",
  54006=>"101100011",
  54007=>"010100011",
  54008=>"001111001",
  54009=>"001110100",
  54010=>"000101111",
  54011=>"000000100",
  54012=>"011011011",
  54013=>"000100101",
  54014=>"101011010",
  54015=>"010100000",
  54016=>"100001010",
  54017=>"010100111",
  54018=>"101100110",
  54019=>"111111000",
  54020=>"100101000",
  54021=>"111000001",
  54022=>"000100100",
  54023=>"001110111",
  54024=>"000110101",
  54025=>"100000111",
  54026=>"101010100",
  54027=>"111000101",
  54028=>"010001001",
  54029=>"101101101",
  54030=>"111100111",
  54031=>"111100000",
  54032=>"010010010",
  54033=>"100100100",
  54034=>"101001101",
  54035=>"000110100",
  54036=>"101000011",
  54037=>"110000100",
  54038=>"011001010",
  54039=>"001010011",
  54040=>"010010000",
  54041=>"110000000",
  54042=>"000000010",
  54043=>"000110001",
  54044=>"010100010",
  54045=>"001110100",
  54046=>"000010001",
  54047=>"010001000",
  54048=>"010110000",
  54049=>"000001111",
  54050=>"101101111",
  54051=>"111101010",
  54052=>"111101010",
  54053=>"000101011",
  54054=>"010001100",
  54055=>"111111111",
  54056=>"011010100",
  54057=>"110111100",
  54058=>"111110000",
  54059=>"111110001",
  54060=>"100111101",
  54061=>"000010100",
  54062=>"000001011",
  54063=>"110110110",
  54064=>"000001111",
  54065=>"001100100",
  54066=>"001101111",
  54067=>"010001001",
  54068=>"100111100",
  54069=>"111010100",
  54070=>"110101110",
  54071=>"011010111",
  54072=>"101001011",
  54073=>"011101111",
  54074=>"111101011",
  54075=>"011010011",
  54076=>"010100000",
  54077=>"010100010",
  54078=>"110001000",
  54079=>"010100010",
  54080=>"001100000",
  54081=>"010001110",
  54082=>"011101001",
  54083=>"000011001",
  54084=>"101001110",
  54085=>"100110010",
  54086=>"110111000",
  54087=>"011100111",
  54088=>"000100101",
  54089=>"110010000",
  54090=>"000100101",
  54091=>"110101011",
  54092=>"011000111",
  54093=>"000010010",
  54094=>"100000000",
  54095=>"101110001",
  54096=>"111101101",
  54097=>"011000000",
  54098=>"011011001",
  54099=>"101000011",
  54100=>"001110010",
  54101=>"001111000",
  54102=>"011001111",
  54103=>"101000101",
  54104=>"111111111",
  54105=>"011100101",
  54106=>"000011111",
  54107=>"001110010",
  54108=>"000010001",
  54109=>"100001100",
  54110=>"101000000",
  54111=>"001011000",
  54112=>"111101111",
  54113=>"100111000",
  54114=>"101010000",
  54115=>"000111010",
  54116=>"111110010",
  54117=>"110011000",
  54118=>"100100010",
  54119=>"001010000",
  54120=>"110101011",
  54121=>"100110100",
  54122=>"010001110",
  54123=>"001010101",
  54124=>"101001001",
  54125=>"000001001",
  54126=>"101111111",
  54127=>"000100010",
  54128=>"101011100",
  54129=>"010011010",
  54130=>"100001011",
  54131=>"101111110",
  54132=>"001000000",
  54133=>"000010011",
  54134=>"100101001",
  54135=>"011111100",
  54136=>"100110111",
  54137=>"011011100",
  54138=>"110111101",
  54139=>"001011001",
  54140=>"100000000",
  54141=>"010011000",
  54142=>"101110101",
  54143=>"010111001",
  54144=>"011011001",
  54145=>"011010001",
  54146=>"001011000",
  54147=>"111110110",
  54148=>"000111100",
  54149=>"100001001",
  54150=>"110111000",
  54151=>"111011110",
  54152=>"000100011",
  54153=>"010110100",
  54154=>"001011000",
  54155=>"101010001",
  54156=>"111011100",
  54157=>"110001111",
  54158=>"010100011",
  54159=>"110101110",
  54160=>"111101101",
  54161=>"100111100",
  54162=>"011011010",
  54163=>"110001100",
  54164=>"100011000",
  54165=>"011001001",
  54166=>"101101101",
  54167=>"110111010",
  54168=>"111010010",
  54169=>"111010100",
  54170=>"100100111",
  54171=>"011001110",
  54172=>"110000101",
  54173=>"100000110",
  54174=>"110011000",
  54175=>"001011000",
  54176=>"101001000",
  54177=>"111011011",
  54178=>"101001011",
  54179=>"101111011",
  54180=>"000010111",
  54181=>"010110101",
  54182=>"001010101",
  54183=>"111111011",
  54184=>"010000000",
  54185=>"111010010",
  54186=>"011110110",
  54187=>"110011110",
  54188=>"110001011",
  54189=>"111100100",
  54190=>"111001001",
  54191=>"011010111",
  54192=>"000011111",
  54193=>"001100101",
  54194=>"000110101",
  54195=>"111001001",
  54196=>"101011010",
  54197=>"100011110",
  54198=>"001011110",
  54199=>"111111001",
  54200=>"011001001",
  54201=>"101001101",
  54202=>"110111001",
  54203=>"011010101",
  54204=>"000001001",
  54205=>"101010000",
  54206=>"111100000",
  54207=>"110101111",
  54208=>"000000000",
  54209=>"101000110",
  54210=>"001000011",
  54211=>"010011001",
  54212=>"000100011",
  54213=>"000111011",
  54214=>"100000101",
  54215=>"110101110",
  54216=>"011100001",
  54217=>"101001100",
  54218=>"011010101",
  54219=>"011100111",
  54220=>"101110000",
  54221=>"101000101",
  54222=>"000110000",
  54223=>"010010100",
  54224=>"100101000",
  54225=>"000010101",
  54226=>"110100000",
  54227=>"011011101",
  54228=>"000110111",
  54229=>"110100100",
  54230=>"001101010",
  54231=>"001001000",
  54232=>"110111010",
  54233=>"000100101",
  54234=>"000111010",
  54235=>"000000111",
  54236=>"100111010",
  54237=>"100011111",
  54238=>"000000110",
  54239=>"110111010",
  54240=>"011000110",
  54241=>"110110100",
  54242=>"001000100",
  54243=>"001000001",
  54244=>"101100100",
  54245=>"111001000",
  54246=>"110110101",
  54247=>"101110101",
  54248=>"100001000",
  54249=>"000010111",
  54250=>"001100001",
  54251=>"000000111",
  54252=>"011100010",
  54253=>"001100110",
  54254=>"000011000",
  54255=>"000110100",
  54256=>"001000000",
  54257=>"000001100",
  54258=>"011111110",
  54259=>"111010100",
  54260=>"101001111",
  54261=>"001011000",
  54262=>"100100100",
  54263=>"111011100",
  54264=>"010011010",
  54265=>"111001001",
  54266=>"000111011",
  54267=>"010101101",
  54268=>"110000100",
  54269=>"111101101",
  54270=>"001010000",
  54271=>"011110100",
  54272=>"100010010",
  54273=>"101010100",
  54274=>"110011100",
  54275=>"101001000",
  54276=>"010101001",
  54277=>"101100100",
  54278=>"101101100",
  54279=>"000111000",
  54280=>"111111101",
  54281=>"000100010",
  54282=>"010001110",
  54283=>"101101111",
  54284=>"011010000",
  54285=>"010111111",
  54286=>"111101100",
  54287=>"110101111",
  54288=>"111101110",
  54289=>"010001100",
  54290=>"000110010",
  54291=>"001101111",
  54292=>"011001000",
  54293=>"001000001",
  54294=>"000101101",
  54295=>"011001001",
  54296=>"010010011",
  54297=>"100011110",
  54298=>"100010010",
  54299=>"101000110",
  54300=>"001010011",
  54301=>"100100010",
  54302=>"010110000",
  54303=>"110100100",
  54304=>"100101001",
  54305=>"100110111",
  54306=>"011001011",
  54307=>"011110000",
  54308=>"100111110",
  54309=>"011110101",
  54310=>"101110111",
  54311=>"111110000",
  54312=>"111100101",
  54313=>"001110100",
  54314=>"101111110",
  54315=>"110110000",
  54316=>"000100100",
  54317=>"011011010",
  54318=>"000011010",
  54319=>"101011011",
  54320=>"110110101",
  54321=>"000111111",
  54322=>"110100100",
  54323=>"000000000",
  54324=>"000001110",
  54325=>"010101010",
  54326=>"000100100",
  54327=>"111111100",
  54328=>"110111011",
  54329=>"011000101",
  54330=>"110000000",
  54331=>"110011011",
  54332=>"010010000",
  54333=>"010000001",
  54334=>"001001000",
  54335=>"010101001",
  54336=>"001111111",
  54337=>"000111001",
  54338=>"000110110",
  54339=>"111001010",
  54340=>"010011011",
  54341=>"100110010",
  54342=>"001110001",
  54343=>"000101001",
  54344=>"100000110",
  54345=>"011001101",
  54346=>"000010000",
  54347=>"001100001",
  54348=>"001101011",
  54349=>"011000111",
  54350=>"010101111",
  54351=>"000101100",
  54352=>"000110111",
  54353=>"010010010",
  54354=>"100100101",
  54355=>"001000100",
  54356=>"101010010",
  54357=>"101101111",
  54358=>"101110000",
  54359=>"111100111",
  54360=>"001110100",
  54361=>"100101110",
  54362=>"000011110",
  54363=>"110010000",
  54364=>"101111001",
  54365=>"000101000",
  54366=>"011100110",
  54367=>"001011111",
  54368=>"010100010",
  54369=>"001110101",
  54370=>"101101000",
  54371=>"010100000",
  54372=>"110010111",
  54373=>"000001101",
  54374=>"100010110",
  54375=>"011100111",
  54376=>"011000100",
  54377=>"000001110",
  54378=>"101011110",
  54379=>"101101110",
  54380=>"011001110",
  54381=>"101100111",
  54382=>"011001000",
  54383=>"011001111",
  54384=>"001000000",
  54385=>"010010101",
  54386=>"000000001",
  54387=>"000011101",
  54388=>"101111110",
  54389=>"111001100",
  54390=>"110110110",
  54391=>"010000000",
  54392=>"100011101",
  54393=>"110100010",
  54394=>"110111111",
  54395=>"010010111",
  54396=>"011000101",
  54397=>"101100111",
  54398=>"111111111",
  54399=>"101110101",
  54400=>"010101111",
  54401=>"011000110",
  54402=>"101011000",
  54403=>"011010111",
  54404=>"110110010",
  54405=>"111101101",
  54406=>"111001101",
  54407=>"010000011",
  54408=>"100111111",
  54409=>"100001001",
  54410=>"100111010",
  54411=>"010000100",
  54412=>"011000000",
  54413=>"111110101",
  54414=>"100111010",
  54415=>"000100101",
  54416=>"110111000",
  54417=>"001001110",
  54418=>"010000010",
  54419=>"101011010",
  54420=>"001010100",
  54421=>"110010000",
  54422=>"010101110",
  54423=>"010111010",
  54424=>"010001111",
  54425=>"111101010",
  54426=>"101100110",
  54427=>"110111101",
  54428=>"110000100",
  54429=>"001010011",
  54430=>"010001011",
  54431=>"011000111",
  54432=>"001101111",
  54433=>"111100110",
  54434=>"101100001",
  54435=>"001111110",
  54436=>"100001110",
  54437=>"111011000",
  54438=>"110011110",
  54439=>"100010011",
  54440=>"011011110",
  54441=>"110111011",
  54442=>"110000010",
  54443=>"110001011",
  54444=>"100110011",
  54445=>"100000001",
  54446=>"100111101",
  54447=>"100000110",
  54448=>"111110001",
  54449=>"010010100",
  54450=>"001001001",
  54451=>"111111000",
  54452=>"110000011",
  54453=>"110001100",
  54454=>"100110000",
  54455=>"110000111",
  54456=>"001000111",
  54457=>"001101100",
  54458=>"111011111",
  54459=>"111110001",
  54460=>"100111001",
  54461=>"011110101",
  54462=>"011011111",
  54463=>"010111001",
  54464=>"001011111",
  54465=>"001010110",
  54466=>"010000000",
  54467=>"000011011",
  54468=>"011010111",
  54469=>"111101011",
  54470=>"001010110",
  54471=>"110101001",
  54472=>"000011001",
  54473=>"100101101",
  54474=>"001010001",
  54475=>"110110110",
  54476=>"110010100",
  54477=>"111001101",
  54478=>"000101011",
  54479=>"010010001",
  54480=>"000110000",
  54481=>"010001010",
  54482=>"000110000",
  54483=>"100111110",
  54484=>"100000000",
  54485=>"010111100",
  54486=>"000011000",
  54487=>"010010110",
  54488=>"001000101",
  54489=>"010111010",
  54490=>"001000010",
  54491=>"100010111",
  54492=>"011001000",
  54493=>"001101110",
  54494=>"000111100",
  54495=>"100001010",
  54496=>"100011111",
  54497=>"001101011",
  54498=>"110000011",
  54499=>"011011010",
  54500=>"101101000",
  54501=>"001011011",
  54502=>"100101010",
  54503=>"000011011",
  54504=>"011000001",
  54505=>"111000010",
  54506=>"000100010",
  54507=>"111111001",
  54508=>"100110010",
  54509=>"100011001",
  54510=>"110100010",
  54511=>"000100010",
  54512=>"000110001",
  54513=>"000001110",
  54514=>"000000101",
  54515=>"010011011",
  54516=>"111000110",
  54517=>"111110101",
  54518=>"111010100",
  54519=>"001010111",
  54520=>"100010011",
  54521=>"010101001",
  54522=>"101110010",
  54523=>"110111010",
  54524=>"010011011",
  54525=>"001111000",
  54526=>"100101010",
  54527=>"110001001",
  54528=>"000001100",
  54529=>"001101101",
  54530=>"101100010",
  54531=>"101111010",
  54532=>"000111000",
  54533=>"000011110",
  54534=>"010110000",
  54535=>"001010110",
  54536=>"110101001",
  54537=>"011110101",
  54538=>"010011001",
  54539=>"000011110",
  54540=>"100010110",
  54541=>"111111011",
  54542=>"100001010",
  54543=>"000010111",
  54544=>"001100000",
  54545=>"100010100",
  54546=>"100101111",
  54547=>"011010100",
  54548=>"110010000",
  54549=>"010000100",
  54550=>"000001000",
  54551=>"010010111",
  54552=>"001101110",
  54553=>"000000000",
  54554=>"001111001",
  54555=>"011101111",
  54556=>"000010101",
  54557=>"101011111",
  54558=>"011111111",
  54559=>"011100000",
  54560=>"100011111",
  54561=>"101000010",
  54562=>"101010010",
  54563=>"110100110",
  54564=>"000101111",
  54565=>"011100110",
  54566=>"001110101",
  54567=>"110001000",
  54568=>"000011110",
  54569=>"000001010",
  54570=>"010000000",
  54571=>"011010011",
  54572=>"011111110",
  54573=>"000010011",
  54574=>"100001100",
  54575=>"111111000",
  54576=>"011000011",
  54577=>"100111111",
  54578=>"001101100",
  54579=>"000110010",
  54580=>"000010011",
  54581=>"101010010",
  54582=>"011111100",
  54583=>"000110110",
  54584=>"001000101",
  54585=>"101001110",
  54586=>"101011001",
  54587=>"101111011",
  54588=>"111001111",
  54589=>"000101111",
  54590=>"010000011",
  54591=>"101011111",
  54592=>"100011011",
  54593=>"100010010",
  54594=>"110111000",
  54595=>"001010000",
  54596=>"000100010",
  54597=>"000101001",
  54598=>"011001011",
  54599=>"101100000",
  54600=>"001110111",
  54601=>"101010001",
  54602=>"100000001",
  54603=>"000000100",
  54604=>"100001010",
  54605=>"011011100",
  54606=>"010000011",
  54607=>"101000001",
  54608=>"000011111",
  54609=>"101111111",
  54610=>"110001001",
  54611=>"010011000",
  54612=>"000100111",
  54613=>"010100010",
  54614=>"101011110",
  54615=>"010100010",
  54616=>"100011100",
  54617=>"111000111",
  54618=>"001111101",
  54619=>"111000111",
  54620=>"000111110",
  54621=>"111100111",
  54622=>"010110111",
  54623=>"100110000",
  54624=>"010011000",
  54625=>"010011010",
  54626=>"110011100",
  54627=>"111110010",
  54628=>"111000000",
  54629=>"111001010",
  54630=>"101000100",
  54631=>"001001100",
  54632=>"000000000",
  54633=>"110100101",
  54634=>"010000001",
  54635=>"001000100",
  54636=>"110001101",
  54637=>"000001100",
  54638=>"000101110",
  54639=>"100110001",
  54640=>"100110101",
  54641=>"101100001",
  54642=>"110111100",
  54643=>"100001111",
  54644=>"001101100",
  54645=>"111011100",
  54646=>"010111001",
  54647=>"011111110",
  54648=>"101110001",
  54649=>"110000001",
  54650=>"001001010",
  54651=>"101010111",
  54652=>"000100000",
  54653=>"000110011",
  54654=>"001011000",
  54655=>"000000001",
  54656=>"101101001",
  54657=>"111011101",
  54658=>"101011011",
  54659=>"000110000",
  54660=>"011111101",
  54661=>"000111110",
  54662=>"100010001",
  54663=>"100010001",
  54664=>"100000101",
  54665=>"101001000",
  54666=>"111100110",
  54667=>"101101100",
  54668=>"100110001",
  54669=>"001000010",
  54670=>"011010110",
  54671=>"100101001",
  54672=>"111110111",
  54673=>"011010110",
  54674=>"011000101",
  54675=>"001110001",
  54676=>"110011110",
  54677=>"000111110",
  54678=>"110101000",
  54679=>"011000110",
  54680=>"100110001",
  54681=>"111000110",
  54682=>"100000110",
  54683=>"011110100",
  54684=>"010001100",
  54685=>"010010111",
  54686=>"111000010",
  54687=>"000000000",
  54688=>"101101100",
  54689=>"001101001",
  54690=>"101111001",
  54691=>"100110111",
  54692=>"000010011",
  54693=>"001100111",
  54694=>"000010010",
  54695=>"111010001",
  54696=>"110010010",
  54697=>"000011111",
  54698=>"011000110",
  54699=>"100111101",
  54700=>"010101011",
  54701=>"111011111",
  54702=>"010010000",
  54703=>"001111001",
  54704=>"100000001",
  54705=>"011000000",
  54706=>"011101101",
  54707=>"001000100",
  54708=>"011101101",
  54709=>"111100011",
  54710=>"001110010",
  54711=>"111110110",
  54712=>"001010110",
  54713=>"000100100",
  54714=>"110101001",
  54715=>"110110000",
  54716=>"111001000",
  54717=>"111110011",
  54718=>"101011100",
  54719=>"111011111",
  54720=>"101011111",
  54721=>"010110101",
  54722=>"010110011",
  54723=>"011111111",
  54724=>"111000001",
  54725=>"001101010",
  54726=>"111001100",
  54727=>"001100001",
  54728=>"000100101",
  54729=>"010111000",
  54730=>"011000010",
  54731=>"100101101",
  54732=>"010101011",
  54733=>"101000010",
  54734=>"001111101",
  54735=>"000000110",
  54736=>"010010101",
  54737=>"101011101",
  54738=>"001010010",
  54739=>"011111100",
  54740=>"100111111",
  54741=>"111011000",
  54742=>"100111111",
  54743=>"111011110",
  54744=>"001100101",
  54745=>"001110000",
  54746=>"110000100",
  54747=>"000111001",
  54748=>"100110101",
  54749=>"110100011",
  54750=>"000110001",
  54751=>"110110101",
  54752=>"010010111",
  54753=>"111000010",
  54754=>"111010111",
  54755=>"101101110",
  54756=>"001110110",
  54757=>"101111100",
  54758=>"111111100",
  54759=>"001000011",
  54760=>"001101111",
  54761=>"011010100",
  54762=>"100000011",
  54763=>"010000110",
  54764=>"110110011",
  54765=>"010010101",
  54766=>"001111111",
  54767=>"101000001",
  54768=>"001011101",
  54769=>"100101000",
  54770=>"110100001",
  54771=>"111011010",
  54772=>"101011100",
  54773=>"100000010",
  54774=>"001111000",
  54775=>"000111100",
  54776=>"011010111",
  54777=>"110000010",
  54778=>"100010010",
  54779=>"110010011",
  54780=>"011100010",
  54781=>"000011111",
  54782=>"100111100",
  54783=>"000111111",
  54784=>"110000110",
  54785=>"101011101",
  54786=>"000100100",
  54787=>"111100011",
  54788=>"110100111",
  54789=>"000111101",
  54790=>"011011101",
  54791=>"000100000",
  54792=>"001000111",
  54793=>"000100111",
  54794=>"111001100",
  54795=>"000001011",
  54796=>"001001000",
  54797=>"000111101",
  54798=>"001000101",
  54799=>"010011101",
  54800=>"110011010",
  54801=>"110100010",
  54802=>"111001101",
  54803=>"001010110",
  54804=>"010010110",
  54805=>"110000010",
  54806=>"100001010",
  54807=>"100101011",
  54808=>"010001101",
  54809=>"100011110",
  54810=>"011001000",
  54811=>"001100010",
  54812=>"110001110",
  54813=>"000100000",
  54814=>"011011110",
  54815=>"010101010",
  54816=>"111110100",
  54817=>"111010000",
  54818=>"010000011",
  54819=>"111101101",
  54820=>"100100000",
  54821=>"110110001",
  54822=>"110100100",
  54823=>"101111010",
  54824=>"001110110",
  54825=>"000111000",
  54826=>"000110110",
  54827=>"010001011",
  54828=>"010110111",
  54829=>"110100010",
  54830=>"101110001",
  54831=>"110001001",
  54832=>"111000010",
  54833=>"100110010",
  54834=>"101001011",
  54835=>"000101001",
  54836=>"011100110",
  54837=>"100010010",
  54838=>"001000011",
  54839=>"110100111",
  54840=>"000000000",
  54841=>"010000000",
  54842=>"110111110",
  54843=>"000100011",
  54844=>"111101111",
  54845=>"000000011",
  54846=>"000001001",
  54847=>"101000011",
  54848=>"110111101",
  54849=>"101010011",
  54850=>"001000111",
  54851=>"011100010",
  54852=>"010000110",
  54853=>"101010010",
  54854=>"110111110",
  54855=>"010011100",
  54856=>"110111101",
  54857=>"011010100",
  54858=>"010111111",
  54859=>"001111111",
  54860=>"101001111",
  54861=>"000110100",
  54862=>"110000010",
  54863=>"111001010",
  54864=>"011100010",
  54865=>"010100111",
  54866=>"011010100",
  54867=>"111110101",
  54868=>"000011100",
  54869=>"001100100",
  54870=>"000011010",
  54871=>"001110011",
  54872=>"111111111",
  54873=>"001101111",
  54874=>"111000101",
  54875=>"000110010",
  54876=>"000110000",
  54877=>"101110000",
  54878=>"010001110",
  54879=>"100011001",
  54880=>"000010000",
  54881=>"100000000",
  54882=>"000110111",
  54883=>"100110111",
  54884=>"001001100",
  54885=>"101001001",
  54886=>"001001011",
  54887=>"111001010",
  54888=>"000101000",
  54889=>"000001101",
  54890=>"111110011",
  54891=>"001000000",
  54892=>"000010110",
  54893=>"110110001",
  54894=>"001010101",
  54895=>"100000111",
  54896=>"011001101",
  54897=>"001000000",
  54898=>"000111000",
  54899=>"110111100",
  54900=>"000100100",
  54901=>"001111011",
  54902=>"101111001",
  54903=>"100000001",
  54904=>"000011001",
  54905=>"011101101",
  54906=>"110100111",
  54907=>"101000010",
  54908=>"011010111",
  54909=>"000001010",
  54910=>"111001010",
  54911=>"001011111",
  54912=>"000011101",
  54913=>"000000001",
  54914=>"011011010",
  54915=>"111000001",
  54916=>"010111001",
  54917=>"011110011",
  54918=>"001011001",
  54919=>"010011001",
  54920=>"110001001",
  54921=>"111010110",
  54922=>"111100101",
  54923=>"100110100",
  54924=>"100001110",
  54925=>"110100110",
  54926=>"010001100",
  54927=>"011111100",
  54928=>"110001001",
  54929=>"111101010",
  54930=>"110010101",
  54931=>"101011000",
  54932=>"100111110",
  54933=>"111111110",
  54934=>"011001011",
  54935=>"111011011",
  54936=>"001010000",
  54937=>"101000111",
  54938=>"010101001",
  54939=>"000001001",
  54940=>"100001010",
  54941=>"101010010",
  54942=>"011101010",
  54943=>"110111000",
  54944=>"110111110",
  54945=>"011010111",
  54946=>"111011010",
  54947=>"011000101",
  54948=>"010010011",
  54949=>"011010110",
  54950=>"010010000",
  54951=>"110000111",
  54952=>"111101000",
  54953=>"001111001",
  54954=>"011001101",
  54955=>"110100100",
  54956=>"001110001",
  54957=>"000101111",
  54958=>"110100111",
  54959=>"001101101",
  54960=>"101000001",
  54961=>"001011111",
  54962=>"111000011",
  54963=>"001110101",
  54964=>"111101101",
  54965=>"111111001",
  54966=>"101001001",
  54967=>"010111100",
  54968=>"110010101",
  54969=>"011100010",
  54970=>"110000100",
  54971=>"110000111",
  54972=>"011101101",
  54973=>"110000110",
  54974=>"100110011",
  54975=>"001100100",
  54976=>"011110010",
  54977=>"001101100",
  54978=>"001111100",
  54979=>"000110001",
  54980=>"010011001",
  54981=>"011000100",
  54982=>"110110001",
  54983=>"010101100",
  54984=>"000000100",
  54985=>"100010111",
  54986=>"011010010",
  54987=>"111100000",
  54988=>"001101101",
  54989=>"000000000",
  54990=>"111011011",
  54991=>"010100110",
  54992=>"111010100",
  54993=>"110011111",
  54994=>"110100011",
  54995=>"101110000",
  54996=>"010110101",
  54997=>"111111111",
  54998=>"001110000",
  54999=>"110000110",
  55000=>"010000001",
  55001=>"101100001",
  55002=>"000000100",
  55003=>"111101010",
  55004=>"010100101",
  55005=>"000011001",
  55006=>"110111110",
  55007=>"010010110",
  55008=>"000010010",
  55009=>"100100111",
  55010=>"111010100",
  55011=>"000010011",
  55012=>"101111001",
  55013=>"101110000",
  55014=>"111111111",
  55015=>"010110110",
  55016=>"001110001",
  55017=>"110101000",
  55018=>"000110101",
  55019=>"100101110",
  55020=>"101110111",
  55021=>"110100111",
  55022=>"111101010",
  55023=>"110001101",
  55024=>"010110100",
  55025=>"001100110",
  55026=>"100011010",
  55027=>"010010111",
  55028=>"100110101",
  55029=>"010000110",
  55030=>"111110110",
  55031=>"011101000",
  55032=>"011110000",
  55033=>"110101110",
  55034=>"010001111",
  55035=>"110001101",
  55036=>"101010001",
  55037=>"001001011",
  55038=>"100100101",
  55039=>"101001101",
  55040=>"010010101",
  55041=>"101011000",
  55042=>"000111111",
  55043=>"110010010",
  55044=>"110000100",
  55045=>"011000001",
  55046=>"111100110",
  55047=>"011001010",
  55048=>"111101111",
  55049=>"101110111",
  55050=>"110111100",
  55051=>"110101001",
  55052=>"111011111",
  55053=>"000101111",
  55054=>"111100010",
  55055=>"101011110",
  55056=>"111110000",
  55057=>"010101100",
  55058=>"000010001",
  55059=>"101101100",
  55060=>"010010011",
  55061=>"011011001",
  55062=>"011001100",
  55063=>"101001110",
  55064=>"110011001",
  55065=>"000111010",
  55066=>"001000100",
  55067=>"010111001",
  55068=>"100101100",
  55069=>"110001111",
  55070=>"010001011",
  55071=>"111011110",
  55072=>"010100110",
  55073=>"101100110",
  55074=>"100011111",
  55075=>"111000010",
  55076=>"011000111",
  55077=>"101000001",
  55078=>"001110101",
  55079=>"110011111",
  55080=>"111100100",
  55081=>"101001101",
  55082=>"011111110",
  55083=>"001100001",
  55084=>"011100011",
  55085=>"001010001",
  55086=>"110000111",
  55087=>"000100100",
  55088=>"100011111",
  55089=>"011001011",
  55090=>"100110010",
  55091=>"010101000",
  55092=>"101011000",
  55093=>"110111000",
  55094=>"110001010",
  55095=>"001101010",
  55096=>"011110101",
  55097=>"000101000",
  55098=>"010000000",
  55099=>"111011100",
  55100=>"010101011",
  55101=>"010011001",
  55102=>"110011101",
  55103=>"111101101",
  55104=>"001000011",
  55105=>"000001101",
  55106=>"001111111",
  55107=>"100000010",
  55108=>"101100111",
  55109=>"101001011",
  55110=>"110101110",
  55111=>"011011000",
  55112=>"101011000",
  55113=>"100101101",
  55114=>"011000000",
  55115=>"111001110",
  55116=>"110101111",
  55117=>"111001011",
  55118=>"010011010",
  55119=>"111010001",
  55120=>"101111011",
  55121=>"100010111",
  55122=>"011000111",
  55123=>"000001111",
  55124=>"010010100",
  55125=>"111101110",
  55126=>"100110010",
  55127=>"111001001",
  55128=>"001011011",
  55129=>"000001001",
  55130=>"100100110",
  55131=>"001101111",
  55132=>"001001010",
  55133=>"001000111",
  55134=>"101010111",
  55135=>"100011011",
  55136=>"101001000",
  55137=>"001100001",
  55138=>"101011001",
  55139=>"000001110",
  55140=>"111101101",
  55141=>"100100001",
  55142=>"011110101",
  55143=>"101010110",
  55144=>"111000000",
  55145=>"110111111",
  55146=>"000100001",
  55147=>"100010101",
  55148=>"111100010",
  55149=>"011010000",
  55150=>"010011100",
  55151=>"111011111",
  55152=>"001000001",
  55153=>"010100010",
  55154=>"000000110",
  55155=>"010110010",
  55156=>"001011101",
  55157=>"100000011",
  55158=>"110101111",
  55159=>"100011000",
  55160=>"110111110",
  55161=>"001111011",
  55162=>"011110001",
  55163=>"010000101",
  55164=>"011101001",
  55165=>"101110001",
  55166=>"001010111",
  55167=>"001011101",
  55168=>"111110000",
  55169=>"011010101",
  55170=>"011101001",
  55171=>"101000011",
  55172=>"010101000",
  55173=>"101000110",
  55174=>"000001001",
  55175=>"011011011",
  55176=>"000110010",
  55177=>"010100010",
  55178=>"011100110",
  55179=>"000100001",
  55180=>"000010000",
  55181=>"111100001",
  55182=>"100001000",
  55183=>"000101010",
  55184=>"001110111",
  55185=>"110111011",
  55186=>"110100001",
  55187=>"111000010",
  55188=>"101001100",
  55189=>"000010010",
  55190=>"010010000",
  55191=>"100111001",
  55192=>"101010011",
  55193=>"001010101",
  55194=>"101010001",
  55195=>"010011010",
  55196=>"110100111",
  55197=>"010111111",
  55198=>"110101010",
  55199=>"000110000",
  55200=>"000001100",
  55201=>"001110101",
  55202=>"111000001",
  55203=>"010000001",
  55204=>"010000011",
  55205=>"110100101",
  55206=>"111110100",
  55207=>"011011011",
  55208=>"011011111",
  55209=>"100011000",
  55210=>"001101100",
  55211=>"111010011",
  55212=>"000000100",
  55213=>"100011010",
  55214=>"101011100",
  55215=>"000010000",
  55216=>"111111001",
  55217=>"010111110",
  55218=>"011010011",
  55219=>"100000101",
  55220=>"101010101",
  55221=>"000101101",
  55222=>"111100110",
  55223=>"000011101",
  55224=>"110100110",
  55225=>"101100111",
  55226=>"100110010",
  55227=>"000101111",
  55228=>"011010110",
  55229=>"011110010",
  55230=>"011100010",
  55231=>"010111110",
  55232=>"000011011",
  55233=>"010100000",
  55234=>"100001100",
  55235=>"100001011",
  55236=>"010011000",
  55237=>"111010001",
  55238=>"110010011",
  55239=>"000000101",
  55240=>"010011111",
  55241=>"111011110",
  55242=>"101101000",
  55243=>"111111100",
  55244=>"111011000",
  55245=>"001101000",
  55246=>"100000110",
  55247=>"100100101",
  55248=>"010001010",
  55249=>"010001101",
  55250=>"100000000",
  55251=>"011010000",
  55252=>"010011100",
  55253=>"010111110",
  55254=>"000010000",
  55255=>"000101011",
  55256=>"011001110",
  55257=>"000001011",
  55258=>"100000100",
  55259=>"100011001",
  55260=>"111100010",
  55261=>"101011101",
  55262=>"100000010",
  55263=>"110111110",
  55264=>"110111100",
  55265=>"000000001",
  55266=>"011010111",
  55267=>"111110011",
  55268=>"111111010",
  55269=>"111101001",
  55270=>"110000111",
  55271=>"011000010",
  55272=>"110110100",
  55273=>"001100000",
  55274=>"100100011",
  55275=>"110001100",
  55276=>"110101010",
  55277=>"100010101",
  55278=>"110001010",
  55279=>"100000010",
  55280=>"110000000",
  55281=>"101111011",
  55282=>"101000100",
  55283=>"011001110",
  55284=>"011110111",
  55285=>"010111011",
  55286=>"110111100",
  55287=>"111111010",
  55288=>"101001101",
  55289=>"110110101",
  55290=>"011000100",
  55291=>"000100101",
  55292=>"001111010",
  55293=>"011011100",
  55294=>"000011111",
  55295=>"100110111",
  55296=>"011100000",
  55297=>"001011111",
  55298=>"000000010",
  55299=>"001110011",
  55300=>"100111000",
  55301=>"010111111",
  55302=>"001000000",
  55303=>"110101010",
  55304=>"110001011",
  55305=>"011011100",
  55306=>"010101101",
  55307=>"001000001",
  55308=>"010001100",
  55309=>"101110001",
  55310=>"111110011",
  55311=>"100101100",
  55312=>"100010011",
  55313=>"001101110",
  55314=>"100010011",
  55315=>"000010100",
  55316=>"100000000",
  55317=>"000010100",
  55318=>"001110001",
  55319=>"110010101",
  55320=>"110011001",
  55321=>"000101001",
  55322=>"101110111",
  55323=>"100111101",
  55324=>"100010010",
  55325=>"000011101",
  55326=>"011011011",
  55327=>"011000000",
  55328=>"011101001",
  55329=>"101001011",
  55330=>"101100100",
  55331=>"111000111",
  55332=>"111010011",
  55333=>"100110010",
  55334=>"000111010",
  55335=>"101011000",
  55336=>"000100110",
  55337=>"011100111",
  55338=>"100101101",
  55339=>"010001011",
  55340=>"011010001",
  55341=>"101010100",
  55342=>"000100000",
  55343=>"000110010",
  55344=>"100111111",
  55345=>"000010010",
  55346=>"000101110",
  55347=>"000010101",
  55348=>"111000010",
  55349=>"110100011",
  55350=>"010101001",
  55351=>"100100011",
  55352=>"010100011",
  55353=>"010010111",
  55354=>"011000110",
  55355=>"101010110",
  55356=>"111000000",
  55357=>"100010001",
  55358=>"110111110",
  55359=>"000100001",
  55360=>"110011011",
  55361=>"000100011",
  55362=>"001100010",
  55363=>"100010010",
  55364=>"110100100",
  55365=>"100110001",
  55366=>"011001111",
  55367=>"010010001",
  55368=>"001000000",
  55369=>"101111101",
  55370=>"100001111",
  55371=>"010101111",
  55372=>"001000000",
  55373=>"010110101",
  55374=>"111001011",
  55375=>"010110101",
  55376=>"011011110",
  55377=>"010100010",
  55378=>"100101001",
  55379=>"100000110",
  55380=>"001110001",
  55381=>"010110100",
  55382=>"101101000",
  55383=>"001000100",
  55384=>"010111000",
  55385=>"101000111",
  55386=>"011000001",
  55387=>"100000100",
  55388=>"010101101",
  55389=>"001101011",
  55390=>"010010101",
  55391=>"110101001",
  55392=>"011000110",
  55393=>"001001010",
  55394=>"000000111",
  55395=>"000000010",
  55396=>"101110101",
  55397=>"100011101",
  55398=>"011000111",
  55399=>"000001001",
  55400=>"011111011",
  55401=>"110110110",
  55402=>"110111001",
  55403=>"111011010",
  55404=>"010111000",
  55405=>"000101111",
  55406=>"011011100",
  55407=>"001001101",
  55408=>"110101101",
  55409=>"101001001",
  55410=>"101110101",
  55411=>"100011101",
  55412=>"011011110",
  55413=>"101011010",
  55414=>"010110100",
  55415=>"110000001",
  55416=>"101010101",
  55417=>"101001001",
  55418=>"001011101",
  55419=>"000011110",
  55420=>"111101100",
  55421=>"101011100",
  55422=>"101001101",
  55423=>"001100000",
  55424=>"001010011",
  55425=>"110000110",
  55426=>"101010000",
  55427=>"000001100",
  55428=>"111101001",
  55429=>"111001011",
  55430=>"001011111",
  55431=>"010000010",
  55432=>"100001010",
  55433=>"111001000",
  55434=>"000101000",
  55435=>"000001010",
  55436=>"010010010",
  55437=>"111110111",
  55438=>"111010000",
  55439=>"111001000",
  55440=>"001001010",
  55441=>"010011011",
  55442=>"011011101",
  55443=>"000100011",
  55444=>"111111110",
  55445=>"001111111",
  55446=>"001001010",
  55447=>"001000110",
  55448=>"000000001",
  55449=>"010001101",
  55450=>"101000110",
  55451=>"000010101",
  55452=>"101011111",
  55453=>"011010011",
  55454=>"010101010",
  55455=>"100011010",
  55456=>"010110111",
  55457=>"111001101",
  55458=>"000110001",
  55459=>"101000100",
  55460=>"101111100",
  55461=>"110100101",
  55462=>"001010101",
  55463=>"010010001",
  55464=>"000001000",
  55465=>"000000000",
  55466=>"010010001",
  55467=>"001100111",
  55468=>"101101010",
  55469=>"001010111",
  55470=>"010010111",
  55471=>"010010111",
  55472=>"111000111",
  55473=>"011110000",
  55474=>"000001111",
  55475=>"110110010",
  55476=>"000101001",
  55477=>"101111100",
  55478=>"101100111",
  55479=>"010000101",
  55480=>"010001100",
  55481=>"111011000",
  55482=>"001101010",
  55483=>"110111101",
  55484=>"001111001",
  55485=>"000010001",
  55486=>"111101111",
  55487=>"011001010",
  55488=>"101000111",
  55489=>"000011000",
  55490=>"110010100",
  55491=>"000111101",
  55492=>"101000001",
  55493=>"001001101",
  55494=>"001101011",
  55495=>"110010000",
  55496=>"011000001",
  55497=>"100010100",
  55498=>"000001001",
  55499=>"011110101",
  55500=>"000100100",
  55501=>"100010100",
  55502=>"011110100",
  55503=>"000001011",
  55504=>"010000100",
  55505=>"101001111",
  55506=>"010000100",
  55507=>"010011000",
  55508=>"010110000",
  55509=>"010001001",
  55510=>"101011011",
  55511=>"011100100",
  55512=>"010000100",
  55513=>"011101101",
  55514=>"010110001",
  55515=>"000100011",
  55516=>"001011000",
  55517=>"001101011",
  55518=>"010101001",
  55519=>"000010001",
  55520=>"010010100",
  55521=>"000000100",
  55522=>"001110110",
  55523=>"000101110",
  55524=>"110001010",
  55525=>"000111100",
  55526=>"000010101",
  55527=>"010111010",
  55528=>"101000101",
  55529=>"010110101",
  55530=>"000111001",
  55531=>"001001011",
  55532=>"001011011",
  55533=>"111110110",
  55534=>"101101010",
  55535=>"111100000",
  55536=>"011010000",
  55537=>"000111101",
  55538=>"010000000",
  55539=>"011001000",
  55540=>"101010000",
  55541=>"111010101",
  55542=>"000110101",
  55543=>"001100101",
  55544=>"001111000",
  55545=>"100101110",
  55546=>"010110110",
  55547=>"000111111",
  55548=>"010010100",
  55549=>"000011001",
  55550=>"111001111",
  55551=>"010010001",
  55552=>"000111111",
  55553=>"100110000",
  55554=>"111101100",
  55555=>"001101000",
  55556=>"100101110",
  55557=>"100100100",
  55558=>"000100111",
  55559=>"110000000",
  55560=>"110010100",
  55561=>"101110111",
  55562=>"010001011",
  55563=>"111111011",
  55564=>"001000010",
  55565=>"110001000",
  55566=>"111100100",
  55567=>"000001001",
  55568=>"111101101",
  55569=>"110110010",
  55570=>"001101100",
  55571=>"001110100",
  55572=>"001010110",
  55573=>"111010100",
  55574=>"100000010",
  55575=>"001111101",
  55576=>"111110100",
  55577=>"101100000",
  55578=>"110001110",
  55579=>"101001110",
  55580=>"000010010",
  55581=>"111101101",
  55582=>"101011111",
  55583=>"111110000",
  55584=>"001111100",
  55585=>"101011111",
  55586=>"111100011",
  55587=>"110100101",
  55588=>"111100011",
  55589=>"011011101",
  55590=>"100100101",
  55591=>"111101101",
  55592=>"101111111",
  55593=>"000000111",
  55594=>"000101110",
  55595=>"010001111",
  55596=>"001010000",
  55597=>"110101101",
  55598=>"111110010",
  55599=>"110101001",
  55600=>"010000000",
  55601=>"001010110",
  55602=>"010111000",
  55603=>"110010101",
  55604=>"011111000",
  55605=>"100101101",
  55606=>"100011000",
  55607=>"111000110",
  55608=>"100010001",
  55609=>"011101001",
  55610=>"101011111",
  55611=>"001001100",
  55612=>"011110111",
  55613=>"010000100",
  55614=>"111100000",
  55615=>"101100101",
  55616=>"010111001",
  55617=>"100110000",
  55618=>"101101001",
  55619=>"111001011",
  55620=>"001001010",
  55621=>"101111010",
  55622=>"010001001",
  55623=>"111010110",
  55624=>"000111011",
  55625=>"101000000",
  55626=>"100010010",
  55627=>"001100011",
  55628=>"100010111",
  55629=>"101010101",
  55630=>"111100100",
  55631=>"100100011",
  55632=>"101000010",
  55633=>"000011111",
  55634=>"000100010",
  55635=>"000010000",
  55636=>"001011111",
  55637=>"110101100",
  55638=>"101010011",
  55639=>"100010100",
  55640=>"110101010",
  55641=>"000000011",
  55642=>"001000001",
  55643=>"101110101",
  55644=>"111110111",
  55645=>"001100100",
  55646=>"101010011",
  55647=>"000011100",
  55648=>"000000101",
  55649=>"101000010",
  55650=>"011001111",
  55651=>"000011010",
  55652=>"111001010",
  55653=>"001001010",
  55654=>"101110010",
  55655=>"000001010",
  55656=>"100010001",
  55657=>"101101111",
  55658=>"101001010",
  55659=>"101011110",
  55660=>"010111111",
  55661=>"101001100",
  55662=>"101101110",
  55663=>"000100001",
  55664=>"110100011",
  55665=>"011000001",
  55666=>"100011011",
  55667=>"000011000",
  55668=>"110111000",
  55669=>"101001101",
  55670=>"110011011",
  55671=>"000111111",
  55672=>"101110100",
  55673=>"000011111",
  55674=>"000100110",
  55675=>"111001001",
  55676=>"010101011",
  55677=>"001101000",
  55678=>"110101111",
  55679=>"110001111",
  55680=>"100100101",
  55681=>"111101100",
  55682=>"101110100",
  55683=>"000000111",
  55684=>"010001100",
  55685=>"100111011",
  55686=>"100110110",
  55687=>"010111000",
  55688=>"101011000",
  55689=>"000110111",
  55690=>"011011011",
  55691=>"011101010",
  55692=>"100001001",
  55693=>"100100111",
  55694=>"011100011",
  55695=>"010011111",
  55696=>"100100000",
  55697=>"111000001",
  55698=>"101100011",
  55699=>"111110101",
  55700=>"111010100",
  55701=>"111101011",
  55702=>"101010001",
  55703=>"100011100",
  55704=>"101111100",
  55705=>"000000101",
  55706=>"110000100",
  55707=>"000100000",
  55708=>"111111001",
  55709=>"111110101",
  55710=>"010000101",
  55711=>"011000100",
  55712=>"100110000",
  55713=>"001100111",
  55714=>"011110110",
  55715=>"010100010",
  55716=>"110110011",
  55717=>"011000101",
  55718=>"011110100",
  55719=>"100101011",
  55720=>"100110110",
  55721=>"010111100",
  55722=>"011010000",
  55723=>"010100111",
  55724=>"010011011",
  55725=>"001101110",
  55726=>"101000001",
  55727=>"000000101",
  55728=>"111011000",
  55729=>"101111100",
  55730=>"000110000",
  55731=>"101100001",
  55732=>"110100100",
  55733=>"110111010",
  55734=>"001100010",
  55735=>"001110010",
  55736=>"010001001",
  55737=>"101001011",
  55738=>"001101001",
  55739=>"001101111",
  55740=>"111111010",
  55741=>"110100110",
  55742=>"101001001",
  55743=>"110010001",
  55744=>"000000001",
  55745=>"110000111",
  55746=>"011001110",
  55747=>"001100010",
  55748=>"100010001",
  55749=>"111100010",
  55750=>"110110111",
  55751=>"100000010",
  55752=>"110000011",
  55753=>"000010110",
  55754=>"110000100",
  55755=>"010111000",
  55756=>"000011101",
  55757=>"000000010",
  55758=>"111111100",
  55759=>"100010001",
  55760=>"111010101",
  55761=>"111000101",
  55762=>"000110110",
  55763=>"000011101",
  55764=>"010011110",
  55765=>"010100111",
  55766=>"011011011",
  55767=>"011001100",
  55768=>"001101101",
  55769=>"100101011",
  55770=>"101010100",
  55771=>"011100111",
  55772=>"011001000",
  55773=>"010100100",
  55774=>"100010110",
  55775=>"110000000",
  55776=>"111010010",
  55777=>"101111011",
  55778=>"011110010",
  55779=>"011110000",
  55780=>"111000101",
  55781=>"001011100",
  55782=>"000111101",
  55783=>"101001101",
  55784=>"010100101",
  55785=>"001110101",
  55786=>"101000000",
  55787=>"100100100",
  55788=>"001100100",
  55789=>"001100100",
  55790=>"011100001",
  55791=>"010110011",
  55792=>"110010101",
  55793=>"100111000",
  55794=>"100000000",
  55795=>"111100110",
  55796=>"111111111",
  55797=>"000011100",
  55798=>"010001110",
  55799=>"000000001",
  55800=>"101010111",
  55801=>"110111011",
  55802=>"010010000",
  55803=>"101100110",
  55804=>"111100101",
  55805=>"001000000",
  55806=>"111010010",
  55807=>"000000010",
  55808=>"010010001",
  55809=>"010100001",
  55810=>"001110000",
  55811=>"001110100",
  55812=>"000011000",
  55813=>"000011100",
  55814=>"010101010",
  55815=>"011101100",
  55816=>"100101001",
  55817=>"000100000",
  55818=>"100101100",
  55819=>"010000001",
  55820=>"010111110",
  55821=>"100001000",
  55822=>"010011010",
  55823=>"111111001",
  55824=>"000001100",
  55825=>"010001101",
  55826=>"011110100",
  55827=>"111011111",
  55828=>"010010000",
  55829=>"111010111",
  55830=>"010100011",
  55831=>"111100010",
  55832=>"000000101",
  55833=>"001100010",
  55834=>"011001100",
  55835=>"011011111",
  55836=>"011001000",
  55837=>"001100110",
  55838=>"000011010",
  55839=>"000110100",
  55840=>"000010111",
  55841=>"010000001",
  55842=>"110011010",
  55843=>"101100010",
  55844=>"011001111",
  55845=>"110001111",
  55846=>"101011100",
  55847=>"101010110",
  55848=>"110101010",
  55849=>"110100001",
  55850=>"000000000",
  55851=>"010100101",
  55852=>"110011000",
  55853=>"010011011",
  55854=>"101101101",
  55855=>"000101000",
  55856=>"000111011",
  55857=>"111001100",
  55858=>"010001101",
  55859=>"001010101",
  55860=>"101010001",
  55861=>"110101011",
  55862=>"101010001",
  55863=>"000001010",
  55864=>"111111101",
  55865=>"000001001",
  55866=>"010000101",
  55867=>"000101000",
  55868=>"001000111",
  55869=>"110111111",
  55870=>"100011101",
  55871=>"100010101",
  55872=>"011110001",
  55873=>"011110000",
  55874=>"110101001",
  55875=>"001011111",
  55876=>"011011111",
  55877=>"001001100",
  55878=>"001000010",
  55879=>"101011011",
  55880=>"011111000",
  55881=>"010000011",
  55882=>"110111100",
  55883=>"110011001",
  55884=>"001011000",
  55885=>"101100101",
  55886=>"110000110",
  55887=>"110011010",
  55888=>"010001011",
  55889=>"011011010",
  55890=>"101100100",
  55891=>"011010001",
  55892=>"000110111",
  55893=>"000000000",
  55894=>"100100011",
  55895=>"001101000",
  55896=>"010001110",
  55897=>"100111000",
  55898=>"010111110",
  55899=>"010000101",
  55900=>"110100001",
  55901=>"000000000",
  55902=>"011001011",
  55903=>"110000111",
  55904=>"111101000",
  55905=>"010010001",
  55906=>"111100011",
  55907=>"000100001",
  55908=>"001100010",
  55909=>"111110011",
  55910=>"110001011",
  55911=>"101001100",
  55912=>"000111011",
  55913=>"011001001",
  55914=>"110101010",
  55915=>"011100110",
  55916=>"110100011",
  55917=>"111011100",
  55918=>"111111001",
  55919=>"001011101",
  55920=>"001100001",
  55921=>"000011000",
  55922=>"111101011",
  55923=>"101100000",
  55924=>"111010011",
  55925=>"010111110",
  55926=>"110011010",
  55927=>"001110001",
  55928=>"110010110",
  55929=>"101111001",
  55930=>"100100111",
  55931=>"101111000",
  55932=>"001100111",
  55933=>"011110000",
  55934=>"000000011",
  55935=>"111001011",
  55936=>"011011010",
  55937=>"011001000",
  55938=>"111000000",
  55939=>"100110010",
  55940=>"101001001",
  55941=>"011111101",
  55942=>"110001101",
  55943=>"100100111",
  55944=>"000101111",
  55945=>"011100001",
  55946=>"110011100",
  55947=>"010111101",
  55948=>"100100000",
  55949=>"101100111",
  55950=>"110100110",
  55951=>"010011101",
  55952=>"110000101",
  55953=>"011010000",
  55954=>"000110011",
  55955=>"110111110",
  55956=>"010110111",
  55957=>"100011010",
  55958=>"000001010",
  55959=>"011110110",
  55960=>"000010010",
  55961=>"001110101",
  55962=>"111000110",
  55963=>"011011001",
  55964=>"000101000",
  55965=>"011110110",
  55966=>"110011101",
  55967=>"111010011",
  55968=>"011110010",
  55969=>"001101101",
  55970=>"111000100",
  55971=>"010101010",
  55972=>"101110100",
  55973=>"110000010",
  55974=>"011110101",
  55975=>"010111110",
  55976=>"100100001",
  55977=>"011100000",
  55978=>"101110000",
  55979=>"101011111",
  55980=>"010000110",
  55981=>"001001110",
  55982=>"011010001",
  55983=>"101101111",
  55984=>"000101101",
  55985=>"001100110",
  55986=>"010011001",
  55987=>"101101000",
  55988=>"111111110",
  55989=>"111000111",
  55990=>"000010001",
  55991=>"011110101",
  55992=>"111110011",
  55993=>"101101101",
  55994=>"010100001",
  55995=>"100111011",
  55996=>"100110011",
  55997=>"010010010",
  55998=>"101001111",
  55999=>"100010100",
  56000=>"010011001",
  56001=>"010111101",
  56002=>"111111010",
  56003=>"100111111",
  56004=>"111001000",
  56005=>"011111000",
  56006=>"011110111",
  56007=>"110100000",
  56008=>"010110010",
  56009=>"100000011",
  56010=>"011010101",
  56011=>"011000100",
  56012=>"001011110",
  56013=>"101101111",
  56014=>"101111000",
  56015=>"111111111",
  56016=>"011001100",
  56017=>"011110101",
  56018=>"010110111",
  56019=>"000000111",
  56020=>"100101110",
  56021=>"101110000",
  56022=>"101111010",
  56023=>"010000000",
  56024=>"000101001",
  56025=>"010000011",
  56026=>"111000101",
  56027=>"110001011",
  56028=>"101001011",
  56029=>"110111000",
  56030=>"111001111",
  56031=>"001000011",
  56032=>"100011101",
  56033=>"111000111",
  56034=>"000010110",
  56035=>"111000101",
  56036=>"000111001",
  56037=>"110001100",
  56038=>"101001000",
  56039=>"010000010",
  56040=>"100010000",
  56041=>"010010000",
  56042=>"101011001",
  56043=>"001100000",
  56044=>"000000111",
  56045=>"010111110",
  56046=>"111111101",
  56047=>"110101001",
  56048=>"011010010",
  56049=>"111001010",
  56050=>"101100010",
  56051=>"001100010",
  56052=>"011011001",
  56053=>"101000110",
  56054=>"000100101",
  56055=>"010010000",
  56056=>"100110000",
  56057=>"110101011",
  56058=>"110010110",
  56059=>"110010000",
  56060=>"010100101",
  56061=>"111100101",
  56062=>"101001000",
  56063=>"101010101",
  56064=>"000111101",
  56065=>"000100110",
  56066=>"010011110",
  56067=>"000011011",
  56068=>"100101101",
  56069=>"100111010",
  56070=>"110101000",
  56071=>"010011111",
  56072=>"100110110",
  56073=>"000111010",
  56074=>"101001011",
  56075=>"101100111",
  56076=>"101001011",
  56077=>"010010111",
  56078=>"101111101",
  56079=>"110111111",
  56080=>"111011100",
  56081=>"100010111",
  56082=>"000101001",
  56083=>"010100100",
  56084=>"010101010",
  56085=>"010001000",
  56086=>"000101001",
  56087=>"110101000",
  56088=>"100100110",
  56089=>"010000111",
  56090=>"001101100",
  56091=>"100110001",
  56092=>"010110000",
  56093=>"000010100",
  56094=>"111101001",
  56095=>"100001111",
  56096=>"000000010",
  56097=>"110001100",
  56098=>"100100111",
  56099=>"111111000",
  56100=>"010011010",
  56101=>"000000000",
  56102=>"100011111",
  56103=>"010100111",
  56104=>"000100011",
  56105=>"010010000",
  56106=>"001010001",
  56107=>"000110001",
  56108=>"110010001",
  56109=>"000011001",
  56110=>"101111111",
  56111=>"111100100",
  56112=>"010001111",
  56113=>"001110001",
  56114=>"010110000",
  56115=>"010011000",
  56116=>"011001011",
  56117=>"000100000",
  56118=>"111010010",
  56119=>"000011001",
  56120=>"001100000",
  56121=>"011000000",
  56122=>"010011111",
  56123=>"011001000",
  56124=>"001100010",
  56125=>"101100011",
  56126=>"100010100",
  56127=>"100101100",
  56128=>"000100001",
  56129=>"101011100",
  56130=>"001111000",
  56131=>"000100110",
  56132=>"001111001",
  56133=>"001101001",
  56134=>"110010000",
  56135=>"100000100",
  56136=>"110001011",
  56137=>"000101001",
  56138=>"001110101",
  56139=>"110101010",
  56140=>"101111111",
  56141=>"110110100",
  56142=>"110010011",
  56143=>"011010001",
  56144=>"000011011",
  56145=>"001101110",
  56146=>"000100001",
  56147=>"000001000",
  56148=>"000011000",
  56149=>"110010010",
  56150=>"000010011",
  56151=>"101010011",
  56152=>"011111111",
  56153=>"011001000",
  56154=>"010001110",
  56155=>"000110101",
  56156=>"101100001",
  56157=>"101010011",
  56158=>"011110111",
  56159=>"110110000",
  56160=>"100001001",
  56161=>"110010100",
  56162=>"101111100",
  56163=>"111100010",
  56164=>"010100001",
  56165=>"001001000",
  56166=>"111000101",
  56167=>"111011101",
  56168=>"100000001",
  56169=>"001011000",
  56170=>"001000101",
  56171=>"010010000",
  56172=>"101101101",
  56173=>"001111010",
  56174=>"110000101",
  56175=>"011010101",
  56176=>"101110101",
  56177=>"001011101",
  56178=>"110110010",
  56179=>"110111111",
  56180=>"100110100",
  56181=>"000010000",
  56182=>"000010100",
  56183=>"011011000",
  56184=>"111101001",
  56185=>"010100100",
  56186=>"111101000",
  56187=>"011000011",
  56188=>"001111001",
  56189=>"110101100",
  56190=>"011110000",
  56191=>"110010011",
  56192=>"100111110",
  56193=>"101101000",
  56194=>"001000101",
  56195=>"000101011",
  56196=>"010101011",
  56197=>"101000110",
  56198=>"101101100",
  56199=>"000101011",
  56200=>"001101100",
  56201=>"101000101",
  56202=>"011100101",
  56203=>"001010000",
  56204=>"100001101",
  56205=>"011111000",
  56206=>"110111000",
  56207=>"100100110",
  56208=>"001010000",
  56209=>"111010101",
  56210=>"000001000",
  56211=>"001110011",
  56212=>"111100000",
  56213=>"001001110",
  56214=>"110110001",
  56215=>"011100101",
  56216=>"010100011",
  56217=>"000110101",
  56218=>"000111110",
  56219=>"100100110",
  56220=>"101101111",
  56221=>"000011010",
  56222=>"101111000",
  56223=>"001000011",
  56224=>"110101100",
  56225=>"000100001",
  56226=>"000001010",
  56227=>"000101010",
  56228=>"000111101",
  56229=>"111111001",
  56230=>"001011001",
  56231=>"010111101",
  56232=>"001111010",
  56233=>"100001110",
  56234=>"101011100",
  56235=>"111001011",
  56236=>"110101001",
  56237=>"000001001",
  56238=>"111101001",
  56239=>"001110010",
  56240=>"000001111",
  56241=>"110000000",
  56242=>"001010100",
  56243=>"101010101",
  56244=>"010011100",
  56245=>"100011011",
  56246=>"011010011",
  56247=>"111111000",
  56248=>"111011001",
  56249=>"000011110",
  56250=>"100111111",
  56251=>"011111011",
  56252=>"101000111",
  56253=>"111011000",
  56254=>"001100111",
  56255=>"111111000",
  56256=>"110101010",
  56257=>"101101100",
  56258=>"000000111",
  56259=>"101001110",
  56260=>"001101000",
  56261=>"011001100",
  56262=>"101100100",
  56263=>"011000000",
  56264=>"010011101",
  56265=>"110100100",
  56266=>"111011100",
  56267=>"101000000",
  56268=>"101000110",
  56269=>"000101100",
  56270=>"010111111",
  56271=>"101101101",
  56272=>"110101010",
  56273=>"100010000",
  56274=>"001000100",
  56275=>"010010111",
  56276=>"010100001",
  56277=>"110101101",
  56278=>"111111110",
  56279=>"001100111",
  56280=>"010001001",
  56281=>"110001011",
  56282=>"011100010",
  56283=>"110000001",
  56284=>"001011000",
  56285=>"101011000",
  56286=>"100111101",
  56287=>"000100001",
  56288=>"001000011",
  56289=>"001010000",
  56290=>"000011000",
  56291=>"001010000",
  56292=>"000001010",
  56293=>"011110011",
  56294=>"111000100",
  56295=>"000110011",
  56296=>"110000111",
  56297=>"000000101",
  56298=>"001000010",
  56299=>"111111010",
  56300=>"111100000",
  56301=>"100000010",
  56302=>"000000000",
  56303=>"011001101",
  56304=>"010000011",
  56305=>"110011001",
  56306=>"101111111",
  56307=>"000011010",
  56308=>"011100000",
  56309=>"011000001",
  56310=>"110011111",
  56311=>"000000011",
  56312=>"110010100",
  56313=>"011000010",
  56314=>"000010011",
  56315=>"100010000",
  56316=>"000101000",
  56317=>"110011011",
  56318=>"110000100",
  56319=>"110110011",
  56320=>"000100101",
  56321=>"000110110",
  56322=>"011001001",
  56323=>"100011111",
  56324=>"101000000",
  56325=>"101000111",
  56326=>"010010110",
  56327=>"011100111",
  56328=>"101110111",
  56329=>"010100101",
  56330=>"011010000",
  56331=>"100010011",
  56332=>"001000001",
  56333=>"000111101",
  56334=>"110011000",
  56335=>"001000001",
  56336=>"100000001",
  56337=>"011100000",
  56338=>"110000001",
  56339=>"001000000",
  56340=>"000010110",
  56341=>"111000000",
  56342=>"101110010",
  56343=>"111010101",
  56344=>"110101110",
  56345=>"110011100",
  56346=>"011011110",
  56347=>"100110111",
  56348=>"100100001",
  56349=>"100100110",
  56350=>"001000100",
  56351=>"011110010",
  56352=>"010011110",
  56353=>"100111110",
  56354=>"110110110",
  56355=>"101011110",
  56356=>"101001001",
  56357=>"011110110",
  56358=>"010000001",
  56359=>"100011111",
  56360=>"101101010",
  56361=>"110111101",
  56362=>"110011110",
  56363=>"101111100",
  56364=>"001110100",
  56365=>"001011100",
  56366=>"110111100",
  56367=>"010111001",
  56368=>"100000100",
  56369=>"101100001",
  56370=>"110100001",
  56371=>"000100001",
  56372=>"100010110",
  56373=>"010000000",
  56374=>"001000100",
  56375=>"111001110",
  56376=>"111001101",
  56377=>"110000101",
  56378=>"010001100",
  56379=>"011110111",
  56380=>"010000000",
  56381=>"001000110",
  56382=>"000100101",
  56383=>"001001101",
  56384=>"100111000",
  56385=>"011001100",
  56386=>"111000001",
  56387=>"110001101",
  56388=>"011011000",
  56389=>"110100000",
  56390=>"110110011",
  56391=>"111011001",
  56392=>"001001101",
  56393=>"110111010",
  56394=>"001111110",
  56395=>"011100011",
  56396=>"111111100",
  56397=>"100110100",
  56398=>"010101010",
  56399=>"101101000",
  56400=>"010111000",
  56401=>"100010100",
  56402=>"010101011",
  56403=>"111001001",
  56404=>"000000011",
  56405=>"110011100",
  56406=>"011011010",
  56407=>"011110010",
  56408=>"110101111",
  56409=>"000001011",
  56410=>"101001110",
  56411=>"110000001",
  56412=>"100011000",
  56413=>"001001100",
  56414=>"000011000",
  56415=>"111111110",
  56416=>"010001000",
  56417=>"010001010",
  56418=>"001010101",
  56419=>"001010011",
  56420=>"001001010",
  56421=>"001001101",
  56422=>"000000111",
  56423=>"001100101",
  56424=>"011111100",
  56425=>"101011110",
  56426=>"110110100",
  56427=>"110100010",
  56428=>"000001000",
  56429=>"000001011",
  56430=>"110111000",
  56431=>"000111001",
  56432=>"100000110",
  56433=>"111000011",
  56434=>"000011000",
  56435=>"110101111",
  56436=>"001110001",
  56437=>"001011110",
  56438=>"001100110",
  56439=>"010011110",
  56440=>"000111011",
  56441=>"111011110",
  56442=>"011111100",
  56443=>"011010111",
  56444=>"111110110",
  56445=>"010101110",
  56446=>"010110000",
  56447=>"011010001",
  56448=>"011001001",
  56449=>"011001110",
  56450=>"011110011",
  56451=>"011011000",
  56452=>"011010100",
  56453=>"010100110",
  56454=>"111111000",
  56455=>"011011111",
  56456=>"111000011",
  56457=>"011111101",
  56458=>"011110010",
  56459=>"000101001",
  56460=>"011100011",
  56461=>"111100111",
  56462=>"000001001",
  56463=>"011011111",
  56464=>"111001011",
  56465=>"000110010",
  56466=>"111111111",
  56467=>"000111000",
  56468=>"000101000",
  56469=>"100100101",
  56470=>"010111011",
  56471=>"001000000",
  56472=>"111000111",
  56473=>"111110000",
  56474=>"111111011",
  56475=>"001101011",
  56476=>"010111001",
  56477=>"101000010",
  56478=>"110101111",
  56479=>"000000011",
  56480=>"001110101",
  56481=>"011001001",
  56482=>"111101100",
  56483=>"100110010",
  56484=>"101110111",
  56485=>"101100000",
  56486=>"111010001",
  56487=>"111011100",
  56488=>"100011100",
  56489=>"100100000",
  56490=>"110110011",
  56491=>"000011101",
  56492=>"001100100",
  56493=>"000011000",
  56494=>"110110000",
  56495=>"110000001",
  56496=>"001100100",
  56497=>"111011010",
  56498=>"110110001",
  56499=>"001000000",
  56500=>"010000011",
  56501=>"111001010",
  56502=>"110000001",
  56503=>"111111011",
  56504=>"000001001",
  56505=>"000100010",
  56506=>"101110100",
  56507=>"101011001",
  56508=>"100011110",
  56509=>"000000010",
  56510=>"010111001",
  56511=>"001010000",
  56512=>"110110011",
  56513=>"110101010",
  56514=>"101111011",
  56515=>"100111010",
  56516=>"000110100",
  56517=>"001100001",
  56518=>"001000110",
  56519=>"110100011",
  56520=>"011000010",
  56521=>"101011111",
  56522=>"110011001",
  56523=>"011110110",
  56524=>"100011111",
  56525=>"111011110",
  56526=>"011000010",
  56527=>"000100001",
  56528=>"101110000",
  56529=>"010001001",
  56530=>"011100100",
  56531=>"001001111",
  56532=>"101101011",
  56533=>"100111000",
  56534=>"100100101",
  56535=>"000011101",
  56536=>"101111101",
  56537=>"111100110",
  56538=>"001010111",
  56539=>"010001110",
  56540=>"111101111",
  56541=>"100001001",
  56542=>"011000001",
  56543=>"000011011",
  56544=>"110001110",
  56545=>"010000100",
  56546=>"111001111",
  56547=>"010011010",
  56548=>"101101001",
  56549=>"000111000",
  56550=>"101111111",
  56551=>"000001001",
  56552=>"111101110",
  56553=>"111111100",
  56554=>"011101010",
  56555=>"001011001",
  56556=>"100011101",
  56557=>"111100000",
  56558=>"110110010",
  56559=>"101111110",
  56560=>"111001111",
  56561=>"000100111",
  56562=>"011010011",
  56563=>"101001101",
  56564=>"001001101",
  56565=>"101111110",
  56566=>"111110110",
  56567=>"011001101",
  56568=>"111111010",
  56569=>"001111000",
  56570=>"010111011",
  56571=>"110000000",
  56572=>"100000110",
  56573=>"000001111",
  56574=>"011010001",
  56575=>"101101000",
  56576=>"100010011",
  56577=>"000010110",
  56578=>"100111010",
  56579=>"001011011",
  56580=>"101011110",
  56581=>"000000110",
  56582=>"001011101",
  56583=>"111110011",
  56584=>"011111111",
  56585=>"111110101",
  56586=>"101111100",
  56587=>"111010010",
  56588=>"000101100",
  56589=>"110110100",
  56590=>"010001000",
  56591=>"110010011",
  56592=>"111011000",
  56593=>"101000010",
  56594=>"001001001",
  56595=>"010110111",
  56596=>"000101100",
  56597=>"111001001",
  56598=>"100000110",
  56599=>"001010110",
  56600=>"001011101",
  56601=>"000100000",
  56602=>"100111111",
  56603=>"101001010",
  56604=>"101101001",
  56605=>"000111000",
  56606=>"101100111",
  56607=>"011001000",
  56608=>"000000000",
  56609=>"011100101",
  56610=>"110101011",
  56611=>"101101010",
  56612=>"001111100",
  56613=>"110110100",
  56614=>"100001101",
  56615=>"000101100",
  56616=>"000000100",
  56617=>"011110110",
  56618=>"000011000",
  56619=>"110011100",
  56620=>"111111110",
  56621=>"111101000",
  56622=>"111010010",
  56623=>"111000110",
  56624=>"011001101",
  56625=>"111111000",
  56626=>"111110010",
  56627=>"111010011",
  56628=>"011100100",
  56629=>"011010010",
  56630=>"100001101",
  56631=>"000110011",
  56632=>"000110111",
  56633=>"011001011",
  56634=>"000011101",
  56635=>"110110000",
  56636=>"000011101",
  56637=>"100100000",
  56638=>"100001010",
  56639=>"110001000",
  56640=>"101001010",
  56641=>"111010110",
  56642=>"100100000",
  56643=>"101000001",
  56644=>"111010010",
  56645=>"001010110",
  56646=>"110010010",
  56647=>"011110010",
  56648=>"101100100",
  56649=>"110000011",
  56650=>"011101111",
  56651=>"101101101",
  56652=>"000110101",
  56653=>"100110100",
  56654=>"110011001",
  56655=>"100100010",
  56656=>"000000000",
  56657=>"011101011",
  56658=>"011110000",
  56659=>"000011001",
  56660=>"001111110",
  56661=>"111011010",
  56662=>"010111101",
  56663=>"000000110",
  56664=>"110111011",
  56665=>"101100000",
  56666=>"111001101",
  56667=>"001011000",
  56668=>"010010111",
  56669=>"001101111",
  56670=>"000010000",
  56671=>"110000011",
  56672=>"111000001",
  56673=>"111100011",
  56674=>"010010100",
  56675=>"000011001",
  56676=>"100101100",
  56677=>"001011011",
  56678=>"011101101",
  56679=>"011011000",
  56680=>"000000000",
  56681=>"101011001",
  56682=>"111100001",
  56683=>"000010100",
  56684=>"000001010",
  56685=>"101010110",
  56686=>"001110011",
  56687=>"010111011",
  56688=>"111011111",
  56689=>"101001100",
  56690=>"100000110",
  56691=>"111110000",
  56692=>"111011001",
  56693=>"001101100",
  56694=>"010001001",
  56695=>"101001111",
  56696=>"001011011",
  56697=>"001010001",
  56698=>"000000000",
  56699=>"000100110",
  56700=>"001001011",
  56701=>"000011111",
  56702=>"110111110",
  56703=>"000000010",
  56704=>"000111101",
  56705=>"010000100",
  56706=>"001000011",
  56707=>"010010010",
  56708=>"100111011",
  56709=>"010110001",
  56710=>"010000000",
  56711=>"110110001",
  56712=>"111100110",
  56713=>"101010011",
  56714=>"100000000",
  56715=>"001111011",
  56716=>"101010101",
  56717=>"000111001",
  56718=>"110110010",
  56719=>"001010000",
  56720=>"010101101",
  56721=>"001011010",
  56722=>"011101111",
  56723=>"110101110",
  56724=>"010111111",
  56725=>"010010101",
  56726=>"111100100",
  56727=>"110101011",
  56728=>"110010011",
  56729=>"001011000",
  56730=>"100101010",
  56731=>"111111110",
  56732=>"011111111",
  56733=>"111110111",
  56734=>"100100111",
  56735=>"111110111",
  56736=>"010100110",
  56737=>"111010000",
  56738=>"110010010",
  56739=>"001001011",
  56740=>"111101000",
  56741=>"010101101",
  56742=>"001000000",
  56743=>"111011101",
  56744=>"100001001",
  56745=>"001000000",
  56746=>"111101110",
  56747=>"010101010",
  56748=>"100000001",
  56749=>"010111100",
  56750=>"001100001",
  56751=>"111001011",
  56752=>"110010111",
  56753=>"000000011",
  56754=>"101111011",
  56755=>"100001111",
  56756=>"100111101",
  56757=>"101011101",
  56758=>"111001110",
  56759=>"010001110",
  56760=>"110110110",
  56761=>"101011101",
  56762=>"001010000",
  56763=>"010110100",
  56764=>"101110110",
  56765=>"010011011",
  56766=>"000110100",
  56767=>"000011000",
  56768=>"110101011",
  56769=>"101110110",
  56770=>"111110001",
  56771=>"001111111",
  56772=>"110111101",
  56773=>"000011011",
  56774=>"011111000",
  56775=>"011100111",
  56776=>"110010000",
  56777=>"001111011",
  56778=>"001101101",
  56779=>"101111110",
  56780=>"000001010",
  56781=>"000100111",
  56782=>"101101101",
  56783=>"011000110",
  56784=>"100010111",
  56785=>"100001010",
  56786=>"101011011",
  56787=>"011011101",
  56788=>"111111001",
  56789=>"100010111",
  56790=>"111000000",
  56791=>"110110011",
  56792=>"101001011",
  56793=>"101011001",
  56794=>"000110110",
  56795=>"101000001",
  56796=>"010000000",
  56797=>"101101000",
  56798=>"010010001",
  56799=>"011100101",
  56800=>"100100111",
  56801=>"011101111",
  56802=>"011101011",
  56803=>"111110100",
  56804=>"110100000",
  56805=>"010100110",
  56806=>"001000001",
  56807=>"011011101",
  56808=>"111101110",
  56809=>"011010000",
  56810=>"101101110",
  56811=>"111101001",
  56812=>"000010001",
  56813=>"010100000",
  56814=>"111100111",
  56815=>"100100011",
  56816=>"010000011",
  56817=>"000111001",
  56818=>"111011010",
  56819=>"111010110",
  56820=>"000100110",
  56821=>"111001011",
  56822=>"111000100",
  56823=>"000000111",
  56824=>"011010111",
  56825=>"111111111",
  56826=>"010010000",
  56827=>"100100010",
  56828=>"010101100",
  56829=>"110010110",
  56830=>"010101010",
  56831=>"000111110",
  56832=>"100011111",
  56833=>"110011110",
  56834=>"010000001",
  56835=>"000110100",
  56836=>"011111010",
  56837=>"101111100",
  56838=>"011001001",
  56839=>"101111111",
  56840=>"001101000",
  56841=>"000100101",
  56842=>"011100111",
  56843=>"111110001",
  56844=>"010100001",
  56845=>"011001111",
  56846=>"111100000",
  56847=>"000010101",
  56848=>"110101111",
  56849=>"011111001",
  56850=>"101100011",
  56851=>"110010001",
  56852=>"010110101",
  56853=>"011111000",
  56854=>"010011101",
  56855=>"001000000",
  56856=>"011010100",
  56857=>"100011011",
  56858=>"001111010",
  56859=>"010000111",
  56860=>"000000000",
  56861=>"111000011",
  56862=>"010010000",
  56863=>"001010001",
  56864=>"101101011",
  56865=>"111110000",
  56866=>"111100100",
  56867=>"011101110",
  56868=>"011001111",
  56869=>"111001101",
  56870=>"011000000",
  56871=>"010001000",
  56872=>"011111111",
  56873=>"000110000",
  56874=>"100000000",
  56875=>"111111110",
  56876=>"000001001",
  56877=>"011101001",
  56878=>"011100101",
  56879=>"111110101",
  56880=>"011100011",
  56881=>"000000100",
  56882=>"101100010",
  56883=>"000110110",
  56884=>"000110011",
  56885=>"001110101",
  56886=>"010011111",
  56887=>"101111010",
  56888=>"011101011",
  56889=>"011100010",
  56890=>"001000101",
  56891=>"101110000",
  56892=>"001101000",
  56893=>"101100110",
  56894=>"101011000",
  56895=>"110100111",
  56896=>"001100010",
  56897=>"111000100",
  56898=>"001111011",
  56899=>"001001000",
  56900=>"100101101",
  56901=>"010100000",
  56902=>"000100010",
  56903=>"000010000",
  56904=>"000100010",
  56905=>"000001100",
  56906=>"000011000",
  56907=>"010001111",
  56908=>"011101010",
  56909=>"100101001",
  56910=>"100000010",
  56911=>"010111010",
  56912=>"001000001",
  56913=>"110100100",
  56914=>"110111111",
  56915=>"110001001",
  56916=>"000001110",
  56917=>"000000101",
  56918=>"000110100",
  56919=>"000011100",
  56920=>"111111010",
  56921=>"100010010",
  56922=>"010000110",
  56923=>"010110100",
  56924=>"000000000",
  56925=>"111011111",
  56926=>"001110011",
  56927=>"001100100",
  56928=>"100110001",
  56929=>"011011101",
  56930=>"000101111",
  56931=>"110000110",
  56932=>"100111010",
  56933=>"010111011",
  56934=>"101000100",
  56935=>"000000010",
  56936=>"000101000",
  56937=>"100101111",
  56938=>"100011011",
  56939=>"100010001",
  56940=>"111010100",
  56941=>"010111011",
  56942=>"101110011",
  56943=>"100011000",
  56944=>"011111010",
  56945=>"010000000",
  56946=>"010000010",
  56947=>"011001100",
  56948=>"000110100",
  56949=>"001000101",
  56950=>"101011111",
  56951=>"011000101",
  56952=>"100001111",
  56953=>"000101100",
  56954=>"011010111",
  56955=>"010010010",
  56956=>"010011001",
  56957=>"110101101",
  56958=>"001101100",
  56959=>"000010111",
  56960=>"000100111",
  56961=>"001101100",
  56962=>"110001101",
  56963=>"011000101",
  56964=>"001111100",
  56965=>"000000100",
  56966=>"101000101",
  56967=>"110001010",
  56968=>"000010000",
  56969=>"111111110",
  56970=>"100100000",
  56971=>"110111000",
  56972=>"110110001",
  56973=>"110011001",
  56974=>"110111111",
  56975=>"001000000",
  56976=>"111111110",
  56977=>"111000000",
  56978=>"111000000",
  56979=>"001001010",
  56980=>"101001100",
  56981=>"110100100",
  56982=>"100111101",
  56983=>"000001001",
  56984=>"000000100",
  56985=>"111100001",
  56986=>"110101111",
  56987=>"110101101",
  56988=>"111001101",
  56989=>"101101011",
  56990=>"111111000",
  56991=>"101001000",
  56992=>"100111111",
  56993=>"011011111",
  56994=>"011101011",
  56995=>"010010110",
  56996=>"001011001",
  56997=>"001110000",
  56998=>"011011001",
  56999=>"000001010",
  57000=>"000100101",
  57001=>"101000100",
  57002=>"111001110",
  57003=>"100011000",
  57004=>"100001000",
  57005=>"101011010",
  57006=>"101010101",
  57007=>"010010111",
  57008=>"100101110",
  57009=>"010010000",
  57010=>"011101110",
  57011=>"010010111",
  57012=>"000110001",
  57013=>"110111110",
  57014=>"011111010",
  57015=>"100011011",
  57016=>"110100111",
  57017=>"101110100",
  57018=>"010001010",
  57019=>"000011110",
  57020=>"101101100",
  57021=>"011000001",
  57022=>"111001111",
  57023=>"100101101",
  57024=>"011111010",
  57025=>"000010101",
  57026=>"010101101",
  57027=>"011001110",
  57028=>"110111000",
  57029=>"010111010",
  57030=>"101110110",
  57031=>"011000100",
  57032=>"010011011",
  57033=>"010001110",
  57034=>"101001110",
  57035=>"010011000",
  57036=>"000101010",
  57037=>"101100111",
  57038=>"001100110",
  57039=>"000001000",
  57040=>"001000001",
  57041=>"000011100",
  57042=>"010000101",
  57043=>"010011001",
  57044=>"000010010",
  57045=>"011100010",
  57046=>"000010010",
  57047=>"110000110",
  57048=>"101001101",
  57049=>"100011110",
  57050=>"100010001",
  57051=>"100100101",
  57052=>"111110011",
  57053=>"001101111",
  57054=>"000100011",
  57055=>"111101010",
  57056=>"110010001",
  57057=>"111111111",
  57058=>"010110101",
  57059=>"111001001",
  57060=>"110001100",
  57061=>"001111000",
  57062=>"001010100",
  57063=>"101000110",
  57064=>"000110101",
  57065=>"001111001",
  57066=>"001110011",
  57067=>"101111000",
  57068=>"000110111",
  57069=>"010000011",
  57070=>"101000000",
  57071=>"001000001",
  57072=>"011100010",
  57073=>"000000011",
  57074=>"011111000",
  57075=>"001010011",
  57076=>"011100111",
  57077=>"010011101",
  57078=>"111001000",
  57079=>"101110100",
  57080=>"101000010",
  57081=>"000100100",
  57082=>"000000110",
  57083=>"111000101",
  57084=>"011010100",
  57085=>"101101001",
  57086=>"101101100",
  57087=>"000111110",
  57088=>"111001100",
  57089=>"111001111",
  57090=>"110100011",
  57091=>"101000001",
  57092=>"010101101",
  57093=>"101111111",
  57094=>"000101111",
  57095=>"101110110",
  57096=>"111101001",
  57097=>"111010110",
  57098=>"100101110",
  57099=>"010101010",
  57100=>"001110100",
  57101=>"111000100",
  57102=>"000001110",
  57103=>"011001010",
  57104=>"001001110",
  57105=>"110011111",
  57106=>"010000010",
  57107=>"010101110",
  57108=>"001101011",
  57109=>"101111010",
  57110=>"001101000",
  57111=>"100111100",
  57112=>"001101100",
  57113=>"000110011",
  57114=>"010000100",
  57115=>"001010110",
  57116=>"101110000",
  57117=>"011001001",
  57118=>"000001001",
  57119=>"000101001",
  57120=>"001000001",
  57121=>"010001111",
  57122=>"000011000",
  57123=>"000110001",
  57124=>"010101011",
  57125=>"101011010",
  57126=>"100101011",
  57127=>"100110010",
  57128=>"110100001",
  57129=>"000000101",
  57130=>"111000101",
  57131=>"110000001",
  57132=>"000111001",
  57133=>"111000011",
  57134=>"001111011",
  57135=>"011000000",
  57136=>"100100100",
  57137=>"010111111",
  57138=>"000010110",
  57139=>"001001111",
  57140=>"111011110",
  57141=>"100001100",
  57142=>"100010100",
  57143=>"110111001",
  57144=>"110001111",
  57145=>"000101001",
  57146=>"101101000",
  57147=>"001100011",
  57148=>"100101101",
  57149=>"100000001",
  57150=>"110010101",
  57151=>"000000111",
  57152=>"000100100",
  57153=>"011100100",
  57154=>"101110000",
  57155=>"111010001",
  57156=>"000001000",
  57157=>"000000001",
  57158=>"110111100",
  57159=>"011111110",
  57160=>"100110000",
  57161=>"111000100",
  57162=>"010011110",
  57163=>"011000110",
  57164=>"001010110",
  57165=>"101110010",
  57166=>"100011101",
  57167=>"011000110",
  57168=>"000101101",
  57169=>"101011011",
  57170=>"111010000",
  57171=>"000001101",
  57172=>"001100001",
  57173=>"001001110",
  57174=>"000101111",
  57175=>"101010000",
  57176=>"111111010",
  57177=>"111001111",
  57178=>"010001110",
  57179=>"011011000",
  57180=>"101100010",
  57181=>"111111101",
  57182=>"001001000",
  57183=>"100010101",
  57184=>"110000010",
  57185=>"100110000",
  57186=>"100001111",
  57187=>"000100000",
  57188=>"000100110",
  57189=>"110011110",
  57190=>"111111111",
  57191=>"100001011",
  57192=>"111111110",
  57193=>"100111011",
  57194=>"000010101",
  57195=>"001010001",
  57196=>"000000011",
  57197=>"101111101",
  57198=>"011010001",
  57199=>"000011101",
  57200=>"101000010",
  57201=>"010001101",
  57202=>"101110000",
  57203=>"000100110",
  57204=>"010101100",
  57205=>"000011011",
  57206=>"001000101",
  57207=>"110010011",
  57208=>"010011101",
  57209=>"100000010",
  57210=>"010110011",
  57211=>"010101001",
  57212=>"001111001",
  57213=>"100110011",
  57214=>"010000011",
  57215=>"010100001",
  57216=>"000110011",
  57217=>"110100111",
  57218=>"000100101",
  57219=>"001000001",
  57220=>"011000001",
  57221=>"110111111",
  57222=>"101000011",
  57223=>"010001100",
  57224=>"001000110",
  57225=>"110110000",
  57226=>"000001011",
  57227=>"010111011",
  57228=>"101101110",
  57229=>"101010111",
  57230=>"010110101",
  57231=>"000001101",
  57232=>"010111010",
  57233=>"001111001",
  57234=>"010001000",
  57235=>"010100011",
  57236=>"000001000",
  57237=>"011000000",
  57238=>"011010111",
  57239=>"001001011",
  57240=>"010011011",
  57241=>"101001101",
  57242=>"001110011",
  57243=>"100101111",
  57244=>"101110111",
  57245=>"011010101",
  57246=>"110111111",
  57247=>"001001010",
  57248=>"111111101",
  57249=>"110010101",
  57250=>"010001111",
  57251=>"111000000",
  57252=>"001000010",
  57253=>"110011111",
  57254=>"110100011",
  57255=>"111110111",
  57256=>"010001010",
  57257=>"100111000",
  57258=>"011111111",
  57259=>"100000011",
  57260=>"110001001",
  57261=>"000110011",
  57262=>"000011100",
  57263=>"101011100",
  57264=>"100110010",
  57265=>"000100000",
  57266=>"110001010",
  57267=>"111111111",
  57268=>"011111111",
  57269=>"001000111",
  57270=>"011101010",
  57271=>"001010110",
  57272=>"101010001",
  57273=>"100001000",
  57274=>"110001101",
  57275=>"000000110",
  57276=>"100010101",
  57277=>"000101001",
  57278=>"100110111",
  57279=>"001001111",
  57280=>"101111101",
  57281=>"000000111",
  57282=>"100111111",
  57283=>"101001010",
  57284=>"100000111",
  57285=>"100010111",
  57286=>"001001100",
  57287=>"111010110",
  57288=>"100010100",
  57289=>"101110001",
  57290=>"011010011",
  57291=>"100001011",
  57292=>"010111110",
  57293=>"100000001",
  57294=>"111000001",
  57295=>"011110000",
  57296=>"101100011",
  57297=>"010001110",
  57298=>"010111011",
  57299=>"101110010",
  57300=>"110001101",
  57301=>"001011101",
  57302=>"100010010",
  57303=>"010010101",
  57304=>"011110001",
  57305=>"010010100",
  57306=>"000010101",
  57307=>"010111011",
  57308=>"100101110",
  57309=>"001111101",
  57310=>"101101110",
  57311=>"101000101",
  57312=>"010001111",
  57313=>"011010000",
  57314=>"111010011",
  57315=>"001111011",
  57316=>"011100111",
  57317=>"111100111",
  57318=>"011110010",
  57319=>"100001110",
  57320=>"000000010",
  57321=>"110110110",
  57322=>"010010101",
  57323=>"010101011",
  57324=>"111111011",
  57325=>"100100111",
  57326=>"101011111",
  57327=>"001000000",
  57328=>"001111101",
  57329=>"101101100",
  57330=>"000010101",
  57331=>"011010101",
  57332=>"000000110",
  57333=>"001000111",
  57334=>"111101110",
  57335=>"000001111",
  57336=>"010101010",
  57337=>"000000010",
  57338=>"111101010",
  57339=>"001110011",
  57340=>"110001001",
  57341=>"010000111",
  57342=>"111110110",
  57343=>"010111111",
  57344=>"111001110",
  57345=>"110110111",
  57346=>"101101010",
  57347=>"111111000",
  57348=>"001001010",
  57349=>"001100101",
  57350=>"000001001",
  57351=>"001110111",
  57352=>"001111100",
  57353=>"100011101",
  57354=>"010001010",
  57355=>"100111100",
  57356=>"111110011",
  57357=>"100101110",
  57358=>"011100001",
  57359=>"111100111",
  57360=>"111010101",
  57361=>"101111101",
  57362=>"111001101",
  57363=>"010110101",
  57364=>"110000010",
  57365=>"001100101",
  57366=>"111011111",
  57367=>"101100011",
  57368=>"101100100",
  57369=>"100100100",
  57370=>"100101110",
  57371=>"010000101",
  57372=>"110100011",
  57373=>"011101101",
  57374=>"000000001",
  57375=>"001000000",
  57376=>"100111100",
  57377=>"011001110",
  57378=>"000001101",
  57379=>"110111000",
  57380=>"011110010",
  57381=>"000010110",
  57382=>"011000011",
  57383=>"100101011",
  57384=>"101001011",
  57385=>"000111110",
  57386=>"011100100",
  57387=>"111011110",
  57388=>"101110111",
  57389=>"100100100",
  57390=>"101101100",
  57391=>"100110100",
  57392=>"010010100",
  57393=>"100111001",
  57394=>"101000001",
  57395=>"100010011",
  57396=>"110110010",
  57397=>"101101101",
  57398=>"110110101",
  57399=>"110111010",
  57400=>"000000101",
  57401=>"110110100",
  57402=>"101000111",
  57403=>"101101010",
  57404=>"111101000",
  57405=>"101011101",
  57406=>"001111100",
  57407=>"011001110",
  57408=>"000101011",
  57409=>"101100001",
  57410=>"010111100",
  57411=>"000000001",
  57412=>"101010110",
  57413=>"000100001",
  57414=>"010000011",
  57415=>"011101101",
  57416=>"000100001",
  57417=>"110111101",
  57418=>"110110111",
  57419=>"111011101",
  57420=>"011000000",
  57421=>"110110000",
  57422=>"111000001",
  57423=>"000101100",
  57424=>"000100101",
  57425=>"110111000",
  57426=>"101001000",
  57427=>"000100101",
  57428=>"101100100",
  57429=>"000100000",
  57430=>"001111101",
  57431=>"001101111",
  57432=>"101110110",
  57433=>"000010001",
  57434=>"000100001",
  57435=>"100111011",
  57436=>"010111101",
  57437=>"001011000",
  57438=>"100000110",
  57439=>"010000110",
  57440=>"010001001",
  57441=>"111001010",
  57442=>"101001111",
  57443=>"010000100",
  57444=>"111000001",
  57445=>"011011110",
  57446=>"001100011",
  57447=>"010111000",
  57448=>"101100011",
  57449=>"011001000",
  57450=>"000010111",
  57451=>"010010000",
  57452=>"110100000",
  57453=>"000001101",
  57454=>"100110101",
  57455=>"111000110",
  57456=>"000100110",
  57457=>"011000001",
  57458=>"110101111",
  57459=>"001011010",
  57460=>"001110101",
  57461=>"111111101",
  57462=>"010001101",
  57463=>"001110111",
  57464=>"000100101",
  57465=>"001011011",
  57466=>"100111111",
  57467=>"100000000",
  57468=>"110101010",
  57469=>"011011111",
  57470=>"101011101",
  57471=>"110001010",
  57472=>"001001110",
  57473=>"101011011",
  57474=>"101110101",
  57475=>"111010111",
  57476=>"111100100",
  57477=>"100010110",
  57478=>"010010011",
  57479=>"111111111",
  57480=>"100110100",
  57481=>"011000011",
  57482=>"110001011",
  57483=>"101111111",
  57484=>"111011100",
  57485=>"011000101",
  57486=>"011011101",
  57487=>"101000000",
  57488=>"001011111",
  57489=>"011001101",
  57490=>"000011111",
  57491=>"011110111",
  57492=>"101110011",
  57493=>"110100000",
  57494=>"101011001",
  57495=>"100000010",
  57496=>"000010011",
  57497=>"110010010",
  57498=>"100011111",
  57499=>"101001011",
  57500=>"011100000",
  57501=>"110101111",
  57502=>"101100001",
  57503=>"001010111",
  57504=>"010011001",
  57505=>"110010100",
  57506=>"101100010",
  57507=>"101101110",
  57508=>"100111111",
  57509=>"010000011",
  57510=>"100111111",
  57511=>"000101100",
  57512=>"100100000",
  57513=>"100101101",
  57514=>"010011111",
  57515=>"000101111",
  57516=>"001100111",
  57517=>"010000000",
  57518=>"001010011",
  57519=>"111111001",
  57520=>"111100101",
  57521=>"111110110",
  57522=>"011111000",
  57523=>"111110010",
  57524=>"101101101",
  57525=>"011010001",
  57526=>"000001110",
  57527=>"010001101",
  57528=>"101001010",
  57529=>"011000000",
  57530=>"000100110",
  57531=>"101011001",
  57532=>"101010011",
  57533=>"000110000",
  57534=>"000110000",
  57535=>"011011110",
  57536=>"000111110",
  57537=>"011101111",
  57538=>"000101010",
  57539=>"011111000",
  57540=>"101111000",
  57541=>"010101110",
  57542=>"101100011",
  57543=>"101110111",
  57544=>"011111011",
  57545=>"100001111",
  57546=>"011001010",
  57547=>"111011011",
  57548=>"110001010",
  57549=>"000101111",
  57550=>"001110100",
  57551=>"001110111",
  57552=>"100101101",
  57553=>"011000101",
  57554=>"100110111",
  57555=>"101111110",
  57556=>"010000001",
  57557=>"000000001",
  57558=>"010100111",
  57559=>"000101010",
  57560=>"110110100",
  57561=>"101100100",
  57562=>"010101010",
  57563=>"100001011",
  57564=>"111111110",
  57565=>"100010110",
  57566=>"010110011",
  57567=>"001000101",
  57568=>"100000110",
  57569=>"101001011",
  57570=>"000100001",
  57571=>"100010111",
  57572=>"001000000",
  57573=>"111010110",
  57574=>"010100100",
  57575=>"010111101",
  57576=>"100001110",
  57577=>"111101000",
  57578=>"000100111",
  57579=>"000001110",
  57580=>"000101011",
  57581=>"000010100",
  57582=>"100101101",
  57583=>"010101111",
  57584=>"001001010",
  57585=>"011110100",
  57586=>"001011101",
  57587=>"101000110",
  57588=>"100010001",
  57589=>"000011000",
  57590=>"111101110",
  57591=>"100000001",
  57592=>"000010101",
  57593=>"111111000",
  57594=>"011010010",
  57595=>"101110111",
  57596=>"001100111",
  57597=>"110110101",
  57598=>"010101010",
  57599=>"111011011",
  57600=>"111011001",
  57601=>"101001111",
  57602=>"001110010",
  57603=>"100111000",
  57604=>"101100111",
  57605=>"001111100",
  57606=>"001110011",
  57607=>"111010000",
  57608=>"011111011",
  57609=>"011101111",
  57610=>"110010001",
  57611=>"000101101",
  57612=>"000111000",
  57613=>"001111011",
  57614=>"010100000",
  57615=>"100011111",
  57616=>"111101101",
  57617=>"100010011",
  57618=>"111100010",
  57619=>"111001011",
  57620=>"011000111",
  57621=>"011100100",
  57622=>"100001111",
  57623=>"101010110",
  57624=>"000001000",
  57625=>"010111110",
  57626=>"000010110",
  57627=>"111000101",
  57628=>"001011010",
  57629=>"010001000",
  57630=>"110100111",
  57631=>"000100100",
  57632=>"101001001",
  57633=>"011101000",
  57634=>"100000101",
  57635=>"100100101",
  57636=>"000111100",
  57637=>"111011011",
  57638=>"011010000",
  57639=>"100100111",
  57640=>"100000101",
  57641=>"111010011",
  57642=>"000100001",
  57643=>"010001001",
  57644=>"000100010",
  57645=>"110101100",
  57646=>"100101000",
  57647=>"111111111",
  57648=>"000101111",
  57649=>"101101000",
  57650=>"010101001",
  57651=>"110000001",
  57652=>"111110111",
  57653=>"010011101",
  57654=>"110000110",
  57655=>"010010010",
  57656=>"000000010",
  57657=>"101100111",
  57658=>"100010110",
  57659=>"110000000",
  57660=>"010011011",
  57661=>"110111010",
  57662=>"110101101",
  57663=>"000100111",
  57664=>"000111100",
  57665=>"100110111",
  57666=>"100110001",
  57667=>"011111010",
  57668=>"111001001",
  57669=>"100101011",
  57670=>"000001001",
  57671=>"101000101",
  57672=>"001000010",
  57673=>"010000010",
  57674=>"000101101",
  57675=>"101110011",
  57676=>"100100011",
  57677=>"001001111",
  57678=>"000010001",
  57679=>"011011010",
  57680=>"011010100",
  57681=>"111000001",
  57682=>"100010001",
  57683=>"100000110",
  57684=>"000100100",
  57685=>"110011001",
  57686=>"001000100",
  57687=>"001010100",
  57688=>"111101000",
  57689=>"100011011",
  57690=>"111001100",
  57691=>"000010010",
  57692=>"110010111",
  57693=>"001111111",
  57694=>"011111001",
  57695=>"010010111",
  57696=>"101001001",
  57697=>"011101101",
  57698=>"101101010",
  57699=>"010110100",
  57700=>"010010111",
  57701=>"010100101",
  57702=>"000010001",
  57703=>"110111001",
  57704=>"111100110",
  57705=>"000100001",
  57706=>"000001101",
  57707=>"011011001",
  57708=>"000001111",
  57709=>"011000000",
  57710=>"111100001",
  57711=>"000110001",
  57712=>"000100000",
  57713=>"000100110",
  57714=>"101111101",
  57715=>"010001011",
  57716=>"101100001",
  57717=>"011111000",
  57718=>"010010011",
  57719=>"101000011",
  57720=>"100011100",
  57721=>"110111011",
  57722=>"101100100",
  57723=>"010101100",
  57724=>"000111111",
  57725=>"101111011",
  57726=>"110011110",
  57727=>"000010100",
  57728=>"011011001",
  57729=>"001101010",
  57730=>"101100001",
  57731=>"110100100",
  57732=>"111100101",
  57733=>"001011011",
  57734=>"010010011",
  57735=>"001101001",
  57736=>"011101111",
  57737=>"011000000",
  57738=>"000000110",
  57739=>"101111001",
  57740=>"010000100",
  57741=>"010000101",
  57742=>"101111001",
  57743=>"011101011",
  57744=>"000111110",
  57745=>"000101001",
  57746=>"000001000",
  57747=>"011000001",
  57748=>"011100011",
  57749=>"101100111",
  57750=>"100101110",
  57751=>"110100010",
  57752=>"011111101",
  57753=>"111001000",
  57754=>"011011101",
  57755=>"111110010",
  57756=>"010010101",
  57757=>"111001011",
  57758=>"111100000",
  57759=>"110111001",
  57760=>"000010100",
  57761=>"001101110",
  57762=>"000011110",
  57763=>"010000000",
  57764=>"100011111",
  57765=>"001001010",
  57766=>"111001100",
  57767=>"100011110",
  57768=>"011011110",
  57769=>"011010011",
  57770=>"011111111",
  57771=>"111111010",
  57772=>"011011000",
  57773=>"010101110",
  57774=>"111100010",
  57775=>"100100110",
  57776=>"010000000",
  57777=>"010000000",
  57778=>"110111011",
  57779=>"101101001",
  57780=>"111011000",
  57781=>"110000101",
  57782=>"001000000",
  57783=>"111001100",
  57784=>"111100010",
  57785=>"001000110",
  57786=>"110001001",
  57787=>"100011101",
  57788=>"101010110",
  57789=>"011010110",
  57790=>"111011000",
  57791=>"111001010",
  57792=>"010101100",
  57793=>"101001110",
  57794=>"110010100",
  57795=>"001111011",
  57796=>"001001111",
  57797=>"101000101",
  57798=>"010001011",
  57799=>"000101011",
  57800=>"100101111",
  57801=>"100101110",
  57802=>"010011010",
  57803=>"100100110",
  57804=>"100100101",
  57805=>"001100111",
  57806=>"111011001",
  57807=>"101010000",
  57808=>"101111000",
  57809=>"001001000",
  57810=>"111101111",
  57811=>"010100011",
  57812=>"010000000",
  57813=>"111100101",
  57814=>"111011000",
  57815=>"011000101",
  57816=>"100000111",
  57817=>"010100010",
  57818=>"000110000",
  57819=>"111110101",
  57820=>"001001000",
  57821=>"011001011",
  57822=>"100001011",
  57823=>"001011010",
  57824=>"100110100",
  57825=>"100101111",
  57826=>"111000001",
  57827=>"111111000",
  57828=>"001100001",
  57829=>"101111011",
  57830=>"110011111",
  57831=>"100001001",
  57832=>"000100110",
  57833=>"000110101",
  57834=>"101011110",
  57835=>"010001001",
  57836=>"011000000",
  57837=>"000010110",
  57838=>"101111010",
  57839=>"100100000",
  57840=>"111001001",
  57841=>"101111111",
  57842=>"110100000",
  57843=>"011110011",
  57844=>"101001011",
  57845=>"010001101",
  57846=>"100001100",
  57847=>"000101111",
  57848=>"011010001",
  57849=>"100110101",
  57850=>"110001100",
  57851=>"011000100",
  57852=>"001001001",
  57853=>"111111111",
  57854=>"100010010",
  57855=>"111100001",
  57856=>"011110001",
  57857=>"101111100",
  57858=>"100010010",
  57859=>"011101010",
  57860=>"111111010",
  57861=>"111101010",
  57862=>"011101011",
  57863=>"100000100",
  57864=>"111100001",
  57865=>"100011001",
  57866=>"101000111",
  57867=>"111101101",
  57868=>"111011011",
  57869=>"010000010",
  57870=>"000100101",
  57871=>"011110011",
  57872=>"000100011",
  57873=>"011101111",
  57874=>"001111000",
  57875=>"111011100",
  57876=>"101001111",
  57877=>"101000101",
  57878=>"110101100",
  57879=>"110010011",
  57880=>"100000101",
  57881=>"101110110",
  57882=>"011111110",
  57883=>"001110000",
  57884=>"011110000",
  57885=>"101011001",
  57886=>"010100010",
  57887=>"100100100",
  57888=>"011000010",
  57889=>"010000000",
  57890=>"010000100",
  57891=>"111010101",
  57892=>"101011010",
  57893=>"101001010",
  57894=>"000100001",
  57895=>"010010011",
  57896=>"100101001",
  57897=>"000010100",
  57898=>"010000010",
  57899=>"111110000",
  57900=>"100001110",
  57901=>"101001100",
  57902=>"110100100",
  57903=>"101010001",
  57904=>"010010001",
  57905=>"110011010",
  57906=>"001101101",
  57907=>"100000011",
  57908=>"101101100",
  57909=>"101001100",
  57910=>"110101011",
  57911=>"000100111",
  57912=>"011111100",
  57913=>"000101110",
  57914=>"111010110",
  57915=>"110000101",
  57916=>"111100110",
  57917=>"111111011",
  57918=>"111100011",
  57919=>"010011101",
  57920=>"001010001",
  57921=>"101101010",
  57922=>"111101100",
  57923=>"101000101",
  57924=>"001100110",
  57925=>"000110110",
  57926=>"000110100",
  57927=>"110101100",
  57928=>"010000110",
  57929=>"101101111",
  57930=>"011001101",
  57931=>"111011001",
  57932=>"010110001",
  57933=>"001001110",
  57934=>"101101101",
  57935=>"011001010",
  57936=>"110101001",
  57937=>"000011001",
  57938=>"000101000",
  57939=>"010010101",
  57940=>"001101011",
  57941=>"110000100",
  57942=>"010100101",
  57943=>"010110101",
  57944=>"010000011",
  57945=>"000010100",
  57946=>"001000000",
  57947=>"001010101",
  57948=>"100111110",
  57949=>"000011110",
  57950=>"000011011",
  57951=>"011010000",
  57952=>"001000110",
  57953=>"110110100",
  57954=>"100011110",
  57955=>"001001010",
  57956=>"110001110",
  57957=>"111001010",
  57958=>"100010101",
  57959=>"000100100",
  57960=>"000010100",
  57961=>"001100101",
  57962=>"110100001",
  57963=>"000110000",
  57964=>"010011011",
  57965=>"001001010",
  57966=>"100101011",
  57967=>"011101001",
  57968=>"111111010",
  57969=>"000000100",
  57970=>"100110100",
  57971=>"001110001",
  57972=>"101101011",
  57973=>"001100001",
  57974=>"011101011",
  57975=>"100010011",
  57976=>"110101111",
  57977=>"100011010",
  57978=>"001000111",
  57979=>"011111101",
  57980=>"011000101",
  57981=>"110111101",
  57982=>"110011000",
  57983=>"011101110",
  57984=>"101110101",
  57985=>"001011001",
  57986=>"010101111",
  57987=>"001101000",
  57988=>"000010011",
  57989=>"111000010",
  57990=>"011100011",
  57991=>"111001100",
  57992=>"101111001",
  57993=>"101010100",
  57994=>"110010000",
  57995=>"110010000",
  57996=>"100101111",
  57997=>"101011111",
  57998=>"111111110",
  57999=>"100101010",
  58000=>"101001011",
  58001=>"100001101",
  58002=>"010110010",
  58003=>"110011110",
  58004=>"001000001",
  58005=>"011101111",
  58006=>"010111110",
  58007=>"110100100",
  58008=>"101101110",
  58009=>"011110100",
  58010=>"001110101",
  58011=>"000100011",
  58012=>"001010000",
  58013=>"000110111",
  58014=>"000110001",
  58015=>"000010100",
  58016=>"011001000",
  58017=>"111101100",
  58018=>"000111000",
  58019=>"011010110",
  58020=>"001100111",
  58021=>"011010010",
  58022=>"110101111",
  58023=>"110000000",
  58024=>"010111111",
  58025=>"000000011",
  58026=>"101111101",
  58027=>"110001001",
  58028=>"111011001",
  58029=>"011011011",
  58030=>"100101100",
  58031=>"110000010",
  58032=>"110101111",
  58033=>"001000000",
  58034=>"101010001",
  58035=>"001001010",
  58036=>"001000100",
  58037=>"111011011",
  58038=>"110011000",
  58039=>"110110111",
  58040=>"110010000",
  58041=>"100111001",
  58042=>"111001000",
  58043=>"110110101",
  58044=>"001000110",
  58045=>"011010011",
  58046=>"111001001",
  58047=>"101001010",
  58048=>"000111011",
  58049=>"101111110",
  58050=>"000000010",
  58051=>"111010011",
  58052=>"001111101",
  58053=>"111010000",
  58054=>"001101110",
  58055=>"100100001",
  58056=>"011001011",
  58057=>"010000011",
  58058=>"110101010",
  58059=>"010111111",
  58060=>"010000010",
  58061=>"110011111",
  58062=>"011010010",
  58063=>"111011010",
  58064=>"011101011",
  58065=>"010011111",
  58066=>"001010011",
  58067=>"001011001",
  58068=>"111010111",
  58069=>"100001010",
  58070=>"100000111",
  58071=>"010010100",
  58072=>"010101000",
  58073=>"010100011",
  58074=>"000010100",
  58075=>"011101110",
  58076=>"101100000",
  58077=>"111010000",
  58078=>"100000000",
  58079=>"010000101",
  58080=>"101000101",
  58081=>"000000001",
  58082=>"110111100",
  58083=>"000100101",
  58084=>"100100010",
  58085=>"000010110",
  58086=>"111111101",
  58087=>"110110100",
  58088=>"001111001",
  58089=>"110100001",
  58090=>"001001010",
  58091=>"010101111",
  58092=>"001111001",
  58093=>"010000001",
  58094=>"001011101",
  58095=>"000110110",
  58096=>"011101011",
  58097=>"100011011",
  58098=>"110001100",
  58099=>"010100101",
  58100=>"001110111",
  58101=>"000000000",
  58102=>"110101011",
  58103=>"111010100",
  58104=>"010111010",
  58105=>"010000110",
  58106=>"010001000",
  58107=>"101101000",
  58108=>"000010001",
  58109=>"000101100",
  58110=>"110101111",
  58111=>"011110111",
  58112=>"000111101",
  58113=>"100101000",
  58114=>"100100110",
  58115=>"010010011",
  58116=>"111001101",
  58117=>"111111100",
  58118=>"100101001",
  58119=>"010100110",
  58120=>"101010001",
  58121=>"000000101",
  58122=>"100011110",
  58123=>"101000011",
  58124=>"000001110",
  58125=>"101110101",
  58126=>"000001010",
  58127=>"100110111",
  58128=>"110111110",
  58129=>"101010101",
  58130=>"111100110",
  58131=>"111010010",
  58132=>"110011001",
  58133=>"010001100",
  58134=>"010011001",
  58135=>"111010011",
  58136=>"010100100",
  58137=>"111001001",
  58138=>"011101000",
  58139=>"111001001",
  58140=>"100000010",
  58141=>"101101101",
  58142=>"000011000",
  58143=>"011110011",
  58144=>"110010100",
  58145=>"110101100",
  58146=>"011110011",
  58147=>"011101000",
  58148=>"001101011",
  58149=>"111001110",
  58150=>"001011010",
  58151=>"100000110",
  58152=>"011011111",
  58153=>"011100000",
  58154=>"111101010",
  58155=>"011101100",
  58156=>"000111001",
  58157=>"101011000",
  58158=>"011010001",
  58159=>"001101110",
  58160=>"101100011",
  58161=>"000101111",
  58162=>"000000000",
  58163=>"000110111",
  58164=>"110011100",
  58165=>"110110101",
  58166=>"110110001",
  58167=>"010111011",
  58168=>"001001010",
  58169=>"101100100",
  58170=>"000001100",
  58171=>"101010000",
  58172=>"101000110",
  58173=>"000001011",
  58174=>"000101010",
  58175=>"100100100",
  58176=>"010011101",
  58177=>"101110110",
  58178=>"101111111",
  58179=>"111011000",
  58180=>"100111001",
  58181=>"010100000",
  58182=>"100001100",
  58183=>"001001010",
  58184=>"111000011",
  58185=>"011110010",
  58186=>"101010011",
  58187=>"101001001",
  58188=>"010000101",
  58189=>"100001101",
  58190=>"010111011",
  58191=>"110001101",
  58192=>"111110010",
  58193=>"010110100",
  58194=>"111010001",
  58195=>"111111111",
  58196=>"110110011",
  58197=>"011100000",
  58198=>"100000000",
  58199=>"011111011",
  58200=>"010000000",
  58201=>"010101010",
  58202=>"110000001",
  58203=>"100111111",
  58204=>"010101100",
  58205=>"101101000",
  58206=>"000001100",
  58207=>"111111101",
  58208=>"001100100",
  58209=>"101110011",
  58210=>"101100110",
  58211=>"000101110",
  58212=>"010111111",
  58213=>"011011100",
  58214=>"011010110",
  58215=>"110011000",
  58216=>"011100000",
  58217=>"111100100",
  58218=>"000000100",
  58219=>"111010100",
  58220=>"010000100",
  58221=>"001000101",
  58222=>"011010110",
  58223=>"111011010",
  58224=>"100001010",
  58225=>"010010111",
  58226=>"010001101",
  58227=>"111011110",
  58228=>"010101100",
  58229=>"100111110",
  58230=>"111110100",
  58231=>"111011000",
  58232=>"001100111",
  58233=>"101101010",
  58234=>"110100111",
  58235=>"000100110",
  58236=>"111000001",
  58237=>"110000101",
  58238=>"110101011",
  58239=>"011001000",
  58240=>"101010111",
  58241=>"101111001",
  58242=>"111110101",
  58243=>"111010111",
  58244=>"011110100",
  58245=>"000001111",
  58246=>"010100101",
  58247=>"101101100",
  58248=>"000001111",
  58249=>"000000000",
  58250=>"101001010",
  58251=>"111111101",
  58252=>"010000111",
  58253=>"100011001",
  58254=>"001011110",
  58255=>"000010110",
  58256=>"100110010",
  58257=>"101101111",
  58258=>"000000100",
  58259=>"101010111",
  58260=>"111011100",
  58261=>"001001010",
  58262=>"110111101",
  58263=>"110011010",
  58264=>"001011010",
  58265=>"101011000",
  58266=>"010001110",
  58267=>"010100100",
  58268=>"010010011",
  58269=>"101100111",
  58270=>"000110100",
  58271=>"000011000",
  58272=>"111000000",
  58273=>"011010001",
  58274=>"111111100",
  58275=>"011000001",
  58276=>"010110011",
  58277=>"100101110",
  58278=>"111110000",
  58279=>"111111111",
  58280=>"110101100",
  58281=>"001110011",
  58282=>"001110010",
  58283=>"100011100",
  58284=>"100100101",
  58285=>"000011100",
  58286=>"000100010",
  58287=>"111100100",
  58288=>"000000010",
  58289=>"011111111",
  58290=>"010001110",
  58291=>"110011000",
  58292=>"111101001",
  58293=>"101000100",
  58294=>"010000100",
  58295=>"010110110",
  58296=>"010110101",
  58297=>"010110001",
  58298=>"010101101",
  58299=>"111001110",
  58300=>"010100110",
  58301=>"000000010",
  58302=>"011101111",
  58303=>"100000100",
  58304=>"110100001",
  58305=>"101010001",
  58306=>"100010011",
  58307=>"001101101",
  58308=>"011100111",
  58309=>"100010011",
  58310=>"101101010",
  58311=>"110001010",
  58312=>"010101101",
  58313=>"111100000",
  58314=>"100101101",
  58315=>"101110000",
  58316=>"001010111",
  58317=>"001110100",
  58318=>"001010011",
  58319=>"110000000",
  58320=>"001001111",
  58321=>"101001011",
  58322=>"010010000",
  58323=>"101011100",
  58324=>"111111011",
  58325=>"011101011",
  58326=>"101011101",
  58327=>"011111001",
  58328=>"111000000",
  58329=>"111101001",
  58330=>"010100010",
  58331=>"100011110",
  58332=>"111010000",
  58333=>"010110000",
  58334=>"111101011",
  58335=>"011011011",
  58336=>"000011101",
  58337=>"110101111",
  58338=>"100000010",
  58339=>"110111100",
  58340=>"010011000",
  58341=>"000000110",
  58342=>"000000010",
  58343=>"000010111",
  58344=>"101100110",
  58345=>"010110100",
  58346=>"010010110",
  58347=>"110100001",
  58348=>"010100110",
  58349=>"000010000",
  58350=>"011011110",
  58351=>"110010100",
  58352=>"011101011",
  58353=>"000010001",
  58354=>"001011001",
  58355=>"100100110",
  58356=>"001110001",
  58357=>"011010111",
  58358=>"001010011",
  58359=>"010011000",
  58360=>"010011000",
  58361=>"010000000",
  58362=>"001100110",
  58363=>"011000100",
  58364=>"000010110",
  58365=>"110111111",
  58366=>"101010101",
  58367=>"110000110",
  58368=>"111111001",
  58369=>"100111111",
  58370=>"011111111",
  58371=>"000001101",
  58372=>"100000000",
  58373=>"100011101",
  58374=>"111101111",
  58375=>"101111100",
  58376=>"010001011",
  58377=>"010000111",
  58378=>"111010100",
  58379=>"101000001",
  58380=>"010100110",
  58381=>"010100111",
  58382=>"100001101",
  58383=>"100111001",
  58384=>"001000100",
  58385=>"111110110",
  58386=>"110011000",
  58387=>"001101010",
  58388=>"000000011",
  58389=>"011000101",
  58390=>"101111110",
  58391=>"001010000",
  58392=>"001101011",
  58393=>"010111110",
  58394=>"100110110",
  58395=>"110011011",
  58396=>"110110110",
  58397=>"001010001",
  58398=>"000111001",
  58399=>"100111111",
  58400=>"010001100",
  58401=>"001111001",
  58402=>"001100100",
  58403=>"001000010",
  58404=>"110111110",
  58405=>"111011011",
  58406=>"000011010",
  58407=>"000110111",
  58408=>"101101010",
  58409=>"101110010",
  58410=>"000110001",
  58411=>"010000111",
  58412=>"010010000",
  58413=>"111001000",
  58414=>"010000001",
  58415=>"111100110",
  58416=>"111101101",
  58417=>"111001100",
  58418=>"111111001",
  58419=>"111010011",
  58420=>"101101101",
  58421=>"111011000",
  58422=>"101100100",
  58423=>"011010101",
  58424=>"011111101",
  58425=>"100001110",
  58426=>"011110001",
  58427=>"100001100",
  58428=>"100001101",
  58429=>"001101101",
  58430=>"001101000",
  58431=>"100011101",
  58432=>"001010111",
  58433=>"000100000",
  58434=>"010000110",
  58435=>"000000010",
  58436=>"011010110",
  58437=>"001111011",
  58438=>"111001010",
  58439=>"111100010",
  58440=>"100110000",
  58441=>"000111000",
  58442=>"001011001",
  58443=>"000111110",
  58444=>"100001000",
  58445=>"111011100",
  58446=>"001011001",
  58447=>"111111111",
  58448=>"000101001",
  58449=>"010101000",
  58450=>"101101010",
  58451=>"000000000",
  58452=>"010010000",
  58453=>"000111110",
  58454=>"111011110",
  58455=>"000100011",
  58456=>"110011000",
  58457=>"011011111",
  58458=>"011111011",
  58459=>"011001001",
  58460=>"010001000",
  58461=>"000001111",
  58462=>"100001000",
  58463=>"110110100",
  58464=>"000101101",
  58465=>"111001000",
  58466=>"010100100",
  58467=>"111110100",
  58468=>"100110101",
  58469=>"100111000",
  58470=>"000110011",
  58471=>"001000110",
  58472=>"100001000",
  58473=>"011101110",
  58474=>"110000100",
  58475=>"000001111",
  58476=>"100100010",
  58477=>"100011010",
  58478=>"111110000",
  58479=>"101111010",
  58480=>"011111111",
  58481=>"100110110",
  58482=>"110101100",
  58483=>"001111000",
  58484=>"001010110",
  58485=>"101100000",
  58486=>"110001100",
  58487=>"000010000",
  58488=>"001100000",
  58489=>"111100010",
  58490=>"101100010",
  58491=>"110111111",
  58492=>"001100011",
  58493=>"110100101",
  58494=>"000010111",
  58495=>"111011011",
  58496=>"111101010",
  58497=>"000111010",
  58498=>"000000001",
  58499=>"000011111",
  58500=>"110101000",
  58501=>"100110100",
  58502=>"111100100",
  58503=>"001111011",
  58504=>"011100000",
  58505=>"001100111",
  58506=>"110110110",
  58507=>"000000011",
  58508=>"001111100",
  58509=>"101010010",
  58510=>"011101100",
  58511=>"110100101",
  58512=>"010000000",
  58513=>"100101101",
  58514=>"110111010",
  58515=>"000010001",
  58516=>"111011010",
  58517=>"110100000",
  58518=>"111111011",
  58519=>"100100001",
  58520=>"001000001",
  58521=>"000011010",
  58522=>"000100010",
  58523=>"001011010",
  58524=>"010000010",
  58525=>"100000001",
  58526=>"010001110",
  58527=>"110101000",
  58528=>"011000000",
  58529=>"011111001",
  58530=>"010111110",
  58531=>"010111010",
  58532=>"101101100",
  58533=>"011111000",
  58534=>"000010001",
  58535=>"110110111",
  58536=>"000011011",
  58537=>"110001000",
  58538=>"010101011",
  58539=>"111110101",
  58540=>"100101101",
  58541=>"101000000",
  58542=>"011111000",
  58543=>"100011001",
  58544=>"001011100",
  58545=>"000101000",
  58546=>"110001011",
  58547=>"000100000",
  58548=>"000011100",
  58549=>"100000101",
  58550=>"110010010",
  58551=>"101000011",
  58552=>"010011110",
  58553=>"111001011",
  58554=>"000000000",
  58555=>"111011100",
  58556=>"110110111",
  58557=>"110001001",
  58558=>"001111010",
  58559=>"000011110",
  58560=>"100011101",
  58561=>"011000101",
  58562=>"000111110",
  58563=>"110010110",
  58564=>"110101100",
  58565=>"000010011",
  58566=>"010001010",
  58567=>"000010100",
  58568=>"110101101",
  58569=>"011101100",
  58570=>"000011000",
  58571=>"111101011",
  58572=>"110111100",
  58573=>"000111010",
  58574=>"000100100",
  58575=>"110100101",
  58576=>"110110100",
  58577=>"111011111",
  58578=>"101000111",
  58579=>"101011100",
  58580=>"100101100",
  58581=>"000001111",
  58582=>"000110100",
  58583=>"001010010",
  58584=>"011101101",
  58585=>"101011001",
  58586=>"110010100",
  58587=>"000011101",
  58588=>"100110011",
  58589=>"101101100",
  58590=>"100000001",
  58591=>"100110001",
  58592=>"010100101",
  58593=>"001001000",
  58594=>"001101101",
  58595=>"000100010",
  58596=>"101011001",
  58597=>"000100001",
  58598=>"101000001",
  58599=>"000101010",
  58600=>"100111100",
  58601=>"100101110",
  58602=>"111000101",
  58603=>"010001100",
  58604=>"000010000",
  58605=>"110101010",
  58606=>"000000111",
  58607=>"000110100",
  58608=>"000100101",
  58609=>"110000101",
  58610=>"000010010",
  58611=>"000111010",
  58612=>"000001101",
  58613=>"101010010",
  58614=>"101010001",
  58615=>"010010001",
  58616=>"000001100",
  58617=>"010110011",
  58618=>"110011100",
  58619=>"000111010",
  58620=>"110000000",
  58621=>"100101100",
  58622=>"110101011",
  58623=>"001011100",
  58624=>"010011001",
  58625=>"100011011",
  58626=>"001101011",
  58627=>"010011000",
  58628=>"110111100",
  58629=>"110010011",
  58630=>"001000010",
  58631=>"000101110",
  58632=>"001001101",
  58633=>"110110001",
  58634=>"101101001",
  58635=>"111001101",
  58636=>"000110111",
  58637=>"000000101",
  58638=>"001001001",
  58639=>"010000100",
  58640=>"110101101",
  58641=>"010100100",
  58642=>"011000101",
  58643=>"001001111",
  58644=>"011110111",
  58645=>"001100011",
  58646=>"100000010",
  58647=>"100101001",
  58648=>"100101001",
  58649=>"000100101",
  58650=>"010110101",
  58651=>"111001010",
  58652=>"110101101",
  58653=>"100001111",
  58654=>"011100100",
  58655=>"011101011",
  58656=>"100100111",
  58657=>"111010000",
  58658=>"010000000",
  58659=>"100101110",
  58660=>"110101010",
  58661=>"011111001",
  58662=>"001101101",
  58663=>"101100010",
  58664=>"110111000",
  58665=>"111110000",
  58666=>"001111111",
  58667=>"111000000",
  58668=>"011111011",
  58669=>"011011111",
  58670=>"101100001",
  58671=>"010110010",
  58672=>"111100100",
  58673=>"001000110",
  58674=>"001111101",
  58675=>"001100011",
  58676=>"100110010",
  58677=>"110000000",
  58678=>"110000001",
  58679=>"111100101",
  58680=>"000010001",
  58681=>"111100101",
  58682=>"010011100",
  58683=>"101101001",
  58684=>"001000110",
  58685=>"110001000",
  58686=>"011111001",
  58687=>"111101001",
  58688=>"111111000",
  58689=>"011010111",
  58690=>"110111101",
  58691=>"000011001",
  58692=>"011011110",
  58693=>"011010011",
  58694=>"110100110",
  58695=>"111000001",
  58696=>"001110010",
  58697=>"011011101",
  58698=>"100010101",
  58699=>"000100010",
  58700=>"101111110",
  58701=>"101001110",
  58702=>"000110100",
  58703=>"000010011",
  58704=>"101011110",
  58705=>"001110001",
  58706=>"000100000",
  58707=>"100100001",
  58708=>"011101010",
  58709=>"010111111",
  58710=>"000111111",
  58711=>"011010101",
  58712=>"101011100",
  58713=>"110000000",
  58714=>"110001010",
  58715=>"000001100",
  58716=>"000010100",
  58717=>"111011001",
  58718=>"101001110",
  58719=>"000111001",
  58720=>"000111010",
  58721=>"111110110",
  58722=>"000010000",
  58723=>"110101110",
  58724=>"100001110",
  58725=>"010010000",
  58726=>"101111011",
  58727=>"001010000",
  58728=>"010101100",
  58729=>"011111001",
  58730=>"000110100",
  58731=>"111101101",
  58732=>"100000100",
  58733=>"101100001",
  58734=>"001010111",
  58735=>"001101100",
  58736=>"100111000",
  58737=>"011101001",
  58738=>"100111001",
  58739=>"100100010",
  58740=>"000101011",
  58741=>"000011001",
  58742=>"110100000",
  58743=>"000110101",
  58744=>"111101101",
  58745=>"110000001",
  58746=>"101010011",
  58747=>"101001001",
  58748=>"001010001",
  58749=>"111010000",
  58750=>"111000010",
  58751=>"101000011",
  58752=>"110110001",
  58753=>"000001010",
  58754=>"110110000",
  58755=>"010001010",
  58756=>"101111011",
  58757=>"010010000",
  58758=>"010000001",
  58759=>"011101001",
  58760=>"000111000",
  58761=>"100110000",
  58762=>"101001110",
  58763=>"100111101",
  58764=>"011000110",
  58765=>"010100000",
  58766=>"000010110",
  58767=>"000010100",
  58768=>"101011010",
  58769=>"000111001",
  58770=>"100100010",
  58771=>"001101101",
  58772=>"001110010",
  58773=>"100011110",
  58774=>"101100000",
  58775=>"001011101",
  58776=>"000101100",
  58777=>"010100011",
  58778=>"000000000",
  58779=>"000101000",
  58780=>"110111100",
  58781=>"001011000",
  58782=>"100100101",
  58783=>"110111100",
  58784=>"111100100",
  58785=>"111101001",
  58786=>"101010000",
  58787=>"000010010",
  58788=>"111101000",
  58789=>"000110001",
  58790=>"000001100",
  58791=>"110000001",
  58792=>"111110110",
  58793=>"001001110",
  58794=>"000100011",
  58795=>"011100100",
  58796=>"001100110",
  58797=>"001000001",
  58798=>"100010011",
  58799=>"101001010",
  58800=>"011100001",
  58801=>"111001100",
  58802=>"011110111",
  58803=>"111111111",
  58804=>"000101001",
  58805=>"000111100",
  58806=>"011010101",
  58807=>"000001001",
  58808=>"000111010",
  58809=>"100011110",
  58810=>"101111010",
  58811=>"100001101",
  58812=>"000100010",
  58813=>"001000101",
  58814=>"001100100",
  58815=>"101010000",
  58816=>"011010100",
  58817=>"010110100",
  58818=>"000011000",
  58819=>"011100101",
  58820=>"100001100",
  58821=>"101000101",
  58822=>"001010101",
  58823=>"101101100",
  58824=>"101000001",
  58825=>"001110111",
  58826=>"000000111",
  58827=>"001100100",
  58828=>"000101101",
  58829=>"100001111",
  58830=>"000001001",
  58831=>"100101011",
  58832=>"100000111",
  58833=>"001101001",
  58834=>"000010010",
  58835=>"100101110",
  58836=>"001000101",
  58837=>"001010111",
  58838=>"110111001",
  58839=>"001011010",
  58840=>"000011100",
  58841=>"011001101",
  58842=>"010111111",
  58843=>"011100111",
  58844=>"101111101",
  58845=>"111001000",
  58846=>"100000111",
  58847=>"111100100",
  58848=>"000010101",
  58849=>"100001000",
  58850=>"101000111",
  58851=>"101011111",
  58852=>"101010110",
  58853=>"100000111",
  58854=>"000001000",
  58855=>"011100111",
  58856=>"111110011",
  58857=>"111001010",
  58858=>"110101100",
  58859=>"111110101",
  58860=>"011101100",
  58861=>"011001101",
  58862=>"010011110",
  58863=>"111111101",
  58864=>"000101111",
  58865=>"001111101",
  58866=>"010110111",
  58867=>"101011010",
  58868=>"101010001",
  58869=>"001101110",
  58870=>"101111011",
  58871=>"111110111",
  58872=>"100110111",
  58873=>"000111011",
  58874=>"010010011",
  58875=>"011001000",
  58876=>"011001010",
  58877=>"010001011",
  58878=>"111101100",
  58879=>"010100111",
  58880=>"001001001",
  58881=>"000100001",
  58882=>"100011000",
  58883=>"010000000",
  58884=>"110111110",
  58885=>"100100101",
  58886=>"100111100",
  58887=>"000101001",
  58888=>"100101011",
  58889=>"000000100",
  58890=>"000010000",
  58891=>"111101000",
  58892=>"001000011",
  58893=>"011010011",
  58894=>"101000111",
  58895=>"101101101",
  58896=>"000110101",
  58897=>"111111010",
  58898=>"010110111",
  58899=>"001101011",
  58900=>"001000100",
  58901=>"110101100",
  58902=>"000100000",
  58903=>"011110110",
  58904=>"010010111",
  58905=>"000100101",
  58906=>"001111001",
  58907=>"010100001",
  58908=>"111010001",
  58909=>"111100111",
  58910=>"111011011",
  58911=>"100011000",
  58912=>"111001001",
  58913=>"000000001",
  58914=>"101110100",
  58915=>"000100001",
  58916=>"011100001",
  58917=>"000000110",
  58918=>"000001010",
  58919=>"000000001",
  58920=>"001100000",
  58921=>"000101001",
  58922=>"011001100",
  58923=>"100010011",
  58924=>"010101001",
  58925=>"100000010",
  58926=>"011111110",
  58927=>"101111101",
  58928=>"001000011",
  58929=>"101000110",
  58930=>"000011000",
  58931=>"100001011",
  58932=>"001011100",
  58933=>"101001111",
  58934=>"010001100",
  58935=>"111111111",
  58936=>"101101000",
  58937=>"001001011",
  58938=>"010001110",
  58939=>"100111001",
  58940=>"010110111",
  58941=>"000001000",
  58942=>"110001110",
  58943=>"001110100",
  58944=>"000101100",
  58945=>"100001010",
  58946=>"001100010",
  58947=>"111101101",
  58948=>"001110101",
  58949=>"010011001",
  58950=>"110101010",
  58951=>"110100110",
  58952=>"011100111",
  58953=>"010011111",
  58954=>"011111111",
  58955=>"001101101",
  58956=>"010100101",
  58957=>"010000010",
  58958=>"101001010",
  58959=>"110000110",
  58960=>"111101111",
  58961=>"001000101",
  58962=>"111101111",
  58963=>"110010100",
  58964=>"001100100",
  58965=>"100110001",
  58966=>"100110001",
  58967=>"011111000",
  58968=>"010110001",
  58969=>"100100110",
  58970=>"100111101",
  58971=>"000101000",
  58972=>"000001000",
  58973=>"111010000",
  58974=>"010000000",
  58975=>"000110001",
  58976=>"001001000",
  58977=>"000010101",
  58978=>"001000000",
  58979=>"011001111",
  58980=>"010111101",
  58981=>"001000000",
  58982=>"001000100",
  58983=>"001011011",
  58984=>"111110111",
  58985=>"111011100",
  58986=>"010001001",
  58987=>"111010010",
  58988=>"111001011",
  58989=>"001110011",
  58990=>"001101111",
  58991=>"101110101",
  58992=>"010111100",
  58993=>"010111111",
  58994=>"000100010",
  58995=>"111111010",
  58996=>"001101100",
  58997=>"011000100",
  58998=>"001100100",
  58999=>"101000010",
  59000=>"110100100",
  59001=>"100101110",
  59002=>"101101100",
  59003=>"100011111",
  59004=>"110010011",
  59005=>"000111011",
  59006=>"000010010",
  59007=>"000101100",
  59008=>"010111100",
  59009=>"101011011",
  59010=>"100011000",
  59011=>"011101101",
  59012=>"100111100",
  59013=>"110011100",
  59014=>"011100101",
  59015=>"110100101",
  59016=>"110100001",
  59017=>"100011111",
  59018=>"000000010",
  59019=>"011000101",
  59020=>"100000000",
  59021=>"010111011",
  59022=>"001110111",
  59023=>"110000111",
  59024=>"000011010",
  59025=>"100111010",
  59026=>"110011001",
  59027=>"000111100",
  59028=>"100000000",
  59029=>"111001010",
  59030=>"101111000",
  59031=>"101010010",
  59032=>"101000001",
  59033=>"101000001",
  59034=>"001110011",
  59035=>"101101101",
  59036=>"101100111",
  59037=>"111011011",
  59038=>"001011001",
  59039=>"011010000",
  59040=>"001011001",
  59041=>"100110011",
  59042=>"100110111",
  59043=>"111011010",
  59044=>"011111111",
  59045=>"010010111",
  59046=>"101101111",
  59047=>"100000110",
  59048=>"111000000",
  59049=>"111010011",
  59050=>"000000000",
  59051=>"110110010",
  59052=>"111001001",
  59053=>"100011111",
  59054=>"101011110",
  59055=>"110011111",
  59056=>"110001010",
  59057=>"010110100",
  59058=>"101010010",
  59059=>"001001101",
  59060=>"011110110",
  59061=>"011101000",
  59062=>"110001111",
  59063=>"001010010",
  59064=>"110110001",
  59065=>"001010001",
  59066=>"001110110",
  59067=>"001010110",
  59068=>"000101111",
  59069=>"101101000",
  59070=>"111110110",
  59071=>"101001010",
  59072=>"100001111",
  59073=>"101001000",
  59074=>"010010110",
  59075=>"110110001",
  59076=>"010110111",
  59077=>"011000000",
  59078=>"001101001",
  59079=>"001011011",
  59080=>"101011111",
  59081=>"101110110",
  59082=>"110100101",
  59083=>"000111011",
  59084=>"110001000",
  59085=>"001100011",
  59086=>"101110100",
  59087=>"000001110",
  59088=>"101110110",
  59089=>"010100101",
  59090=>"000011000",
  59091=>"011100111",
  59092=>"000101100",
  59093=>"011101111",
  59094=>"011111111",
  59095=>"111000001",
  59096=>"001001101",
  59097=>"100001001",
  59098=>"110011110",
  59099=>"100010010",
  59100=>"110011100",
  59101=>"000111101",
  59102=>"111111001",
  59103=>"000111100",
  59104=>"101111101",
  59105=>"101001100",
  59106=>"101011011",
  59107=>"101111000",
  59108=>"000111110",
  59109=>"010000010",
  59110=>"101010001",
  59111=>"000010001",
  59112=>"001001010",
  59113=>"100110101",
  59114=>"100101111",
  59115=>"001001000",
  59116=>"111101101",
  59117=>"111110100",
  59118=>"000100100",
  59119=>"111101101",
  59120=>"111111110",
  59121=>"001111010",
  59122=>"001110100",
  59123=>"001000000",
  59124=>"111000101",
  59125=>"100111010",
  59126=>"111110010",
  59127=>"111011100",
  59128=>"011101011",
  59129=>"100010011",
  59130=>"001010010",
  59131=>"110111010",
  59132=>"010110000",
  59133=>"111011011",
  59134=>"001111011",
  59135=>"000001100",
  59136=>"000000000",
  59137=>"110000010",
  59138=>"100101011",
  59139=>"111111000",
  59140=>"011100110",
  59141=>"000101000",
  59142=>"101101011",
  59143=>"100011000",
  59144=>"101000001",
  59145=>"110001111",
  59146=>"100000001",
  59147=>"010110110",
  59148=>"100001001",
  59149=>"101011101",
  59150=>"110000111",
  59151=>"100110100",
  59152=>"010000110",
  59153=>"000001101",
  59154=>"111011100",
  59155=>"000011110",
  59156=>"010101010",
  59157=>"100110001",
  59158=>"010010100",
  59159=>"100111000",
  59160=>"111010000",
  59161=>"110010000",
  59162=>"110000001",
  59163=>"000001000",
  59164=>"111100001",
  59165=>"011101001",
  59166=>"010011011",
  59167=>"000011101",
  59168=>"110101110",
  59169=>"001000110",
  59170=>"000100010",
  59171=>"101100100",
  59172=>"110000101",
  59173=>"000100111",
  59174=>"000011010",
  59175=>"011110111",
  59176=>"010110100",
  59177=>"010010000",
  59178=>"001101000",
  59179=>"101000001",
  59180=>"011101111",
  59181=>"001111000",
  59182=>"111001110",
  59183=>"100010101",
  59184=>"000100011",
  59185=>"100101000",
  59186=>"110010100",
  59187=>"111101110",
  59188=>"111011111",
  59189=>"101001111",
  59190=>"011011101",
  59191=>"011010000",
  59192=>"011011011",
  59193=>"100101110",
  59194=>"000110100",
  59195=>"010110111",
  59196=>"101111100",
  59197=>"111000100",
  59198=>"011000100",
  59199=>"110100010",
  59200=>"111001011",
  59201=>"100101110",
  59202=>"001000011",
  59203=>"110110101",
  59204=>"000010011",
  59205=>"111111011",
  59206=>"101001001",
  59207=>"111100010",
  59208=>"101011100",
  59209=>"000100000",
  59210=>"001110111",
  59211=>"010100100",
  59212=>"100110001",
  59213=>"010010110",
  59214=>"001110011",
  59215=>"100000001",
  59216=>"000101010",
  59217=>"110111011",
  59218=>"110000000",
  59219=>"000011110",
  59220=>"011100000",
  59221=>"001000000",
  59222=>"101100001",
  59223=>"100000101",
  59224=>"001001011",
  59225=>"110011111",
  59226=>"110110001",
  59227=>"000111111",
  59228=>"111001101",
  59229=>"000011001",
  59230=>"101011010",
  59231=>"111001010",
  59232=>"100111110",
  59233=>"111000010",
  59234=>"001011010",
  59235=>"101010001",
  59236=>"001101010",
  59237=>"011010001",
  59238=>"001001001",
  59239=>"110101000",
  59240=>"111100100",
  59241=>"111100111",
  59242=>"101011101",
  59243=>"101100110",
  59244=>"011101001",
  59245=>"110011000",
  59246=>"011011010",
  59247=>"101111110",
  59248=>"001011000",
  59249=>"100000101",
  59250=>"111110111",
  59251=>"001111011",
  59252=>"110100011",
  59253=>"000000111",
  59254=>"100111101",
  59255=>"101001000",
  59256=>"010111011",
  59257=>"000001000",
  59258=>"110101111",
  59259=>"000101000",
  59260=>"001110011",
  59261=>"100001010",
  59262=>"001111010",
  59263=>"010111000",
  59264=>"010111110",
  59265=>"100101000",
  59266=>"101111000",
  59267=>"101001101",
  59268=>"100011110",
  59269=>"001101101",
  59270=>"000101101",
  59271=>"011110001",
  59272=>"001011100",
  59273=>"000000010",
  59274=>"100111011",
  59275=>"011010111",
  59276=>"110100010",
  59277=>"010101110",
  59278=>"111111000",
  59279=>"000011011",
  59280=>"111010001",
  59281=>"000101011",
  59282=>"111100101",
  59283=>"110000111",
  59284=>"011111010",
  59285=>"101101110",
  59286=>"110000011",
  59287=>"110010101",
  59288=>"101001111",
  59289=>"111101100",
  59290=>"111100111",
  59291=>"010110011",
  59292=>"011010100",
  59293=>"111011000",
  59294=>"000000001",
  59295=>"111101100",
  59296=>"010000011",
  59297=>"110001011",
  59298=>"100110000",
  59299=>"100101010",
  59300=>"111011110",
  59301=>"001011011",
  59302=>"111111100",
  59303=>"111110101",
  59304=>"111111101",
  59305=>"000010001",
  59306=>"100111111",
  59307=>"101111011",
  59308=>"101110010",
  59309=>"011011011",
  59310=>"000111001",
  59311=>"100000010",
  59312=>"001010110",
  59313=>"101001111",
  59314=>"000000001",
  59315=>"001001110",
  59316=>"000000001",
  59317=>"001111011",
  59318=>"000001110",
  59319=>"010111100",
  59320=>"000001101",
  59321=>"100110111",
  59322=>"101010110",
  59323=>"000010101",
  59324=>"110010000",
  59325=>"101000101",
  59326=>"111011010",
  59327=>"110000000",
  59328=>"110101010",
  59329=>"100101101",
  59330=>"011100010",
  59331=>"011001000",
  59332=>"100100010",
  59333=>"011111000",
  59334=>"101010101",
  59335=>"101001010",
  59336=>"010011011",
  59337=>"100101101",
  59338=>"100010010",
  59339=>"000000111",
  59340=>"010101011",
  59341=>"101001011",
  59342=>"001000000",
  59343=>"101001101",
  59344=>"011001111",
  59345=>"101101001",
  59346=>"011101100",
  59347=>"111001100",
  59348=>"001001111",
  59349=>"000111010",
  59350=>"011000001",
  59351=>"101010101",
  59352=>"111100100",
  59353=>"101111010",
  59354=>"111111000",
  59355=>"101101010",
  59356=>"010000000",
  59357=>"011000000",
  59358=>"111100101",
  59359=>"000000010",
  59360=>"100100111",
  59361=>"011010001",
  59362=>"111010001",
  59363=>"110101001",
  59364=>"100010100",
  59365=>"000000100",
  59366=>"010001101",
  59367=>"110101011",
  59368=>"001010110",
  59369=>"011010001",
  59370=>"011101111",
  59371=>"100011001",
  59372=>"101001001",
  59373=>"110010010",
  59374=>"000001011",
  59375=>"000000000",
  59376=>"111000010",
  59377=>"101000101",
  59378=>"011101111",
  59379=>"010111110",
  59380=>"101001110",
  59381=>"000110000",
  59382=>"101001100",
  59383=>"111110000",
  59384=>"001000001",
  59385=>"001100110",
  59386=>"001010001",
  59387=>"001000010",
  59388=>"000111110",
  59389=>"101100010",
  59390=>"011100100",
  59391=>"101000101",
  59392=>"100100111",
  59393=>"000000100",
  59394=>"001001011",
  59395=>"011000010",
  59396=>"100110011",
  59397=>"010010010",
  59398=>"010101111",
  59399=>"110010101",
  59400=>"111010000",
  59401=>"010010110",
  59402=>"001111001",
  59403=>"010011100",
  59404=>"001000110",
  59405=>"001101011",
  59406=>"101001000",
  59407=>"001001101",
  59408=>"010011111",
  59409=>"111011000",
  59410=>"110011000",
  59411=>"100100110",
  59412=>"101011010",
  59413=>"111010110",
  59414=>"000110011",
  59415=>"011001000",
  59416=>"100001110",
  59417=>"001010100",
  59418=>"011100111",
  59419=>"101001000",
  59420=>"000101010",
  59421=>"110011010",
  59422=>"111001000",
  59423=>"110110001",
  59424=>"000100110",
  59425=>"111110000",
  59426=>"111100101",
  59427=>"010110011",
  59428=>"100100111",
  59429=>"101010101",
  59430=>"101100100",
  59431=>"001100010",
  59432=>"001000001",
  59433=>"110010100",
  59434=>"010001011",
  59435=>"001000010",
  59436=>"000110100",
  59437=>"100000010",
  59438=>"010010100",
  59439=>"000001100",
  59440=>"000001001",
  59441=>"111010110",
  59442=>"000111110",
  59443=>"011001111",
  59444=>"011100110",
  59445=>"101010001",
  59446=>"010100000",
  59447=>"001100101",
  59448=>"111100000",
  59449=>"000000100",
  59450=>"011110111",
  59451=>"111101111",
  59452=>"000000111",
  59453=>"001111100",
  59454=>"100011110",
  59455=>"001110000",
  59456=>"111010001",
  59457=>"100011000",
  59458=>"000100101",
  59459=>"111001000",
  59460=>"010000110",
  59461=>"001111010",
  59462=>"000111111",
  59463=>"100101010",
  59464=>"100010101",
  59465=>"100111001",
  59466=>"000000011",
  59467=>"000101001",
  59468=>"101110011",
  59469=>"100000000",
  59470=>"110101111",
  59471=>"101111011",
  59472=>"111001010",
  59473=>"010010000",
  59474=>"100000110",
  59475=>"101111100",
  59476=>"111001101",
  59477=>"011101000",
  59478=>"001101101",
  59479=>"101111111",
  59480=>"111010011",
  59481=>"000111000",
  59482=>"100111010",
  59483=>"100100001",
  59484=>"100100110",
  59485=>"001111101",
  59486=>"010110111",
  59487=>"111000111",
  59488=>"010001010",
  59489=>"111100010",
  59490=>"011010111",
  59491=>"100110111",
  59492=>"010110100",
  59493=>"000010111",
  59494=>"010101010",
  59495=>"010100001",
  59496=>"110111001",
  59497=>"000101010",
  59498=>"100101100",
  59499=>"010101001",
  59500=>"101001000",
  59501=>"000110111",
  59502=>"010010000",
  59503=>"010111111",
  59504=>"101110001",
  59505=>"001010001",
  59506=>"110111010",
  59507=>"100101101",
  59508=>"110111000",
  59509=>"110001110",
  59510=>"000111000",
  59511=>"100111101",
  59512=>"011001011",
  59513=>"111111100",
  59514=>"001001101",
  59515=>"100001010",
  59516=>"101100011",
  59517=>"100100111",
  59518=>"110000011",
  59519=>"100001010",
  59520=>"011101000",
  59521=>"110101101",
  59522=>"101001101",
  59523=>"111110011",
  59524=>"010000000",
  59525=>"011111101",
  59526=>"001010010",
  59527=>"000100011",
  59528=>"101101001",
  59529=>"110000010",
  59530=>"111000011",
  59531=>"000110111",
  59532=>"111100010",
  59533=>"100010010",
  59534=>"011100101",
  59535=>"001100011",
  59536=>"111101111",
  59537=>"010010111",
  59538=>"111111011",
  59539=>"101000011",
  59540=>"010010001",
  59541=>"010111011",
  59542=>"001010111",
  59543=>"010000110",
  59544=>"111000010",
  59545=>"000000010",
  59546=>"000101010",
  59547=>"111011000",
  59548=>"010110111",
  59549=>"010111110",
  59550=>"100111111",
  59551=>"111110101",
  59552=>"010101010",
  59553=>"001000111",
  59554=>"111100000",
  59555=>"010000000",
  59556=>"000011001",
  59557=>"010000110",
  59558=>"001011111",
  59559=>"101000001",
  59560=>"111100001",
  59561=>"000110001",
  59562=>"111011110",
  59563=>"101101010",
  59564=>"111001011",
  59565=>"101110100",
  59566=>"000100011",
  59567=>"110011110",
  59568=>"101001011",
  59569=>"100110000",
  59570=>"010110010",
  59571=>"010000101",
  59572=>"111101111",
  59573=>"010011111",
  59574=>"010010110",
  59575=>"011010000",
  59576=>"101001010",
  59577=>"001110001",
  59578=>"011001001",
  59579=>"100111010",
  59580=>"101000100",
  59581=>"100100011",
  59582=>"001100010",
  59583=>"100101101",
  59584=>"101110010",
  59585=>"100001001",
  59586=>"001110111",
  59587=>"001011011",
  59588=>"001111111",
  59589=>"001000101",
  59590=>"111001000",
  59591=>"000100111",
  59592=>"001111110",
  59593=>"111111001",
  59594=>"101001000",
  59595=>"001001000",
  59596=>"110011101",
  59597=>"111010110",
  59598=>"001111111",
  59599=>"011111101",
  59600=>"010101100",
  59601=>"100010110",
  59602=>"111000001",
  59603=>"001101100",
  59604=>"011100010",
  59605=>"011110011",
  59606=>"001001000",
  59607=>"000010010",
  59608=>"101100101",
  59609=>"101100010",
  59610=>"000011001",
  59611=>"001011100",
  59612=>"110100101",
  59613=>"000000110",
  59614=>"001001000",
  59615=>"101100111",
  59616=>"001010001",
  59617=>"000001100",
  59618=>"111101011",
  59619=>"110000000",
  59620=>"010110101",
  59621=>"011011101",
  59622=>"101000000",
  59623=>"101110000",
  59624=>"010110001",
  59625=>"110111001",
  59626=>"000010111",
  59627=>"110110111",
  59628=>"111111000",
  59629=>"011101101",
  59630=>"010100001",
  59631=>"000000101",
  59632=>"100001101",
  59633=>"110001101",
  59634=>"101001110",
  59635=>"100100101",
  59636=>"101111111",
  59637=>"101000000",
  59638=>"001000000",
  59639=>"001110000",
  59640=>"100101101",
  59641=>"110000011",
  59642=>"011111010",
  59643=>"001000010",
  59644=>"011100101",
  59645=>"000100100",
  59646=>"111110110",
  59647=>"000111001",
  59648=>"011000101",
  59649=>"111100000",
  59650=>"010100110",
  59651=>"110000000",
  59652=>"001011111",
  59653=>"101111101",
  59654=>"000000101",
  59655=>"101010111",
  59656=>"011000011",
  59657=>"110011101",
  59658=>"110011000",
  59659=>"010110000",
  59660=>"111100110",
  59661=>"100110100",
  59662=>"000100001",
  59663=>"000111000",
  59664=>"101111011",
  59665=>"100010001",
  59666=>"001010111",
  59667=>"110111001",
  59668=>"000000011",
  59669=>"010101100",
  59670=>"101000000",
  59671=>"110001000",
  59672=>"001011011",
  59673=>"100000111",
  59674=>"110100000",
  59675=>"100011000",
  59676=>"001000000",
  59677=>"111011010",
  59678=>"001000110",
  59679=>"010011011",
  59680=>"100100100",
  59681=>"111100111",
  59682=>"001011110",
  59683=>"001010000",
  59684=>"001111010",
  59685=>"101110010",
  59686=>"111011000",
  59687=>"011110001",
  59688=>"011010001",
  59689=>"010001001",
  59690=>"000101011",
  59691=>"000000111",
  59692=>"111000111",
  59693=>"100000011",
  59694=>"001000011",
  59695=>"011011111",
  59696=>"001001010",
  59697=>"100110111",
  59698=>"011100101",
  59699=>"101010011",
  59700=>"010111110",
  59701=>"101101000",
  59702=>"110001110",
  59703=>"011101011",
  59704=>"110000011",
  59705=>"001011100",
  59706=>"011101110",
  59707=>"001010010",
  59708=>"100000000",
  59709=>"000010000",
  59710=>"110100101",
  59711=>"101101010",
  59712=>"011001000",
  59713=>"000111111",
  59714=>"100110111",
  59715=>"110100000",
  59716=>"001010111",
  59717=>"100100100",
  59718=>"011101011",
  59719=>"000100001",
  59720=>"100111101",
  59721=>"010011000",
  59722=>"110100110",
  59723=>"001001010",
  59724=>"000000011",
  59725=>"011110110",
  59726=>"010011011",
  59727=>"100000101",
  59728=>"110100000",
  59729=>"111010000",
  59730=>"100001001",
  59731=>"100111100",
  59732=>"110110010",
  59733=>"000101110",
  59734=>"011110000",
  59735=>"101001010",
  59736=>"101000010",
  59737=>"001000000",
  59738=>"111011010",
  59739=>"101101101",
  59740=>"010001010",
  59741=>"101010101",
  59742=>"111011110",
  59743=>"100011111",
  59744=>"001110000",
  59745=>"011010111",
  59746=>"110101100",
  59747=>"100100110",
  59748=>"100110011",
  59749=>"011001001",
  59750=>"000110010",
  59751=>"000011110",
  59752=>"110100001",
  59753=>"011101001",
  59754=>"000101010",
  59755=>"000001110",
  59756=>"100001001",
  59757=>"001111100",
  59758=>"111111001",
  59759=>"010001010",
  59760=>"010110011",
  59761=>"000011010",
  59762=>"110010011",
  59763=>"000000000",
  59764=>"100100010",
  59765=>"101011100",
  59766=>"100000111",
  59767=>"000000011",
  59768=>"001011001",
  59769=>"111010001",
  59770=>"011011001",
  59771=>"011011011",
  59772=>"001101101",
  59773=>"111110110",
  59774=>"010001010",
  59775=>"110110111",
  59776=>"001100000",
  59777=>"110101000",
  59778=>"001101111",
  59779=>"000001000",
  59780=>"110001001",
  59781=>"000010000",
  59782=>"010011100",
  59783=>"011010111",
  59784=>"011011000",
  59785=>"110000000",
  59786=>"011000000",
  59787=>"010001010",
  59788=>"110001110",
  59789=>"100100110",
  59790=>"110000011",
  59791=>"110110100",
  59792=>"110101000",
  59793=>"011011110",
  59794=>"011011000",
  59795=>"001100001",
  59796=>"100111010",
  59797=>"010100101",
  59798=>"000111011",
  59799=>"111110101",
  59800=>"011111101",
  59801=>"000100001",
  59802=>"111000101",
  59803=>"110100110",
  59804=>"111001011",
  59805=>"000011111",
  59806=>"001100010",
  59807=>"011100000",
  59808=>"110100100",
  59809=>"101001101",
  59810=>"001111101",
  59811=>"000001101",
  59812=>"000000001",
  59813=>"100000010",
  59814=>"010101010",
  59815=>"110101011",
  59816=>"011000001",
  59817=>"101100001",
  59818=>"100100000",
  59819=>"100011000",
  59820=>"010111000",
  59821=>"100001110",
  59822=>"010101001",
  59823=>"111110011",
  59824=>"100111001",
  59825=>"001011010",
  59826=>"001100110",
  59827=>"010000000",
  59828=>"000101010",
  59829=>"001011110",
  59830=>"011110110",
  59831=>"001010101",
  59832=>"111111110",
  59833=>"010010100",
  59834=>"001011001",
  59835=>"110110110",
  59836=>"100001011",
  59837=>"100101110",
  59838=>"001100011",
  59839=>"010010101",
  59840=>"000100011",
  59841=>"100111010",
  59842=>"110100011",
  59843=>"101010000",
  59844=>"111101011",
  59845=>"111100001",
  59846=>"001011001",
  59847=>"011111010",
  59848=>"001101111",
  59849=>"101100110",
  59850=>"110101101",
  59851=>"001100000",
  59852=>"010011011",
  59853=>"000001100",
  59854=>"100010001",
  59855=>"000110000",
  59856=>"001011000",
  59857=>"000011100",
  59858=>"101110110",
  59859=>"011010011",
  59860=>"000110100",
  59861=>"010111101",
  59862=>"111001000",
  59863=>"010110010",
  59864=>"000111000",
  59865=>"100100010",
  59866=>"011011000",
  59867=>"111100010",
  59868=>"011011111",
  59869=>"010111100",
  59870=>"011101111",
  59871=>"101001111",
  59872=>"000011011",
  59873=>"100011101",
  59874=>"101001001",
  59875=>"110001000",
  59876=>"001000111",
  59877=>"010100000",
  59878=>"100100100",
  59879=>"010101000",
  59880=>"011010110",
  59881=>"110010111",
  59882=>"101000000",
  59883=>"001111001",
  59884=>"010000010",
  59885=>"001010000",
  59886=>"110101110",
  59887=>"110100110",
  59888=>"000111010",
  59889=>"000001101",
  59890=>"011011101",
  59891=>"001100101",
  59892=>"000101011",
  59893=>"101101010",
  59894=>"011010101",
  59895=>"100011101",
  59896=>"000001100",
  59897=>"111011010",
  59898=>"010111000",
  59899=>"011111010",
  59900=>"110011111",
  59901=>"010000111",
  59902=>"001100100",
  59903=>"110101110",
  59904=>"100010100",
  59905=>"000110110",
  59906=>"000011101",
  59907=>"000010000",
  59908=>"000101100",
  59909=>"110100100",
  59910=>"110110100",
  59911=>"011000101",
  59912=>"011111001",
  59913=>"100111001",
  59914=>"100001010",
  59915=>"000110101",
  59916=>"101101000",
  59917=>"001101000",
  59918=>"000010000",
  59919=>"110001000",
  59920=>"100001001",
  59921=>"000001110",
  59922=>"000001110",
  59923=>"111111000",
  59924=>"100001011",
  59925=>"111111001",
  59926=>"111100001",
  59927=>"010100000",
  59928=>"100100011",
  59929=>"011011111",
  59930=>"101111101",
  59931=>"001110010",
  59932=>"010000101",
  59933=>"111011010",
  59934=>"111011111",
  59935=>"010010010",
  59936=>"010000101",
  59937=>"101100101",
  59938=>"000000000",
  59939=>"000110001",
  59940=>"110001101",
  59941=>"011001101",
  59942=>"100001010",
  59943=>"000110110",
  59944=>"011110110",
  59945=>"110101101",
  59946=>"001111011",
  59947=>"000110110",
  59948=>"101010001",
  59949=>"010001110",
  59950=>"100000001",
  59951=>"010010010",
  59952=>"100110110",
  59953=>"110010011",
  59954=>"000000101",
  59955=>"001110001",
  59956=>"001101000",
  59957=>"000010100",
  59958=>"100101011",
  59959=>"100101101",
  59960=>"101010001",
  59961=>"110110010",
  59962=>"100110101",
  59963=>"011110011",
  59964=>"001010010",
  59965=>"011011000",
  59966=>"110001000",
  59967=>"011000000",
  59968=>"111111111",
  59969=>"011101111",
  59970=>"100110101",
  59971=>"101101101",
  59972=>"110011001",
  59973=>"101100001",
  59974=>"111011100",
  59975=>"001010001",
  59976=>"100111100",
  59977=>"110100101",
  59978=>"111100100",
  59979=>"100101111",
  59980=>"010000011",
  59981=>"001000000",
  59982=>"111100111",
  59983=>"110111010",
  59984=>"100011001",
  59985=>"101000111",
  59986=>"011100111",
  59987=>"011100110",
  59988=>"100100111",
  59989=>"110000001",
  59990=>"110101100",
  59991=>"100011100",
  59992=>"011110100",
  59993=>"111100111",
  59994=>"001101111",
  59995=>"001000110",
  59996=>"111100011",
  59997=>"111011010",
  59998=>"100000001",
  59999=>"110101110",
  60000=>"100101001",
  60001=>"111011110",
  60002=>"001110010",
  60003=>"000101011",
  60004=>"110111010",
  60005=>"111001101",
  60006=>"001011110",
  60007=>"001111101",
  60008=>"111110110",
  60009=>"110011111",
  60010=>"110010011",
  60011=>"110001011",
  60012=>"000101010",
  60013=>"100101000",
  60014=>"000100010",
  60015=>"000110000",
  60016=>"111000000",
  60017=>"000111001",
  60018=>"111000111",
  60019=>"110111000",
  60020=>"000011011",
  60021=>"111110100",
  60022=>"111101101",
  60023=>"111100011",
  60024=>"001111111",
  60025=>"001100101",
  60026=>"110011100",
  60027=>"010110010",
  60028=>"000010010",
  60029=>"101010001",
  60030=>"000101101",
  60031=>"111110111",
  60032=>"100111111",
  60033=>"011000110",
  60034=>"111000100",
  60035=>"101101001",
  60036=>"101101111",
  60037=>"100011010",
  60038=>"110011100",
  60039=>"111111010",
  60040=>"011100010",
  60041=>"100001100",
  60042=>"100001111",
  60043=>"001111100",
  60044=>"101100000",
  60045=>"101100101",
  60046=>"110001010",
  60047=>"111001001",
  60048=>"101010000",
  60049=>"000111011",
  60050=>"101001001",
  60051=>"010100110",
  60052=>"101111111",
  60053=>"101001001",
  60054=>"110110010",
  60055=>"001110000",
  60056=>"000110000",
  60057=>"011111000",
  60058=>"011110001",
  60059=>"110011111",
  60060=>"111010011",
  60061=>"100111101",
  60062=>"110101010",
  60063=>"001100100",
  60064=>"110101000",
  60065=>"000101110",
  60066=>"001100010",
  60067=>"101000101",
  60068=>"010011001",
  60069=>"011011011",
  60070=>"011010101",
  60071=>"011000010",
  60072=>"110010000",
  60073=>"101001011",
  60074=>"001001101",
  60075=>"000101111",
  60076=>"011100111",
  60077=>"110000000",
  60078=>"100010011",
  60079=>"001011011",
  60080=>"010001001",
  60081=>"100100001",
  60082=>"110001101",
  60083=>"101000110",
  60084=>"011000000",
  60085=>"011101001",
  60086=>"001110111",
  60087=>"001101110",
  60088=>"101010011",
  60089=>"110110110",
  60090=>"100000111",
  60091=>"100001110",
  60092=>"010110000",
  60093=>"111100100",
  60094=>"000101000",
  60095=>"111001000",
  60096=>"101110101",
  60097=>"000001101",
  60098=>"101111100",
  60099=>"010101000",
  60100=>"101001010",
  60101=>"000010000",
  60102=>"101110001",
  60103=>"100000100",
  60104=>"111110100",
  60105=>"101001101",
  60106=>"000001001",
  60107=>"001110110",
  60108=>"000001100",
  60109=>"110011111",
  60110=>"000010110",
  60111=>"010011111",
  60112=>"111111010",
  60113=>"110110011",
  60114=>"010111000",
  60115=>"110000001",
  60116=>"100001001",
  60117=>"101010110",
  60118=>"010110001",
  60119=>"010101010",
  60120=>"000010111",
  60121=>"000011100",
  60122=>"000010011",
  60123=>"101101100",
  60124=>"000100011",
  60125=>"110010110",
  60126=>"011011110",
  60127=>"111011010",
  60128=>"000011101",
  60129=>"110101101",
  60130=>"100110111",
  60131=>"111001011",
  60132=>"101001001",
  60133=>"000110011",
  60134=>"111011111",
  60135=>"110000010",
  60136=>"111111111",
  60137=>"000111110",
  60138=>"011100011",
  60139=>"010011011",
  60140=>"101110100",
  60141=>"101101101",
  60142=>"110000111",
  60143=>"011111100",
  60144=>"001011010",
  60145=>"101110100",
  60146=>"101100010",
  60147=>"101001110",
  60148=>"110000100",
  60149=>"111010100",
  60150=>"111110011",
  60151=>"010000011",
  60152=>"101101000",
  60153=>"010001000",
  60154=>"011100011",
  60155=>"000110000",
  60156=>"011011101",
  60157=>"001000000",
  60158=>"011011001",
  60159=>"110010100",
  60160=>"010001100",
  60161=>"011100001",
  60162=>"010100100",
  60163=>"001101111",
  60164=>"110111001",
  60165=>"011010111",
  60166=>"000000111",
  60167=>"000010001",
  60168=>"110000000",
  60169=>"001101111",
  60170=>"000111011",
  60171=>"100011101",
  60172=>"110011111",
  60173=>"000011111",
  60174=>"011111111",
  60175=>"110010110",
  60176=>"001110111",
  60177=>"100010001",
  60178=>"001100101",
  60179=>"100101111",
  60180=>"110001010",
  60181=>"101000110",
  60182=>"011111001",
  60183=>"101010101",
  60184=>"011000010",
  60185=>"110110111",
  60186=>"000000100",
  60187=>"010001010",
  60188=>"111111010",
  60189=>"011101110",
  60190=>"000010000",
  60191=>"010001000",
  60192=>"101101101",
  60193=>"000001001",
  60194=>"011111101",
  60195=>"111101000",
  60196=>"111011110",
  60197=>"000010000",
  60198=>"101100001",
  60199=>"111111000",
  60200=>"010011111",
  60201=>"101101111",
  60202=>"100101100",
  60203=>"000110011",
  60204=>"010101111",
  60205=>"001000010",
  60206=>"000011100",
  60207=>"010011100",
  60208=>"011000111",
  60209=>"010001111",
  60210=>"010011111",
  60211=>"111110110",
  60212=>"111011101",
  60213=>"110010001",
  60214=>"111010101",
  60215=>"110010001",
  60216=>"101111010",
  60217=>"001011010",
  60218=>"000100101",
  60219=>"111011000",
  60220=>"111101010",
  60221=>"111001000",
  60222=>"000000101",
  60223=>"110010100",
  60224=>"000100000",
  60225=>"010110010",
  60226=>"111101011",
  60227=>"011111101",
  60228=>"110000010",
  60229=>"001110111",
  60230=>"011011100",
  60231=>"110111110",
  60232=>"000110010",
  60233=>"111000000",
  60234=>"100100010",
  60235=>"001010010",
  60236=>"101110111",
  60237=>"010010010",
  60238=>"110111101",
  60239=>"010001000",
  60240=>"101101101",
  60241=>"110010111",
  60242=>"010111010",
  60243=>"101101111",
  60244=>"100001011",
  60245=>"001000001",
  60246=>"101000110",
  60247=>"111001101",
  60248=>"110001011",
  60249=>"000001001",
  60250=>"111100111",
  60251=>"100100000",
  60252=>"100111111",
  60253=>"000011110",
  60254=>"000111101",
  60255=>"000000000",
  60256=>"010101101",
  60257=>"101001111",
  60258=>"011100111",
  60259=>"101001000",
  60260=>"100100100",
  60261=>"010111110",
  60262=>"011111000",
  60263=>"000001010",
  60264=>"100010010",
  60265=>"010001000",
  60266=>"011001101",
  60267=>"111110010",
  60268=>"001101111",
  60269=>"100010110",
  60270=>"110100001",
  60271=>"011001010",
  60272=>"100100101",
  60273=>"011011110",
  60274=>"100110010",
  60275=>"111010010",
  60276=>"110000000",
  60277=>"001101110",
  60278=>"111011011",
  60279=>"010000001",
  60280=>"010011101",
  60281=>"110111010",
  60282=>"010101110",
  60283=>"010001101",
  60284=>"001010000",
  60285=>"010111010",
  60286=>"101010010",
  60287=>"101111010",
  60288=>"110010011",
  60289=>"110111111",
  60290=>"111010000",
  60291=>"011111111",
  60292=>"010011111",
  60293=>"010011011",
  60294=>"111000110",
  60295=>"001001111",
  60296=>"101010111",
  60297=>"100000100",
  60298=>"011101110",
  60299=>"010100010",
  60300=>"001010000",
  60301=>"001101011",
  60302=>"001100101",
  60303=>"010010010",
  60304=>"000110111",
  60305=>"011000111",
  60306=>"011110011",
  60307=>"011101001",
  60308=>"010000000",
  60309=>"000101000",
  60310=>"001000001",
  60311=>"101111101",
  60312=>"000000111",
  60313=>"100010100",
  60314=>"000001011",
  60315=>"111110000",
  60316=>"010001000",
  60317=>"100010011",
  60318=>"100010011",
  60319=>"011101011",
  60320=>"100011101",
  60321=>"010001111",
  60322=>"010011110",
  60323=>"011011011",
  60324=>"011101001",
  60325=>"111111101",
  60326=>"100100111",
  60327=>"101111101",
  60328=>"001110110",
  60329=>"111101101",
  60330=>"011010101",
  60331=>"010111010",
  60332=>"001000110",
  60333=>"010000101",
  60334=>"101101101",
  60335=>"000011001",
  60336=>"011000100",
  60337=>"100010011",
  60338=>"011111101",
  60339=>"000000110",
  60340=>"100000000",
  60341=>"010010010",
  60342=>"110101101",
  60343=>"100011011",
  60344=>"110001011",
  60345=>"110101011",
  60346=>"110100001",
  60347=>"101000101",
  60348=>"111010001",
  60349=>"010101010",
  60350=>"001011101",
  60351=>"110101100",
  60352=>"111000101",
  60353=>"000000000",
  60354=>"111110100",
  60355=>"100011100",
  60356=>"000100111",
  60357=>"101111001",
  60358=>"000011011",
  60359=>"010011000",
  60360=>"000010000",
  60361=>"001111001",
  60362=>"001101000",
  60363=>"011100011",
  60364=>"110011011",
  60365=>"111100000",
  60366=>"110000110",
  60367=>"001001110",
  60368=>"010010101",
  60369=>"010111011",
  60370=>"001010010",
  60371=>"100001110",
  60372=>"100000011",
  60373=>"010000100",
  60374=>"111000010",
  60375=>"110001110",
  60376=>"100000110",
  60377=>"111101010",
  60378=>"001110011",
  60379=>"000001010",
  60380=>"000010001",
  60381=>"000111011",
  60382=>"100001101",
  60383=>"100010001",
  60384=>"110101111",
  60385=>"100000010",
  60386=>"101100000",
  60387=>"001010000",
  60388=>"001010010",
  60389=>"111000111",
  60390=>"001111011",
  60391=>"000010011",
  60392=>"001111110",
  60393=>"010100010",
  60394=>"111101101",
  60395=>"111000000",
  60396=>"011011001",
  60397=>"101000010",
  60398=>"111101010",
  60399=>"011000011",
  60400=>"000011110",
  60401=>"000101101",
  60402=>"011100111",
  60403=>"010000010",
  60404=>"101010000",
  60405=>"111000001",
  60406=>"110110100",
  60407=>"101010101",
  60408=>"001000011",
  60409=>"101111101",
  60410=>"011010010",
  60411=>"011000100",
  60412=>"000000010",
  60413=>"100110101",
  60414=>"101111011",
  60415=>"110001001",
  60416=>"000001000",
  60417=>"100111001",
  60418=>"010110110",
  60419=>"010000000",
  60420=>"010110111",
  60421=>"111001110",
  60422=>"111001000",
  60423=>"100010100",
  60424=>"011101001",
  60425=>"110110010",
  60426=>"000011111",
  60427=>"100101001",
  60428=>"111001101",
  60429=>"110100000",
  60430=>"111100100",
  60431=>"000000001",
  60432=>"101111111",
  60433=>"010110100",
  60434=>"101000100",
  60435=>"111001001",
  60436=>"010000001",
  60437=>"001111100",
  60438=>"111010101",
  60439=>"000001110",
  60440=>"110000000",
  60441=>"000100010",
  60442=>"100101000",
  60443=>"000010100",
  60444=>"010010101",
  60445=>"010001100",
  60446=>"001111111",
  60447=>"111011101",
  60448=>"110101000",
  60449=>"001000001",
  60450=>"111000110",
  60451=>"000100100",
  60452=>"101011100",
  60453=>"001100101",
  60454=>"010001011",
  60455=>"111100010",
  60456=>"000111011",
  60457=>"000000110",
  60458=>"100011001",
  60459=>"100101001",
  60460=>"000100011",
  60461=>"111001010",
  60462=>"101111011",
  60463=>"011111110",
  60464=>"000011000",
  60465=>"101000100",
  60466=>"101001101",
  60467=>"101101111",
  60468=>"111110111",
  60469=>"001001100",
  60470=>"110001100",
  60471=>"101011011",
  60472=>"100011001",
  60473=>"010000110",
  60474=>"010100100",
  60475=>"110111111",
  60476=>"001101000",
  60477=>"000100011",
  60478=>"101001000",
  60479=>"001001100",
  60480=>"001110000",
  60481=>"000011001",
  60482=>"110110110",
  60483=>"111101010",
  60484=>"100111011",
  60485=>"111000001",
  60486=>"110000110",
  60487=>"000010111",
  60488=>"010010111",
  60489=>"110100010",
  60490=>"000010000",
  60491=>"001010011",
  60492=>"011101010",
  60493=>"011110100",
  60494=>"000010010",
  60495=>"001010010",
  60496=>"100110110",
  60497=>"000001110",
  60498=>"110111111",
  60499=>"101010111",
  60500=>"111110010",
  60501=>"111000101",
  60502=>"010010100",
  60503=>"110111010",
  60504=>"010111010",
  60505=>"100110010",
  60506=>"110001001",
  60507=>"110000011",
  60508=>"001000110",
  60509=>"101111110",
  60510=>"100011111",
  60511=>"101101000",
  60512=>"010000000",
  60513=>"101100011",
  60514=>"001001111",
  60515=>"111101110",
  60516=>"010010010",
  60517=>"010000100",
  60518=>"010010000",
  60519=>"101110110",
  60520=>"001111111",
  60521=>"001111110",
  60522=>"111011111",
  60523=>"000010001",
  60524=>"110111010",
  60525=>"000000011",
  60526=>"100001110",
  60527=>"110110000",
  60528=>"011000111",
  60529=>"100100111",
  60530=>"000100001",
  60531=>"111110110",
  60532=>"001100011",
  60533=>"110100111",
  60534=>"001000101",
  60535=>"010110011",
  60536=>"010100110",
  60537=>"011101000",
  60538=>"100101111",
  60539=>"000100001",
  60540=>"000100000",
  60541=>"010001100",
  60542=>"011000000",
  60543=>"101111000",
  60544=>"000101001",
  60545=>"011010001",
  60546=>"001111111",
  60547=>"010010110",
  60548=>"001110010",
  60549=>"100001010",
  60550=>"000101110",
  60551=>"001110010",
  60552=>"010010101",
  60553=>"001101001",
  60554=>"100000011",
  60555=>"111010001",
  60556=>"011000111",
  60557=>"111011010",
  60558=>"111110010",
  60559=>"001111111",
  60560=>"011111010",
  60561=>"100111011",
  60562=>"111111010",
  60563=>"010110001",
  60564=>"110101000",
  60565=>"111100000",
  60566=>"101010101",
  60567=>"110001111",
  60568=>"100101100",
  60569=>"000000101",
  60570=>"010011010",
  60571=>"001110011",
  60572=>"001010111",
  60573=>"101011100",
  60574=>"000100100",
  60575=>"001101100",
  60576=>"001110100",
  60577=>"010100011",
  60578=>"000000001",
  60579=>"100010101",
  60580=>"010001001",
  60581=>"100110101",
  60582=>"010010011",
  60583=>"001001110",
  60584=>"001100010",
  60585=>"111000000",
  60586=>"011000101",
  60587=>"101001101",
  60588=>"001011110",
  60589=>"010001100",
  60590=>"011001101",
  60591=>"001000000",
  60592=>"101101010",
  60593=>"011010110",
  60594=>"111001001",
  60595=>"100100111",
  60596=>"110011101",
  60597=>"110000100",
  60598=>"011000001",
  60599=>"000100000",
  60600=>"010100111",
  60601=>"101010101",
  60602=>"000111001",
  60603=>"010011010",
  60604=>"111000110",
  60605=>"000100001",
  60606=>"100010111",
  60607=>"011010110",
  60608=>"000010011",
  60609=>"110101110",
  60610=>"101100110",
  60611=>"101010011",
  60612=>"101110100",
  60613=>"101101100",
  60614=>"011010111",
  60615=>"110100010",
  60616=>"111010001",
  60617=>"111011110",
  60618=>"111110111",
  60619=>"101111110",
  60620=>"011110111",
  60621=>"011110000",
  60622=>"101111100",
  60623=>"011111100",
  60624=>"110101111",
  60625=>"010011100",
  60626=>"111000001",
  60627=>"111011000",
  60628=>"011111001",
  60629=>"011001001",
  60630=>"011011100",
  60631=>"111110110",
  60632=>"101000001",
  60633=>"000110010",
  60634=>"010101011",
  60635=>"000101010",
  60636=>"111001000",
  60637=>"000011100",
  60638=>"010001111",
  60639=>"110100011",
  60640=>"110001010",
  60641=>"010100100",
  60642=>"011001001",
  60643=>"000010000",
  60644=>"000101000",
  60645=>"010000000",
  60646=>"110101100",
  60647=>"101011110",
  60648=>"000010100",
  60649=>"100001110",
  60650=>"011111110",
  60651=>"001100110",
  60652=>"010001011",
  60653=>"101010111",
  60654=>"001110000",
  60655=>"100101000",
  60656=>"101110011",
  60657=>"101011010",
  60658=>"101011011",
  60659=>"110011100",
  60660=>"011000100",
  60661=>"001000100",
  60662=>"100000101",
  60663=>"000110111",
  60664=>"001000010",
  60665=>"000111101",
  60666=>"111101111",
  60667=>"100000010",
  60668=>"001010001",
  60669=>"100110110",
  60670=>"000100110",
  60671=>"110010000",
  60672=>"001011111",
  60673=>"010101101",
  60674=>"101111000",
  60675=>"000111010",
  60676=>"101100111",
  60677=>"011001001",
  60678=>"001110001",
  60679=>"100000111",
  60680=>"101100001",
  60681=>"101011010",
  60682=>"010011110",
  60683=>"001000111",
  60684=>"011000111",
  60685=>"101011100",
  60686=>"010011001",
  60687=>"111000100",
  60688=>"111100111",
  60689=>"100011111",
  60690=>"001011111",
  60691=>"111110111",
  60692=>"101101111",
  60693=>"110000000",
  60694=>"100111000",
  60695=>"010100100",
  60696=>"111000111",
  60697=>"110011000",
  60698=>"010100110",
  60699=>"111000100",
  60700=>"010011000",
  60701=>"101010000",
  60702=>"100101001",
  60703=>"000110110",
  60704=>"000100000",
  60705=>"110000100",
  60706=>"001001100",
  60707=>"110101110",
  60708=>"000000101",
  60709=>"001111000",
  60710=>"011110000",
  60711=>"101010100",
  60712=>"110000011",
  60713=>"111101110",
  60714=>"101010111",
  60715=>"011101101",
  60716=>"100100110",
  60717=>"111111111",
  60718=>"000001000",
  60719=>"100010010",
  60720=>"110010111",
  60721=>"001100001",
  60722=>"010000100",
  60723=>"100011101",
  60724=>"110000111",
  60725=>"111101000",
  60726=>"101111101",
  60727=>"011011011",
  60728=>"111010101",
  60729=>"110000100",
  60730=>"000010011",
  60731=>"001111101",
  60732=>"011110110",
  60733=>"001001101",
  60734=>"111011111",
  60735=>"101001100",
  60736=>"110011101",
  60737=>"110101111",
  60738=>"001001010",
  60739=>"100000100",
  60740=>"100000010",
  60741=>"000010111",
  60742=>"110010101",
  60743=>"001000110",
  60744=>"100010000",
  60745=>"101001001",
  60746=>"101101000",
  60747=>"100101011",
  60748=>"100100110",
  60749=>"101001010",
  60750=>"001110011",
  60751=>"010011001",
  60752=>"100011000",
  60753=>"001000100",
  60754=>"101011111",
  60755=>"011100111",
  60756=>"001010011",
  60757=>"011011000",
  60758=>"011111010",
  60759=>"101010011",
  60760=>"001101010",
  60761=>"000100100",
  60762=>"111100011",
  60763=>"011101000",
  60764=>"000110111",
  60765=>"110101110",
  60766=>"001111110",
  60767=>"010101101",
  60768=>"111100110",
  60769=>"110011010",
  60770=>"101011111",
  60771=>"000111011",
  60772=>"110111110",
  60773=>"100100110",
  60774=>"000000010",
  60775=>"101101111",
  60776=>"010101100",
  60777=>"000010000",
  60778=>"100111111",
  60779=>"001001100",
  60780=>"101000010",
  60781=>"111101011",
  60782=>"010011011",
  60783=>"110010111",
  60784=>"010101111",
  60785=>"111101110",
  60786=>"100101100",
  60787=>"101100011",
  60788=>"111100101",
  60789=>"010011001",
  60790=>"000110010",
  60791=>"111000101",
  60792=>"011101100",
  60793=>"111101111",
  60794=>"011110001",
  60795=>"100100100",
  60796=>"000110000",
  60797=>"011111001",
  60798=>"001101010",
  60799=>"000011000",
  60800=>"110110101",
  60801=>"011010111",
  60802=>"111001111",
  60803=>"101001000",
  60804=>"110000001",
  60805=>"101011111",
  60806=>"111001101",
  60807=>"000010100",
  60808=>"101111101",
  60809=>"011000110",
  60810=>"100111111",
  60811=>"110011111",
  60812=>"101111001",
  60813=>"110111101",
  60814=>"111101001",
  60815=>"000100111",
  60816=>"000100111",
  60817=>"011110010",
  60818=>"000100001",
  60819=>"010011110",
  60820=>"101001111",
  60821=>"001101101",
  60822=>"011111010",
  60823=>"011010100",
  60824=>"111010110",
  60825=>"000011010",
  60826=>"100000100",
  60827=>"110110100",
  60828=>"111110010",
  60829=>"100000010",
  60830=>"001110110",
  60831=>"110100101",
  60832=>"000001000",
  60833=>"001111111",
  60834=>"000001001",
  60835=>"011110000",
  60836=>"011001101",
  60837=>"110010110",
  60838=>"011000010",
  60839=>"000101111",
  60840=>"010100010",
  60841=>"011111011",
  60842=>"011101110",
  60843=>"111111111",
  60844=>"011100011",
  60845=>"001011101",
  60846=>"101110000",
  60847=>"111100000",
  60848=>"010000101",
  60849=>"100010001",
  60850=>"100100110",
  60851=>"001101011",
  60852=>"110110111",
  60853=>"111101001",
  60854=>"011010111",
  60855=>"010001001",
  60856=>"101011010",
  60857=>"111101101",
  60858=>"100011001",
  60859=>"010110110",
  60860=>"010100000",
  60861=>"101111101",
  60862=>"011010000",
  60863=>"111100010",
  60864=>"001011001",
  60865=>"111101000",
  60866=>"111101001",
  60867=>"110110100",
  60868=>"101001011",
  60869=>"000000010",
  60870=>"101010101",
  60871=>"011011001",
  60872=>"100100010",
  60873=>"000100001",
  60874=>"101101000",
  60875=>"010001100",
  60876=>"100100100",
  60877=>"011101011",
  60878=>"010100111",
  60879=>"101100111",
  60880=>"011010001",
  60881=>"010010100",
  60882=>"101010000",
  60883=>"110101100",
  60884=>"011110010",
  60885=>"101111100",
  60886=>"001001001",
  60887=>"000011000",
  60888=>"010100000",
  60889=>"010111000",
  60890=>"001111110",
  60891=>"111001001",
  60892=>"101100000",
  60893=>"101110001",
  60894=>"001101101",
  60895=>"011000000",
  60896=>"100011110",
  60897=>"101011001",
  60898=>"100001000",
  60899=>"110100010",
  60900=>"100000001",
  60901=>"110000110",
  60902=>"100110111",
  60903=>"010100111",
  60904=>"100111100",
  60905=>"011101001",
  60906=>"000100110",
  60907=>"001100010",
  60908=>"010010001",
  60909=>"001101000",
  60910=>"011101100",
  60911=>"111110000",
  60912=>"000000111",
  60913=>"111101101",
  60914=>"010111000",
  60915=>"111011110",
  60916=>"111001101",
  60917=>"011001001",
  60918=>"000101000",
  60919=>"010111010",
  60920=>"010100100",
  60921=>"100001100",
  60922=>"001011010",
  60923=>"010001100",
  60924=>"111011110",
  60925=>"111111111",
  60926=>"000000100",
  60927=>"010000100",
  60928=>"100001100",
  60929=>"011011001",
  60930=>"010110100",
  60931=>"001111010",
  60932=>"101101011",
  60933=>"001000000",
  60934=>"111111100",
  60935=>"100010010",
  60936=>"001100011",
  60937=>"100010111",
  60938=>"011110111",
  60939=>"100001110",
  60940=>"001100100",
  60941=>"100011000",
  60942=>"010011111",
  60943=>"011010011",
  60944=>"110100111",
  60945=>"110000110",
  60946=>"011011001",
  60947=>"111011111",
  60948=>"111101111",
  60949=>"100111100",
  60950=>"101111001",
  60951=>"111110001",
  60952=>"001000110",
  60953=>"110010100",
  60954=>"010000101",
  60955=>"000111101",
  60956=>"111100100",
  60957=>"010000000",
  60958=>"101101101",
  60959=>"011000101",
  60960=>"000000111",
  60961=>"101010111",
  60962=>"000000011",
  60963=>"110110101",
  60964=>"110000010",
  60965=>"001100011",
  60966=>"101110100",
  60967=>"001100101",
  60968=>"100011110",
  60969=>"001100111",
  60970=>"010110000",
  60971=>"011110000",
  60972=>"011011011",
  60973=>"011011001",
  60974=>"100010011",
  60975=>"101101111",
  60976=>"011000110",
  60977=>"111010000",
  60978=>"011000000",
  60979=>"111101000",
  60980=>"001110000",
  60981=>"101110101",
  60982=>"100000000",
  60983=>"100110000",
  60984=>"110011010",
  60985=>"001000100",
  60986=>"100101001",
  60987=>"010110111",
  60988=>"010101011",
  60989=>"010101001",
  60990=>"000111101",
  60991=>"000000101",
  60992=>"001011110",
  60993=>"010011101",
  60994=>"000010101",
  60995=>"010001011",
  60996=>"000110100",
  60997=>"101110110",
  60998=>"000010110",
  60999=>"110101111",
  61000=>"010000001",
  61001=>"001011110",
  61002=>"111000111",
  61003=>"010010000",
  61004=>"000010001",
  61005=>"001100011",
  61006=>"000110010",
  61007=>"001111100",
  61008=>"111111101",
  61009=>"010110110",
  61010=>"111011111",
  61011=>"000101100",
  61012=>"010110110",
  61013=>"001010000",
  61014=>"011100000",
  61015=>"110010001",
  61016=>"110110000",
  61017=>"101111101",
  61018=>"000001100",
  61019=>"110010100",
  61020=>"000001000",
  61021=>"011110111",
  61022=>"000000001",
  61023=>"100101011",
  61024=>"111101110",
  61025=>"111100100",
  61026=>"001110010",
  61027=>"100101000",
  61028=>"011000000",
  61029=>"010101110",
  61030=>"111010001",
  61031=>"110011111",
  61032=>"011100000",
  61033=>"111001000",
  61034=>"100110111",
  61035=>"111010111",
  61036=>"011001101",
  61037=>"010101010",
  61038=>"000101001",
  61039=>"110101001",
  61040=>"000010000",
  61041=>"110111111",
  61042=>"001111110",
  61043=>"101100001",
  61044=>"010111111",
  61045=>"100010010",
  61046=>"001000010",
  61047=>"001101010",
  61048=>"010101110",
  61049=>"001001011",
  61050=>"011111010",
  61051=>"110001110",
  61052=>"110010101",
  61053=>"101110101",
  61054=>"111111111",
  61055=>"100101001",
  61056=>"011110001",
  61057=>"011010101",
  61058=>"011110011",
  61059=>"000111111",
  61060=>"001101101",
  61061=>"100100001",
  61062=>"100100110",
  61063=>"011111010",
  61064=>"111111101",
  61065=>"001101011",
  61066=>"011000000",
  61067=>"001001110",
  61068=>"011001001",
  61069=>"001010000",
  61070=>"101111100",
  61071=>"000010000",
  61072=>"000101110",
  61073=>"111000101",
  61074=>"101001011",
  61075=>"011111110",
  61076=>"010100011",
  61077=>"110000011",
  61078=>"010110010",
  61079=>"000111111",
  61080=>"101110101",
  61081=>"110111101",
  61082=>"010010100",
  61083=>"001001111",
  61084=>"011010001",
  61085=>"110101101",
  61086=>"011000000",
  61087=>"000110111",
  61088=>"110111100",
  61089=>"010010000",
  61090=>"111001100",
  61091=>"010101010",
  61092=>"100000010",
  61093=>"001101011",
  61094=>"001100101",
  61095=>"101000101",
  61096=>"100001010",
  61097=>"101001100",
  61098=>"010111111",
  61099=>"101001111",
  61100=>"100101000",
  61101=>"011000110",
  61102=>"011001001",
  61103=>"100111001",
  61104=>"010011100",
  61105=>"000011011",
  61106=>"100101010",
  61107=>"011110100",
  61108=>"101011001",
  61109=>"101101001",
  61110=>"101101001",
  61111=>"101000101",
  61112=>"100001111",
  61113=>"101110011",
  61114=>"100000001",
  61115=>"100111101",
  61116=>"000100110",
  61117=>"000001011",
  61118=>"100111100",
  61119=>"011111011",
  61120=>"110011001",
  61121=>"100101110",
  61122=>"000001101",
  61123=>"000000100",
  61124=>"000000101",
  61125=>"000101100",
  61126=>"100011111",
  61127=>"011011101",
  61128=>"000100000",
  61129=>"101111000",
  61130=>"101001110",
  61131=>"000000010",
  61132=>"101111111",
  61133=>"111101111",
  61134=>"000110111",
  61135=>"011101011",
  61136=>"100001100",
  61137=>"011000111",
  61138=>"011101011",
  61139=>"111010110",
  61140=>"111001111",
  61141=>"001000110",
  61142=>"000000000",
  61143=>"101011110",
  61144=>"000010101",
  61145=>"111100100",
  61146=>"101010101",
  61147=>"111101001",
  61148=>"101101101",
  61149=>"111000011",
  61150=>"010001000",
  61151=>"100001101",
  61152=>"011111101",
  61153=>"101101110",
  61154=>"110100010",
  61155=>"010100000",
  61156=>"110100101",
  61157=>"011111110",
  61158=>"111011110",
  61159=>"011011100",
  61160=>"110101001",
  61161=>"110110110",
  61162=>"110011100",
  61163=>"111111110",
  61164=>"000000101",
  61165=>"011111111",
  61166=>"111001010",
  61167=>"000001101",
  61168=>"111111010",
  61169=>"100000101",
  61170=>"111010110",
  61171=>"101000001",
  61172=>"110101111",
  61173=>"110101100",
  61174=>"000000111",
  61175=>"100110111",
  61176=>"111101010",
  61177=>"110111110",
  61178=>"000000011",
  61179=>"000001110",
  61180=>"000010101",
  61181=>"101110110",
  61182=>"100111011",
  61183=>"000010100",
  61184=>"001010101",
  61185=>"100000000",
  61186=>"101000111",
  61187=>"000110101",
  61188=>"000111010",
  61189=>"000010100",
  61190=>"101110101",
  61191=>"001100001",
  61192=>"110010010",
  61193=>"011101000",
  61194=>"101000000",
  61195=>"001100000",
  61196=>"110011100",
  61197=>"101011010",
  61198=>"000001100",
  61199=>"101100101",
  61200=>"000000100",
  61201=>"111001000",
  61202=>"000011111",
  61203=>"100110010",
  61204=>"111101101",
  61205=>"010111100",
  61206=>"011011001",
  61207=>"000010100",
  61208=>"010011001",
  61209=>"011001010",
  61210=>"001100010",
  61211=>"001001010",
  61212=>"000100111",
  61213=>"001001000",
  61214=>"110011010",
  61215=>"011011110",
  61216=>"001000011",
  61217=>"100111001",
  61218=>"000000110",
  61219=>"100101111",
  61220=>"101011111",
  61221=>"010101000",
  61222=>"001010111",
  61223=>"101101011",
  61224=>"100110010",
  61225=>"010101001",
  61226=>"100101011",
  61227=>"011111001",
  61228=>"010011101",
  61229=>"111111111",
  61230=>"000010111",
  61231=>"000010011",
  61232=>"010000001",
  61233=>"101000100",
  61234=>"011000001",
  61235=>"001011111",
  61236=>"000000000",
  61237=>"011101011",
  61238=>"010011001",
  61239=>"100110001",
  61240=>"101000001",
  61241=>"100110101",
  61242=>"001001001",
  61243=>"110000001",
  61244=>"100001110",
  61245=>"010111011",
  61246=>"000011000",
  61247=>"100110101",
  61248=>"100111001",
  61249=>"110110101",
  61250=>"001001011",
  61251=>"100100101",
  61252=>"101001011",
  61253=>"001000111",
  61254=>"100101111",
  61255=>"110110111",
  61256=>"000110111",
  61257=>"001101010",
  61258=>"101101110",
  61259=>"000000001",
  61260=>"110011011",
  61261=>"111000011",
  61262=>"111111000",
  61263=>"011011000",
  61264=>"000001100",
  61265=>"000001100",
  61266=>"001000101",
  61267=>"010110000",
  61268=>"101010000",
  61269=>"101011111",
  61270=>"000011011",
  61271=>"011010111",
  61272=>"010010111",
  61273=>"011111101",
  61274=>"100110101",
  61275=>"111011101",
  61276=>"011001111",
  61277=>"011010000",
  61278=>"010011101",
  61279=>"100110100",
  61280=>"010101000",
  61281=>"011001000",
  61282=>"111011111",
  61283=>"001010001",
  61284=>"010001011",
  61285=>"110001111",
  61286=>"100000011",
  61287=>"100110101",
  61288=>"000010000",
  61289=>"101111000",
  61290=>"010001011",
  61291=>"111011111",
  61292=>"110110110",
  61293=>"011100101",
  61294=>"111000110",
  61295=>"101001000",
  61296=>"111101111",
  61297=>"010001010",
  61298=>"010101010",
  61299=>"001100100",
  61300=>"010110001",
  61301=>"101110000",
  61302=>"011001111",
  61303=>"110011011",
  61304=>"011111001",
  61305=>"011011101",
  61306=>"110100100",
  61307=>"010010100",
  61308=>"111111000",
  61309=>"000010100",
  61310=>"101111110",
  61311=>"011000111",
  61312=>"001101111",
  61313=>"000010010",
  61314=>"101000101",
  61315=>"111100011",
  61316=>"010011101",
  61317=>"010011011",
  61318=>"111101111",
  61319=>"000010000",
  61320=>"011110001",
  61321=>"101111100",
  61322=>"010001110",
  61323=>"011010100",
  61324=>"111111111",
  61325=>"010100101",
  61326=>"101001110",
  61327=>"001100001",
  61328=>"000010000",
  61329=>"000100101",
  61330=>"000110110",
  61331=>"100001001",
  61332=>"111011011",
  61333=>"110001001",
  61334=>"011100010",
  61335=>"011100000",
  61336=>"110101101",
  61337=>"001011000",
  61338=>"000111110",
  61339=>"000010110",
  61340=>"101001011",
  61341=>"010101100",
  61342=>"110110010",
  61343=>"101111000",
  61344=>"101111101",
  61345=>"111011001",
  61346=>"001011100",
  61347=>"110111000",
  61348=>"010111100",
  61349=>"111110101",
  61350=>"010111000",
  61351=>"110010110",
  61352=>"011100000",
  61353=>"010100001",
  61354=>"000100000",
  61355=>"001011100",
  61356=>"000001101",
  61357=>"110100110",
  61358=>"101100111",
  61359=>"101000110",
  61360=>"001000011",
  61361=>"010111111",
  61362=>"100001000",
  61363=>"111000101",
  61364=>"000110011",
  61365=>"100101011",
  61366=>"110110110",
  61367=>"111010101",
  61368=>"111100110",
  61369=>"011000100",
  61370=>"101010100",
  61371=>"111110100",
  61372=>"110010001",
  61373=>"111000010",
  61374=>"111101100",
  61375=>"110011010",
  61376=>"011010010",
  61377=>"011000001",
  61378=>"111111111",
  61379=>"001111010",
  61380=>"010110101",
  61381=>"111001100",
  61382=>"010001100",
  61383=>"110101011",
  61384=>"011010001",
  61385=>"011001001",
  61386=>"100011010",
  61387=>"011100110",
  61388=>"000001101",
  61389=>"000010101",
  61390=>"100100101",
  61391=>"001101110",
  61392=>"100101110",
  61393=>"100101101",
  61394=>"010000111",
  61395=>"110001011",
  61396=>"100000100",
  61397=>"111111111",
  61398=>"110001010",
  61399=>"101010100",
  61400=>"111000100",
  61401=>"011100011",
  61402=>"111001111",
  61403=>"011101110",
  61404=>"000011110",
  61405=>"011010110",
  61406=>"111110111",
  61407=>"000001001",
  61408=>"010010111",
  61409=>"011100110",
  61410=>"101110100",
  61411=>"101110000",
  61412=>"000101010",
  61413=>"111100111",
  61414=>"111110100",
  61415=>"111111011",
  61416=>"111000000",
  61417=>"011000011",
  61418=>"000101000",
  61419=>"100100011",
  61420=>"011100001",
  61421=>"000000101",
  61422=>"100101010",
  61423=>"001111010",
  61424=>"101010111",
  61425=>"101011110",
  61426=>"110110110",
  61427=>"110110011",
  61428=>"111001101",
  61429=>"100110101",
  61430=>"001011010",
  61431=>"110111111",
  61432=>"100010111",
  61433=>"100100010",
  61434=>"001111100",
  61435=>"001111100",
  61436=>"111000111",
  61437=>"010000000",
  61438=>"110001111",
  61439=>"011110101",
  61440=>"101001110",
  61441=>"000000100",
  61442=>"110000011",
  61443=>"111001010",
  61444=>"100100010",
  61445=>"110010110",
  61446=>"010011010",
  61447=>"110000010",
  61448=>"011001010",
  61449=>"100110011",
  61450=>"110010000",
  61451=>"001000111",
  61452=>"100110101",
  61453=>"101101010",
  61454=>"000001000",
  61455=>"001010010",
  61456=>"101100011",
  61457=>"000110001",
  61458=>"101011010",
  61459=>"011010101",
  61460=>"011101110",
  61461=>"010110101",
  61462=>"000110100",
  61463=>"101000111",
  61464=>"010100110",
  61465=>"001111000",
  61466=>"111111111",
  61467=>"010100010",
  61468=>"000100000",
  61469=>"110000101",
  61470=>"011010111",
  61471=>"010011110",
  61472=>"010010101",
  61473=>"110000110",
  61474=>"011111001",
  61475=>"100000101",
  61476=>"001111000",
  61477=>"100001001",
  61478=>"101000100",
  61479=>"101100111",
  61480=>"001101000",
  61481=>"100100100",
  61482=>"011111101",
  61483=>"011000100",
  61484=>"110101001",
  61485=>"000100001",
  61486=>"010010110",
  61487=>"111001101",
  61488=>"011001011",
  61489=>"000010011",
  61490=>"010110011",
  61491=>"111111111",
  61492=>"010000100",
  61493=>"000101000",
  61494=>"110011010",
  61495=>"000010010",
  61496=>"011110111",
  61497=>"100111000",
  61498=>"100001010",
  61499=>"101101011",
  61500=>"000011010",
  61501=>"001101001",
  61502=>"110000100",
  61503=>"100010100",
  61504=>"010110000",
  61505=>"000000011",
  61506=>"100011001",
  61507=>"001000001",
  61508=>"110101110",
  61509=>"000011001",
  61510=>"011111100",
  61511=>"111101000",
  61512=>"011111101",
  61513=>"110011100",
  61514=>"101010111",
  61515=>"001000000",
  61516=>"010011010",
  61517=>"111101001",
  61518=>"011111000",
  61519=>"000100000",
  61520=>"010110101",
  61521=>"000000010",
  61522=>"010001110",
  61523=>"111011000",
  61524=>"010000100",
  61525=>"100001010",
  61526=>"001101101",
  61527=>"001001101",
  61528=>"110011011",
  61529=>"001010101",
  61530=>"111000010",
  61531=>"110111010",
  61532=>"101000001",
  61533=>"100010100",
  61534=>"001001110",
  61535=>"010100101",
  61536=>"100100110",
  61537=>"110111101",
  61538=>"010100111",
  61539=>"000101011",
  61540=>"011000100",
  61541=>"010000110",
  61542=>"110101110",
  61543=>"111011101",
  61544=>"000010111",
  61545=>"000010110",
  61546=>"010010011",
  61547=>"110101010",
  61548=>"010110000",
  61549=>"111010001",
  61550=>"001001011",
  61551=>"001000000",
  61552=>"010100010",
  61553=>"010001111",
  61554=>"001101110",
  61555=>"101011110",
  61556=>"111011010",
  61557=>"011001110",
  61558=>"101010000",
  61559=>"011011011",
  61560=>"001000000",
  61561=>"100000010",
  61562=>"100100011",
  61563=>"110101000",
  61564=>"010101110",
  61565=>"011001011",
  61566=>"000010101",
  61567=>"010001100",
  61568=>"010010000",
  61569=>"010000100",
  61570=>"010100001",
  61571=>"101011001",
  61572=>"111010010",
  61573=>"111111111",
  61574=>"011111101",
  61575=>"110001001",
  61576=>"110010011",
  61577=>"100100000",
  61578=>"000110100",
  61579=>"111001110",
  61580=>"111010111",
  61581=>"010010110",
  61582=>"100001000",
  61583=>"100011001",
  61584=>"000100011",
  61585=>"011110110",
  61586=>"101011011",
  61587=>"001100101",
  61588=>"001110100",
  61589=>"100100100",
  61590=>"010110100",
  61591=>"001010110",
  61592=>"000111110",
  61593=>"101110110",
  61594=>"111111011",
  61595=>"011101011",
  61596=>"000001100",
  61597=>"001100100",
  61598=>"111101111",
  61599=>"110011101",
  61600=>"010100010",
  61601=>"101100111",
  61602=>"000101111",
  61603=>"111111100",
  61604=>"110110111",
  61605=>"100011111",
  61606=>"101010001",
  61607=>"100011011",
  61608=>"101100001",
  61609=>"110101011",
  61610=>"110010010",
  61611=>"001011110",
  61612=>"111110111",
  61613=>"101111111",
  61614=>"000011110",
  61615=>"101111010",
  61616=>"001001110",
  61617=>"000111011",
  61618=>"101111001",
  61619=>"100001101",
  61620=>"101010111",
  61621=>"100111001",
  61622=>"000011100",
  61623=>"001010000",
  61624=>"011010011",
  61625=>"000110010",
  61626=>"001000110",
  61627=>"010010000",
  61628=>"010110011",
  61629=>"110011100",
  61630=>"011110110",
  61631=>"101100101",
  61632=>"111101000",
  61633=>"110100111",
  61634=>"011000000",
  61635=>"011011110",
  61636=>"010000101",
  61637=>"100101111",
  61638=>"101001110",
  61639=>"111111000",
  61640=>"100001011",
  61641=>"010101110",
  61642=>"001100110",
  61643=>"011001001",
  61644=>"111101000",
  61645=>"111100110",
  61646=>"000001000",
  61647=>"110110110",
  61648=>"110100000",
  61649=>"101000011",
  61650=>"011011010",
  61651=>"011100111",
  61652=>"110000111",
  61653=>"010110100",
  61654=>"100011000",
  61655=>"000001000",
  61656=>"001101001",
  61657=>"101110010",
  61658=>"010001000",
  61659=>"010000111",
  61660=>"100010011",
  61661=>"011111000",
  61662=>"000000010",
  61663=>"110000010",
  61664=>"101101100",
  61665=>"000011111",
  61666=>"010010111",
  61667=>"010001010",
  61668=>"100001100",
  61669=>"101001110",
  61670=>"100001001",
  61671=>"011001111",
  61672=>"000101001",
  61673=>"110011011",
  61674=>"101100011",
  61675=>"001010000",
  61676=>"000100000",
  61677=>"111001000",
  61678=>"101110011",
  61679=>"001001001",
  61680=>"101100001",
  61681=>"010011000",
  61682=>"001111000",
  61683=>"010000010",
  61684=>"101001000",
  61685=>"000011001",
  61686=>"011010010",
  61687=>"100000111",
  61688=>"100101111",
  61689=>"101101001",
  61690=>"010101110",
  61691=>"001000011",
  61692=>"000100001",
  61693=>"010101010",
  61694=>"001010010",
  61695=>"000111100",
  61696=>"011100010",
  61697=>"010001001",
  61698=>"101010111",
  61699=>"001101011",
  61700=>"100000011",
  61701=>"111110100",
  61702=>"001111101",
  61703=>"111001100",
  61704=>"000100100",
  61705=>"000111011",
  61706=>"001000100",
  61707=>"101100101",
  61708=>"000111000",
  61709=>"000111111",
  61710=>"111010111",
  61711=>"001000001",
  61712=>"101000001",
  61713=>"011110111",
  61714=>"000110101",
  61715=>"111110111",
  61716=>"000001110",
  61717=>"100111111",
  61718=>"001000011",
  61719=>"001000101",
  61720=>"101101111",
  61721=>"110011000",
  61722=>"000011011",
  61723=>"000110011",
  61724=>"010100000",
  61725=>"110110101",
  61726=>"001010010",
  61727=>"011100000",
  61728=>"000010000",
  61729=>"100111010",
  61730=>"110101000",
  61731=>"100011100",
  61732=>"011001110",
  61733=>"001110101",
  61734=>"111110111",
  61735=>"111101101",
  61736=>"011010101",
  61737=>"000010110",
  61738=>"111101101",
  61739=>"011011001",
  61740=>"000110010",
  61741=>"101100000",
  61742=>"000100110",
  61743=>"010010011",
  61744=>"010101000",
  61745=>"111011110",
  61746=>"111001000",
  61747=>"110001101",
  61748=>"111000111",
  61749=>"000101100",
  61750=>"011100111",
  61751=>"111000101",
  61752=>"000111001",
  61753=>"010001111",
  61754=>"000110110",
  61755=>"111100100",
  61756=>"100000110",
  61757=>"111110001",
  61758=>"011111110",
  61759=>"110100001",
  61760=>"101110101",
  61761=>"000000110",
  61762=>"101100110",
  61763=>"001011110",
  61764=>"101111011",
  61765=>"010101000",
  61766=>"100110011",
  61767=>"011110001",
  61768=>"010101000",
  61769=>"000010010",
  61770=>"101011010",
  61771=>"001100011",
  61772=>"101010100",
  61773=>"000111000",
  61774=>"111011011",
  61775=>"111110101",
  61776=>"111010100",
  61777=>"011010110",
  61778=>"110101101",
  61779=>"101101111",
  61780=>"101001100",
  61781=>"000000011",
  61782=>"001000011",
  61783=>"100001001",
  61784=>"010000101",
  61785=>"110000000",
  61786=>"000101011",
  61787=>"100000110",
  61788=>"001100111",
  61789=>"110010001",
  61790=>"001001000",
  61791=>"011100010",
  61792=>"111110111",
  61793=>"000101111",
  61794=>"110000000",
  61795=>"010101000",
  61796=>"011010000",
  61797=>"101101010",
  61798=>"000100101",
  61799=>"111101110",
  61800=>"111011110",
  61801=>"010100001",
  61802=>"011000100",
  61803=>"001001011",
  61804=>"110000011",
  61805=>"011101100",
  61806=>"101001010",
  61807=>"101101101",
  61808=>"101111011",
  61809=>"101101000",
  61810=>"100110000",
  61811=>"011110101",
  61812=>"101011011",
  61813=>"111010011",
  61814=>"100100101",
  61815=>"111110010",
  61816=>"001111100",
  61817=>"100110111",
  61818=>"100111111",
  61819=>"010010010",
  61820=>"110001000",
  61821=>"100001010",
  61822=>"010111011",
  61823=>"101000101",
  61824=>"011110100",
  61825=>"010101110",
  61826=>"100111001",
  61827=>"011111101",
  61828=>"101011011",
  61829=>"000001101",
  61830=>"001110110",
  61831=>"111000111",
  61832=>"111010100",
  61833=>"111100011",
  61834=>"100010101",
  61835=>"000111011",
  61836=>"011111101",
  61837=>"111010110",
  61838=>"110110111",
  61839=>"011101101",
  61840=>"111101010",
  61841=>"000001111",
  61842=>"101110011",
  61843=>"011101011",
  61844=>"100011001",
  61845=>"010011100",
  61846=>"010111111",
  61847=>"011010001",
  61848=>"010110001",
  61849=>"010010010",
  61850=>"111011110",
  61851=>"100101001",
  61852=>"011010100",
  61853=>"101100001",
  61854=>"100100001",
  61855=>"000100111",
  61856=>"000100011",
  61857=>"100010111",
  61858=>"011001000",
  61859=>"010000100",
  61860=>"000100100",
  61861=>"010000000",
  61862=>"011010100",
  61863=>"111010100",
  61864=>"100101011",
  61865=>"001100010",
  61866=>"100001000",
  61867=>"011101010",
  61868=>"101101110",
  61869=>"101100110",
  61870=>"000001110",
  61871=>"101101111",
  61872=>"101100010",
  61873=>"111101000",
  61874=>"100101011",
  61875=>"100111111",
  61876=>"101110111",
  61877=>"000100100",
  61878=>"000101101",
  61879=>"100010110",
  61880=>"001110000",
  61881=>"000110100",
  61882=>"001010011",
  61883=>"111000110",
  61884=>"001001101",
  61885=>"101011011",
  61886=>"000010110",
  61887=>"010010101",
  61888=>"110010101",
  61889=>"101011110",
  61890=>"010011101",
  61891=>"011101001",
  61892=>"001110011",
  61893=>"010100111",
  61894=>"111011111",
  61895=>"110000000",
  61896=>"001111000",
  61897=>"000011101",
  61898=>"011000111",
  61899=>"011010011",
  61900=>"110100101",
  61901=>"100010100",
  61902=>"011100001",
  61903=>"101000011",
  61904=>"111110110",
  61905=>"110000100",
  61906=>"011000110",
  61907=>"000110101",
  61908=>"101010011",
  61909=>"111001000",
  61910=>"001101111",
  61911=>"010110011",
  61912=>"101100001",
  61913=>"011011101",
  61914=>"111111100",
  61915=>"011101101",
  61916=>"010011001",
  61917=>"010010011",
  61918=>"110110011",
  61919=>"001000000",
  61920=>"000100000",
  61921=>"001010010",
  61922=>"001110111",
  61923=>"110011010",
  61924=>"001010010",
  61925=>"101111000",
  61926=>"011110010",
  61927=>"100001010",
  61928=>"110100011",
  61929=>"001001111",
  61930=>"000101100",
  61931=>"011101100",
  61932=>"110110111",
  61933=>"011001111",
  61934=>"011100101",
  61935=>"001000110",
  61936=>"100001110",
  61937=>"111001110",
  61938=>"000000010",
  61939=>"001100110",
  61940=>"100101100",
  61941=>"001101001",
  61942=>"110101111",
  61943=>"111100100",
  61944=>"110110101",
  61945=>"110101011",
  61946=>"110111001",
  61947=>"000111111",
  61948=>"001110010",
  61949=>"100010110",
  61950=>"010001011",
  61951=>"000111101",
  61952=>"100000000",
  61953=>"111101111",
  61954=>"110011011",
  61955=>"100011100",
  61956=>"011101010",
  61957=>"011100000",
  61958=>"011010110",
  61959=>"010111101",
  61960=>"001110011",
  61961=>"011100110",
  61962=>"101001000",
  61963=>"010000111",
  61964=>"000111001",
  61965=>"100100101",
  61966=>"010110000",
  61967=>"111011110",
  61968=>"011011010",
  61969=>"110000111",
  61970=>"100001111",
  61971=>"100100110",
  61972=>"010001111",
  61973=>"101100101",
  61974=>"101110111",
  61975=>"000010001",
  61976=>"000000110",
  61977=>"011010100",
  61978=>"101001000",
  61979=>"111011110",
  61980=>"011101100",
  61981=>"011011100",
  61982=>"110100010",
  61983=>"000111010",
  61984=>"010111011",
  61985=>"010010101",
  61986=>"000001011",
  61987=>"000001010",
  61988=>"000111010",
  61989=>"111010011",
  61990=>"000110011",
  61991=>"001101101",
  61992=>"110101101",
  61993=>"110111110",
  61994=>"110000111",
  61995=>"100111010",
  61996=>"000101111",
  61997=>"100100100",
  61998=>"001010000",
  61999=>"011010101",
  62000=>"000011110",
  62001=>"111011011",
  62002=>"100100111",
  62003=>"001100011",
  62004=>"010011101",
  62005=>"010101000",
  62006=>"010011110",
  62007=>"010100000",
  62008=>"000100000",
  62009=>"101010110",
  62010=>"111010111",
  62011=>"100010000",
  62012=>"000101011",
  62013=>"000010000",
  62014=>"110011010",
  62015=>"001110101",
  62016=>"100010101",
  62017=>"000111011",
  62018=>"101000101",
  62019=>"101010000",
  62020=>"010001001",
  62021=>"001001110",
  62022=>"100000000",
  62023=>"110000101",
  62024=>"011001100",
  62025=>"010111001",
  62026=>"110011010",
  62027=>"110000100",
  62028=>"101110100",
  62029=>"011010010",
  62030=>"011000111",
  62031=>"001000101",
  62032=>"010110011",
  62033=>"101000010",
  62034=>"001100110",
  62035=>"110000110",
  62036=>"100000001",
  62037=>"000101101",
  62038=>"001100000",
  62039=>"000100110",
  62040=>"000110011",
  62041=>"110110011",
  62042=>"110001001",
  62043=>"101100011",
  62044=>"111110100",
  62045=>"101001010",
  62046=>"110100001",
  62047=>"011011000",
  62048=>"010011100",
  62049=>"101101011",
  62050=>"100010111",
  62051=>"011011101",
  62052=>"101110100",
  62053=>"010011100",
  62054=>"111101111",
  62055=>"111111101",
  62056=>"100010111",
  62057=>"001011001",
  62058=>"001110111",
  62059=>"110000011",
  62060=>"100110110",
  62061=>"001001100",
  62062=>"000110001",
  62063=>"011101000",
  62064=>"001100001",
  62065=>"001001101",
  62066=>"011001100",
  62067=>"000011000",
  62068=>"011111111",
  62069=>"110011011",
  62070=>"011010101",
  62071=>"001011110",
  62072=>"101001011",
  62073=>"000110111",
  62074=>"110011000",
  62075=>"101100110",
  62076=>"010101010",
  62077=>"000001101",
  62078=>"001100010",
  62079=>"111011011",
  62080=>"001010000",
  62081=>"001101110",
  62082=>"011001001",
  62083=>"100101001",
  62084=>"011110110",
  62085=>"111111100",
  62086=>"000100000",
  62087=>"100010001",
  62088=>"000100101",
  62089=>"000000001",
  62090=>"001100110",
  62091=>"011101010",
  62092=>"110100101",
  62093=>"010000111",
  62094=>"010111010",
  62095=>"010111100",
  62096=>"101000010",
  62097=>"111010111",
  62098=>"010000111",
  62099=>"000011100",
  62100=>"100001101",
  62101=>"110110010",
  62102=>"001011101",
  62103=>"000010100",
  62104=>"110110100",
  62105=>"001011000",
  62106=>"001001011",
  62107=>"001000110",
  62108=>"110010100",
  62109=>"110010101",
  62110=>"000101111",
  62111=>"101100000",
  62112=>"000010111",
  62113=>"001010111",
  62114=>"010011110",
  62115=>"101101010",
  62116=>"010000001",
  62117=>"000010111",
  62118=>"101101000",
  62119=>"000101111",
  62120=>"111100001",
  62121=>"010001101",
  62122=>"001111100",
  62123=>"100101011",
  62124=>"100101010",
  62125=>"100000111",
  62126=>"110010101",
  62127=>"010011011",
  62128=>"000001000",
  62129=>"001011000",
  62130=>"011101010",
  62131=>"110001111",
  62132=>"111101101",
  62133=>"011111101",
  62134=>"111100111",
  62135=>"100000010",
  62136=>"100010010",
  62137=>"101110011",
  62138=>"000101110",
  62139=>"010000110",
  62140=>"111000000",
  62141=>"100011000",
  62142=>"000100011",
  62143=>"000001000",
  62144=>"110110011",
  62145=>"010000101",
  62146=>"000111011",
  62147=>"101001100",
  62148=>"011011000",
  62149=>"101000000",
  62150=>"101000000",
  62151=>"000000000",
  62152=>"010000001",
  62153=>"011000010",
  62154=>"011111000",
  62155=>"000010000",
  62156=>"100000010",
  62157=>"011011011",
  62158=>"100111000",
  62159=>"010101011",
  62160=>"010010000",
  62161=>"000000010",
  62162=>"000001111",
  62163=>"010100010",
  62164=>"000011110",
  62165=>"001000110",
  62166=>"000000100",
  62167=>"100010110",
  62168=>"100101111",
  62169=>"000010010",
  62170=>"111111110",
  62171=>"011001010",
  62172=>"000101100",
  62173=>"100010000",
  62174=>"010100010",
  62175=>"100001010",
  62176=>"100001001",
  62177=>"001010100",
  62178=>"111011010",
  62179=>"010001111",
  62180=>"001011010",
  62181=>"111100101",
  62182=>"100110101",
  62183=>"010101100",
  62184=>"000011111",
  62185=>"010001101",
  62186=>"111001000",
  62187=>"110001000",
  62188=>"000100011",
  62189=>"101111110",
  62190=>"000000101",
  62191=>"010111110",
  62192=>"011011001",
  62193=>"110011111",
  62194=>"110111011",
  62195=>"110110011",
  62196=>"010111010",
  62197=>"100101101",
  62198=>"100011111",
  62199=>"011001000",
  62200=>"000011110",
  62201=>"100010100",
  62202=>"111101111",
  62203=>"100000110",
  62204=>"111111101",
  62205=>"011010101",
  62206=>"000001000",
  62207=>"100111001",
  62208=>"101001010",
  62209=>"101011110",
  62210=>"111100011",
  62211=>"100010001",
  62212=>"000001001",
  62213=>"000001100",
  62214=>"010101011",
  62215=>"101100000",
  62216=>"101101101",
  62217=>"100000100",
  62218=>"010101100",
  62219=>"100000101",
  62220=>"101010100",
  62221=>"111001110",
  62222=>"000000000",
  62223=>"100110100",
  62224=>"100100101",
  62225=>"101101110",
  62226=>"010001110",
  62227=>"101011111",
  62228=>"110000000",
  62229=>"001001110",
  62230=>"000100000",
  62231=>"010000010",
  62232=>"001100111",
  62233=>"001110110",
  62234=>"000101100",
  62235=>"010000000",
  62236=>"000111101",
  62237=>"100100011",
  62238=>"010101110",
  62239=>"110000001",
  62240=>"010101101",
  62241=>"011101110",
  62242=>"110100011",
  62243=>"101100110",
  62244=>"111011111",
  62245=>"000101000",
  62246=>"000101011",
  62247=>"011101101",
  62248=>"000111010",
  62249=>"111100001",
  62250=>"011001111",
  62251=>"110001110",
  62252=>"101110110",
  62253=>"101010010",
  62254=>"110100110",
  62255=>"100110110",
  62256=>"101100110",
  62257=>"101011110",
  62258=>"100010010",
  62259=>"001010010",
  62260=>"100110100",
  62261=>"111010010",
  62262=>"111001010",
  62263=>"000110100",
  62264=>"110001100",
  62265=>"100100001",
  62266=>"000100100",
  62267=>"111010010",
  62268=>"001101001",
  62269=>"000011000",
  62270=>"100100001",
  62271=>"111010100",
  62272=>"000011000",
  62273=>"100110011",
  62274=>"010001110",
  62275=>"101010111",
  62276=>"010110110",
  62277=>"001111010",
  62278=>"111110011",
  62279=>"000011000",
  62280=>"101010001",
  62281=>"100000011",
  62282=>"001011110",
  62283=>"101011010",
  62284=>"010111001",
  62285=>"001101000",
  62286=>"000100000",
  62287=>"010110110",
  62288=>"110101000",
  62289=>"101111011",
  62290=>"100001000",
  62291=>"011111011",
  62292=>"111000100",
  62293=>"100100101",
  62294=>"001101101",
  62295=>"000000011",
  62296=>"001100110",
  62297=>"001010000",
  62298=>"100111110",
  62299=>"001111111",
  62300=>"111011111",
  62301=>"111010011",
  62302=>"001011101",
  62303=>"010010110",
  62304=>"100000000",
  62305=>"011110011",
  62306=>"110110001",
  62307=>"110100010",
  62308=>"111101100",
  62309=>"110100000",
  62310=>"000111010",
  62311=>"010100101",
  62312=>"011000100",
  62313=>"110110011",
  62314=>"101000101",
  62315=>"000111010",
  62316=>"000001000",
  62317=>"001001110",
  62318=>"111010000",
  62319=>"010111100",
  62320=>"111000010",
  62321=>"100010000",
  62322=>"010100010",
  62323=>"111001110",
  62324=>"010000111",
  62325=>"101100100",
  62326=>"100001100",
  62327=>"101101010",
  62328=>"010000101",
  62329=>"111111010",
  62330=>"100011100",
  62331=>"110110001",
  62332=>"000001100",
  62333=>"100110000",
  62334=>"111001000",
  62335=>"110111111",
  62336=>"110000100",
  62337=>"000001010",
  62338=>"111000101",
  62339=>"001010100",
  62340=>"110110101",
  62341=>"110011110",
  62342=>"100100110",
  62343=>"000010001",
  62344=>"100111000",
  62345=>"010011111",
  62346=>"000111010",
  62347=>"001001001",
  62348=>"001100100",
  62349=>"110001110",
  62350=>"010101001",
  62351=>"010111110",
  62352=>"010100010",
  62353=>"110000010",
  62354=>"000000000",
  62355=>"011000001",
  62356=>"000110100",
  62357=>"111101100",
  62358=>"010010010",
  62359=>"000011101",
  62360=>"001100101",
  62361=>"101111000",
  62362=>"000111010",
  62363=>"100001001",
  62364=>"111000000",
  62365=>"110001101",
  62366=>"101100000",
  62367=>"110000101",
  62368=>"011000011",
  62369=>"011100000",
  62370=>"011010110",
  62371=>"111010011",
  62372=>"100100000",
  62373=>"101111101",
  62374=>"111110010",
  62375=>"100010111",
  62376=>"101010111",
  62377=>"111001101",
  62378=>"000010010",
  62379=>"101101100",
  62380=>"111001010",
  62381=>"010101110",
  62382=>"111111001",
  62383=>"100010001",
  62384=>"111101011",
  62385=>"110110001",
  62386=>"100100010",
  62387=>"010110010",
  62388=>"111001000",
  62389=>"010011100",
  62390=>"011011110",
  62391=>"000111100",
  62392=>"010100010",
  62393=>"101100111",
  62394=>"101011000",
  62395=>"011001111",
  62396=>"010010111",
  62397=>"000100000",
  62398=>"011110011",
  62399=>"110010101",
  62400=>"010110010",
  62401=>"100101110",
  62402=>"001111100",
  62403=>"010010110",
  62404=>"101010001",
  62405=>"000100100",
  62406=>"010000100",
  62407=>"111111110",
  62408=>"001110001",
  62409=>"101011001",
  62410=>"110110111",
  62411=>"101010011",
  62412=>"011010010",
  62413=>"110101000",
  62414=>"000001000",
  62415=>"001011110",
  62416=>"111111110",
  62417=>"110001001",
  62418=>"110010111",
  62419=>"111100000",
  62420=>"011110010",
  62421=>"100111100",
  62422=>"010100001",
  62423=>"101011010",
  62424=>"111000110",
  62425=>"000100000",
  62426=>"111010010",
  62427=>"111100100",
  62428=>"110011010",
  62429=>"010101000",
  62430=>"000001100",
  62431=>"001010110",
  62432=>"101100111",
  62433=>"111110011",
  62434=>"111011001",
  62435=>"111111111",
  62436=>"001101001",
  62437=>"100000110",
  62438=>"110010101",
  62439=>"111010000",
  62440=>"101011101",
  62441=>"000010101",
  62442=>"110000000",
  62443=>"100000111",
  62444=>"000100010",
  62445=>"000110001",
  62446=>"111000000",
  62447=>"011110111",
  62448=>"000010100",
  62449=>"110111010",
  62450=>"001100110",
  62451=>"101101011",
  62452=>"001100010",
  62453=>"100110001",
  62454=>"101010101",
  62455=>"001000000",
  62456=>"100010010",
  62457=>"001001101",
  62458=>"100111011",
  62459=>"011111111",
  62460=>"010001101",
  62461=>"110010001",
  62462=>"111010000",
  62463=>"101100000",
  62464=>"000000000",
  62465=>"001000000",
  62466=>"111111001",
  62467=>"000101001",
  62468=>"011000000",
  62469=>"001100111",
  62470=>"000011010",
  62471=>"000010100",
  62472=>"011110000",
  62473=>"100101110",
  62474=>"011000100",
  62475=>"001000110",
  62476=>"100111100",
  62477=>"011101011",
  62478=>"101101010",
  62479=>"101000111",
  62480=>"010000010",
  62481=>"101010011",
  62482=>"100111100",
  62483=>"010111101",
  62484=>"100001100",
  62485=>"010100100",
  62486=>"000100101",
  62487=>"110011100",
  62488=>"011110001",
  62489=>"001111110",
  62490=>"100110000",
  62491=>"000000001",
  62492=>"000111101",
  62493=>"010111111",
  62494=>"010010001",
  62495=>"000011110",
  62496=>"000010110",
  62497=>"111110110",
  62498=>"101010101",
  62499=>"110000110",
  62500=>"110100000",
  62501=>"110101110",
  62502=>"100100011",
  62503=>"101011010",
  62504=>"110001001",
  62505=>"110001000",
  62506=>"001011101",
  62507=>"000101100",
  62508=>"110000011",
  62509=>"001111111",
  62510=>"111101100",
  62511=>"100011111",
  62512=>"100110011",
  62513=>"011110100",
  62514=>"101101001",
  62515=>"011111100",
  62516=>"011100100",
  62517=>"111001001",
  62518=>"000110001",
  62519=>"110011110",
  62520=>"000001010",
  62521=>"101100011",
  62522=>"011011001",
  62523=>"001000110",
  62524=>"000110111",
  62525=>"000000100",
  62526=>"110010111",
  62527=>"000101001",
  62528=>"001011011",
  62529=>"110101000",
  62530=>"000001110",
  62531=>"010000100",
  62532=>"010011010",
  62533=>"111011001",
  62534=>"111111010",
  62535=>"101000000",
  62536=>"001000100",
  62537=>"010010011",
  62538=>"010110011",
  62539=>"000101110",
  62540=>"011101110",
  62541=>"001000011",
  62542=>"111101101",
  62543=>"111010100",
  62544=>"001011010",
  62545=>"110101110",
  62546=>"011011110",
  62547=>"111111101",
  62548=>"100011000",
  62549=>"010000001",
  62550=>"011110011",
  62551=>"101000001",
  62552=>"001101111",
  62553=>"111100000",
  62554=>"101010110",
  62555=>"100101010",
  62556=>"000100001",
  62557=>"100100110",
  62558=>"110110100",
  62559=>"010101010",
  62560=>"100000001",
  62561=>"100100101",
  62562=>"110010000",
  62563=>"110000010",
  62564=>"011000101",
  62565=>"001001000",
  62566=>"111010111",
  62567=>"000110000",
  62568=>"011011010",
  62569=>"101100111",
  62570=>"000101010",
  62571=>"100110110",
  62572=>"010000101",
  62573=>"010111011",
  62574=>"101011111",
  62575=>"100001010",
  62576=>"111011110",
  62577=>"000000000",
  62578=>"000010111",
  62579=>"101011100",
  62580=>"010001010",
  62581=>"011110100",
  62582=>"100100000",
  62583=>"010010100",
  62584=>"101111010",
  62585=>"011111000",
  62586=>"100110110",
  62587=>"110100101",
  62588=>"000010110",
  62589=>"111101010",
  62590=>"100111110",
  62591=>"011011101",
  62592=>"111110000",
  62593=>"011110100",
  62594=>"111000100",
  62595=>"100100101",
  62596=>"011001011",
  62597=>"011001000",
  62598=>"101110100",
  62599=>"000000110",
  62600=>"110111010",
  62601=>"001010111",
  62602=>"100001110",
  62603=>"010000100",
  62604=>"110010111",
  62605=>"010111010",
  62606=>"010011110",
  62607=>"010011010",
  62608=>"011010010",
  62609=>"110001001",
  62610=>"110101100",
  62611=>"000101110",
  62612=>"010000110",
  62613=>"010010110",
  62614=>"101011010",
  62615=>"000101110",
  62616=>"100101011",
  62617=>"110001100",
  62618=>"110010000",
  62619=>"100010011",
  62620=>"101110110",
  62621=>"011101100",
  62622=>"010100110",
  62623=>"000100000",
  62624=>"000111101",
  62625=>"000111101",
  62626=>"111001010",
  62627=>"000111100",
  62628=>"101110101",
  62629=>"010011100",
  62630=>"001110001",
  62631=>"100010001",
  62632=>"000000010",
  62633=>"000010010",
  62634=>"011111101",
  62635=>"001001010",
  62636=>"011010010",
  62637=>"110010111",
  62638=>"101010000",
  62639=>"001110000",
  62640=>"111011111",
  62641=>"111111111",
  62642=>"000110110",
  62643=>"010010000",
  62644=>"100011000",
  62645=>"110110101",
  62646=>"101101000",
  62647=>"000001001",
  62648=>"011100100",
  62649=>"000101111",
  62650=>"100000111",
  62651=>"011010011",
  62652=>"101110011",
  62653=>"000100100",
  62654=>"110101111",
  62655=>"000101110",
  62656=>"001100001",
  62657=>"100111110",
  62658=>"111000010",
  62659=>"010011000",
  62660=>"011100111",
  62661=>"100111101",
  62662=>"001010010",
  62663=>"001100011",
  62664=>"111000010",
  62665=>"110101001",
  62666=>"101100011",
  62667=>"000101101",
  62668=>"001010000",
  62669=>"110001110",
  62670=>"110001101",
  62671=>"001000010",
  62672=>"100100010",
  62673=>"001001110",
  62674=>"100000010",
  62675=>"001010111",
  62676=>"111100101",
  62677=>"100110000",
  62678=>"001101111",
  62679=>"100111010",
  62680=>"001000111",
  62681=>"000010000",
  62682=>"000000101",
  62683=>"111100000",
  62684=>"010000001",
  62685=>"100001010",
  62686=>"000001101",
  62687=>"000000010",
  62688=>"100110001",
  62689=>"101010010",
  62690=>"111111100",
  62691=>"100111001",
  62692=>"111011110",
  62693=>"010011001",
  62694=>"000110000",
  62695=>"110100001",
  62696=>"010110111",
  62697=>"111011101",
  62698=>"000001111",
  62699=>"110001100",
  62700=>"100111101",
  62701=>"110001101",
  62702=>"110010100",
  62703=>"100001010",
  62704=>"000010000",
  62705=>"111101010",
  62706=>"111011011",
  62707=>"100001011",
  62708=>"101011110",
  62709=>"110101100",
  62710=>"110100001",
  62711=>"110110110",
  62712=>"010101100",
  62713=>"110011100",
  62714=>"101100010",
  62715=>"110001000",
  62716=>"000010001",
  62717=>"010000110",
  62718=>"100100010",
  62719=>"101001100",
  62720=>"011110011",
  62721=>"001011010",
  62722=>"110010110",
  62723=>"001100001",
  62724=>"100110010",
  62725=>"111101011",
  62726=>"010011011",
  62727=>"000101011",
  62728=>"011000001",
  62729=>"111010000",
  62730=>"111110011",
  62731=>"010010110",
  62732=>"011010111",
  62733=>"101100110",
  62734=>"001110010",
  62735=>"001010010",
  62736=>"011010010",
  62737=>"000100001",
  62738=>"100001010",
  62739=>"000001011",
  62740=>"001010111",
  62741=>"100110001",
  62742=>"100110001",
  62743=>"000011001",
  62744=>"000010110",
  62745=>"111001001",
  62746=>"011110011",
  62747=>"101111000",
  62748=>"011110011",
  62749=>"010110111",
  62750=>"011010100",
  62751=>"000100110",
  62752=>"000111000",
  62753=>"011001000",
  62754=>"001010011",
  62755=>"001110111",
  62756=>"111001011",
  62757=>"110100110",
  62758=>"111110100",
  62759=>"001010001",
  62760=>"100110110",
  62761=>"110000111",
  62762=>"001011111",
  62763=>"011101111",
  62764=>"011011100",
  62765=>"111111011",
  62766=>"010000011",
  62767=>"111110001",
  62768=>"000010000",
  62769=>"010101110",
  62770=>"010011001",
  62771=>"000110000",
  62772=>"101100111",
  62773=>"110010111",
  62774=>"111110110",
  62775=>"110000101",
  62776=>"001000100",
  62777=>"101000010",
  62778=>"110111110",
  62779=>"001111000",
  62780=>"110011101",
  62781=>"111100101",
  62782=>"111111110",
  62783=>"011010110",
  62784=>"111010111",
  62785=>"001101011",
  62786=>"010110100",
  62787=>"001010001",
  62788=>"110110111",
  62789=>"000001001",
  62790=>"011001001",
  62791=>"000100010",
  62792=>"110011111",
  62793=>"000110110",
  62794=>"111000011",
  62795=>"100011011",
  62796=>"100001111",
  62797=>"010000010",
  62798=>"110100111",
  62799=>"110000011",
  62800=>"111100011",
  62801=>"010110100",
  62802=>"101110111",
  62803=>"001100110",
  62804=>"000110001",
  62805=>"010011000",
  62806=>"000001101",
  62807=>"010111100",
  62808=>"010010001",
  62809=>"100010011",
  62810=>"111111101",
  62811=>"000001101",
  62812=>"110110110",
  62813=>"011111100",
  62814=>"001111100",
  62815=>"101011110",
  62816=>"101011001",
  62817=>"001000001",
  62818=>"000100000",
  62819=>"001000001",
  62820=>"000100111",
  62821=>"001100010",
  62822=>"001011000",
  62823=>"010011011",
  62824=>"101011001",
  62825=>"001010100",
  62826=>"100111011",
  62827=>"110100111",
  62828=>"000001111",
  62829=>"001000010",
  62830=>"111000100",
  62831=>"110110100",
  62832=>"101000010",
  62833=>"001111110",
  62834=>"111111111",
  62835=>"011001000",
  62836=>"011101111",
  62837=>"011100110",
  62838=>"011011000",
  62839=>"111001111",
  62840=>"101110001",
  62841=>"011101010",
  62842=>"011010011",
  62843=>"110111100",
  62844=>"101111010",
  62845=>"111000010",
  62846=>"110011101",
  62847=>"110011101",
  62848=>"100100010",
  62849=>"101011010",
  62850=>"000110001",
  62851=>"100011000",
  62852=>"010010010",
  62853=>"100101000",
  62854=>"101011110",
  62855=>"101111001",
  62856=>"100000001",
  62857=>"101001101",
  62858=>"101111110",
  62859=>"011111001",
  62860=>"110000110",
  62861=>"110000001",
  62862=>"011111100",
  62863=>"110101100",
  62864=>"001101111",
  62865=>"100100001",
  62866=>"100101011",
  62867=>"000110011",
  62868=>"100001111",
  62869=>"100101100",
  62870=>"011010010",
  62871=>"101110100",
  62872=>"110101001",
  62873=>"010001101",
  62874=>"101011111",
  62875=>"011011110",
  62876=>"011000000",
  62877=>"010011100",
  62878=>"110011000",
  62879=>"111010111",
  62880=>"111101111",
  62881=>"111101101",
  62882=>"011010110",
  62883=>"001101001",
  62884=>"011111001",
  62885=>"110011000",
  62886=>"001010000",
  62887=>"010010111",
  62888=>"010111011",
  62889=>"100000000",
  62890=>"110110111",
  62891=>"101100101",
  62892=>"101101100",
  62893=>"111101011",
  62894=>"010011000",
  62895=>"110111100",
  62896=>"100010101",
  62897=>"100001110",
  62898=>"100110011",
  62899=>"000000000",
  62900=>"011100000",
  62901=>"110010010",
  62902=>"111010011",
  62903=>"111011100",
  62904=>"101000001",
  62905=>"000010000",
  62906=>"110001010",
  62907=>"111101000",
  62908=>"110011101",
  62909=>"110101110",
  62910=>"011110010",
  62911=>"001000111",
  62912=>"100001010",
  62913=>"011001000",
  62914=>"110010000",
  62915=>"101010000",
  62916=>"110111000",
  62917=>"111010110",
  62918=>"001011101",
  62919=>"010001101",
  62920=>"000100000",
  62921=>"100100000",
  62922=>"000100110",
  62923=>"101110000",
  62924=>"011100000",
  62925=>"101100101",
  62926=>"100001010",
  62927=>"001111100",
  62928=>"110111111",
  62929=>"000010100",
  62930=>"000110111",
  62931=>"100011010",
  62932=>"000110000",
  62933=>"010100000",
  62934=>"101101101",
  62935=>"110100100",
  62936=>"100011010",
  62937=>"111111001",
  62938=>"011100001",
  62939=>"110111011",
  62940=>"011010111",
  62941=>"011000101",
  62942=>"001111111",
  62943=>"011010111",
  62944=>"111101001",
  62945=>"110111101",
  62946=>"100000101",
  62947=>"101101010",
  62948=>"110010000",
  62949=>"101110110",
  62950=>"110110111",
  62951=>"000100011",
  62952=>"011001011",
  62953=>"111110000",
  62954=>"111001011",
  62955=>"011000101",
  62956=>"000001101",
  62957=>"001101111",
  62958=>"110100011",
  62959=>"011110001",
  62960=>"111101000",
  62961=>"000000111",
  62962=>"001110100",
  62963=>"100100010",
  62964=>"001111110",
  62965=>"010111100",
  62966=>"011111110",
  62967=>"010100001",
  62968=>"001001101",
  62969=>"110011101",
  62970=>"100101110",
  62971=>"010000000",
  62972=>"111010110",
  62973=>"010010111",
  62974=>"010010101",
  62975=>"001011010",
  62976=>"100111111",
  62977=>"000111001",
  62978=>"011100111",
  62979=>"001110001",
  62980=>"000111001",
  62981=>"101111011",
  62982=>"100011010",
  62983=>"011110011",
  62984=>"010111100",
  62985=>"110101111",
  62986=>"100100100",
  62987=>"011000011",
  62988=>"000101010",
  62989=>"011100001",
  62990=>"111001011",
  62991=>"001000001",
  62992=>"001011011",
  62993=>"011111100",
  62994=>"001000010",
  62995=>"001100001",
  62996=>"100001000",
  62997=>"011001000",
  62998=>"001111111",
  62999=>"110110101",
  63000=>"010111100",
  63001=>"100011110",
  63002=>"001010001",
  63003=>"000111111",
  63004=>"101110101",
  63005=>"111101001",
  63006=>"100110101",
  63007=>"100011101",
  63008=>"001010111",
  63009=>"001001101",
  63010=>"000100001",
  63011=>"110111010",
  63012=>"101011100",
  63013=>"110100101",
  63014=>"101100011",
  63015=>"110111100",
  63016=>"111111001",
  63017=>"001000011",
  63018=>"000110010",
  63019=>"100000111",
  63020=>"100001011",
  63021=>"011101001",
  63022=>"101100111",
  63023=>"100100011",
  63024=>"111100010",
  63025=>"101011100",
  63026=>"011010000",
  63027=>"101100010",
  63028=>"110011100",
  63029=>"100100100",
  63030=>"101100100",
  63031=>"110010101",
  63032=>"000011111",
  63033=>"101010111",
  63034=>"100011111",
  63035=>"111111111",
  63036=>"001101001",
  63037=>"110010110",
  63038=>"000001110",
  63039=>"101110010",
  63040=>"001010100",
  63041=>"111010010",
  63042=>"100100110",
  63043=>"101000001",
  63044=>"000000001",
  63045=>"000111111",
  63046=>"000100101",
  63047=>"110110110",
  63048=>"011100001",
  63049=>"000110100",
  63050=>"010111001",
  63051=>"100110111",
  63052=>"101010011",
  63053=>"101111110",
  63054=>"111010101",
  63055=>"110101111",
  63056=>"100001101",
  63057=>"111101101",
  63058=>"111010101",
  63059=>"001110000",
  63060=>"000110110",
  63061=>"010101000",
  63062=>"100100100",
  63063=>"100101001",
  63064=>"010011100",
  63065=>"111011011",
  63066=>"001100010",
  63067=>"000101111",
  63068=>"100101011",
  63069=>"001010010",
  63070=>"001100111",
  63071=>"111010000",
  63072=>"011011101",
  63073=>"000001010",
  63074=>"011001010",
  63075=>"000110010",
  63076=>"010111011",
  63077=>"111111110",
  63078=>"111111011",
  63079=>"100111101",
  63080=>"011010000",
  63081=>"111110110",
  63082=>"010101011",
  63083=>"010111100",
  63084=>"101110101",
  63085=>"111001001",
  63086=>"101110000",
  63087=>"100010111",
  63088=>"100100001",
  63089=>"111000000",
  63090=>"001101101",
  63091=>"110110001",
  63092=>"010111100",
  63093=>"010001111",
  63094=>"111001001",
  63095=>"100000001",
  63096=>"010011101",
  63097=>"010011110",
  63098=>"100110111",
  63099=>"110010001",
  63100=>"011101001",
  63101=>"000001110",
  63102=>"101101111",
  63103=>"101101101",
  63104=>"110110110",
  63105=>"001100101",
  63106=>"110111110",
  63107=>"010011100",
  63108=>"010101111",
  63109=>"010111111",
  63110=>"011001000",
  63111=>"111010110",
  63112=>"000001001",
  63113=>"110000000",
  63114=>"101110001",
  63115=>"110000001",
  63116=>"011001101",
  63117=>"101100110",
  63118=>"100111010",
  63119=>"100010010",
  63120=>"111100100",
  63121=>"110100000",
  63122=>"000011000",
  63123=>"101001010",
  63124=>"010101100",
  63125=>"001000101",
  63126=>"011010010",
  63127=>"101101001",
  63128=>"011100011",
  63129=>"001000100",
  63130=>"110000001",
  63131=>"101000010",
  63132=>"010000001",
  63133=>"101101101",
  63134=>"011100000",
  63135=>"100110100",
  63136=>"001101110",
  63137=>"111010000",
  63138=>"000111110",
  63139=>"011101111",
  63140=>"111100000",
  63141=>"111110001",
  63142=>"111000100",
  63143=>"110111000",
  63144=>"111000111",
  63145=>"010110010",
  63146=>"101001110",
  63147=>"010010010",
  63148=>"010111110",
  63149=>"000000001",
  63150=>"010001010",
  63151=>"110110111",
  63152=>"110011000",
  63153=>"111110111",
  63154=>"010100100",
  63155=>"101110110",
  63156=>"001010100",
  63157=>"000111100",
  63158=>"100110111",
  63159=>"001111101",
  63160=>"001100111",
  63161=>"011011101",
  63162=>"101101101",
  63163=>"111010101",
  63164=>"111000011",
  63165=>"000100011",
  63166=>"111001100",
  63167=>"001111001",
  63168=>"010011011",
  63169=>"011000000",
  63170=>"101001000",
  63171=>"001010111",
  63172=>"000010111",
  63173=>"011110011",
  63174=>"111010011",
  63175=>"001011110",
  63176=>"011111110",
  63177=>"110000110",
  63178=>"110101010",
  63179=>"100010100",
  63180=>"011100110",
  63181=>"111001100",
  63182=>"001100001",
  63183=>"000010001",
  63184=>"101111000",
  63185=>"010011011",
  63186=>"010010101",
  63187=>"100000011",
  63188=>"001101110",
  63189=>"011000110",
  63190=>"100101111",
  63191=>"100101000",
  63192=>"000110000",
  63193=>"010111000",
  63194=>"000110000",
  63195=>"011001000",
  63196=>"010100000",
  63197=>"110111010",
  63198=>"011001111",
  63199=>"100111110",
  63200=>"110111010",
  63201=>"111111011",
  63202=>"010100100",
  63203=>"110100001",
  63204=>"011000001",
  63205=>"111111011",
  63206=>"001100001",
  63207=>"000000110",
  63208=>"001000010",
  63209=>"101101011",
  63210=>"101110001",
  63211=>"001101101",
  63212=>"101000000",
  63213=>"100100111",
  63214=>"100110000",
  63215=>"010011011",
  63216=>"000101111",
  63217=>"000011010",
  63218=>"011011100",
  63219=>"100101001",
  63220=>"111110100",
  63221=>"000001011",
  63222=>"111101000",
  63223=>"011100010",
  63224=>"000000011",
  63225=>"011000001",
  63226=>"011010110",
  63227=>"010010101",
  63228=>"001010111",
  63229=>"110111001",
  63230=>"010000000",
  63231=>"000100000",
  63232=>"001000011",
  63233=>"010101010",
  63234=>"001001110",
  63235=>"001110010",
  63236=>"110111111",
  63237=>"110100001",
  63238=>"101011000",
  63239=>"000111101",
  63240=>"100110000",
  63241=>"111001110",
  63242=>"110100000",
  63243=>"100111010",
  63244=>"111100011",
  63245=>"010000001",
  63246=>"001001011",
  63247=>"000001000",
  63248=>"111100011",
  63249=>"100010100",
  63250=>"000001000",
  63251=>"111111101",
  63252=>"010001001",
  63253=>"000010111",
  63254=>"011010111",
  63255=>"000011011",
  63256=>"000100000",
  63257=>"001100010",
  63258=>"011010001",
  63259=>"011010010",
  63260=>"111100011",
  63261=>"001011110",
  63262=>"100110010",
  63263=>"101011011",
  63264=>"101001000",
  63265=>"000001110",
  63266=>"110110110",
  63267=>"111100000",
  63268=>"011011101",
  63269=>"111110110",
  63270=>"101011111",
  63271=>"110010100",
  63272=>"100110001",
  63273=>"100101100",
  63274=>"100100000",
  63275=>"001011110",
  63276=>"011010111",
  63277=>"011001110",
  63278=>"110000100",
  63279=>"000110001",
  63280=>"111110100",
  63281=>"111101111",
  63282=>"000000101",
  63283=>"011001110",
  63284=>"110110111",
  63285=>"110000111",
  63286=>"111111111",
  63287=>"000110110",
  63288=>"101110101",
  63289=>"011110111",
  63290=>"101001111",
  63291=>"110001100",
  63292=>"111011010",
  63293=>"111001111",
  63294=>"001000001",
  63295=>"101010000",
  63296=>"101011001",
  63297=>"110101001",
  63298=>"110010010",
  63299=>"100111001",
  63300=>"100100001",
  63301=>"010011010",
  63302=>"100000100",
  63303=>"100100101",
  63304=>"110011010",
  63305=>"001001100",
  63306=>"000001111",
  63307=>"000001010",
  63308=>"001101010",
  63309=>"111101011",
  63310=>"111110110",
  63311=>"000010000",
  63312=>"100100100",
  63313=>"111100011",
  63314=>"011110111",
  63315=>"111000001",
  63316=>"101110000",
  63317=>"001000011",
  63318=>"011101001",
  63319=>"011101101",
  63320=>"111111101",
  63321=>"001100101",
  63322=>"010110110",
  63323=>"111000000",
  63324=>"100101111",
  63325=>"011011001",
  63326=>"100000111",
  63327=>"111100000",
  63328=>"110111000",
  63329=>"001101100",
  63330=>"011111100",
  63331=>"110000000",
  63332=>"110101011",
  63333=>"111111010",
  63334=>"010011110",
  63335=>"110001001",
  63336=>"111110001",
  63337=>"011100101",
  63338=>"000000100",
  63339=>"111000011",
  63340=>"010010110",
  63341=>"111000110",
  63342=>"110101110",
  63343=>"010011001",
  63344=>"110101110",
  63345=>"101110000",
  63346=>"001100100",
  63347=>"110001010",
  63348=>"001001011",
  63349=>"000100010",
  63350=>"101010000",
  63351=>"010011001",
  63352=>"001011001",
  63353=>"100001101",
  63354=>"001110100",
  63355=>"100001110",
  63356=>"010100000",
  63357=>"111010001",
  63358=>"101110010",
  63359=>"110111110",
  63360=>"011001110",
  63361=>"011110101",
  63362=>"001011100",
  63363=>"111001100",
  63364=>"101101100",
  63365=>"111000110",
  63366=>"101000000",
  63367=>"101111101",
  63368=>"000110100",
  63369=>"101010001",
  63370=>"001111010",
  63371=>"101111111",
  63372=>"101101111",
  63373=>"011001011",
  63374=>"001110010",
  63375=>"111110111",
  63376=>"100110110",
  63377=>"100000110",
  63378=>"001000100",
  63379=>"001000000",
  63380=>"101111100",
  63381=>"101100101",
  63382=>"100100010",
  63383=>"011110001",
  63384=>"001001010",
  63385=>"010111100",
  63386=>"101011010",
  63387=>"001101111",
  63388=>"111110111",
  63389=>"000011000",
  63390=>"111010110",
  63391=>"000011101",
  63392=>"101101011",
  63393=>"100111110",
  63394=>"110010001",
  63395=>"110010011",
  63396=>"011001011",
  63397=>"011100000",
  63398=>"110100111",
  63399=>"010111011",
  63400=>"000101110",
  63401=>"001110111",
  63402=>"110010111",
  63403=>"001110010",
  63404=>"000000100",
  63405=>"001111000",
  63406=>"010010101",
  63407=>"110110010",
  63408=>"011110111",
  63409=>"010101100",
  63410=>"001100101",
  63411=>"111000010",
  63412=>"011001001",
  63413=>"111001111",
  63414=>"000101011",
  63415=>"111101001",
  63416=>"101101001",
  63417=>"101100100",
  63418=>"100010100",
  63419=>"101001010",
  63420=>"010011010",
  63421=>"010101110",
  63422=>"111011100",
  63423=>"100101111",
  63424=>"001000010",
  63425=>"010011111",
  63426=>"011000000",
  63427=>"010110100",
  63428=>"110110011",
  63429=>"000100101",
  63430=>"101000000",
  63431=>"110001000",
  63432=>"001010111",
  63433=>"101000011",
  63434=>"011111111",
  63435=>"110101110",
  63436=>"001110101",
  63437=>"101101000",
  63438=>"100010110",
  63439=>"001000001",
  63440=>"000100100",
  63441=>"111010001",
  63442=>"010111100",
  63443=>"101111101",
  63444=>"010111010",
  63445=>"010000111",
  63446=>"011000110",
  63447=>"111011010",
  63448=>"011100100",
  63449=>"100111101",
  63450=>"001011111",
  63451=>"000001110",
  63452=>"011101100",
  63453=>"011000001",
  63454=>"001101101",
  63455=>"111010101",
  63456=>"011000000",
  63457=>"001001110",
  63458=>"111010111",
  63459=>"111001010",
  63460=>"010100010",
  63461=>"010000101",
  63462=>"111101001",
  63463=>"101100100",
  63464=>"101010011",
  63465=>"000001010",
  63466=>"100100001",
  63467=>"000001100",
  63468=>"011100000",
  63469=>"010110100",
  63470=>"010011001",
  63471=>"010001101",
  63472=>"100001001",
  63473=>"110100010",
  63474=>"000000010",
  63475=>"100101100",
  63476=>"111010001",
  63477=>"011011111",
  63478=>"101010000",
  63479=>"011000101",
  63480=>"110001111",
  63481=>"011011111",
  63482=>"001101101",
  63483=>"010001110",
  63484=>"101001000",
  63485=>"100000011",
  63486=>"011001000",
  63487=>"011001000",
  63488=>"000101110",
  63489=>"001000000",
  63490=>"111110101",
  63491=>"010111001",
  63492=>"111101100",
  63493=>"011110001",
  63494=>"111101100",
  63495=>"000011011",
  63496=>"000001101",
  63497=>"100101110",
  63498=>"010001000",
  63499=>"010011000",
  63500=>"010111101",
  63501=>"111000100",
  63502=>"001100011",
  63503=>"100010101",
  63504=>"100100000",
  63505=>"000111011",
  63506=>"110110011",
  63507=>"100100101",
  63508=>"101010001",
  63509=>"010100001",
  63510=>"111100110",
  63511=>"100001000",
  63512=>"011001100",
  63513=>"101010000",
  63514=>"000101111",
  63515=>"110010010",
  63516=>"110101010",
  63517=>"011101011",
  63518=>"110100000",
  63519=>"010110100",
  63520=>"100010100",
  63521=>"111000101",
  63522=>"100001110",
  63523=>"100000001",
  63524=>"000011000",
  63525=>"010000011",
  63526=>"100100000",
  63527=>"010010000",
  63528=>"010011000",
  63529=>"100100100",
  63530=>"101000110",
  63531=>"000000100",
  63532=>"100000000",
  63533=>"111001110",
  63534=>"011001011",
  63535=>"111110110",
  63536=>"111000111",
  63537=>"111111001",
  63538=>"000100101",
  63539=>"010010010",
  63540=>"101110101",
  63541=>"010111000",
  63542=>"000001000",
  63543=>"000101110",
  63544=>"011010011",
  63545=>"111010110",
  63546=>"111000000",
  63547=>"100001100",
  63548=>"011111110",
  63549=>"101100001",
  63550=>"111101000",
  63551=>"001110100",
  63552=>"100111111",
  63553=>"001010111",
  63554=>"101010101",
  63555=>"000010010",
  63556=>"011110110",
  63557=>"101000011",
  63558=>"111011111",
  63559=>"101100100",
  63560=>"011011000",
  63561=>"001001010",
  63562=>"001000101",
  63563=>"000001111",
  63564=>"111101101",
  63565=>"010001000",
  63566=>"010010011",
  63567=>"010100100",
  63568=>"110010100",
  63569=>"000010010",
  63570=>"000100001",
  63571=>"111000000",
  63572=>"111101001",
  63573=>"111011000",
  63574=>"100010110",
  63575=>"001001001",
  63576=>"010100011",
  63577=>"011010011",
  63578=>"011100110",
  63579=>"000001000",
  63580=>"000000010",
  63581=>"011100101",
  63582=>"110011110",
  63583=>"010101100",
  63584=>"001011010",
  63585=>"100100001",
  63586=>"110101000",
  63587=>"010001000",
  63588=>"011010000",
  63589=>"101101001",
  63590=>"000000110",
  63591=>"000100111",
  63592=>"110000100",
  63593=>"000011010",
  63594=>"000100001",
  63595=>"100101100",
  63596=>"110001100",
  63597=>"111101110",
  63598=>"001111101",
  63599=>"010001000",
  63600=>"001010010",
  63601=>"001001001",
  63602=>"011100110",
  63603=>"100000011",
  63604=>"000101010",
  63605=>"110011110",
  63606=>"010000111",
  63607=>"100111001",
  63608=>"110000011",
  63609=>"001010011",
  63610=>"100001110",
  63611=>"110000100",
  63612=>"110100100",
  63613=>"110000110",
  63614=>"010000010",
  63615=>"100100110",
  63616=>"010001000",
  63617=>"111010110",
  63618=>"110011000",
  63619=>"010010100",
  63620=>"100101110",
  63621=>"010001011",
  63622=>"111100010",
  63623=>"010111100",
  63624=>"010010111",
  63625=>"010100011",
  63626=>"100100011",
  63627=>"000000111",
  63628=>"100101000",
  63629=>"110000000",
  63630=>"100110111",
  63631=>"100000111",
  63632=>"101100100",
  63633=>"001000011",
  63634=>"000101111",
  63635=>"001001000",
  63636=>"101001100",
  63637=>"001111001",
  63638=>"100000001",
  63639=>"100110101",
  63640=>"101001000",
  63641=>"000001010",
  63642=>"110111011",
  63643=>"001001011",
  63644=>"001100000",
  63645=>"110110011",
  63646=>"000111011",
  63647=>"011001111",
  63648=>"110101100",
  63649=>"110111001",
  63650=>"010010100",
  63651=>"000011001",
  63652=>"001100001",
  63653=>"000001010",
  63654=>"100110101",
  63655=>"010111011",
  63656=>"111100111",
  63657=>"000011111",
  63658=>"111110110",
  63659=>"010010101",
  63660=>"000110010",
  63661=>"111010001",
  63662=>"101110001",
  63663=>"000100001",
  63664=>"111001111",
  63665=>"010111111",
  63666=>"011011010",
  63667=>"110100110",
  63668=>"001111010",
  63669=>"101000000",
  63670=>"111101011",
  63671=>"001100001",
  63672=>"000010001",
  63673=>"101110110",
  63674=>"001001110",
  63675=>"100111110",
  63676=>"010000110",
  63677=>"100110110",
  63678=>"110000000",
  63679=>"111101010",
  63680=>"000111110",
  63681=>"110001100",
  63682=>"011001011",
  63683=>"110010000",
  63684=>"110010101",
  63685=>"010100001",
  63686=>"110011110",
  63687=>"011111110",
  63688=>"101111111",
  63689=>"101010111",
  63690=>"001101010",
  63691=>"011110100",
  63692=>"011101001",
  63693=>"010000111",
  63694=>"101111100",
  63695=>"011010001",
  63696=>"111100101",
  63697=>"010011010",
  63698=>"100011110",
  63699=>"011111110",
  63700=>"100000110",
  63701=>"111010001",
  63702=>"000100110",
  63703=>"000001110",
  63704=>"011011111",
  63705=>"100110110",
  63706=>"101000010",
  63707=>"010000011",
  63708=>"111011000",
  63709=>"111111111",
  63710=>"111001111",
  63711=>"101101011",
  63712=>"011000011",
  63713=>"101101101",
  63714=>"100010111",
  63715=>"100011011",
  63716=>"111110000",
  63717=>"011011101",
  63718=>"100011101",
  63719=>"001001110",
  63720=>"100010110",
  63721=>"111001111",
  63722=>"011101111",
  63723=>"011101000",
  63724=>"000011100",
  63725=>"010110110",
  63726=>"001111110",
  63727=>"111111111",
  63728=>"111101000",
  63729=>"000001100",
  63730=>"000101111",
  63731=>"011011110",
  63732=>"110001010",
  63733=>"111001100",
  63734=>"010110111",
  63735=>"111100111",
  63736=>"011011000",
  63737=>"011100101",
  63738=>"011000111",
  63739=>"100111001",
  63740=>"001011101",
  63741=>"101101001",
  63742=>"101010011",
  63743=>"110111000",
  63744=>"000111110",
  63745=>"011001100",
  63746=>"001001111",
  63747=>"101111001",
  63748=>"111000110",
  63749=>"110011011",
  63750=>"111001110",
  63751=>"100100101",
  63752=>"000000110",
  63753=>"110011011",
  63754=>"100001011",
  63755=>"011010001",
  63756=>"011000111",
  63757=>"011011100",
  63758=>"001111000",
  63759=>"111111001",
  63760=>"111101001",
  63761=>"001000001",
  63762=>"111111101",
  63763=>"001001011",
  63764=>"111001001",
  63765=>"010011001",
  63766=>"101010011",
  63767=>"100110000",
  63768=>"111011000",
  63769=>"100000011",
  63770=>"111111001",
  63771=>"110001111",
  63772=>"101111000",
  63773=>"001010010",
  63774=>"101110111",
  63775=>"010001101",
  63776=>"001100011",
  63777=>"011111110",
  63778=>"000111110",
  63779=>"010100111",
  63780=>"011011100",
  63781=>"111110010",
  63782=>"100001000",
  63783=>"100101000",
  63784=>"101010010",
  63785=>"111111010",
  63786=>"000010101",
  63787=>"001000101",
  63788=>"010000111",
  63789=>"100100000",
  63790=>"110001111",
  63791=>"000011010",
  63792=>"010000100",
  63793=>"001101111",
  63794=>"110101111",
  63795=>"110100111",
  63796=>"001000010",
  63797=>"001111001",
  63798=>"000001100",
  63799=>"111001001",
  63800=>"010011001",
  63801=>"010011011",
  63802=>"001001011",
  63803=>"100101001",
  63804=>"111011101",
  63805=>"000001110",
  63806=>"110100101",
  63807=>"100101111",
  63808=>"101000101",
  63809=>"110010011",
  63810=>"110110110",
  63811=>"111000011",
  63812=>"111000100",
  63813=>"110111101",
  63814=>"001011001",
  63815=>"111001101",
  63816=>"110110001",
  63817=>"101001000",
  63818=>"111101001",
  63819=>"110101101",
  63820=>"111000010",
  63821=>"000110000",
  63822=>"101010001",
  63823=>"001110101",
  63824=>"101001101",
  63825=>"101001111",
  63826=>"110001001",
  63827=>"001000101",
  63828=>"110110111",
  63829=>"100110000",
  63830=>"100010010",
  63831=>"010000011",
  63832=>"110010100",
  63833=>"010110010",
  63834=>"001100010",
  63835=>"001001010",
  63836=>"101000100",
  63837=>"001011011",
  63838=>"111101100",
  63839=>"111110111",
  63840=>"010011000",
  63841=>"001101011",
  63842=>"010001001",
  63843=>"010110010",
  63844=>"000000001",
  63845=>"000101010",
  63846=>"011100001",
  63847=>"000000001",
  63848=>"110010110",
  63849=>"011010011",
  63850=>"011110101",
  63851=>"011100111",
  63852=>"011011100",
  63853=>"001000110",
  63854=>"000101010",
  63855=>"100111011",
  63856=>"110001110",
  63857=>"101100000",
  63858=>"110001000",
  63859=>"110011110",
  63860=>"101100101",
  63861=>"100001111",
  63862=>"100001010",
  63863=>"011100010",
  63864=>"000100001",
  63865=>"000001110",
  63866=>"101000010",
  63867=>"001010100",
  63868=>"010111100",
  63869=>"100000111",
  63870=>"100111000",
  63871=>"111110000",
  63872=>"101011101",
  63873=>"110110111",
  63874=>"001010010",
  63875=>"110011101",
  63876=>"101110011",
  63877=>"000001110",
  63878=>"000010111",
  63879=>"011000010",
  63880=>"001001100",
  63881=>"001100101",
  63882=>"001100111",
  63883=>"110100101",
  63884=>"110100111",
  63885=>"110111000",
  63886=>"100010111",
  63887=>"001011111",
  63888=>"101000110",
  63889=>"000101000",
  63890=>"101000001",
  63891=>"111110111",
  63892=>"010011110",
  63893=>"000110101",
  63894=>"100100010",
  63895=>"101100110",
  63896=>"011000100",
  63897=>"000011011",
  63898=>"110011111",
  63899=>"101100110",
  63900=>"000100100",
  63901=>"010011011",
  63902=>"011111101",
  63903=>"101011110",
  63904=>"100110000",
  63905=>"111010101",
  63906=>"000111111",
  63907=>"000101101",
  63908=>"101100001",
  63909=>"000011001",
  63910=>"001001100",
  63911=>"101101000",
  63912=>"110101011",
  63913=>"011101000",
  63914=>"010000001",
  63915=>"110110011",
  63916=>"100000010",
  63917=>"001010100",
  63918=>"000101111",
  63919=>"010110110",
  63920=>"100000110",
  63921=>"000111101",
  63922=>"101001110",
  63923=>"001011010",
  63924=>"011001111",
  63925=>"101101011",
  63926=>"101100110",
  63927=>"110111101",
  63928=>"111001110",
  63929=>"101110011",
  63930=>"111100100",
  63931=>"100110111",
  63932=>"100100111",
  63933=>"100100011",
  63934=>"010000111",
  63935=>"111000101",
  63936=>"011111001",
  63937=>"001111110",
  63938=>"101101000",
  63939=>"000011100",
  63940=>"100101100",
  63941=>"010011010",
  63942=>"010000011",
  63943=>"110111011",
  63944=>"000000111",
  63945=>"010110001",
  63946=>"101011110",
  63947=>"001001010",
  63948=>"010011101",
  63949=>"110001111",
  63950=>"010010000",
  63951=>"000101101",
  63952=>"111101111",
  63953=>"011000010",
  63954=>"000011001",
  63955=>"000110111",
  63956=>"000000000",
  63957=>"010011011",
  63958=>"100110000",
  63959=>"001110010",
  63960=>"100111000",
  63961=>"001000011",
  63962=>"001101010",
  63963=>"010000001",
  63964=>"100110101",
  63965=>"001111011",
  63966=>"000010111",
  63967=>"100111110",
  63968=>"010101100",
  63969=>"011110000",
  63970=>"110000001",
  63971=>"110100110",
  63972=>"000101101",
  63973=>"001011001",
  63974=>"100011011",
  63975=>"011100111",
  63976=>"001010001",
  63977=>"101110100",
  63978=>"100101101",
  63979=>"111100110",
  63980=>"100101100",
  63981=>"001001000",
  63982=>"000110101",
  63983=>"010000001",
  63984=>"011010100",
  63985=>"111100001",
  63986=>"001111011",
  63987=>"000001111",
  63988=>"101100110",
  63989=>"011001110",
  63990=>"100010000",
  63991=>"010000001",
  63992=>"101100001",
  63993=>"000010000",
  63994=>"110100100",
  63995=>"011101110",
  63996=>"010101100",
  63997=>"000000010",
  63998=>"001100110",
  63999=>"011001111",
  64000=>"010010101",
  64001=>"100011111",
  64002=>"111011001",
  64003=>"111110010",
  64004=>"100111111",
  64005=>"111111011",
  64006=>"111111111",
  64007=>"110010000",
  64008=>"000011000",
  64009=>"101111001",
  64010=>"110001011",
  64011=>"001101101",
  64012=>"001110101",
  64013=>"001110001",
  64014=>"011101010",
  64015=>"011101110",
  64016=>"100001000",
  64017=>"011011000",
  64018=>"110000101",
  64019=>"110111000",
  64020=>"100000001",
  64021=>"101001001",
  64022=>"100010111",
  64023=>"011110001",
  64024=>"001001100",
  64025=>"010101110",
  64026=>"001111101",
  64027=>"101110010",
  64028=>"011110110",
  64029=>"010111100",
  64030=>"001100111",
  64031=>"101110101",
  64032=>"101010011",
  64033=>"110001101",
  64034=>"011000000",
  64035=>"100110000",
  64036=>"010000010",
  64037=>"101110001",
  64038=>"110110000",
  64039=>"110111000",
  64040=>"001100011",
  64041=>"100001110",
  64042=>"101010010",
  64043=>"010010011",
  64044=>"011110000",
  64045=>"000000000",
  64046=>"110111101",
  64047=>"000000100",
  64048=>"000101001",
  64049=>"101010010",
  64050=>"101011110",
  64051=>"001010111",
  64052=>"010001101",
  64053=>"011001100",
  64054=>"001110000",
  64055=>"010101000",
  64056=>"000101011",
  64057=>"100011100",
  64058=>"000110011",
  64059=>"110101001",
  64060=>"100001100",
  64061=>"001110010",
  64062=>"111001101",
  64063=>"100100001",
  64064=>"101000111",
  64065=>"000001100",
  64066=>"011001111",
  64067=>"000000011",
  64068=>"011001001",
  64069=>"101111111",
  64070=>"001001011",
  64071=>"101111001",
  64072=>"011000111",
  64073=>"000000011",
  64074=>"000101111",
  64075=>"011111101",
  64076=>"001101010",
  64077=>"011000100",
  64078=>"111001001",
  64079=>"111010000",
  64080=>"100000000",
  64081=>"010000000",
  64082=>"100010001",
  64083=>"000000101",
  64084=>"011001101",
  64085=>"110000111",
  64086=>"111010110",
  64087=>"010011101",
  64088=>"110011101",
  64089=>"111000010",
  64090=>"001100100",
  64091=>"110000100",
  64092=>"000001010",
  64093=>"110101100",
  64094=>"101110011",
  64095=>"011001100",
  64096=>"110000010",
  64097=>"000001000",
  64098=>"101011001",
  64099=>"111010011",
  64100=>"011100010",
  64101=>"111001000",
  64102=>"101001011",
  64103=>"010001110",
  64104=>"101001111",
  64105=>"110101011",
  64106=>"100011110",
  64107=>"111100110",
  64108=>"111111100",
  64109=>"000101011",
  64110=>"101010011",
  64111=>"001000111",
  64112=>"110110011",
  64113=>"010111111",
  64114=>"111111101",
  64115=>"111010010",
  64116=>"111101000",
  64117=>"111111001",
  64118=>"101011000",
  64119=>"011011001",
  64120=>"011111100",
  64121=>"000011111",
  64122=>"001111100",
  64123=>"000110101",
  64124=>"000010010",
  64125=>"111000100",
  64126=>"111111100",
  64127=>"110101010",
  64128=>"011111111",
  64129=>"111000011",
  64130=>"100101000",
  64131=>"001001000",
  64132=>"110011100",
  64133=>"010010000",
  64134=>"111011100",
  64135=>"000110100",
  64136=>"111100001",
  64137=>"110000101",
  64138=>"100111111",
  64139=>"111000100",
  64140=>"101011111",
  64141=>"111111111",
  64142=>"000001100",
  64143=>"000010101",
  64144=>"110001100",
  64145=>"110100011",
  64146=>"011011000",
  64147=>"111111000",
  64148=>"100010010",
  64149=>"010011010",
  64150=>"100001010",
  64151=>"111100000",
  64152=>"010111101",
  64153=>"010101000",
  64154=>"111001100",
  64155=>"001110101",
  64156=>"000000101",
  64157=>"110011010",
  64158=>"110101100",
  64159=>"011001100",
  64160=>"101010001",
  64161=>"001100101",
  64162=>"100011110",
  64163=>"101011101",
  64164=>"011111101",
  64165=>"101011010",
  64166=>"011011101",
  64167=>"111101100",
  64168=>"110101110",
  64169=>"000111001",
  64170=>"001111101",
  64171=>"100111010",
  64172=>"110000010",
  64173=>"000100000",
  64174=>"000010000",
  64175=>"010001001",
  64176=>"011011000",
  64177=>"110101000",
  64178=>"101100111",
  64179=>"101100001",
  64180=>"010010110",
  64181=>"010001010",
  64182=>"111110001",
  64183=>"111111101",
  64184=>"010101110",
  64185=>"110111111",
  64186=>"011100110",
  64187=>"001001001",
  64188=>"001011000",
  64189=>"001110101",
  64190=>"011111000",
  64191=>"000010111",
  64192=>"110111110",
  64193=>"101011000",
  64194=>"111110001",
  64195=>"010100110",
  64196=>"011110100",
  64197=>"110100101",
  64198=>"100010111",
  64199=>"101101101",
  64200=>"010001101",
  64201=>"011000100",
  64202=>"110011001",
  64203=>"001111011",
  64204=>"101010001",
  64205=>"000111111",
  64206=>"010110011",
  64207=>"110110101",
  64208=>"100100101",
  64209=>"111010010",
  64210=>"000001011",
  64211=>"001000011",
  64212=>"011001101",
  64213=>"010010010",
  64214=>"000011111",
  64215=>"101010000",
  64216=>"010011010",
  64217=>"100000000",
  64218=>"110111110",
  64219=>"100011111",
  64220=>"000110011",
  64221=>"100000111",
  64222=>"101001001",
  64223=>"111001100",
  64224=>"101000000",
  64225=>"010110111",
  64226=>"111000100",
  64227=>"111110100",
  64228=>"111000010",
  64229=>"101001101",
  64230=>"110110111",
  64231=>"100001100",
  64232=>"000110101",
  64233=>"001011011",
  64234=>"000011011",
  64235=>"011100111",
  64236=>"100010010",
  64237=>"011101100",
  64238=>"010111001",
  64239=>"011001100",
  64240=>"000011100",
  64241=>"001101110",
  64242=>"101110001",
  64243=>"011110100",
  64244=>"110110111",
  64245=>"001111001",
  64246=>"110101111",
  64247=>"100101001",
  64248=>"110001110",
  64249=>"011011011",
  64250=>"000001001",
  64251=>"001001100",
  64252=>"010100111",
  64253=>"101010110",
  64254=>"001100110",
  64255=>"010100100",
  64256=>"000100011",
  64257=>"001111000",
  64258=>"000100101",
  64259=>"100000011",
  64260=>"100011000",
  64261=>"000111010",
  64262=>"101001110",
  64263=>"100010111",
  64264=>"001000010",
  64265=>"101011111",
  64266=>"001011010",
  64267=>"110010000",
  64268=>"001000000",
  64269=>"110100010",
  64270=>"000111100",
  64271=>"101111101",
  64272=>"000001110",
  64273=>"001011101",
  64274=>"011111000",
  64275=>"001000111",
  64276=>"100111010",
  64277=>"110010010",
  64278=>"001111000",
  64279=>"011110000",
  64280=>"111001001",
  64281=>"001001101",
  64282=>"000110111",
  64283=>"110000110",
  64284=>"111100001",
  64285=>"010101000",
  64286=>"011010010",
  64287=>"110000110",
  64288=>"001101011",
  64289=>"100100011",
  64290=>"001011011",
  64291=>"011111000",
  64292=>"111000000",
  64293=>"101110011",
  64294=>"011010111",
  64295=>"101100101",
  64296=>"111010110",
  64297=>"000001111",
  64298=>"110111101",
  64299=>"101101010",
  64300=>"111101100",
  64301=>"000010011",
  64302=>"100001011",
  64303=>"110010101",
  64304=>"101011001",
  64305=>"100101111",
  64306=>"010010110",
  64307=>"111010010",
  64308=>"110010101",
  64309=>"100010101",
  64310=>"011110111",
  64311=>"011010100",
  64312=>"101011000",
  64313=>"101110111",
  64314=>"101011010",
  64315=>"100110011",
  64316=>"000001010",
  64317=>"111101010",
  64318=>"101110111",
  64319=>"101101111",
  64320=>"000011000",
  64321=>"100010100",
  64322=>"010110111",
  64323=>"010110000",
  64324=>"011001001",
  64325=>"000101100",
  64326=>"000001001",
  64327=>"010111001",
  64328=>"110101010",
  64329=>"111101111",
  64330=>"011001010",
  64331=>"011001101",
  64332=>"000011101",
  64333=>"110001101",
  64334=>"111100111",
  64335=>"001010100",
  64336=>"000010010",
  64337=>"011010100",
  64338=>"010000000",
  64339=>"001010100",
  64340=>"000110011",
  64341=>"101001001",
  64342=>"111000111",
  64343=>"001110100",
  64344=>"110001111",
  64345=>"110111011",
  64346=>"000010011",
  64347=>"111000111",
  64348=>"001100010",
  64349=>"111000000",
  64350=>"010001001",
  64351=>"000101001",
  64352=>"101110011",
  64353=>"110001101",
  64354=>"010100001",
  64355=>"101111001",
  64356=>"010010000",
  64357=>"011101110",
  64358=>"010010000",
  64359=>"101011000",
  64360=>"101111000",
  64361=>"000100001",
  64362=>"100011001",
  64363=>"011110111",
  64364=>"010100111",
  64365=>"011110010",
  64366=>"001101110",
  64367=>"011101001",
  64368=>"001001000",
  64369=>"001111010",
  64370=>"100011010",
  64371=>"110101111",
  64372=>"000011010",
  64373=>"000001000",
  64374=>"001001100",
  64375=>"101101111",
  64376=>"111011001",
  64377=>"101000011",
  64378=>"010000110",
  64379=>"111000010",
  64380=>"000000000",
  64381=>"011011010",
  64382=>"010111000",
  64383=>"110111001",
  64384=>"000111101",
  64385=>"000010101",
  64386=>"110010010",
  64387=>"000110110",
  64388=>"110001110",
  64389=>"101101101",
  64390=>"111111100",
  64391=>"000110001",
  64392=>"111011111",
  64393=>"110111011",
  64394=>"101011011",
  64395=>"010111101",
  64396=>"110111101",
  64397=>"011101010",
  64398=>"100001111",
  64399=>"001000010",
  64400=>"011110011",
  64401=>"100010101",
  64402=>"010100001",
  64403=>"001001101",
  64404=>"000101001",
  64405=>"101011111",
  64406=>"110010000",
  64407=>"100001101",
  64408=>"000110101",
  64409=>"100010000",
  64410=>"010001110",
  64411=>"000011110",
  64412=>"001000101",
  64413=>"010011000",
  64414=>"101110001",
  64415=>"101010000",
  64416=>"011100011",
  64417=>"001001000",
  64418=>"001011100",
  64419=>"100000000",
  64420=>"101000011",
  64421=>"010100100",
  64422=>"000011111",
  64423=>"101000111",
  64424=>"011000010",
  64425=>"001001011",
  64426=>"111000000",
  64427=>"100111011",
  64428=>"011100111",
  64429=>"010010111",
  64430=>"001100111",
  64431=>"100000000",
  64432=>"101011000",
  64433=>"010100110",
  64434=>"000100010",
  64435=>"001011001",
  64436=>"111011001",
  64437=>"101000010",
  64438=>"000000100",
  64439=>"100001000",
  64440=>"000001111",
  64441=>"011011110",
  64442=>"111111010",
  64443=>"100101001",
  64444=>"000000110",
  64445=>"100111010",
  64446=>"111000000",
  64447=>"011111000",
  64448=>"010110110",
  64449=>"010011110",
  64450=>"001000100",
  64451=>"100110001",
  64452=>"001100110",
  64453=>"101111010",
  64454=>"110101000",
  64455=>"100011101",
  64456=>"000010000",
  64457=>"011000001",
  64458=>"110100011",
  64459=>"110110001",
  64460=>"000100111",
  64461=>"010011010",
  64462=>"111110101",
  64463=>"011100011",
  64464=>"010000001",
  64465=>"001010101",
  64466=>"010111111",
  64467=>"011100100",
  64468=>"101101010",
  64469=>"111111110",
  64470=>"001001000",
  64471=>"110010010",
  64472=>"000111101",
  64473=>"100011011",
  64474=>"100101111",
  64475=>"010101110",
  64476=>"101000011",
  64477=>"000111110",
  64478=>"101101001",
  64479=>"111001010",
  64480=>"011000111",
  64481=>"011010001",
  64482=>"010001111",
  64483=>"100100111",
  64484=>"001111100",
  64485=>"111010111",
  64486=>"000001001",
  64487=>"011010011",
  64488=>"101000100",
  64489=>"000101011",
  64490=>"110100010",
  64491=>"111011110",
  64492=>"011011111",
  64493=>"000000001",
  64494=>"110100001",
  64495=>"000111111",
  64496=>"001001100",
  64497=>"011100011",
  64498=>"011101010",
  64499=>"101010001",
  64500=>"110001100",
  64501=>"111011101",
  64502=>"110100110",
  64503=>"110110111",
  64504=>"010001101",
  64505=>"100001001",
  64506=>"101110101",
  64507=>"111001100",
  64508=>"001111110",
  64509=>"111101110",
  64510=>"101000000",
  64511=>"011101000",
  64512=>"101111101",
  64513=>"011110000",
  64514=>"100110100",
  64515=>"111101110",
  64516=>"000000010",
  64517=>"000011111",
  64518=>"001001001",
  64519=>"001011100",
  64520=>"101001010",
  64521=>"010111001",
  64522=>"000001010",
  64523=>"110110111",
  64524=>"110101011",
  64525=>"000001110",
  64526=>"110011010",
  64527=>"001011110",
  64528=>"111001110",
  64529=>"100001001",
  64530=>"010001000",
  64531=>"000010001",
  64532=>"110001010",
  64533=>"101000110",
  64534=>"101011100",
  64535=>"101000101",
  64536=>"111111000",
  64537=>"010010110",
  64538=>"000100001",
  64539=>"101110001",
  64540=>"011011010",
  64541=>"111110010",
  64542=>"001010101",
  64543=>"000011100",
  64544=>"110101101",
  64545=>"100011110",
  64546=>"111110010",
  64547=>"110001110",
  64548=>"000000000",
  64549=>"000011110",
  64550=>"010011101",
  64551=>"111110101",
  64552=>"111011101",
  64553=>"010101100",
  64554=>"110001011",
  64555=>"101001100",
  64556=>"010000100",
  64557=>"000010100",
  64558=>"110101111",
  64559=>"101011101",
  64560=>"110101011",
  64561=>"010101010",
  64562=>"011011101",
  64563=>"111000101",
  64564=>"011110110",
  64565=>"101001111",
  64566=>"101000101",
  64567=>"010000101",
  64568=>"100010100",
  64569=>"100010010",
  64570=>"111101111",
  64571=>"001101001",
  64572=>"100110001",
  64573=>"111101001",
  64574=>"110101111",
  64575=>"001001010",
  64576=>"111010011",
  64577=>"000000001",
  64578=>"111001001",
  64579=>"011100111",
  64580=>"110110001",
  64581=>"100001101",
  64582=>"100110000",
  64583=>"100101010",
  64584=>"111011111",
  64585=>"011000100",
  64586=>"101011000",
  64587=>"001111101",
  64588=>"110100101",
  64589=>"111110111",
  64590=>"110111100",
  64591=>"101010110",
  64592=>"101101010",
  64593=>"111010110",
  64594=>"100010110",
  64595=>"010110001",
  64596=>"110101001",
  64597=>"000111000",
  64598=>"110000011",
  64599=>"101000100",
  64600=>"110101110",
  64601=>"100110010",
  64602=>"000110101",
  64603=>"001100101",
  64604=>"011001101",
  64605=>"000011101",
  64606=>"110110011",
  64607=>"111111000",
  64608=>"011010100",
  64609=>"101110101",
  64610=>"100101111",
  64611=>"011100000",
  64612=>"100101011",
  64613=>"011110000",
  64614=>"010101010",
  64615=>"001111000",
  64616=>"110001011",
  64617=>"001100000",
  64618=>"010000010",
  64619=>"010110001",
  64620=>"101011101",
  64621=>"010110110",
  64622=>"011001110",
  64623=>"011110101",
  64624=>"110101010",
  64625=>"010011001",
  64626=>"111001111",
  64627=>"010110111",
  64628=>"010111001",
  64629=>"101101001",
  64630=>"000100000",
  64631=>"110001001",
  64632=>"001100100",
  64633=>"100011010",
  64634=>"111001001",
  64635=>"011110111",
  64636=>"101100100",
  64637=>"111100111",
  64638=>"111001111",
  64639=>"010101001",
  64640=>"110000100",
  64641=>"000010010",
  64642=>"000011000",
  64643=>"011111000",
  64644=>"001101111",
  64645=>"100001010",
  64646=>"001111000",
  64647=>"101101000",
  64648=>"111110111",
  64649=>"001101010",
  64650=>"110011110",
  64651=>"111110011",
  64652=>"000010001",
  64653=>"111111001",
  64654=>"110000110",
  64655=>"101110110",
  64656=>"010001111",
  64657=>"111011011",
  64658=>"111000101",
  64659=>"011101101",
  64660=>"100010011",
  64661=>"101100000",
  64662=>"001000101",
  64663=>"010111001",
  64664=>"000010100",
  64665=>"111001110",
  64666=>"100000100",
  64667=>"000110100",
  64668=>"010010100",
  64669=>"101110011",
  64670=>"101100011",
  64671=>"110100001",
  64672=>"000000001",
  64673=>"011100001",
  64674=>"011000010",
  64675=>"010011010",
  64676=>"000001000",
  64677=>"101011111",
  64678=>"000000001",
  64679=>"001011000",
  64680=>"100101010",
  64681=>"000000110",
  64682=>"011110110",
  64683=>"101001100",
  64684=>"011010000",
  64685=>"111101101",
  64686=>"010111011",
  64687=>"100101010",
  64688=>"001111101",
  64689=>"000101010",
  64690=>"010110010",
  64691=>"101010101",
  64692=>"100010101",
  64693=>"010110111",
  64694=>"011001000",
  64695=>"001010000",
  64696=>"111000001",
  64697=>"010000000",
  64698=>"100000010",
  64699=>"000110111",
  64700=>"101110001",
  64701=>"100100110",
  64702=>"011000001",
  64703=>"111111011",
  64704=>"111110010",
  64705=>"110101000",
  64706=>"110010100",
  64707=>"111001101",
  64708=>"101010000",
  64709=>"001111100",
  64710=>"111010011",
  64711=>"011001111",
  64712=>"100010101",
  64713=>"111111111",
  64714=>"110001010",
  64715=>"001100101",
  64716=>"000110100",
  64717=>"011111111",
  64718=>"101101101",
  64719=>"100001110",
  64720=>"001110000",
  64721=>"010100001",
  64722=>"011011001",
  64723=>"011000010",
  64724=>"101100000",
  64725=>"110011110",
  64726=>"100000011",
  64727=>"010001100",
  64728=>"100001101",
  64729=>"001011100",
  64730=>"000000000",
  64731=>"111010000",
  64732=>"011001111",
  64733=>"100101110",
  64734=>"000110110",
  64735=>"001111011",
  64736=>"001010101",
  64737=>"100000110",
  64738=>"110010100",
  64739=>"010010101",
  64740=>"011001100",
  64741=>"110011001",
  64742=>"110110110",
  64743=>"001010010",
  64744=>"100000010",
  64745=>"110100101",
  64746=>"100011100",
  64747=>"100001001",
  64748=>"100001110",
  64749=>"000001011",
  64750=>"000000111",
  64751=>"011111011",
  64752=>"111010111",
  64753=>"100001010",
  64754=>"101011110",
  64755=>"110111100",
  64756=>"100010001",
  64757=>"011010000",
  64758=>"001111011",
  64759=>"000100101",
  64760=>"000010111",
  64761=>"001001101",
  64762=>"101100100",
  64763=>"000100011",
  64764=>"011111110",
  64765=>"010011000",
  64766=>"100100001",
  64767=>"000100100",
  64768=>"111101010",
  64769=>"101111000",
  64770=>"000100111",
  64771=>"011000001",
  64772=>"100001100",
  64773=>"000000110",
  64774=>"010001010",
  64775=>"110001101",
  64776=>"100111101",
  64777=>"011101011",
  64778=>"110111000",
  64779=>"101111101",
  64780=>"001011011",
  64781=>"010110000",
  64782=>"010100010",
  64783=>"000000000",
  64784=>"111111010",
  64785=>"111000100",
  64786=>"111001111",
  64787=>"001001000",
  64788=>"111111111",
  64789=>"001100101",
  64790=>"000101110",
  64791=>"010010011",
  64792=>"101111100",
  64793=>"001001001",
  64794=>"100110000",
  64795=>"001010001",
  64796=>"100100100",
  64797=>"111001100",
  64798=>"011111111",
  64799=>"100010000",
  64800=>"001010101",
  64801=>"101000010",
  64802=>"000101011",
  64803=>"000110000",
  64804=>"111010010",
  64805=>"000111000",
  64806=>"100011101",
  64807=>"011111010",
  64808=>"010001000",
  64809=>"101000010",
  64810=>"111111011",
  64811=>"001111110",
  64812=>"000011000",
  64813=>"100110101",
  64814=>"010011100",
  64815=>"000001010",
  64816=>"000101110",
  64817=>"111111011",
  64818=>"101011000",
  64819=>"100111011",
  64820=>"111010001",
  64821=>"000000001",
  64822=>"011000101",
  64823=>"011100111",
  64824=>"010001010",
  64825=>"000101110",
  64826=>"101001001",
  64827=>"001111100",
  64828=>"000110110",
  64829=>"111011100",
  64830=>"000001100",
  64831=>"110101110",
  64832=>"011001110",
  64833=>"100110111",
  64834=>"010100010",
  64835=>"110110111",
  64836=>"010111000",
  64837=>"101100101",
  64838=>"000001100",
  64839=>"101011000",
  64840=>"000000101",
  64841=>"001100010",
  64842=>"110100011",
  64843=>"000101110",
  64844=>"000010001",
  64845=>"000101110",
  64846=>"000111100",
  64847=>"101110011",
  64848=>"100010111",
  64849=>"101001010",
  64850=>"110111110",
  64851=>"100100111",
  64852=>"000100000",
  64853=>"010111100",
  64854=>"101110100",
  64855=>"110111110",
  64856=>"001100000",
  64857=>"100011101",
  64858=>"101001011",
  64859=>"111000111",
  64860=>"101100001",
  64861=>"000001011",
  64862=>"100111011",
  64863=>"011000001",
  64864=>"001011100",
  64865=>"001001111",
  64866=>"100110101",
  64867=>"001000011",
  64868=>"000000101",
  64869=>"011110101",
  64870=>"010110111",
  64871=>"111111011",
  64872=>"001010110",
  64873=>"000000001",
  64874=>"000001110",
  64875=>"000000110",
  64876=>"010011010",
  64877=>"110001101",
  64878=>"011101110",
  64879=>"000001000",
  64880=>"100010100",
  64881=>"000101100",
  64882=>"001101111",
  64883=>"010111011",
  64884=>"000011010",
  64885=>"000010001",
  64886=>"101111110",
  64887=>"010101011",
  64888=>"010001111",
  64889=>"010010110",
  64890=>"011111010",
  64891=>"001100011",
  64892=>"100110110",
  64893=>"111100010",
  64894=>"100111000",
  64895=>"100000111",
  64896=>"001000110",
  64897=>"000101111",
  64898=>"010101111",
  64899=>"000011111",
  64900=>"011011101",
  64901=>"100100010",
  64902=>"110111010",
  64903=>"001100100",
  64904=>"011001111",
  64905=>"101000111",
  64906=>"000101100",
  64907=>"000111111",
  64908=>"101001100",
  64909=>"100110111",
  64910=>"101111001",
  64911=>"100011011",
  64912=>"110010000",
  64913=>"001000010",
  64914=>"000110100",
  64915=>"101001110",
  64916=>"011100010",
  64917=>"100110000",
  64918=>"100111000",
  64919=>"011111101",
  64920=>"111110101",
  64921=>"010000111",
  64922=>"101111110",
  64923=>"100111000",
  64924=>"111111100",
  64925=>"010011000",
  64926=>"111111011",
  64927=>"110101000",
  64928=>"010000001",
  64929=>"100010001",
  64930=>"011110011",
  64931=>"111101100",
  64932=>"110110100",
  64933=>"101001000",
  64934=>"010100110",
  64935=>"011010100",
  64936=>"010010001",
  64937=>"010011000",
  64938=>"001111001",
  64939=>"000000110",
  64940=>"000001110",
  64941=>"001101101",
  64942=>"001101010",
  64943=>"111110010",
  64944=>"001001010",
  64945=>"000011001",
  64946=>"000001000",
  64947=>"000001011",
  64948=>"001001111",
  64949=>"101000110",
  64950=>"100001110",
  64951=>"011011000",
  64952=>"010110011",
  64953=>"000000101",
  64954=>"101111101",
  64955=>"001101100",
  64956=>"001110011",
  64957=>"111100011",
  64958=>"100111010",
  64959=>"100011011",
  64960=>"000101101",
  64961=>"011010000",
  64962=>"011001110",
  64963=>"011010011",
  64964=>"010111111",
  64965=>"100100001",
  64966=>"001110011",
  64967=>"101000100",
  64968=>"110011011",
  64969=>"100110011",
  64970=>"011011000",
  64971=>"110010001",
  64972=>"000001000",
  64973=>"011101010",
  64974=>"101111010",
  64975=>"010001101",
  64976=>"110101111",
  64977=>"010110011",
  64978=>"011001011",
  64979=>"111100101",
  64980=>"110110001",
  64981=>"011111111",
  64982=>"011000001",
  64983=>"001001000",
  64984=>"100111011",
  64985=>"111101000",
  64986=>"111001000",
  64987=>"110111001",
  64988=>"001100001",
  64989=>"111000111",
  64990=>"111101001",
  64991=>"001100000",
  64992=>"111000010",
  64993=>"100011010",
  64994=>"010110010",
  64995=>"100011100",
  64996=>"111001001",
  64997=>"110010000",
  64998=>"000010110",
  64999=>"000001000",
  65000=>"000100001",
  65001=>"000100100",
  65002=>"000000001",
  65003=>"000111110",
  65004=>"111101001",
  65005=>"111101101",
  65006=>"010000001",
  65007=>"100001000",
  65008=>"000010000",
  65009=>"000110010",
  65010=>"010010011",
  65011=>"000010110",
  65012=>"101001000",
  65013=>"001111011",
  65014=>"110001110",
  65015=>"000011111",
  65016=>"000011000",
  65017=>"011101110",
  65018=>"101101100",
  65019=>"010001111",
  65020=>"000000010",
  65021=>"010000101",
  65022=>"110101010",
  65023=>"001101010",
  65024=>"001001000",
  65025=>"110110111",
  65026=>"111110110",
  65027=>"011100111",
  65028=>"001101110",
  65029=>"111001011",
  65030=>"010100010",
  65031=>"101011000",
  65032=>"111010100",
  65033=>"001110100",
  65034=>"010010110",
  65035=>"100110100",
  65036=>"110101111",
  65037=>"001100101",
  65038=>"001011111",
  65039=>"111101001",
  65040=>"101000000",
  65041=>"010000011",
  65042=>"111001011",
  65043=>"010110001",
  65044=>"101110101",
  65045=>"110100100",
  65046=>"110010111",
  65047=>"110000000",
  65048=>"000000100",
  65049=>"000010000",
  65050=>"011010100",
  65051=>"110001000",
  65052=>"111100001",
  65053=>"111111000",
  65054=>"110101000",
  65055=>"110110110",
  65056=>"111010000",
  65057=>"110011000",
  65058=>"000110100",
  65059=>"010010001",
  65060=>"001000011",
  65061=>"001110000",
  65062=>"000000111",
  65063=>"010000100",
  65064=>"110000010",
  65065=>"100001010",
  65066=>"101111111",
  65067=>"110000011",
  65068=>"101101000",
  65069=>"101110100",
  65070=>"110011100",
  65071=>"100110010",
  65072=>"010001001",
  65073=>"110000010",
  65074=>"000101101",
  65075=>"100111111",
  65076=>"100101000",
  65077=>"011000011",
  65078=>"001101110",
  65079=>"111110100",
  65080=>"111110001",
  65081=>"111000001",
  65082=>"101011000",
  65083=>"001000101",
  65084=>"110100011",
  65085=>"000000110",
  65086=>"010010001",
  65087=>"001110000",
  65088=>"001010101",
  65089=>"010000100",
  65090=>"000011010",
  65091=>"111100111",
  65092=>"010001100",
  65093=>"101110010",
  65094=>"111001001",
  65095=>"000100100",
  65096=>"111010111",
  65097=>"011010100",
  65098=>"100000101",
  65099=>"100001101",
  65100=>"010100111",
  65101=>"000011101",
  65102=>"000110101",
  65103=>"111001101",
  65104=>"010001101",
  65105=>"001001000",
  65106=>"001111001",
  65107=>"011000111",
  65108=>"011101100",
  65109=>"010000110",
  65110=>"100100000",
  65111=>"000111111",
  65112=>"111101111",
  65113=>"000001001",
  65114=>"101101011",
  65115=>"000001001",
  65116=>"100000100",
  65117=>"010000100",
  65118=>"000011110",
  65119=>"000000101",
  65120=>"010100000",
  65121=>"001110100",
  65122=>"010100100",
  65123=>"011100101",
  65124=>"101000001",
  65125=>"110001000",
  65126=>"100000100",
  65127=>"010111100",
  65128=>"110110111",
  65129=>"001101010",
  65130=>"000110000",
  65131=>"010000100",
  65132=>"000110110",
  65133=>"111100011",
  65134=>"001001111",
  65135=>"110000100",
  65136=>"010010000",
  65137=>"000110101",
  65138=>"111010000",
  65139=>"110010001",
  65140=>"100011111",
  65141=>"011000100",
  65142=>"110011101",
  65143=>"100001100",
  65144=>"001000000",
  65145=>"100111101",
  65146=>"110100010",
  65147=>"101101110",
  65148=>"010110100",
  65149=>"100101101",
  65150=>"000010010",
  65151=>"011101100",
  65152=>"001011010",
  65153=>"011011101",
  65154=>"001101011",
  65155=>"111101001",
  65156=>"000111010",
  65157=>"001111101",
  65158=>"001111110",
  65159=>"101001111",
  65160=>"101100001",
  65161=>"110111111",
  65162=>"111101010",
  65163=>"010110101",
  65164=>"101000100",
  65165=>"111100000",
  65166=>"101101100",
  65167=>"010101011",
  65168=>"101111110",
  65169=>"110011000",
  65170=>"111111100",
  65171=>"010001101",
  65172=>"000001100",
  65173=>"010101000",
  65174=>"101111010",
  65175=>"001101101",
  65176=>"100111100",
  65177=>"101111110",
  65178=>"111110010",
  65179=>"001001010",
  65180=>"001011100",
  65181=>"000011001",
  65182=>"010010001",
  65183=>"000110001",
  65184=>"110000000",
  65185=>"001011001",
  65186=>"101010101",
  65187=>"111101011",
  65188=>"000010010",
  65189=>"000011000",
  65190=>"000100111",
  65191=>"010011000",
  65192=>"110110101",
  65193=>"001001000",
  65194=>"001001011",
  65195=>"110001101",
  65196=>"111101110",
  65197=>"011010001",
  65198=>"110101110",
  65199=>"000000011",
  65200=>"000100111",
  65201=>"110011100",
  65202=>"101010010",
  65203=>"101011010",
  65204=>"100100111",
  65205=>"110000111",
  65206=>"001011110",
  65207=>"000110001",
  65208=>"001000101",
  65209=>"110101000",
  65210=>"000111111",
  65211=>"011010100",
  65212=>"110100000",
  65213=>"011110011",
  65214=>"100000100",
  65215=>"100001010",
  65216=>"111100101",
  65217=>"100111000",
  65218=>"010111001",
  65219=>"001010011",
  65220=>"001000110",
  65221=>"000010010",
  65222=>"100100010",
  65223=>"111001000",
  65224=>"011000011",
  65225=>"011011001",
  65226=>"111100111",
  65227=>"101111100",
  65228=>"001011000",
  65229=>"111110001",
  65230=>"100111011",
  65231=>"001010101",
  65232=>"100100011",
  65233=>"000000010",
  65234=>"001101000",
  65235=>"000011001",
  65236=>"011101000",
  65237=>"010010001",
  65238=>"100011010",
  65239=>"001110001",
  65240=>"000111100",
  65241=>"100011101",
  65242=>"100000101",
  65243=>"000110101",
  65244=>"101100000",
  65245=>"000100010",
  65246=>"000011110",
  65247=>"111111100",
  65248=>"110100110",
  65249=>"010001110",
  65250=>"100100111",
  65251=>"000000110",
  65252=>"110000010",
  65253=>"110000101",
  65254=>"011100000",
  65255=>"110110110",
  65256=>"110011000",
  65257=>"101001001",
  65258=>"000010101",
  65259=>"101010000",
  65260=>"000000011",
  65261=>"011000111",
  65262=>"111110111",
  65263=>"010111011",
  65264=>"101001000",
  65265=>"011110111",
  65266=>"010000011",
  65267=>"101111100",
  65268=>"111111110",
  65269=>"110011110",
  65270=>"110010010",
  65271=>"100011101",
  65272=>"010000111",
  65273=>"010100110",
  65274=>"011010111",
  65275=>"010110001",
  65276=>"011001110",
  65277=>"111111101",
  65278=>"101110110",
  65279=>"001101111",
  65280=>"001011010",
  65281=>"000101011",
  65282=>"111010111",
  65283=>"000000110",
  65284=>"010101010",
  65285=>"001001000",
  65286=>"001010010",
  65287=>"110000100",
  65288=>"000000000",
  65289=>"100010010",
  65290=>"100101010",
  65291=>"000101110",
  65292=>"111110100",
  65293=>"111110110",
  65294=>"111010000",
  65295=>"111111011",
  65296=>"101100101",
  65297=>"000000001",
  65298=>"001101100",
  65299=>"110011001",
  65300=>"100000110",
  65301=>"001111100",
  65302=>"101010001",
  65303=>"000011001",
  65304=>"001001110",
  65305=>"011101010",
  65306=>"000111110",
  65307=>"010010110",
  65308=>"100001111",
  65309=>"101111011",
  65310=>"110010111",
  65311=>"111011011",
  65312=>"011001100",
  65313=>"110001010",
  65314=>"111001100",
  65315=>"111010000",
  65316=>"000110101",
  65317=>"000000111",
  65318=>"010001011",
  65319=>"111110001",
  65320=>"000111011",
  65321=>"000001001",
  65322=>"010000000",
  65323=>"000010010",
  65324=>"011110111",
  65325=>"000001010",
  65326=>"010101100",
  65327=>"111111000",
  65328=>"100011110",
  65329=>"011001111",
  65330=>"001110001",
  65331=>"100000101",
  65332=>"010011000",
  65333=>"111001000",
  65334=>"010111011",
  65335=>"000111101",
  65336=>"100111000",
  65337=>"100011010",
  65338=>"000011011",
  65339=>"001111111",
  65340=>"110011110",
  65341=>"001110010",
  65342=>"001000100",
  65343=>"101011010",
  65344=>"100010110",
  65345=>"000000000",
  65346=>"001111001",
  65347=>"101100101",
  65348=>"001101100",
  65349=>"000001010",
  65350=>"000100100",
  65351=>"111100000",
  65352=>"110011111",
  65353=>"001110110",
  65354=>"000110101",
  65355=>"101011011",
  65356=>"100111100",
  65357=>"011001110",
  65358=>"001100001",
  65359=>"011110011",
  65360=>"100110101",
  65361=>"011010000",
  65362=>"001101000",
  65363=>"000000101",
  65364=>"011111001",
  65365=>"000100111",
  65366=>"001010000",
  65367=>"010001010",
  65368=>"100001101",
  65369=>"111111001",
  65370=>"011001101",
  65371=>"101101010",
  65372=>"101101001",
  65373=>"010100110",
  65374=>"111001000",
  65375=>"000001111",
  65376=>"100001101",
  65377=>"011000010",
  65378=>"000010101",
  65379=>"010011010",
  65380=>"010011100",
  65381=>"100010011",
  65382=>"101011110",
  65383=>"100110100",
  65384=>"111110011",
  65385=>"000010010",
  65386=>"011100011",
  65387=>"011101001",
  65388=>"111011001",
  65389=>"011100110",
  65390=>"110101110",
  65391=>"110101111",
  65392=>"001101011",
  65393=>"011100001",
  65394=>"110010100",
  65395=>"011010010",
  65396=>"110100011",
  65397=>"011011001",
  65398=>"011100000",
  65399=>"110111100",
  65400=>"001011010",
  65401=>"001101100",
  65402=>"111000000",
  65403=>"000001010",
  65404=>"000111101",
  65405=>"000111011",
  65406=>"001101000",
  65407=>"111111110",
  65408=>"100010010",
  65409=>"010000001",
  65410=>"001100011",
  65411=>"110101111",
  65412=>"000110110",
  65413=>"010111100",
  65414=>"001011011",
  65415=>"111011010",
  65416=>"100101001",
  65417=>"001000110",
  65418=>"101111011",
  65419=>"000010110",
  65420=>"101001000",
  65421=>"101011000",
  65422=>"110011000",
  65423=>"100000011",
  65424=>"011010110",
  65425=>"111010111",
  65426=>"010111001",
  65427=>"110011000",
  65428=>"001011100",
  65429=>"111111011",
  65430=>"111000000",
  65431=>"110110001",
  65432=>"100011011",
  65433=>"110110000",
  65434=>"001100101",
  65435=>"001011001",
  65436=>"101111110",
  65437=>"011000000",
  65438=>"010010000",
  65439=>"001001111",
  65440=>"000001000",
  65441=>"010110000",
  65442=>"000110111",
  65443=>"000111001",
  65444=>"010000100",
  65445=>"101011111",
  65446=>"100011111",
  65447=>"110010101",
  65448=>"011111111",
  65449=>"001101111",
  65450=>"001011101",
  65451=>"111000111",
  65452=>"101011000",
  65453=>"101011001",
  65454=>"110110110",
  65455=>"010001001",
  65456=>"001000101",
  65457=>"110011111",
  65458=>"010101100",
  65459=>"101001001",
  65460=>"000011011",
  65461=>"110000110",
  65462=>"111000110",
  65463=>"111100101",
  65464=>"101000010",
  65465=>"000111010",
  65466=>"010001111",
  65467=>"110010011",
  65468=>"000111100",
  65469=>"100000010",
  65470=>"011010001",
  65471=>"101010111",
  65472=>"001101111",
  65473=>"011101101",
  65474=>"000001011",
  65475=>"010111011",
  65476=>"010000110",
  65477=>"111010100",
  65478=>"001101111",
  65479=>"100000100",
  65480=>"100011000",
  65481=>"111101110",
  65482=>"011100011",
  65483=>"001110111",
  65484=>"100011011",
  65485=>"011000011",
  65486=>"110000110",
  65487=>"011100011",
  65488=>"000000110",
  65489=>"010000100",
  65490=>"100010001",
  65491=>"000001110",
  65492=>"001010111",
  65493=>"110010111",
  65494=>"110001100",
  65495=>"011010101",
  65496=>"010010001",
  65497=>"111101001",
  65498=>"101001101",
  65499=>"110110000",
  65500=>"100001000",
  65501=>"101101100",
  65502=>"111010011",
  65503=>"000110001",
  65504=>"100000100",
  65505=>"111100011",
  65506=>"001011011",
  65507=>"111110111",
  65508=>"011001001",
  65509=>"000010000",
  65510=>"000100111",
  65511=>"011111100",
  65512=>"001001000",
  65513=>"011010110",
  65514=>"100101101",
  65515=>"001110001",
  65516=>"011110100",
  65517=>"101010110",
  65518=>"001010001",
  65519=>"001011111",
  65520=>"000101001",
  65521=>"100010000",
  65522=>"000010011",
  65523=>"100100111",
  65524=>"010110100",
  65525=>"000111011",
  65526=>"010001001",
  65527=>"001011000",
  65528=>"000110001",
  65529=>"011111111",
  65530=>"100011010",
  65531=>"001010011",
  65532=>"110111101",
  65533=>"001010001",
  65534=>"101101101",
  65535=>"010001001");

BEGIN
  weight <= ROM_content(to_integer(address));
END RTL;