LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L8_4_WROM IS
  PORT (
    weight : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
    address : IN unsigned(weightsbitsAddress(8)-1 DOWNTO 0));
END L8_4_WROM;

ARCHITECTURE RTL OF L8_4_WROM IS

  TYPE ROM_mem IS ARRAY (0 TO 65535) OF STD_LOGIC_VECTOR(8 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem := (0=>"000100100",
  1=>"100110011",
  2=>"001101011",
  3=>"001010001",
  4=>"100100111",
  5=>"001111010",
  6=>"010100101",
  7=>"100000010",
  8=>"111111011",
  9=>"001001001",
  10=>"101110101",
  11=>"011110100",
  12=>"111010111",
  13=>"101011101",
  14=>"010100001",
  15=>"000101111",
  16=>"110000001",
  17=>"001111011",
  18=>"011011101",
  19=>"010111010",
  20=>"000001000",
  21=>"101111100",
  22=>"001111010",
  23=>"010010100",
  24=>"000111011",
  25=>"001000101",
  26=>"110110101",
  27=>"010000110",
  28=>"101001101",
  29=>"100111010",
  30=>"010010000",
  31=>"001010010",
  32=>"010001001",
  33=>"100001101",
  34=>"101010001",
  35=>"001000100",
  36=>"111011010",
  37=>"000000101",
  38=>"000100100",
  39=>"001110111",
  40=>"101111111",
  41=>"000110111",
  42=>"111010101",
  43=>"001010111",
  44=>"101110100",
  45=>"001100110",
  46=>"101011011",
  47=>"011011111",
  48=>"001110001",
  49=>"110011100",
  50=>"101010111",
  51=>"111011100",
  52=>"011111010",
  53=>"100010000",
  54=>"111100010",
  55=>"011110010",
  56=>"011010010",
  57=>"100000001",
  58=>"111010110",
  59=>"000101100",
  60=>"110110000",
  61=>"101010000",
  62=>"011100100",
  63=>"111011111",
  64=>"100010000",
  65=>"000000101",
  66=>"101011001",
  67=>"010011000",
  68=>"100111110",
  69=>"101101111",
  70=>"000000111",
  71=>"000110000",
  72=>"100101100",
  73=>"011000011",
  74=>"001011110",
  75=>"011110101",
  76=>"001000010",
  77=>"111000110",
  78=>"111111100",
  79=>"010100010",
  80=>"101001001",
  81=>"101111111",
  82=>"110110010",
  83=>"100111101",
  84=>"000010000",
  85=>"111001101",
  86=>"010110010",
  87=>"110011100",
  88=>"100100101",
  89=>"010101011",
  90=>"010111111",
  91=>"001100001",
  92=>"011001101",
  93=>"000110000",
  94=>"011000110",
  95=>"010000010",
  96=>"001100001",
  97=>"111111110",
  98=>"111011000",
  99=>"001011100",
  100=>"011110110",
  101=>"100101110",
  102=>"101110110",
  103=>"111011110",
  104=>"000001000",
  105=>"011101100",
  106=>"010011011",
  107=>"100011110",
  108=>"001011111",
  109=>"000101110",
  110=>"110010000",
  111=>"010101000",
  112=>"101101100",
  113=>"111001011",
  114=>"101011011",
  115=>"100100001",
  116=>"101011100",
  117=>"111010010",
  118=>"111100110",
  119=>"101101100",
  120=>"001110111",
  121=>"101101111",
  122=>"101000000",
  123=>"100010000",
  124=>"110110010",
  125=>"001001001",
  126=>"011000110",
  127=>"000001000",
  128=>"111000001",
  129=>"001011001",
  130=>"111101011",
  131=>"101011011",
  132=>"110001000",
  133=>"111110011",
  134=>"110110100",
  135=>"100011000",
  136=>"011101011",
  137=>"000000011",
  138=>"110000000",
  139=>"010011010",
  140=>"000110001",
  141=>"010010010",
  142=>"001110001",
  143=>"011010011",
  144=>"011110010",
  145=>"000010101",
  146=>"001000100",
  147=>"001111111",
  148=>"100000011",
  149=>"111100100",
  150=>"001000001",
  151=>"110011110",
  152=>"100101011",
  153=>"111111111",
  154=>"001011100",
  155=>"110011001",
  156=>"000011010",
  157=>"000100000",
  158=>"001101010",
  159=>"101110011",
  160=>"011110000",
  161=>"110001111",
  162=>"010010000",
  163=>"011010000",
  164=>"111101101",
  165=>"100000110",
  166=>"011000010",
  167=>"111100000",
  168=>"001111010",
  169=>"011111000",
  170=>"101110111",
  171=>"101101001",
  172=>"001010100",
  173=>"100110010",
  174=>"100100001",
  175=>"111111110",
  176=>"111011001",
  177=>"000111111",
  178=>"000100001",
  179=>"011100000",
  180=>"000001110",
  181=>"010111001",
  182=>"011000101",
  183=>"010000101",
  184=>"011100001",
  185=>"100001010",
  186=>"000010000",
  187=>"111111011",
  188=>"011000011",
  189=>"011000111",
  190=>"110000111",
  191=>"101000001",
  192=>"110111000",
  193=>"011011110",
  194=>"010010010",
  195=>"000101011",
  196=>"000111011",
  197=>"001011010",
  198=>"010111111",
  199=>"000001010",
  200=>"000000100",
  201=>"001110100",
  202=>"001011111",
  203=>"001101100",
  204=>"000111001",
  205=>"111100011",
  206=>"100111000",
  207=>"101101011",
  208=>"110000001",
  209=>"110001100",
  210=>"011001111",
  211=>"010110001",
  212=>"110001100",
  213=>"111110001",
  214=>"110101000",
  215=>"001001011",
  216=>"010000010",
  217=>"000000111",
  218=>"001000000",
  219=>"111011111",
  220=>"111100011",
  221=>"000100111",
  222=>"100001000",
  223=>"100100000",
  224=>"101011010",
  225=>"101100101",
  226=>"011001010",
  227=>"000110110",
  228=>"101100111",
  229=>"100000011",
  230=>"001011101",
  231=>"001010010",
  232=>"100000011",
  233=>"110110010",
  234=>"011111110",
  235=>"011000010",
  236=>"111110110",
  237=>"001000101",
  238=>"010111100",
  239=>"011111100",
  240=>"000010010",
  241=>"110000101",
  242=>"010110011",
  243=>"101101100",
  244=>"100010000",
  245=>"001011100",
  246=>"001011100",
  247=>"101001101",
  248=>"100110011",
  249=>"001110011",
  250=>"010011111",
  251=>"101000111",
  252=>"111100101",
  253=>"111101010",
  254=>"100001111",
  255=>"100101001",
  256=>"010010011",
  257=>"010101101",
  258=>"000100111",
  259=>"101111001",
  260=>"000010010",
  261=>"111010000",
  262=>"101010001",
  263=>"001000000",
  264=>"000110101",
  265=>"000101111",
  266=>"100001001",
  267=>"011101001",
  268=>"011000110",
  269=>"110000010",
  270=>"000111110",
  271=>"011001000",
  272=>"000111110",
  273=>"100100111",
  274=>"000110000",
  275=>"000010001",
  276=>"001000010",
  277=>"000111001",
  278=>"001110111",
  279=>"000011111",
  280=>"110001010",
  281=>"000101100",
  282=>"001001000",
  283=>"101101011",
  284=>"101000000",
  285=>"011111010",
  286=>"000001010",
  287=>"111111101",
  288=>"110011111",
  289=>"111111000",
  290=>"001011010",
  291=>"100111101",
  292=>"110100000",
  293=>"010111001",
  294=>"000000110",
  295=>"110100001",
  296=>"000011100",
  297=>"011111001",
  298=>"110010101",
  299=>"101010001",
  300=>"011100011",
  301=>"101001010",
  302=>"100001010",
  303=>"000001111",
  304=>"001101111",
  305=>"100011001",
  306=>"101001011",
  307=>"001001011",
  308=>"000111001",
  309=>"000000100",
  310=>"110100010",
  311=>"010001100",
  312=>"100001000",
  313=>"001010101",
  314=>"111000111",
  315=>"011100011",
  316=>"000001110",
  317=>"001011100",
  318=>"011110011",
  319=>"010101111",
  320=>"010000001",
  321=>"001001010",
  322=>"101000101",
  323=>"011010100",
  324=>"011111100",
  325=>"001110101",
  326=>"011000100",
  327=>"100000001",
  328=>"011001001",
  329=>"001101001",
  330=>"101111000",
  331=>"010010110",
  332=>"101101000",
  333=>"110011101",
  334=>"111100100",
  335=>"100000010",
  336=>"011000111",
  337=>"100001000",
  338=>"111110001",
  339=>"000110011",
  340=>"010000001",
  341=>"001101101",
  342=>"101000010",
  343=>"001111101",
  344=>"000001101",
  345=>"100010011",
  346=>"111101100",
  347=>"011101000",
  348=>"101101100",
  349=>"110100110",
  350=>"110110010",
  351=>"011110010",
  352=>"001100110",
  353=>"100111011",
  354=>"000110111",
  355=>"000101111",
  356=>"100010110",
  357=>"100011110",
  358=>"101111010",
  359=>"001011011",
  360=>"101111011",
  361=>"000100101",
  362=>"000001000",
  363=>"000001100",
  364=>"100011000",
  365=>"111001101",
  366=>"010101001",
  367=>"101001110",
  368=>"001111001",
  369=>"011001001",
  370=>"111101111",
  371=>"100001110",
  372=>"000000001",
  373=>"000001100",
  374=>"100100100",
  375=>"010100011",
  376=>"010001100",
  377=>"100011001",
  378=>"111111010",
  379=>"011101011",
  380=>"000000100",
  381=>"000011011",
  382=>"010010011",
  383=>"100101100",
  384=>"010001110",
  385=>"011011001",
  386=>"101011100",
  387=>"000100101",
  388=>"011111111",
  389=>"111101000",
  390=>"011011101",
  391=>"000110011",
  392=>"001001011",
  393=>"101001111",
  394=>"100000000",
  395=>"110010001",
  396=>"100101001",
  397=>"101000011",
  398=>"001000000",
  399=>"100010110",
  400=>"111001010",
  401=>"000011011",
  402=>"001110100",
  403=>"001111000",
  404=>"010101100",
  405=>"100110100",
  406=>"100101101",
  407=>"010111111",
  408=>"001100001",
  409=>"000000101",
  410=>"001011011",
  411=>"110001010",
  412=>"010000011",
  413=>"101010001",
  414=>"001110010",
  415=>"010001100",
  416=>"111000010",
  417=>"000000000",
  418=>"001001110",
  419=>"010100010",
  420=>"100010001",
  421=>"001100111",
  422=>"111100011",
  423=>"001101101",
  424=>"011101111",
  425=>"100111010",
  426=>"010000011",
  427=>"101000000",
  428=>"000101111",
  429=>"110101111",
  430=>"011110111",
  431=>"010000010",
  432=>"001101101",
  433=>"010100000",
  434=>"011010000",
  435=>"011110100",
  436=>"110000010",
  437=>"101110010",
  438=>"110101111",
  439=>"001001100",
  440=>"000100011",
  441=>"010100100",
  442=>"100001000",
  443=>"110010010",
  444=>"000010000",
  445=>"101001011",
  446=>"010011111",
  447=>"110001010",
  448=>"001010010",
  449=>"001111010",
  450=>"000100000",
  451=>"100010101",
  452=>"101010101",
  453=>"000101001",
  454=>"010100110",
  455=>"110111110",
  456=>"100001100",
  457=>"101000101",
  458=>"000010011",
  459=>"010010000",
  460=>"010000111",
  461=>"101101011",
  462=>"001100001",
  463=>"110111100",
  464=>"001000011",
  465=>"010101101",
  466=>"000000011",
  467=>"010010000",
  468=>"000000010",
  469=>"110110111",
  470=>"100100000",
  471=>"010100010",
  472=>"010101001",
  473=>"101101101",
  474=>"100010000",
  475=>"010111100",
  476=>"011111101",
  477=>"001100001",
  478=>"000110100",
  479=>"001111011",
  480=>"111100000",
  481=>"001110101",
  482=>"111100001",
  483=>"001000010",
  484=>"100101110",
  485=>"101011110",
  486=>"000001111",
  487=>"001111010",
  488=>"001110000",
  489=>"001001101",
  490=>"010000010",
  491=>"001011101",
  492=>"001000110",
  493=>"011101011",
  494=>"000100001",
  495=>"000000001",
  496=>"011100001",
  497=>"100100010",
  498=>"001010000",
  499=>"101100001",
  500=>"101000010",
  501=>"100010010",
  502=>"000100011",
  503=>"110011001",
  504=>"011111111",
  505=>"010001011",
  506=>"110100101",
  507=>"110011000",
  508=>"010100100",
  509=>"111011101",
  510=>"100111100",
  511=>"001101011",
  512=>"010111100",
  513=>"011001011",
  514=>"111011111",
  515=>"010000010",
  516=>"010111010",
  517=>"000100100",
  518=>"001011111",
  519=>"100000011",
  520=>"011000000",
  521=>"111111100",
  522=>"000110010",
  523=>"000000000",
  524=>"011100000",
  525=>"110110010",
  526=>"101000111",
  527=>"100011100",
  528=>"100111011",
  529=>"110101000",
  530=>"110011000",
  531=>"011011111",
  532=>"000010011",
  533=>"110010000",
  534=>"110010100",
  535=>"110000100",
  536=>"111001100",
  537=>"110010111",
  538=>"101111001",
  539=>"011100000",
  540=>"111010111",
  541=>"101101101",
  542=>"001111101",
  543=>"011101011",
  544=>"110100000",
  545=>"010011111",
  546=>"001011000",
  547=>"111001010",
  548=>"000101101",
  549=>"100111010",
  550=>"000001011",
  551=>"011111010",
  552=>"100101010",
  553=>"100001001",
  554=>"101110110",
  555=>"111111010",
  556=>"111001001",
  557=>"010110010",
  558=>"101001101",
  559=>"000101000",
  560=>"011001011",
  561=>"101110110",
  562=>"000100001",
  563=>"110001001",
  564=>"001110001",
  565=>"101101000",
  566=>"110000010",
  567=>"010001001",
  568=>"010000010",
  569=>"101110001",
  570=>"110110010",
  571=>"000111101",
  572=>"011101000",
  573=>"110000110",
  574=>"110110010",
  575=>"100111000",
  576=>"011101001",
  577=>"010001110",
  578=>"110011000",
  579=>"000100101",
  580=>"001110001",
  581=>"110010000",
  582=>"001111110",
  583=>"100000100",
  584=>"010110010",
  585=>"100111001",
  586=>"011011010",
  587=>"101111000",
  588=>"010001110",
  589=>"001101000",
  590=>"111010001",
  591=>"100011010",
  592=>"101100110",
  593=>"101111100",
  594=>"101100001",
  595=>"001011010",
  596=>"010100100",
  597=>"110111111",
  598=>"110110000",
  599=>"000000100",
  600=>"110100001",
  601=>"010100000",
  602=>"000100111",
  603=>"100001100",
  604=>"110010100",
  605=>"101111000",
  606=>"100100110",
  607=>"000111100",
  608=>"111110000",
  609=>"011000111",
  610=>"100010101",
  611=>"001100101",
  612=>"001010010",
  613=>"001100110",
  614=>"001111110",
  615=>"001101110",
  616=>"010101101",
  617=>"100101010",
  618=>"001110010",
  619=>"110001000",
  620=>"110110010",
  621=>"110001000",
  622=>"011111110",
  623=>"110101101",
  624=>"000001101",
  625=>"001111110",
  626=>"001101110",
  627=>"100001011",
  628=>"010101001",
  629=>"011001011",
  630=>"111110001",
  631=>"100010010",
  632=>"101010110",
  633=>"110101001",
  634=>"001100010",
  635=>"111000101",
  636=>"011000001",
  637=>"110010111",
  638=>"001000100",
  639=>"001100010",
  640=>"000010000",
  641=>"110110110",
  642=>"011110010",
  643=>"100001000",
  644=>"101001010",
  645=>"010110100",
  646=>"001110101",
  647=>"101010100",
  648=>"000011101",
  649=>"101100111",
  650=>"110110110",
  651=>"100001100",
  652=>"000111011",
  653=>"101101100",
  654=>"011001101",
  655=>"010000100",
  656=>"101110001",
  657=>"001000111",
  658=>"001111110",
  659=>"011001010",
  660=>"101001001",
  661=>"100001000",
  662=>"010101110",
  663=>"111100110",
  664=>"011001100",
  665=>"110110000",
  666=>"101110110",
  667=>"001001001",
  668=>"111000110",
  669=>"011011011",
  670=>"010110000",
  671=>"111100010",
  672=>"111111001",
  673=>"000101001",
  674=>"001101001",
  675=>"011001011",
  676=>"100001100",
  677=>"110011110",
  678=>"010001101",
  679=>"101000111",
  680=>"001110100",
  681=>"101000101",
  682=>"111010011",
  683=>"011000000",
  684=>"000000001",
  685=>"101011010",
  686=>"100100010",
  687=>"011001010",
  688=>"111111001",
  689=>"000100011",
  690=>"000100000",
  691=>"110000101",
  692=>"110001011",
  693=>"111101110",
  694=>"100000001",
  695=>"001010000",
  696=>"100111000",
  697=>"111010100",
  698=>"110011100",
  699=>"001101101",
  700=>"100101111",
  701=>"100010100",
  702=>"011000011",
  703=>"110111111",
  704=>"101101101",
  705=>"111011001",
  706=>"100001011",
  707=>"100111001",
  708=>"111111000",
  709=>"101000110",
  710=>"100000010",
  711=>"001111100",
  712=>"011100110",
  713=>"111101010",
  714=>"001101101",
  715=>"010100101",
  716=>"111000001",
  717=>"001011010",
  718=>"000000100",
  719=>"110110011",
  720=>"100000010",
  721=>"011011000",
  722=>"010100001",
  723=>"101010000",
  724=>"101101100",
  725=>"111000111",
  726=>"111110111",
  727=>"011010111",
  728=>"010000101",
  729=>"010011000",
  730=>"000111111",
  731=>"110101111",
  732=>"100010011",
  733=>"010100010",
  734=>"100001110",
  735=>"001000101",
  736=>"111101011",
  737=>"110101110",
  738=>"100101101",
  739=>"110110100",
  740=>"000111101",
  741=>"110001000",
  742=>"100100111",
  743=>"001000010",
  744=>"111110011",
  745=>"100000010",
  746=>"110010011",
  747=>"101100000",
  748=>"101110110",
  749=>"100011000",
  750=>"000111000",
  751=>"110110110",
  752=>"100001000",
  753=>"111010111",
  754=>"000111010",
  755=>"101101001",
  756=>"100001110",
  757=>"100110000",
  758=>"110010101",
  759=>"110001001",
  760=>"100001000",
  761=>"110010011",
  762=>"100111101",
  763=>"010001001",
  764=>"011111110",
  765=>"001100110",
  766=>"000011010",
  767=>"000110100",
  768=>"100100110",
  769=>"111110001",
  770=>"111110101",
  771=>"101010010",
  772=>"010011011",
  773=>"011001100",
  774=>"001110111",
  775=>"000000110",
  776=>"001010010",
  777=>"110010110",
  778=>"000111011",
  779=>"000011000",
  780=>"100101011",
  781=>"110011110",
  782=>"010001101",
  783=>"111101101",
  784=>"111000111",
  785=>"010100000",
  786=>"100101011",
  787=>"010011101",
  788=>"111101101",
  789=>"010001001",
  790=>"111111110",
  791=>"010010011",
  792=>"100101101",
  793=>"111011010",
  794=>"111000111",
  795=>"010110101",
  796=>"000011001",
  797=>"100001101",
  798=>"110000110",
  799=>"010101100",
  800=>"111011010",
  801=>"000100010",
  802=>"100111000",
  803=>"100010101",
  804=>"100101001",
  805=>"111101101",
  806=>"101001011",
  807=>"111010111",
  808=>"000011001",
  809=>"000101100",
  810=>"010010010",
  811=>"001011010",
  812=>"001101111",
  813=>"001111001",
  814=>"001110011",
  815=>"000100010",
  816=>"000011011",
  817=>"011000000",
  818=>"001111011",
  819=>"001111011",
  820=>"110100011",
  821=>"101100100",
  822=>"000000100",
  823=>"101101011",
  824=>"001001010",
  825=>"111011010",
  826=>"100101010",
  827=>"010100110",
  828=>"010001101",
  829=>"010110001",
  830=>"110010011",
  831=>"000011001",
  832=>"010000001",
  833=>"101101000",
  834=>"000110100",
  835=>"110001110",
  836=>"110110011",
  837=>"011100111",
  838=>"110111101",
  839=>"010110101",
  840=>"011010110",
  841=>"000101010",
  842=>"100010101",
  843=>"100111010",
  844=>"111110100",
  845=>"110001110",
  846=>"101111111",
  847=>"010101100",
  848=>"111110110",
  849=>"101100011",
  850=>"111110110",
  851=>"110110001",
  852=>"111100101",
  853=>"110111001",
  854=>"000010100",
  855=>"010000101",
  856=>"011010001",
  857=>"000101010",
  858=>"111111111",
  859=>"001101010",
  860=>"110111110",
  861=>"100111100",
  862=>"000001110",
  863=>"000011001",
  864=>"100010010",
  865=>"101011000",
  866=>"001010110",
  867=>"010111110",
  868=>"110011101",
  869=>"101111111",
  870=>"001010101",
  871=>"011110100",
  872=>"000011110",
  873=>"110001000",
  874=>"111110000",
  875=>"110100100",
  876=>"101011001",
  877=>"101000110",
  878=>"111001000",
  879=>"010011010",
  880=>"011110100",
  881=>"011101110",
  882=>"111000111",
  883=>"001100110",
  884=>"010100111",
  885=>"010100001",
  886=>"100111001",
  887=>"010000010",
  888=>"111101111",
  889=>"000111010",
  890=>"111000001",
  891=>"110111110",
  892=>"010100110",
  893=>"101110011",
  894=>"111001110",
  895=>"100100100",
  896=>"100010101",
  897=>"001100100",
  898=>"001010100",
  899=>"110111101",
  900=>"100101001",
  901=>"111101100",
  902=>"100010000",
  903=>"001101110",
  904=>"110100100",
  905=>"101101101",
  906=>"010110001",
  907=>"001000110",
  908=>"011111101",
  909=>"000010001",
  910=>"111110000",
  911=>"001100110",
  912=>"000001101",
  913=>"010010100",
  914=>"101000111",
  915=>"111111011",
  916=>"010100011",
  917=>"100111010",
  918=>"100011101",
  919=>"000011100",
  920=>"111001111",
  921=>"001111111",
  922=>"001111010",
  923=>"101110100",
  924=>"110110010",
  925=>"100001100",
  926=>"110000100",
  927=>"011011101",
  928=>"101100000",
  929=>"000011001",
  930=>"110000101",
  931=>"011101101",
  932=>"110010000",
  933=>"110111011",
  934=>"000010100",
  935=>"101110100",
  936=>"001000010",
  937=>"011010111",
  938=>"110100000",
  939=>"100001100",
  940=>"001010010",
  941=>"100111111",
  942=>"110011010",
  943=>"011100011",
  944=>"011001111",
  945=>"000100001",
  946=>"110110000",
  947=>"010001010",
  948=>"100000101",
  949=>"101101000",
  950=>"001101111",
  951=>"110001101",
  952=>"110011011",
  953=>"011110111",
  954=>"000101010",
  955=>"000000110",
  956=>"001101100",
  957=>"101010000",
  958=>"110110100",
  959=>"000000001",
  960=>"101010111",
  961=>"010101101",
  962=>"100000011",
  963=>"110000010",
  964=>"001011100",
  965=>"101101111",
  966=>"010011010",
  967=>"000000010",
  968=>"111111001",
  969=>"100100011",
  970=>"011001110",
  971=>"000110111",
  972=>"101000110",
  973=>"000100010",
  974=>"000110000",
  975=>"010000001",
  976=>"001100111",
  977=>"100010000",
  978=>"011010100",
  979=>"001101011",
  980=>"101000110",
  981=>"001000110",
  982=>"100010110",
  983=>"011010000",
  984=>"011001110",
  985=>"001000001",
  986=>"010000000",
  987=>"100110101",
  988=>"000001001",
  989=>"010101010",
  990=>"010001101",
  991=>"011101110",
  992=>"011000010",
  993=>"001011100",
  994=>"000100100",
  995=>"011101011",
  996=>"011000001",
  997=>"111100000",
  998=>"010000001",
  999=>"000010100",
  1000=>"010100101",
  1001=>"111011000",
  1002=>"100000001",
  1003=>"000110111",
  1004=>"000111001",
  1005=>"001000101",
  1006=>"110100111",
  1007=>"100110100",
  1008=>"110001111",
  1009=>"010101100",
  1010=>"011010011",
  1011=>"100010101",
  1012=>"100101100",
  1013=>"110000100",
  1014=>"011011101",
  1015=>"110110101",
  1016=>"101101101",
  1017=>"110100101",
  1018=>"110100111",
  1019=>"111100100",
  1020=>"010010010",
  1021=>"000011110",
  1022=>"100000011",
  1023=>"001001101",
  1024=>"110001011",
  1025=>"000111001",
  1026=>"001111101",
  1027=>"001101000",
  1028=>"011100010",
  1029=>"100101001",
  1030=>"010100110",
  1031=>"001101101",
  1032=>"100100000",
  1033=>"011001001",
  1034=>"110000100",
  1035=>"011100101",
  1036=>"011101101",
  1037=>"111011100",
  1038=>"011100011",
  1039=>"110001100",
  1040=>"101011011",
  1041=>"000100001",
  1042=>"111000100",
  1043=>"101111100",
  1044=>"111000111",
  1045=>"000111110",
  1046=>"101010011",
  1047=>"110100100",
  1048=>"001000000",
  1049=>"011011101",
  1050=>"101110010",
  1051=>"011111000",
  1052=>"100110011",
  1053=>"011111111",
  1054=>"110000100",
  1055=>"110101100",
  1056=>"100011010",
  1057=>"001010100",
  1058=>"111101010",
  1059=>"111011001",
  1060=>"110001101",
  1061=>"111000001",
  1062=>"111100001",
  1063=>"010101011",
  1064=>"100001100",
  1065=>"001100001",
  1066=>"010011010",
  1067=>"110101001",
  1068=>"000101011",
  1069=>"110001000",
  1070=>"101100001",
  1071=>"100100110",
  1072=>"100111111",
  1073=>"001010011",
  1074=>"101000111",
  1075=>"011101010",
  1076=>"001000010",
  1077=>"011110100",
  1078=>"110010111",
  1079=>"010010001",
  1080=>"000000001",
  1081=>"001111000",
  1082=>"011010100",
  1083=>"001101010",
  1084=>"111000100",
  1085=>"100111101",
  1086=>"011110111",
  1087=>"010000100",
  1088=>"011000110",
  1089=>"010000001",
  1090=>"011101101",
  1091=>"000101001",
  1092=>"111111110",
  1093=>"111110000",
  1094=>"101101011",
  1095=>"100110001",
  1096=>"011010110",
  1097=>"000010001",
  1098=>"011001001",
  1099=>"101111011",
  1100=>"010110000",
  1101=>"111110011",
  1102=>"000111100",
  1103=>"010101110",
  1104=>"011011100",
  1105=>"010001000",
  1106=>"011110111",
  1107=>"110010001",
  1108=>"101001011",
  1109=>"101000010",
  1110=>"000000010",
  1111=>"010010011",
  1112=>"110111111",
  1113=>"011100001",
  1114=>"010000101",
  1115=>"100000101",
  1116=>"111001101",
  1117=>"010100001",
  1118=>"000001111",
  1119=>"110111000",
  1120=>"101000000",
  1121=>"101001001",
  1122=>"110111101",
  1123=>"001111010",
  1124=>"100111100",
  1125=>"001001010",
  1126=>"010000000",
  1127=>"010000100",
  1128=>"010001001",
  1129=>"101100110",
  1130=>"011111000",
  1131=>"110100010",
  1132=>"111101000",
  1133=>"111011000",
  1134=>"100110010",
  1135=>"011111000",
  1136=>"010110110",
  1137=>"011110000",
  1138=>"011011010",
  1139=>"100100101",
  1140=>"001111000",
  1141=>"101010110",
  1142=>"001101000",
  1143=>"101001000",
  1144=>"101111110",
  1145=>"110100010",
  1146=>"001110000",
  1147=>"010100001",
  1148=>"011000101",
  1149=>"111111101",
  1150=>"000111101",
  1151=>"100101110",
  1152=>"000101010",
  1153=>"010111110",
  1154=>"000010011",
  1155=>"001000111",
  1156=>"111111101",
  1157=>"010000100",
  1158=>"011010100",
  1159=>"101010100",
  1160=>"110100111",
  1161=>"000111111",
  1162=>"111110111",
  1163=>"100001111",
  1164=>"000111100",
  1165=>"100011110",
  1166=>"010100101",
  1167=>"100101100",
  1168=>"111000010",
  1169=>"001110111",
  1170=>"000100011",
  1171=>"101001100",
  1172=>"000001110",
  1173=>"011110010",
  1174=>"111110011",
  1175=>"010110111",
  1176=>"111110110",
  1177=>"001111000",
  1178=>"110011111",
  1179=>"011110110",
  1180=>"010000010",
  1181=>"111001011",
  1182=>"001100001",
  1183=>"101100100",
  1184=>"001001101",
  1185=>"111111011",
  1186=>"011010100",
  1187=>"001010010",
  1188=>"101101010",
  1189=>"010100110",
  1190=>"101001111",
  1191=>"101010000",
  1192=>"101001000",
  1193=>"101101000",
  1194=>"111011101",
  1195=>"101100101",
  1196=>"110100110",
  1197=>"110101100",
  1198=>"110000001",
  1199=>"111011011",
  1200=>"100110010",
  1201=>"000110011",
  1202=>"100000010",
  1203=>"101111011",
  1204=>"010000000",
  1205=>"001110100",
  1206=>"000000110",
  1207=>"101001000",
  1208=>"111011101",
  1209=>"001100101",
  1210=>"001101011",
  1211=>"000100001",
  1212=>"000110100",
  1213=>"101111010",
  1214=>"101110110",
  1215=>"011111111",
  1216=>"111101010",
  1217=>"000011010",
  1218=>"011111001",
  1219=>"100011010",
  1220=>"000110110",
  1221=>"001100100",
  1222=>"001001111",
  1223=>"100111100",
  1224=>"101111100",
  1225=>"001011101",
  1226=>"111001110",
  1227=>"001001100",
  1228=>"111000110",
  1229=>"100111001",
  1230=>"011001111",
  1231=>"110011110",
  1232=>"010011001",
  1233=>"001100011",
  1234=>"011010001",
  1235=>"001000111",
  1236=>"111010010",
  1237=>"100100001",
  1238=>"110011010",
  1239=>"011000110",
  1240=>"110000101",
  1241=>"100011100",
  1242=>"000011011",
  1243=>"110100011",
  1244=>"011111101",
  1245=>"111101100",
  1246=>"010001010",
  1247=>"000001100",
  1248=>"101010000",
  1249=>"001100100",
  1250=>"110000001",
  1251=>"000010001",
  1252=>"100111101",
  1253=>"000110111",
  1254=>"001000011",
  1255=>"010001100",
  1256=>"110110000",
  1257=>"100011011",
  1258=>"001000011",
  1259=>"101001001",
  1260=>"100001100",
  1261=>"100110011",
  1262=>"100110000",
  1263=>"010111101",
  1264=>"011100111",
  1265=>"001100100",
  1266=>"000001110",
  1267=>"111010001",
  1268=>"101101101",
  1269=>"010011001",
  1270=>"001110011",
  1271=>"000000000",
  1272=>"110101111",
  1273=>"010110001",
  1274=>"101011100",
  1275=>"001000000",
  1276=>"111011111",
  1277=>"101010000",
  1278=>"110101011",
  1279=>"001101011",
  1280=>"000111100",
  1281=>"110110010",
  1282=>"111001011",
  1283=>"010011101",
  1284=>"011100001",
  1285=>"011111000",
  1286=>"001100001",
  1287=>"111000010",
  1288=>"100000010",
  1289=>"001000001",
  1290=>"001010101",
  1291=>"101011100",
  1292=>"011001000",
  1293=>"010100100",
  1294=>"101111001",
  1295=>"000000110",
  1296=>"111101001",
  1297=>"111111001",
  1298=>"000101111",
  1299=>"011001011",
  1300=>"010001100",
  1301=>"110101010",
  1302=>"011010100",
  1303=>"010000001",
  1304=>"000001011",
  1305=>"111001101",
  1306=>"110000010",
  1307=>"000011011",
  1308=>"000000100",
  1309=>"111011010",
  1310=>"111100001",
  1311=>"100011101",
  1312=>"010101001",
  1313=>"110100110",
  1314=>"101110001",
  1315=>"111111110",
  1316=>"111010101",
  1317=>"100011110",
  1318=>"110100010",
  1319=>"010000111",
  1320=>"100000100",
  1321=>"001100011",
  1322=>"111101001",
  1323=>"011011000",
  1324=>"101111111",
  1325=>"000110000",
  1326=>"101000000",
  1327=>"011001101",
  1328=>"010011100",
  1329=>"010100001",
  1330=>"101001111",
  1331=>"101011100",
  1332=>"110110111",
  1333=>"111010000",
  1334=>"100100010",
  1335=>"100010101",
  1336=>"110110110",
  1337=>"110011001",
  1338=>"101100010",
  1339=>"000000011",
  1340=>"111111110",
  1341=>"101111111",
  1342=>"001100010",
  1343=>"000010100",
  1344=>"000010110",
  1345=>"011100110",
  1346=>"010000101",
  1347=>"100011101",
  1348=>"010000000",
  1349=>"011111101",
  1350=>"100110000",
  1351=>"000101000",
  1352=>"010101001",
  1353=>"110010010",
  1354=>"110110011",
  1355=>"010000000",
  1356=>"001001010",
  1357=>"100101101",
  1358=>"100000111",
  1359=>"111100011",
  1360=>"111000010",
  1361=>"010101001",
  1362=>"110110101",
  1363=>"110111100",
  1364=>"000111010",
  1365=>"010110000",
  1366=>"111010110",
  1367=>"100110010",
  1368=>"011011111",
  1369=>"001001011",
  1370=>"000011110",
  1371=>"000000101",
  1372=>"101010011",
  1373=>"110000010",
  1374=>"100000000",
  1375=>"001010001",
  1376=>"000110011",
  1377=>"111101001",
  1378=>"000111111",
  1379=>"111001001",
  1380=>"100010111",
  1381=>"110101101",
  1382=>"110010001",
  1383=>"001111010",
  1384=>"011111101",
  1385=>"101010000",
  1386=>"110110000",
  1387=>"101010000",
  1388=>"000111010",
  1389=>"010001010",
  1390=>"110110101",
  1391=>"010010100",
  1392=>"000000101",
  1393=>"111000100",
  1394=>"111010000",
  1395=>"111001011",
  1396=>"111000111",
  1397=>"010101011",
  1398=>"100100100",
  1399=>"010001110",
  1400=>"011010011",
  1401=>"000011011",
  1402=>"001010000",
  1403=>"000011000",
  1404=>"100000101",
  1405=>"011111100",
  1406=>"001111100",
  1407=>"000101110",
  1408=>"100110001",
  1409=>"001000000",
  1410=>"110011011",
  1411=>"000000101",
  1412=>"100100111",
  1413=>"001001011",
  1414=>"110111100",
  1415=>"010010000",
  1416=>"000101111",
  1417=>"000100010",
  1418=>"100110001",
  1419=>"011011100",
  1420=>"100111100",
  1421=>"110111001",
  1422=>"011010110",
  1423=>"111001110",
  1424=>"011100101",
  1425=>"100011001",
  1426=>"000010000",
  1427=>"111110110",
  1428=>"111110110",
  1429=>"010100010",
  1430=>"011111110",
  1431=>"101001100",
  1432=>"000000000",
  1433=>"100010101",
  1434=>"000111101",
  1435=>"100000000",
  1436=>"011111011",
  1437=>"010010110",
  1438=>"110010011",
  1439=>"100000101",
  1440=>"101010100",
  1441=>"110101111",
  1442=>"010110111",
  1443=>"110101111",
  1444=>"101011000",
  1445=>"001111010",
  1446=>"110101111",
  1447=>"100000000",
  1448=>"011100110",
  1449=>"001111000",
  1450=>"100100010",
  1451=>"001010010",
  1452=>"100110000",
  1453=>"011000000",
  1454=>"100010100",
  1455=>"000111000",
  1456=>"111010001",
  1457=>"011100111",
  1458=>"011010110",
  1459=>"011110011",
  1460=>"101100101",
  1461=>"110011001",
  1462=>"010000100",
  1463=>"110110101",
  1464=>"000010100",
  1465=>"001010111",
  1466=>"011111110",
  1467=>"001111010",
  1468=>"000101000",
  1469=>"100011001",
  1470=>"000001010",
  1471=>"110001101",
  1472=>"000100110",
  1473=>"110111101",
  1474=>"000100101",
  1475=>"101000100",
  1476=>"101001111",
  1477=>"100111101",
  1478=>"001101000",
  1479=>"001111100",
  1480=>"001000001",
  1481=>"100001011",
  1482=>"000110010",
  1483=>"100111010",
  1484=>"000000111",
  1485=>"001111001",
  1486=>"000110101",
  1487=>"111100000",
  1488=>"111010111",
  1489=>"000100010",
  1490=>"000000100",
  1491=>"100010000",
  1492=>"010000100",
  1493=>"000000011",
  1494=>"001000101",
  1495=>"011011011",
  1496=>"000110001",
  1497=>"000111111",
  1498=>"110111110",
  1499=>"000011010",
  1500=>"110000111",
  1501=>"111000111",
  1502=>"011110111",
  1503=>"100001011",
  1504=>"101100011",
  1505=>"100101100",
  1506=>"110011101",
  1507=>"001000000",
  1508=>"001101011",
  1509=>"100010100",
  1510=>"110111000",
  1511=>"000111011",
  1512=>"011011101",
  1513=>"011000100",
  1514=>"100101100",
  1515=>"101111010",
  1516=>"010110000",
  1517=>"110010111",
  1518=>"011000011",
  1519=>"011000010",
  1520=>"101100101",
  1521=>"110010110",
  1522=>"110110100",
  1523=>"001010000",
  1524=>"101010100",
  1525=>"101001011",
  1526=>"001011010",
  1527=>"001101011",
  1528=>"001100000",
  1529=>"001110111",
  1530=>"001000000",
  1531=>"000111110",
  1532=>"100101100",
  1533=>"010111101",
  1534=>"100000000",
  1535=>"010010001",
  1536=>"001101011",
  1537=>"011000100",
  1538=>"011011000",
  1539=>"110010011",
  1540=>"010101110",
  1541=>"101001011",
  1542=>"101001011",
  1543=>"110001010",
  1544=>"011100111",
  1545=>"011011001",
  1546=>"110100111",
  1547=>"101110111",
  1548=>"000100010",
  1549=>"010011100",
  1550=>"001010101",
  1551=>"111110100",
  1552=>"111111010",
  1553=>"111011101",
  1554=>"111111000",
  1555=>"000000001",
  1556=>"101100101",
  1557=>"101011111",
  1558=>"010100010",
  1559=>"010000101",
  1560=>"001111111",
  1561=>"000100110",
  1562=>"000000000",
  1563=>"101001001",
  1564=>"011110000",
  1565=>"001101110",
  1566=>"101011000",
  1567=>"010111001",
  1568=>"000111000",
  1569=>"001011101",
  1570=>"100111010",
  1571=>"001111000",
  1572=>"101111111",
  1573=>"110101100",
  1574=>"110010111",
  1575=>"101110111",
  1576=>"011010000",
  1577=>"101011011",
  1578=>"000110110",
  1579=>"110111010",
  1580=>"001111110",
  1581=>"110011111",
  1582=>"010000101",
  1583=>"101101001",
  1584=>"110001001",
  1585=>"111111000",
  1586=>"000010001",
  1587=>"011110011",
  1588=>"010011011",
  1589=>"110100011",
  1590=>"110000001",
  1591=>"100110111",
  1592=>"110111100",
  1593=>"011001010",
  1594=>"010111000",
  1595=>"111010001",
  1596=>"011100101",
  1597=>"010001100",
  1598=>"000010001",
  1599=>"011001010",
  1600=>"000001010",
  1601=>"100011111",
  1602=>"111100001",
  1603=>"000011111",
  1604=>"011111110",
  1605=>"000100110",
  1606=>"001100110",
  1607=>"100110001",
  1608=>"001101100",
  1609=>"111011110",
  1610=>"111000001",
  1611=>"010110001",
  1612=>"001001001",
  1613=>"000001001",
  1614=>"000001100",
  1615=>"111101111",
  1616=>"010110100",
  1617=>"000000001",
  1618=>"011110100",
  1619=>"110001011",
  1620=>"110101101",
  1621=>"000100101",
  1622=>"010100110",
  1623=>"001010001",
  1624=>"000010110",
  1625=>"101101101",
  1626=>"011001010",
  1627=>"100001110",
  1628=>"100101011",
  1629=>"110110000",
  1630=>"100010101",
  1631=>"101101110",
  1632=>"001011010",
  1633=>"001101000",
  1634=>"011010111",
  1635=>"100111101",
  1636=>"010110010",
  1637=>"111001000",
  1638=>"101000110",
  1639=>"010111100",
  1640=>"010100000",
  1641=>"011000100",
  1642=>"011000010",
  1643=>"111000110",
  1644=>"001100011",
  1645=>"110110110",
  1646=>"001001011",
  1647=>"011100011",
  1648=>"100011101",
  1649=>"001101110",
  1650=>"011011011",
  1651=>"000111000",
  1652=>"011101100",
  1653=>"101110100",
  1654=>"101011001",
  1655=>"010110011",
  1656=>"001100010",
  1657=>"111101100",
  1658=>"111110111",
  1659=>"011101010",
  1660=>"101011001",
  1661=>"001111011",
  1662=>"100010000",
  1663=>"110000110",
  1664=>"001100100",
  1665=>"101010001",
  1666=>"001101000",
  1667=>"101010100",
  1668=>"001010111",
  1669=>"100010000",
  1670=>"011111110",
  1671=>"111111001",
  1672=>"001010011",
  1673=>"000010100",
  1674=>"001111011",
  1675=>"011001101",
  1676=>"100000001",
  1677=>"000010000",
  1678=>"111000000",
  1679=>"101100111",
  1680=>"010000110",
  1681=>"100000110",
  1682=>"011111100",
  1683=>"001001010",
  1684=>"100100011",
  1685=>"110111110",
  1686=>"000110010",
  1687=>"001110101",
  1688=>"111000000",
  1689=>"101010101",
  1690=>"010000010",
  1691=>"111100011",
  1692=>"010010001",
  1693=>"010100000",
  1694=>"010100001",
  1695=>"100011111",
  1696=>"101000111",
  1697=>"100111000",
  1698=>"000101010",
  1699=>"010110111",
  1700=>"000101110",
  1701=>"110001100",
  1702=>"001111110",
  1703=>"010111101",
  1704=>"111001101",
  1705=>"000011000",
  1706=>"100100001",
  1707=>"110011011",
  1708=>"101010100",
  1709=>"011001100",
  1710=>"001010001",
  1711=>"000001111",
  1712=>"000011001",
  1713=>"100100000",
  1714=>"010011101",
  1715=>"110001111",
  1716=>"011010000",
  1717=>"110001111",
  1718=>"011001010",
  1719=>"010100101",
  1720=>"110010010",
  1721=>"000011010",
  1722=>"000111101",
  1723=>"100000001",
  1724=>"000101011",
  1725=>"100001010",
  1726=>"111001100",
  1727=>"110101100",
  1728=>"100100100",
  1729=>"110101111",
  1730=>"100111100",
  1731=>"000001111",
  1732=>"100000000",
  1733=>"111111101",
  1734=>"100111011",
  1735=>"100101000",
  1736=>"010111001",
  1737=>"001010001",
  1738=>"111010000",
  1739=>"011010001",
  1740=>"000110111",
  1741=>"110111011",
  1742=>"001100010",
  1743=>"000001001",
  1744=>"101100011",
  1745=>"001101110",
  1746=>"111101011",
  1747=>"101010110",
  1748=>"011000111",
  1749=>"101100001",
  1750=>"000000110",
  1751=>"001111001",
  1752=>"010001100",
  1753=>"110100101",
  1754=>"000001000",
  1755=>"000010111",
  1756=>"100100110",
  1757=>"110110111",
  1758=>"001101000",
  1759=>"001110100",
  1760=>"101100001",
  1761=>"101010011",
  1762=>"111001010",
  1763=>"000001000",
  1764=>"000011001",
  1765=>"000100110",
  1766=>"011100010",
  1767=>"010001110",
  1768=>"111011100",
  1769=>"111100111",
  1770=>"101000001",
  1771=>"001100100",
  1772=>"110110000",
  1773=>"100111001",
  1774=>"110101101",
  1775=>"110100011",
  1776=>"100000110",
  1777=>"000000011",
  1778=>"001001011",
  1779=>"001010000",
  1780=>"011101001",
  1781=>"111010010",
  1782=>"000011110",
  1783=>"101011100",
  1784=>"101100000",
  1785=>"011110011",
  1786=>"111011010",
  1787=>"111000110",
  1788=>"101110110",
  1789=>"000110001",
  1790=>"101010110",
  1791=>"010001011",
  1792=>"101001001",
  1793=>"011000101",
  1794=>"101011000",
  1795=>"111100001",
  1796=>"010101100",
  1797=>"101111000",
  1798=>"101101101",
  1799=>"010010010",
  1800=>"001101011",
  1801=>"010111011",
  1802=>"100001110",
  1803=>"000010000",
  1804=>"111111100",
  1805=>"011000011",
  1806=>"010011100",
  1807=>"101000000",
  1808=>"110001011",
  1809=>"001100010",
  1810=>"100101000",
  1811=>"111111111",
  1812=>"111110011",
  1813=>"000000101",
  1814=>"111001111",
  1815=>"011010000",
  1816=>"000101010",
  1817=>"110011010",
  1818=>"110101111",
  1819=>"011100110",
  1820=>"001010101",
  1821=>"111100101",
  1822=>"111011001",
  1823=>"001111001",
  1824=>"111100101",
  1825=>"000000010",
  1826=>"010101110",
  1827=>"000000011",
  1828=>"110011101",
  1829=>"110110010",
  1830=>"000010101",
  1831=>"001110001",
  1832=>"111010100",
  1833=>"011010100",
  1834=>"000100000",
  1835=>"000110101",
  1836=>"100100110",
  1837=>"100100000",
  1838=>"001000100",
  1839=>"010011011",
  1840=>"111100000",
  1841=>"101001000",
  1842=>"111101101",
  1843=>"010011101",
  1844=>"101000100",
  1845=>"111101111",
  1846=>"000111111",
  1847=>"001000001",
  1848=>"000110010",
  1849=>"111111100",
  1850=>"111000010",
  1851=>"111001111",
  1852=>"000111011",
  1853=>"000100001",
  1854=>"110100010",
  1855=>"001011101",
  1856=>"010011001",
  1857=>"111010001",
  1858=>"000000011",
  1859=>"010111011",
  1860=>"000011001",
  1861=>"110001111",
  1862=>"101100000",
  1863=>"011110110",
  1864=>"110100110",
  1865=>"000000100",
  1866=>"000110100",
  1867=>"100011011",
  1868=>"001001100",
  1869=>"100111100",
  1870=>"011001001",
  1871=>"000001110",
  1872=>"101111011",
  1873=>"101110111",
  1874=>"101001000",
  1875=>"001010100",
  1876=>"111101000",
  1877=>"111000110",
  1878=>"101111101",
  1879=>"100111100",
  1880=>"010000001",
  1881=>"001111101",
  1882=>"111001101",
  1883=>"000111001",
  1884=>"111111011",
  1885=>"100011000",
  1886=>"111101101",
  1887=>"011000110",
  1888=>"011000001",
  1889=>"100001110",
  1890=>"100111101",
  1891=>"110010101",
  1892=>"001000000",
  1893=>"001000011",
  1894=>"001011111",
  1895=>"011011011",
  1896=>"001001001",
  1897=>"010001000",
  1898=>"110011111",
  1899=>"111101101",
  1900=>"110010110",
  1901=>"000011001",
  1902=>"011011101",
  1903=>"000011111",
  1904=>"100111110",
  1905=>"101111010",
  1906=>"010100011",
  1907=>"111000011",
  1908=>"111001100",
  1909=>"000011010",
  1910=>"111100010",
  1911=>"010011010",
  1912=>"111010111",
  1913=>"011000010",
  1914=>"000110100",
  1915=>"100111101",
  1916=>"110100000",
  1917=>"111001010",
  1918=>"000001001",
  1919=>"011101000",
  1920=>"011011111",
  1921=>"101000110",
  1922=>"000101100",
  1923=>"111100101",
  1924=>"101011011",
  1925=>"000010111",
  1926=>"100001111",
  1927=>"110101010",
  1928=>"110001110",
  1929=>"111110110",
  1930=>"000001110",
  1931=>"011011011",
  1932=>"111010101",
  1933=>"101110110",
  1934=>"100110111",
  1935=>"001000001",
  1936=>"100110011",
  1937=>"011110111",
  1938=>"001100000",
  1939=>"101101011",
  1940=>"001010101",
  1941=>"000001000",
  1942=>"010111111",
  1943=>"011000101",
  1944=>"010110011",
  1945=>"110100001",
  1946=>"011001111",
  1947=>"000101100",
  1948=>"011011011",
  1949=>"111001000",
  1950=>"101000111",
  1951=>"011001110",
  1952=>"101011001",
  1953=>"011011001",
  1954=>"011111100",
  1955=>"011101111",
  1956=>"111011001",
  1957=>"001011111",
  1958=>"101110011",
  1959=>"001110100",
  1960=>"100001000",
  1961=>"101011101",
  1962=>"010010110",
  1963=>"100000111",
  1964=>"011110111",
  1965=>"010110010",
  1966=>"101100100",
  1967=>"001100101",
  1968=>"111100001",
  1969=>"000010001",
  1970=>"011101110",
  1971=>"111110100",
  1972=>"110010011",
  1973=>"110000010",
  1974=>"000101001",
  1975=>"010101010",
  1976=>"010010010",
  1977=>"100101001",
  1978=>"000111100",
  1979=>"001110001",
  1980=>"011101000",
  1981=>"110110100",
  1982=>"101110010",
  1983=>"100010001",
  1984=>"110001010",
  1985=>"110100000",
  1986=>"010001111",
  1987=>"111110111",
  1988=>"000010001",
  1989=>"010111100",
  1990=>"100010011",
  1991=>"101111010",
  1992=>"100100000",
  1993=>"101011001",
  1994=>"010010100",
  1995=>"110110001",
  1996=>"001101011",
  1997=>"101010010",
  1998=>"110101111",
  1999=>"101010001",
  2000=>"011101110",
  2001=>"011000001",
  2002=>"010111100",
  2003=>"001000101",
  2004=>"110111110",
  2005=>"000010011",
  2006=>"110111111",
  2007=>"110001000",
  2008=>"010111100",
  2009=>"000001010",
  2010=>"111111111",
  2011=>"100100000",
  2012=>"101000010",
  2013=>"110001100",
  2014=>"101001100",
  2015=>"000000100",
  2016=>"011010011",
  2017=>"000010011",
  2018=>"010011110",
  2019=>"111010001",
  2020=>"110100000",
  2021=>"110001111",
  2022=>"000000110",
  2023=>"000100010",
  2024=>"111010011",
  2025=>"001110011",
  2026=>"011111010",
  2027=>"000011100",
  2028=>"010111110",
  2029=>"100011101",
  2030=>"101101110",
  2031=>"110110010",
  2032=>"001100101",
  2033=>"100110011",
  2034=>"000000100",
  2035=>"100011011",
  2036=>"001100110",
  2037=>"010001000",
  2038=>"100100100",
  2039=>"001100101",
  2040=>"000011010",
  2041=>"001001011",
  2042=>"110000100",
  2043=>"001110111",
  2044=>"100000110",
  2045=>"101000101",
  2046=>"100001010",
  2047=>"010011110",
  2048=>"011101011",
  2049=>"110100010",
  2050=>"110000101",
  2051=>"101000110",
  2052=>"100101110",
  2053=>"101001100",
  2054=>"111111111",
  2055=>"001101101",
  2056=>"111101101",
  2057=>"100111000",
  2058=>"101000000",
  2059=>"010011111",
  2060=>"111100101",
  2061=>"100001000",
  2062=>"010110111",
  2063=>"011000100",
  2064=>"100111000",
  2065=>"001001101",
  2066=>"110100101",
  2067=>"101000100",
  2068=>"110010101",
  2069=>"011011111",
  2070=>"100101111",
  2071=>"101100101",
  2072=>"010101011",
  2073=>"000100110",
  2074=>"001100111",
  2075=>"111111100",
  2076=>"111110000",
  2077=>"000111001",
  2078=>"111010000",
  2079=>"001101010",
  2080=>"100001110",
  2081=>"000000011",
  2082=>"000111010",
  2083=>"101000100",
  2084=>"110001011",
  2085=>"111001110",
  2086=>"101110100",
  2087=>"110010111",
  2088=>"001111001",
  2089=>"001011111",
  2090=>"011100001",
  2091=>"111111010",
  2092=>"101101001",
  2093=>"110110001",
  2094=>"101111011",
  2095=>"110010100",
  2096=>"001110101",
  2097=>"000101111",
  2098=>"001111100",
  2099=>"011010001",
  2100=>"001001011",
  2101=>"101011001",
  2102=>"001011110",
  2103=>"111000110",
  2104=>"010011000",
  2105=>"100001010",
  2106=>"100000010",
  2107=>"001000110",
  2108=>"010001000",
  2109=>"000111110",
  2110=>"111011100",
  2111=>"000110000",
  2112=>"110100111",
  2113=>"001000000",
  2114=>"001011101",
  2115=>"011011001",
  2116=>"000010100",
  2117=>"001000111",
  2118=>"110011010",
  2119=>"101111011",
  2120=>"110111010",
  2121=>"010011011",
  2122=>"110001100",
  2123=>"101000100",
  2124=>"010101111",
  2125=>"110011110",
  2126=>"010011000",
  2127=>"111010011",
  2128=>"011100101",
  2129=>"010010100",
  2130=>"101100100",
  2131=>"001001111",
  2132=>"001010100",
  2133=>"010101001",
  2134=>"111101100",
  2135=>"001111101",
  2136=>"001101100",
  2137=>"000000111",
  2138=>"110100100",
  2139=>"011001010",
  2140=>"110001111",
  2141=>"001001101",
  2142=>"111101001",
  2143=>"011000111",
  2144=>"110000101",
  2145=>"011011111",
  2146=>"010000101",
  2147=>"001010000",
  2148=>"111111101",
  2149=>"001001010",
  2150=>"010011101",
  2151=>"111001111",
  2152=>"010110111",
  2153=>"001010001",
  2154=>"000101100",
  2155=>"010001111",
  2156=>"001111000",
  2157=>"101000000",
  2158=>"101111101",
  2159=>"111011110",
  2160=>"101110001",
  2161=>"010101100",
  2162=>"010001101",
  2163=>"100100101",
  2164=>"010011010",
  2165=>"110110100",
  2166=>"111001010",
  2167=>"000000010",
  2168=>"010001000",
  2169=>"101011111",
  2170=>"100110101",
  2171=>"000110101",
  2172=>"111001001",
  2173=>"000011011",
  2174=>"101010111",
  2175=>"111001010",
  2176=>"100001000",
  2177=>"100000110",
  2178=>"111101111",
  2179=>"010000000",
  2180=>"000000101",
  2181=>"101100111",
  2182=>"000001111",
  2183=>"111101011",
  2184=>"111011110",
  2185=>"101000010",
  2186=>"001101000",
  2187=>"111000001",
  2188=>"010000001",
  2189=>"000111000",
  2190=>"010001011",
  2191=>"011010011",
  2192=>"100101011",
  2193=>"000011010",
  2194=>"100111001",
  2195=>"111100101",
  2196=>"100001000",
  2197=>"010111110",
  2198=>"000001100",
  2199=>"000011101",
  2200=>"110001000",
  2201=>"010001110",
  2202=>"100110000",
  2203=>"110100011",
  2204=>"110010101",
  2205=>"010101100",
  2206=>"111000111",
  2207=>"110010101",
  2208=>"010101010",
  2209=>"111000110",
  2210=>"000101011",
  2211=>"001011001",
  2212=>"001011001",
  2213=>"010010011",
  2214=>"010111110",
  2215=>"000000010",
  2216=>"110010100",
  2217=>"001011111",
  2218=>"000000001",
  2219=>"111110000",
  2220=>"000001110",
  2221=>"110010101",
  2222=>"110001101",
  2223=>"001000110",
  2224=>"000100110",
  2225=>"000101111",
  2226=>"101110101",
  2227=>"110001010",
  2228=>"111010010",
  2229=>"011110101",
  2230=>"010011010",
  2231=>"101001100",
  2232=>"101111000",
  2233=>"001000110",
  2234=>"110010011",
  2235=>"100000000",
  2236=>"101100011",
  2237=>"100011011",
  2238=>"110011000",
  2239=>"100101101",
  2240=>"101001101",
  2241=>"001000000",
  2242=>"101111001",
  2243=>"001010101",
  2244=>"011000110",
  2245=>"001000011",
  2246=>"100100110",
  2247=>"001011000",
  2248=>"001010100",
  2249=>"100101101",
  2250=>"001111001",
  2251=>"111000001",
  2252=>"011111100",
  2253=>"010000111",
  2254=>"001011101",
  2255=>"000101000",
  2256=>"101000101",
  2257=>"000010110",
  2258=>"000011000",
  2259=>"010100011",
  2260=>"110000100",
  2261=>"010001100",
  2262=>"011001110",
  2263=>"000101111",
  2264=>"110001100",
  2265=>"100011100",
  2266=>"111100011",
  2267=>"111110100",
  2268=>"100010010",
  2269=>"010000110",
  2270=>"100000011",
  2271=>"110000101",
  2272=>"110011000",
  2273=>"010110100",
  2274=>"101100111",
  2275=>"101000100",
  2276=>"111001110",
  2277=>"000011110",
  2278=>"000101001",
  2279=>"110011110",
  2280=>"011001100",
  2281=>"100010111",
  2282=>"011011011",
  2283=>"001010011",
  2284=>"000101101",
  2285=>"101000000",
  2286=>"001110000",
  2287=>"111101010",
  2288=>"011101110",
  2289=>"011011111",
  2290=>"011010100",
  2291=>"000100000",
  2292=>"010001001",
  2293=>"100011111",
  2294=>"000011101",
  2295=>"110010001",
  2296=>"001011000",
  2297=>"111110000",
  2298=>"100111101",
  2299=>"001001001",
  2300=>"111011001",
  2301=>"011000100",
  2302=>"110111011",
  2303=>"010111111",
  2304=>"010101110",
  2305=>"100100010",
  2306=>"010011010",
  2307=>"011111111",
  2308=>"100101101",
  2309=>"000011110",
  2310=>"011010000",
  2311=>"100100101",
  2312=>"110011000",
  2313=>"111011000",
  2314=>"010111110",
  2315=>"010110101",
  2316=>"000110110",
  2317=>"010011011",
  2318=>"011011011",
  2319=>"001001011",
  2320=>"111101000",
  2321=>"110101111",
  2322=>"111100101",
  2323=>"111010111",
  2324=>"011111001",
  2325=>"110011000",
  2326=>"111011110",
  2327=>"011100110",
  2328=>"010010011",
  2329=>"010000111",
  2330=>"010000010",
  2331=>"110100001",
  2332=>"011010011",
  2333=>"111000000",
  2334=>"011110010",
  2335=>"011100001",
  2336=>"010110100",
  2337=>"101111000",
  2338=>"111110010",
  2339=>"010000101",
  2340=>"011110100",
  2341=>"001010111",
  2342=>"100011110",
  2343=>"100101111",
  2344=>"101101001",
  2345=>"101101011",
  2346=>"000111110",
  2347=>"100000110",
  2348=>"101100011",
  2349=>"111101001",
  2350=>"100001011",
  2351=>"101100100",
  2352=>"100001010",
  2353=>"011011101",
  2354=>"000001110",
  2355=>"100001011",
  2356=>"110000100",
  2357=>"000001001",
  2358=>"001010011",
  2359=>"100010000",
  2360=>"101011110",
  2361=>"011100000",
  2362=>"100000100",
  2363=>"111011010",
  2364=>"101101000",
  2365=>"111000110",
  2366=>"001111001",
  2367=>"100110011",
  2368=>"001001010",
  2369=>"001101111",
  2370=>"011011001",
  2371=>"100011010",
  2372=>"001011110",
  2373=>"101011010",
  2374=>"101110001",
  2375=>"011011010",
  2376=>"111100010",
  2377=>"110010100",
  2378=>"111010110",
  2379=>"000001110",
  2380=>"001010101",
  2381=>"110111000",
  2382=>"001010010",
  2383=>"010110000",
  2384=>"110000001",
  2385=>"000010001",
  2386=>"111101111",
  2387=>"111101011",
  2388=>"001001001",
  2389=>"001011011",
  2390=>"100001000",
  2391=>"101101011",
  2392=>"011100111",
  2393=>"010011011",
  2394=>"001011100",
  2395=>"110101110",
  2396=>"111101001",
  2397=>"111010000",
  2398=>"001011101",
  2399=>"011000101",
  2400=>"100101111",
  2401=>"110110100",
  2402=>"111100110",
  2403=>"111001001",
  2404=>"010001011",
  2405=>"101110111",
  2406=>"001010111",
  2407=>"111111110",
  2408=>"100111000",
  2409=>"011001101",
  2410=>"110000100",
  2411=>"101111101",
  2412=>"001001000",
  2413=>"011110001",
  2414=>"001000001",
  2415=>"011100110",
  2416=>"110100010",
  2417=>"110010100",
  2418=>"111011111",
  2419=>"010000100",
  2420=>"000100011",
  2421=>"001101101",
  2422=>"000110010",
  2423=>"011100011",
  2424=>"010001100",
  2425=>"000111000",
  2426=>"010100111",
  2427=>"000100001",
  2428=>"001010111",
  2429=>"000111110",
  2430=>"100110100",
  2431=>"101101110",
  2432=>"100111011",
  2433=>"001011110",
  2434=>"011101101",
  2435=>"010111011",
  2436=>"110011111",
  2437=>"101110001",
  2438=>"001111000",
  2439=>"111000011",
  2440=>"011011110",
  2441=>"101100111",
  2442=>"000011001",
  2443=>"001000000",
  2444=>"001001000",
  2445=>"110000110",
  2446=>"010001111",
  2447=>"110010111",
  2448=>"101101001",
  2449=>"011010100",
  2450=>"011111001",
  2451=>"010110110",
  2452=>"110101001",
  2453=>"100001101",
  2454=>"001011011",
  2455=>"010000000",
  2456=>"011010010",
  2457=>"011101111",
  2458=>"101001111",
  2459=>"011110110",
  2460=>"110001110",
  2461=>"110000101",
  2462=>"101100001",
  2463=>"101011101",
  2464=>"111101100",
  2465=>"011000101",
  2466=>"110110100",
  2467=>"000000101",
  2468=>"111111011",
  2469=>"110001101",
  2470=>"001010100",
  2471=>"111101110",
  2472=>"001010000",
  2473=>"011111101",
  2474=>"011011010",
  2475=>"101110111",
  2476=>"011011111",
  2477=>"001001111",
  2478=>"110100100",
  2479=>"101101000",
  2480=>"000100101",
  2481=>"100111000",
  2482=>"101011000",
  2483=>"111011010",
  2484=>"111001000",
  2485=>"101111001",
  2486=>"000011111",
  2487=>"000100010",
  2488=>"111101111",
  2489=>"101101110",
  2490=>"011101000",
  2491=>"000100100",
  2492=>"000111010",
  2493=>"000101001",
  2494=>"111101000",
  2495=>"111111011",
  2496=>"100000000",
  2497=>"101101111",
  2498=>"101110100",
  2499=>"010001101",
  2500=>"011010110",
  2501=>"011001100",
  2502=>"011000000",
  2503=>"001000000",
  2504=>"100011010",
  2505=>"000010100",
  2506=>"101011101",
  2507=>"010110011",
  2508=>"000001101",
  2509=>"111010111",
  2510=>"000010111",
  2511=>"010010000",
  2512=>"011111110",
  2513=>"100111001",
  2514=>"011110010",
  2515=>"000100111",
  2516=>"001101111",
  2517=>"101100000",
  2518=>"001111011",
  2519=>"001011100",
  2520=>"100010011",
  2521=>"111100111",
  2522=>"010101000",
  2523=>"111111100",
  2524=>"000101101",
  2525=>"101001111",
  2526=>"111101010",
  2527=>"100010110",
  2528=>"010011101",
  2529=>"001010110",
  2530=>"111010100",
  2531=>"001011110",
  2532=>"100110010",
  2533=>"011111110",
  2534=>"010111000",
  2535=>"010000100",
  2536=>"010001100",
  2537=>"000010110",
  2538=>"000000001",
  2539=>"001000101",
  2540=>"000010110",
  2541=>"111001000",
  2542=>"101001001",
  2543=>"110100100",
  2544=>"010011011",
  2545=>"011001100",
  2546=>"010010000",
  2547=>"000000010",
  2548=>"100101011",
  2549=>"000000101",
  2550=>"110001100",
  2551=>"010110001",
  2552=>"001000100",
  2553=>"110110010",
  2554=>"001100111",
  2555=>"001110001",
  2556=>"111111011",
  2557=>"010100110",
  2558=>"110110110",
  2559=>"111000001",
  2560=>"011110010",
  2561=>"000011010",
  2562=>"101001110",
  2563=>"101100010",
  2564=>"011001101",
  2565=>"010101111",
  2566=>"000010001",
  2567=>"110010000",
  2568=>"111100000",
  2569=>"111011111",
  2570=>"110001110",
  2571=>"110010101",
  2572=>"101000010",
  2573=>"001110100",
  2574=>"000100001",
  2575=>"110010010",
  2576=>"001101001",
  2577=>"100010100",
  2578=>"111111001",
  2579=>"001010011",
  2580=>"010100000",
  2581=>"010100001",
  2582=>"001110111",
  2583=>"101101000",
  2584=>"100100001",
  2585=>"001010001",
  2586=>"011101101",
  2587=>"001101001",
  2588=>"111001000",
  2589=>"011010100",
  2590=>"101010011",
  2591=>"101011111",
  2592=>"000001010",
  2593=>"101010110",
  2594=>"010010001",
  2595=>"001101100",
  2596=>"011110111",
  2597=>"111011001",
  2598=>"000000010",
  2599=>"001010100",
  2600=>"101000000",
  2601=>"111111111",
  2602=>"000001001",
  2603=>"100100100",
  2604=>"001001111",
  2605=>"101000100",
  2606=>"101000111",
  2607=>"000001010",
  2608=>"000101110",
  2609=>"111001111",
  2610=>"110011100",
  2611=>"111110111",
  2612=>"111100011",
  2613=>"011100011",
  2614=>"010001110",
  2615=>"111000101",
  2616=>"110100000",
  2617=>"111010010",
  2618=>"010001000",
  2619=>"000111011",
  2620=>"101111101",
  2621=>"110110010",
  2622=>"111100001",
  2623=>"000101100",
  2624=>"011100001",
  2625=>"110100100",
  2626=>"011011100",
  2627=>"000101000",
  2628=>"011101000",
  2629=>"100001111",
  2630=>"001000110",
  2631=>"101100001",
  2632=>"011111110",
  2633=>"101000011",
  2634=>"011111010",
  2635=>"011101000",
  2636=>"010010000",
  2637=>"000000001",
  2638=>"110010011",
  2639=>"001111100",
  2640=>"000111000",
  2641=>"101001011",
  2642=>"010001110",
  2643=>"000001101",
  2644=>"111001100",
  2645=>"100000100",
  2646=>"000101000",
  2647=>"101110010",
  2648=>"011010101",
  2649=>"110000000",
  2650=>"001010100",
  2651=>"000000011",
  2652=>"101001110",
  2653=>"100000100",
  2654=>"001110110",
  2655=>"001100110",
  2656=>"011011010",
  2657=>"111011110",
  2658=>"010010110",
  2659=>"111001000",
  2660=>"010001001",
  2661=>"000000011",
  2662=>"110000010",
  2663=>"010010110",
  2664=>"011011010",
  2665=>"101010111",
  2666=>"110010111",
  2667=>"101001111",
  2668=>"101111110",
  2669=>"100000101",
  2670=>"101111000",
  2671=>"101110110",
  2672=>"000110100",
  2673=>"001011001",
  2674=>"101001111",
  2675=>"010001001",
  2676=>"111001101",
  2677=>"111011010",
  2678=>"001110011",
  2679=>"101001001",
  2680=>"101000001",
  2681=>"011011111",
  2682=>"000111001",
  2683=>"001000110",
  2684=>"111001101",
  2685=>"111000110",
  2686=>"010101101",
  2687=>"010010000",
  2688=>"100000111",
  2689=>"110111110",
  2690=>"110110101",
  2691=>"000000111",
  2692=>"010101101",
  2693=>"101100010",
  2694=>"010001010",
  2695=>"111011111",
  2696=>"111110010",
  2697=>"110011110",
  2698=>"001000010",
  2699=>"100011000",
  2700=>"111000101",
  2701=>"111101111",
  2702=>"110001010",
  2703=>"111000110",
  2704=>"111000100",
  2705=>"111110010",
  2706=>"110011010",
  2707=>"001110101",
  2708=>"000110010",
  2709=>"001101001",
  2710=>"010011111",
  2711=>"001001101",
  2712=>"101011011",
  2713=>"110011111",
  2714=>"010100110",
  2715=>"001001101",
  2716=>"100001111",
  2717=>"000110001",
  2718=>"000001111",
  2719=>"111100010",
  2720=>"110111111",
  2721=>"010001111",
  2722=>"000110111",
  2723=>"110010100",
  2724=>"111101101",
  2725=>"010111011",
  2726=>"101000010",
  2727=>"000001011",
  2728=>"111011101",
  2729=>"101100001",
  2730=>"101110001",
  2731=>"110000001",
  2732=>"010100010",
  2733=>"011101000",
  2734=>"000010100",
  2735=>"111011111",
  2736=>"000100101",
  2737=>"101001101",
  2738=>"010000010",
  2739=>"111000111",
  2740=>"011100010",
  2741=>"011010001",
  2742=>"111110001",
  2743=>"100101010",
  2744=>"000111010",
  2745=>"010000100",
  2746=>"010111101",
  2747=>"011110111",
  2748=>"000010111",
  2749=>"111111010",
  2750=>"101110000",
  2751=>"110000001",
  2752=>"011110111",
  2753=>"011000000",
  2754=>"010000000",
  2755=>"101001000",
  2756=>"011001100",
  2757=>"000010111",
  2758=>"100010100",
  2759=>"000110110",
  2760=>"001001100",
  2761=>"011011010",
  2762=>"010100101",
  2763=>"110001111",
  2764=>"010010110",
  2765=>"000101100",
  2766=>"010000100",
  2767=>"011000110",
  2768=>"101111100",
  2769=>"101010101",
  2770=>"111101100",
  2771=>"011010110",
  2772=>"110010110",
  2773=>"000100100",
  2774=>"111011101",
  2775=>"011010100",
  2776=>"000111001",
  2777=>"001101101",
  2778=>"001101001",
  2779=>"001010111",
  2780=>"010100110",
  2781=>"110000011",
  2782=>"110001011",
  2783=>"010110111",
  2784=>"010101101",
  2785=>"001001000",
  2786=>"010011111",
  2787=>"010001011",
  2788=>"010000100",
  2789=>"111101001",
  2790=>"000100000",
  2791=>"110111011",
  2792=>"000001100",
  2793=>"110111000",
  2794=>"000001000",
  2795=>"000011110",
  2796=>"010001010",
  2797=>"101111110",
  2798=>"100001011",
  2799=>"010001111",
  2800=>"111111111",
  2801=>"011101000",
  2802=>"011101101",
  2803=>"111001001",
  2804=>"111100001",
  2805=>"000000010",
  2806=>"111110000",
  2807=>"001000111",
  2808=>"101000111",
  2809=>"111010100",
  2810=>"111111110",
  2811=>"010000101",
  2812=>"011010110",
  2813=>"010001111",
  2814=>"100110101",
  2815=>"100100001",
  2816=>"101100001",
  2817=>"100011001",
  2818=>"011011010",
  2819=>"010000001",
  2820=>"110001000",
  2821=>"001100000",
  2822=>"011000100",
  2823=>"101100101",
  2824=>"111110101",
  2825=>"011100101",
  2826=>"001011011",
  2827=>"101011010",
  2828=>"001110110",
  2829=>"111010000",
  2830=>"100001001",
  2831=>"111111011",
  2832=>"111100111",
  2833=>"000010000",
  2834=>"100011001",
  2835=>"011100101",
  2836=>"111101100",
  2837=>"010101010",
  2838=>"011010111",
  2839=>"000000110",
  2840=>"010110010",
  2841=>"100011111",
  2842=>"000000100",
  2843=>"010000100",
  2844=>"101000000",
  2845=>"000001111",
  2846=>"111011001",
  2847=>"111110110",
  2848=>"000001010",
  2849=>"010100100",
  2850=>"000000001",
  2851=>"111001000",
  2852=>"000000101",
  2853=>"111100000",
  2854=>"010000101",
  2855=>"100010001",
  2856=>"101011011",
  2857=>"100001110",
  2858=>"110111010",
  2859=>"000000110",
  2860=>"000101100",
  2861=>"001100100",
  2862=>"000101001",
  2863=>"101100110",
  2864=>"000101101",
  2865=>"011001000",
  2866=>"010011100",
  2867=>"101010100",
  2868=>"010110001",
  2869=>"010010110",
  2870=>"101100001",
  2871=>"100101111",
  2872=>"111110010",
  2873=>"000000001",
  2874=>"011000110",
  2875=>"010011000",
  2876=>"111111000",
  2877=>"000101100",
  2878=>"110001000",
  2879=>"010011000",
  2880=>"111100001",
  2881=>"010111100",
  2882=>"111010011",
  2883=>"100001101",
  2884=>"000000011",
  2885=>"110001101",
  2886=>"000001011",
  2887=>"001001000",
  2888=>"000001101",
  2889=>"000101010",
  2890=>"011000110",
  2891=>"001001100",
  2892=>"110100111",
  2893=>"110100010",
  2894=>"000111001",
  2895=>"000000110",
  2896=>"010100011",
  2897=>"110001000",
  2898=>"010000011",
  2899=>"001000010",
  2900=>"111101010",
  2901=>"101111100",
  2902=>"010101000",
  2903=>"000110001",
  2904=>"000001011",
  2905=>"001000101",
  2906=>"100111110",
  2907=>"111010100",
  2908=>"010011111",
  2909=>"011100000",
  2910=>"101000011",
  2911=>"010001010",
  2912=>"110010010",
  2913=>"000000100",
  2914=>"111010011",
  2915=>"100010110",
  2916=>"100000111",
  2917=>"111100001",
  2918=>"001101100",
  2919=>"001000000",
  2920=>"111000000",
  2921=>"000101001",
  2922=>"100000100",
  2923=>"111010110",
  2924=>"000000100",
  2925=>"110000100",
  2926=>"001101100",
  2927=>"101000111",
  2928=>"111100111",
  2929=>"010110110",
  2930=>"000000011",
  2931=>"000010011",
  2932=>"000010011",
  2933=>"111100000",
  2934=>"100110010",
  2935=>"001001010",
  2936=>"101010011",
  2937=>"000111011",
  2938=>"011101100",
  2939=>"010101011",
  2940=>"110000010",
  2941=>"001101000",
  2942=>"100010000",
  2943=>"111100110",
  2944=>"000000011",
  2945=>"000001000",
  2946=>"010011001",
  2947=>"010110100",
  2948=>"010001010",
  2949=>"111100010",
  2950=>"000110000",
  2951=>"100001110",
  2952=>"111111010",
  2953=>"110110011",
  2954=>"000010001",
  2955=>"101110101",
  2956=>"111100111",
  2957=>"101101110",
  2958=>"101111000",
  2959=>"011001011",
  2960=>"111011100",
  2961=>"111111000",
  2962=>"000100001",
  2963=>"111100011",
  2964=>"001011110",
  2965=>"110101001",
  2966=>"010010100",
  2967=>"111100101",
  2968=>"000110111",
  2969=>"011001100",
  2970=>"100101110",
  2971=>"100101001",
  2972=>"110000110",
  2973=>"111000100",
  2974=>"001010111",
  2975=>"111100001",
  2976=>"000100110",
  2977=>"000100110",
  2978=>"010110111",
  2979=>"001010110",
  2980=>"000000111",
  2981=>"011110010",
  2982=>"000001101",
  2983=>"100101101",
  2984=>"000110010",
  2985=>"111000001",
  2986=>"001101111",
  2987=>"100000000",
  2988=>"101101011",
  2989=>"010000101",
  2990=>"010100011",
  2991=>"111100100",
  2992=>"110000100",
  2993=>"010100100",
  2994=>"001110101",
  2995=>"000011100",
  2996=>"010011111",
  2997=>"001000101",
  2998=>"010001110",
  2999=>"010011101",
  3000=>"100000101",
  3001=>"100011110",
  3002=>"001100011",
  3003=>"010100011",
  3004=>"110110110",
  3005=>"010001011",
  3006=>"011010110",
  3007=>"110100110",
  3008=>"000011010",
  3009=>"110101001",
  3010=>"011111011",
  3011=>"001101100",
  3012=>"100011000",
  3013=>"001101110",
  3014=>"000010100",
  3015=>"101101100",
  3016=>"101000100",
  3017=>"010001000",
  3018=>"101101101",
  3019=>"001111000",
  3020=>"110010111",
  3021=>"011000110",
  3022=>"010000000",
  3023=>"010000101",
  3024=>"110101011",
  3025=>"011101111",
  3026=>"010111101",
  3027=>"010110000",
  3028=>"011011101",
  3029=>"110111101",
  3030=>"000000101",
  3031=>"110011010",
  3032=>"111000111",
  3033=>"010011000",
  3034=>"111010010",
  3035=>"100011110",
  3036=>"101101111",
  3037=>"101111111",
  3038=>"011101010",
  3039=>"100000001",
  3040=>"111001010",
  3041=>"111011110",
  3042=>"111110011",
  3043=>"111001011",
  3044=>"111010100",
  3045=>"011100100",
  3046=>"001110001",
  3047=>"000000001",
  3048=>"011100111",
  3049=>"010111010",
  3050=>"101101111",
  3051=>"111101011",
  3052=>"100111100",
  3053=>"000111010",
  3054=>"111111100",
  3055=>"111101111",
  3056=>"000000010",
  3057=>"101001010",
  3058=>"100111011",
  3059=>"001100101",
  3060=>"111101101",
  3061=>"000001110",
  3062=>"000001101",
  3063=>"011110010",
  3064=>"101000110",
  3065=>"110101001",
  3066=>"111001110",
  3067=>"011111000",
  3068=>"001011001",
  3069=>"100101000",
  3070=>"111000011",
  3071=>"110000101",
  3072=>"000001000",
  3073=>"011010101",
  3074=>"000000000",
  3075=>"111101111",
  3076=>"111000100",
  3077=>"101011110",
  3078=>"100010001",
  3079=>"101001000",
  3080=>"111011001",
  3081=>"001001011",
  3082=>"010100110",
  3083=>"111110001",
  3084=>"000111111",
  3085=>"110001000",
  3086=>"111100000",
  3087=>"101000101",
  3088=>"000010001",
  3089=>"000000111",
  3090=>"100010101",
  3091=>"000111110",
  3092=>"010111001",
  3093=>"101010011",
  3094=>"110111100",
  3095=>"001000110",
  3096=>"001001110",
  3097=>"100110000",
  3098=>"101111001",
  3099=>"111101001",
  3100=>"011111001",
  3101=>"110111000",
  3102=>"000100010",
  3103=>"111000000",
  3104=>"001111000",
  3105=>"101111101",
  3106=>"001010101",
  3107=>"011110110",
  3108=>"011011000",
  3109=>"010011001",
  3110=>"000001000",
  3111=>"011011010",
  3112=>"111000100",
  3113=>"111001000",
  3114=>"000110100",
  3115=>"001100000",
  3116=>"010101111",
  3117=>"000010001",
  3118=>"101110100",
  3119=>"110000000",
  3120=>"111110111",
  3121=>"000000000",
  3122=>"011000111",
  3123=>"111111110",
  3124=>"101111111",
  3125=>"001111000",
  3126=>"001011100",
  3127=>"110110011",
  3128=>"100001001",
  3129=>"110000010",
  3130=>"100011110",
  3131=>"110010000",
  3132=>"001000000",
  3133=>"000000110",
  3134=>"110101000",
  3135=>"011100000",
  3136=>"001110011",
  3137=>"000001010",
  3138=>"001100011",
  3139=>"011101100",
  3140=>"100011011",
  3141=>"011111010",
  3142=>"010100110",
  3143=>"011111101",
  3144=>"111101100",
  3145=>"110111010",
  3146=>"000001100",
  3147=>"100010011",
  3148=>"001011011",
  3149=>"101011011",
  3150=>"100010101",
  3151=>"101110010",
  3152=>"000000001",
  3153=>"000001001",
  3154=>"010011101",
  3155=>"001001001",
  3156=>"011000100",
  3157=>"000001111",
  3158=>"000100011",
  3159=>"110100100",
  3160=>"100110111",
  3161=>"101111100",
  3162=>"111010001",
  3163=>"000110011",
  3164=>"101110101",
  3165=>"101100101",
  3166=>"000100101",
  3167=>"100010000",
  3168=>"010111110",
  3169=>"011011010",
  3170=>"100001011",
  3171=>"000011100",
  3172=>"101101100",
  3173=>"110100111",
  3174=>"011101110",
  3175=>"010101101",
  3176=>"010100100",
  3177=>"010011110",
  3178=>"000001010",
  3179=>"010010100",
  3180=>"001110010",
  3181=>"010100101",
  3182=>"111100110",
  3183=>"011111000",
  3184=>"100001011",
  3185=>"110101111",
  3186=>"111100010",
  3187=>"001101000",
  3188=>"111111111",
  3189=>"001011111",
  3190=>"001101111",
  3191=>"100110100",
  3192=>"010010110",
  3193=>"011000110",
  3194=>"010000100",
  3195=>"000001000",
  3196=>"100000010",
  3197=>"011001000",
  3198=>"101101011",
  3199=>"110000001",
  3200=>"011010101",
  3201=>"111100000",
  3202=>"001001000",
  3203=>"100101111",
  3204=>"101000000",
  3205=>"010011011",
  3206=>"000100101",
  3207=>"000010010",
  3208=>"101000011",
  3209=>"011101000",
  3210=>"101111000",
  3211=>"110110100",
  3212=>"111110111",
  3213=>"011110100",
  3214=>"011010011",
  3215=>"111101100",
  3216=>"001110110",
  3217=>"000011110",
  3218=>"000011101",
  3219=>"011100000",
  3220=>"000001101",
  3221=>"011111100",
  3222=>"001011001",
  3223=>"011011001",
  3224=>"110111001",
  3225=>"101011100",
  3226=>"001011111",
  3227=>"100110101",
  3228=>"000000010",
  3229=>"000011011",
  3230=>"110000110",
  3231=>"101110010",
  3232=>"100001010",
  3233=>"100011101",
  3234=>"001101001",
  3235=>"000110110",
  3236=>"000100110",
  3237=>"000011101",
  3238=>"111111101",
  3239=>"101001000",
  3240=>"111100000",
  3241=>"110001110",
  3242=>"111110010",
  3243=>"001011001",
  3244=>"110101100",
  3245=>"100001110",
  3246=>"000100010",
  3247=>"000101001",
  3248=>"000011011",
  3249=>"111011011",
  3250=>"001001100",
  3251=>"100100100",
  3252=>"010011111",
  3253=>"000000101",
  3254=>"101110011",
  3255=>"110100001",
  3256=>"011111011",
  3257=>"110100100",
  3258=>"100000000",
  3259=>"101000000",
  3260=>"110011100",
  3261=>"010101010",
  3262=>"000011111",
  3263=>"100111100",
  3264=>"111100011",
  3265=>"001001011",
  3266=>"100101010",
  3267=>"111100000",
  3268=>"111111011",
  3269=>"000111001",
  3270=>"111010100",
  3271=>"011000101",
  3272=>"001101000",
  3273=>"101010110",
  3274=>"001110011",
  3275=>"011110011",
  3276=>"111000111",
  3277=>"011000111",
  3278=>"011100110",
  3279=>"111010101",
  3280=>"001000110",
  3281=>"000100000",
  3282=>"111100000",
  3283=>"111101000",
  3284=>"001100000",
  3285=>"011100010",
  3286=>"000100011",
  3287=>"001010101",
  3288=>"010011101",
  3289=>"001010011",
  3290=>"010001101",
  3291=>"000001010",
  3292=>"111010010",
  3293=>"111111011",
  3294=>"110000000",
  3295=>"000111110",
  3296=>"001000001",
  3297=>"001111111",
  3298=>"101000010",
  3299=>"011011011",
  3300=>"000011011",
  3301=>"100001010",
  3302=>"001100000",
  3303=>"000110000",
  3304=>"001101000",
  3305=>"001101111",
  3306=>"010001101",
  3307=>"111111110",
  3308=>"100100100",
  3309=>"110110100",
  3310=>"110011111",
  3311=>"101111011",
  3312=>"111100011",
  3313=>"011001111",
  3314=>"001010001",
  3315=>"011100000",
  3316=>"000111110",
  3317=>"101101111",
  3318=>"111100001",
  3319=>"000100101",
  3320=>"101011110",
  3321=>"110100000",
  3322=>"000011000",
  3323=>"000101101",
  3324=>"101100011",
  3325=>"001110000",
  3326=>"001010100",
  3327=>"101001000",
  3328=>"101010110",
  3329=>"000001100",
  3330=>"101011110",
  3331=>"101111111",
  3332=>"110010001",
  3333=>"010010101",
  3334=>"000010100",
  3335=>"110011011",
  3336=>"101001001",
  3337=>"010000110",
  3338=>"001111101",
  3339=>"001011001",
  3340=>"000010010",
  3341=>"000110000",
  3342=>"100111001",
  3343=>"011111011",
  3344=>"000101111",
  3345=>"001111100",
  3346=>"010010110",
  3347=>"100010001",
  3348=>"110001011",
  3349=>"001001001",
  3350=>"101101100",
  3351=>"100101110",
  3352=>"101100110",
  3353=>"101011101",
  3354=>"111110101",
  3355=>"101101000",
  3356=>"101111000",
  3357=>"000110101",
  3358=>"010010101",
  3359=>"111111101",
  3360=>"000111010",
  3361=>"000010110",
  3362=>"011011000",
  3363=>"101010110",
  3364=>"001110000",
  3365=>"100000111",
  3366=>"000111010",
  3367=>"000100010",
  3368=>"101000001",
  3369=>"010000010",
  3370=>"111110110",
  3371=>"000000001",
  3372=>"101011001",
  3373=>"110000111",
  3374=>"001110100",
  3375=>"110001101",
  3376=>"001001001",
  3377=>"101110001",
  3378=>"001011111",
  3379=>"011110110",
  3380=>"011000000",
  3381=>"000011101",
  3382=>"011101010",
  3383=>"110100111",
  3384=>"011000100",
  3385=>"110010011",
  3386=>"110100100",
  3387=>"000101111",
  3388=>"111111010",
  3389=>"001111010",
  3390=>"010110001",
  3391=>"011100001",
  3392=>"001001001",
  3393=>"011000100",
  3394=>"100100001",
  3395=>"111110101",
  3396=>"010010100",
  3397=>"011001101",
  3398=>"001100100",
  3399=>"110101101",
  3400=>"101010111",
  3401=>"111000111",
  3402=>"011010000",
  3403=>"001000001",
  3404=>"111001011",
  3405=>"001011100",
  3406=>"011101111",
  3407=>"101011010",
  3408=>"111100011",
  3409=>"100011000",
  3410=>"010110101",
  3411=>"111011101",
  3412=>"011011000",
  3413=>"010001011",
  3414=>"111011111",
  3415=>"110011100",
  3416=>"101011101",
  3417=>"001011000",
  3418=>"011000010",
  3419=>"011100101",
  3420=>"001000000",
  3421=>"011110001",
  3422=>"111000001",
  3423=>"000001001",
  3424=>"011110001",
  3425=>"110110010",
  3426=>"010000000",
  3427=>"011100010",
  3428=>"000011100",
  3429=>"100010100",
  3430=>"111110000",
  3431=>"010000110",
  3432=>"100000000",
  3433=>"110001100",
  3434=>"000101010",
  3435=>"111100000",
  3436=>"011101110",
  3437=>"000110001",
  3438=>"111100010",
  3439=>"110011000",
  3440=>"000011010",
  3441=>"111110011",
  3442=>"100000011",
  3443=>"010110100",
  3444=>"100101101",
  3445=>"010100011",
  3446=>"110000000",
  3447=>"110101001",
  3448=>"101010011",
  3449=>"110000100",
  3450=>"100011110",
  3451=>"010011101",
  3452=>"110011111",
  3453=>"100000110",
  3454=>"010000110",
  3455=>"100001101",
  3456=>"100111100",
  3457=>"111001111",
  3458=>"110101101",
  3459=>"110000011",
  3460=>"111101111",
  3461=>"010100001",
  3462=>"111010011",
  3463=>"001010010",
  3464=>"101101100",
  3465=>"110000111",
  3466=>"000011111",
  3467=>"100000011",
  3468=>"101010101",
  3469=>"010001101",
  3470=>"001111001",
  3471=>"100001101",
  3472=>"000010100",
  3473=>"111101101",
  3474=>"111001100",
  3475=>"100001111",
  3476=>"011101010",
  3477=>"111000010",
  3478=>"000001010",
  3479=>"001110111",
  3480=>"011011100",
  3481=>"001100000",
  3482=>"011100011",
  3483=>"100010000",
  3484=>"011001100",
  3485=>"011001001",
  3486=>"111010110",
  3487=>"000101000",
  3488=>"100100010",
  3489=>"101000011",
  3490=>"100111111",
  3491=>"100111001",
  3492=>"010100011",
  3493=>"011100000",
  3494=>"101011100",
  3495=>"111111010",
  3496=>"111101010",
  3497=>"000110100",
  3498=>"001110110",
  3499=>"010100010",
  3500=>"100010000",
  3501=>"111101001",
  3502=>"110001000",
  3503=>"000100001",
  3504=>"111001011",
  3505=>"001101110",
  3506=>"010101100",
  3507=>"000101110",
  3508=>"010010011",
  3509=>"101010101",
  3510=>"001000101",
  3511=>"111011010",
  3512=>"011110011",
  3513=>"110000010",
  3514=>"011011111",
  3515=>"111010001",
  3516=>"011100111",
  3517=>"010100101",
  3518=>"010011101",
  3519=>"100100000",
  3520=>"110100110",
  3521=>"000100010",
  3522=>"000100011",
  3523=>"001101001",
  3524=>"000101000",
  3525=>"000100000",
  3526=>"100011111",
  3527=>"110111001",
  3528=>"001100100",
  3529=>"100010111",
  3530=>"010010010",
  3531=>"101100110",
  3532=>"100111100",
  3533=>"000001111",
  3534=>"000001011",
  3535=>"000011100",
  3536=>"001111001",
  3537=>"100100010",
  3538=>"110111110",
  3539=>"001111011",
  3540=>"111111010",
  3541=>"001111111",
  3542=>"001000001",
  3543=>"000101010",
  3544=>"010001010",
  3545=>"111001110",
  3546=>"011101010",
  3547=>"001001110",
  3548=>"101111001",
  3549=>"100001111",
  3550=>"100101010",
  3551=>"010000000",
  3552=>"101101001",
  3553=>"101001100",
  3554=>"110100111",
  3555=>"001010010",
  3556=>"101001010",
  3557=>"011100101",
  3558=>"000000110",
  3559=>"010000000",
  3560=>"101000101",
  3561=>"001111011",
  3562=>"001111101",
  3563=>"000011010",
  3564=>"110010101",
  3565=>"101100011",
  3566=>"011011101",
  3567=>"111100011",
  3568=>"100100010",
  3569=>"001000010",
  3570=>"110111000",
  3571=>"011000101",
  3572=>"110101101",
  3573=>"011010101",
  3574=>"100101110",
  3575=>"001001101",
  3576=>"010011100",
  3577=>"001111010",
  3578=>"111000000",
  3579=>"110010110",
  3580=>"110011111",
  3581=>"000000010",
  3582=>"010000011",
  3583=>"101111000",
  3584=>"010000100",
  3585=>"000011001",
  3586=>"111001001",
  3587=>"111111001",
  3588=>"101100111",
  3589=>"101111001",
  3590=>"000000011",
  3591=>"100100001",
  3592=>"000110001",
  3593=>"010011011",
  3594=>"111011010",
  3595=>"111011111",
  3596=>"000000011",
  3597=>"111101110",
  3598=>"111110100",
  3599=>"101000011",
  3600=>"101001111",
  3601=>"000000000",
  3602=>"110000101",
  3603=>"001010000",
  3604=>"111100101",
  3605=>"011000111",
  3606=>"000101101",
  3607=>"000101011",
  3608=>"110000101",
  3609=>"010101010",
  3610=>"011011000",
  3611=>"011101011",
  3612=>"010110010",
  3613=>"111001001",
  3614=>"000000001",
  3615=>"110100110",
  3616=>"111011011",
  3617=>"001000001",
  3618=>"000101011",
  3619=>"111111011",
  3620=>"000000001",
  3621=>"010001101",
  3622=>"111111000",
  3623=>"010100101",
  3624=>"010100010",
  3625=>"000011001",
  3626=>"010111101",
  3627=>"010111111",
  3628=>"011001111",
  3629=>"100011011",
  3630=>"100111100",
  3631=>"000001110",
  3632=>"100110111",
  3633=>"001010000",
  3634=>"000111100",
  3635=>"100010010",
  3636=>"101111011",
  3637=>"100101010",
  3638=>"100000000",
  3639=>"011011001",
  3640=>"010100000",
  3641=>"101000000",
  3642=>"001111101",
  3643=>"000100101",
  3644=>"111110110",
  3645=>"011000101",
  3646=>"010010011",
  3647=>"100111010",
  3648=>"000101000",
  3649=>"101110110",
  3650=>"000100110",
  3651=>"100010011",
  3652=>"001110001",
  3653=>"101001100",
  3654=>"110010011",
  3655=>"110010000",
  3656=>"001000100",
  3657=>"110100111",
  3658=>"000111001",
  3659=>"101010111",
  3660=>"110000101",
  3661=>"110010110",
  3662=>"101001001",
  3663=>"011010011",
  3664=>"011001110",
  3665=>"000010000",
  3666=>"000110100",
  3667=>"111100001",
  3668=>"011100011",
  3669=>"111110010",
  3670=>"111110110",
  3671=>"010110111",
  3672=>"101110111",
  3673=>"101010110",
  3674=>"111111011",
  3675=>"000100000",
  3676=>"011011011",
  3677=>"000110011",
  3678=>"100100101",
  3679=>"000010001",
  3680=>"000001101",
  3681=>"100100100",
  3682=>"100101110",
  3683=>"000101110",
  3684=>"000001110",
  3685=>"101000001",
  3686=>"101001101",
  3687=>"110001101",
  3688=>"110011110",
  3689=>"001101110",
  3690=>"100011001",
  3691=>"110000110",
  3692=>"100100001",
  3693=>"000011101",
  3694=>"101101110",
  3695=>"011010001",
  3696=>"001001011",
  3697=>"001000011",
  3698=>"001001000",
  3699=>"010101100",
  3700=>"111110110",
  3701=>"001100111",
  3702=>"010001101",
  3703=>"111111101",
  3704=>"010101011",
  3705=>"110010000",
  3706=>"101110110",
  3707=>"110000110",
  3708=>"010010101",
  3709=>"010110011",
  3710=>"110101001",
  3711=>"001100000",
  3712=>"000011011",
  3713=>"010000000",
  3714=>"101111010",
  3715=>"101111101",
  3716=>"110100101",
  3717=>"100000000",
  3718=>"010111000",
  3719=>"001001111",
  3720=>"111110111",
  3721=>"011001000",
  3722=>"011000010",
  3723=>"111110001",
  3724=>"001010010",
  3725=>"001100011",
  3726=>"010101010",
  3727=>"111111011",
  3728=>"110111010",
  3729=>"100111100",
  3730=>"010111000",
  3731=>"010111011",
  3732=>"000000110",
  3733=>"000110010",
  3734=>"000101101",
  3735=>"010110010",
  3736=>"110010010",
  3737=>"001110101",
  3738=>"110001100",
  3739=>"110011011",
  3740=>"110101110",
  3741=>"110010101",
  3742=>"010001111",
  3743=>"010111101",
  3744=>"011111010",
  3745=>"100110001",
  3746=>"101000001",
  3747=>"110100000",
  3748=>"011101100",
  3749=>"001110001",
  3750=>"111101101",
  3751=>"101110001",
  3752=>"101101011",
  3753=>"101011111",
  3754=>"001010011",
  3755=>"000000000",
  3756=>"000110000",
  3757=>"110000100",
  3758=>"101100100",
  3759=>"101000100",
  3760=>"010111111",
  3761=>"000111011",
  3762=>"000100001",
  3763=>"110101110",
  3764=>"111110101",
  3765=>"001111110",
  3766=>"001011101",
  3767=>"010101011",
  3768=>"101010011",
  3769=>"000010110",
  3770=>"000010111",
  3771=>"010101110",
  3772=>"111010101",
  3773=>"111100001",
  3774=>"010101000",
  3775=>"011111010",
  3776=>"110000011",
  3777=>"111001101",
  3778=>"000111000",
  3779=>"100001110",
  3780=>"101111101",
  3781=>"010001000",
  3782=>"101110101",
  3783=>"110000000",
  3784=>"110000110",
  3785=>"010000111",
  3786=>"011111000",
  3787=>"111100011",
  3788=>"000000001",
  3789=>"101100011",
  3790=>"000111000",
  3791=>"101100010",
  3792=>"101011100",
  3793=>"000000011",
  3794=>"101111100",
  3795=>"001110111",
  3796=>"011110111",
  3797=>"111111011",
  3798=>"001000000",
  3799=>"011100110",
  3800=>"001001110",
  3801=>"101000001",
  3802=>"010011011",
  3803=>"111110111",
  3804=>"110000000",
  3805=>"000010000",
  3806=>"000011111",
  3807=>"111101101",
  3808=>"001010111",
  3809=>"001000101",
  3810=>"101100010",
  3811=>"000101000",
  3812=>"110001011",
  3813=>"000011111",
  3814=>"101000011",
  3815=>"101011111",
  3816=>"100111000",
  3817=>"100110101",
  3818=>"000001110",
  3819=>"000101111",
  3820=>"000011111",
  3821=>"000111110",
  3822=>"001101011",
  3823=>"101011000",
  3824=>"000111000",
  3825=>"001000000",
  3826=>"000011110",
  3827=>"111011000",
  3828=>"011001010",
  3829=>"010110000",
  3830=>"110001011",
  3831=>"100010000",
  3832=>"111011101",
  3833=>"100000111",
  3834=>"000101011",
  3835=>"001000001",
  3836=>"010111011",
  3837=>"001110011",
  3838=>"010100101",
  3839=>"101111011",
  3840=>"100111000",
  3841=>"010111001",
  3842=>"000101101",
  3843=>"100001000",
  3844=>"000111110",
  3845=>"101001111",
  3846=>"001000000",
  3847=>"010001010",
  3848=>"111000100",
  3849=>"100111000",
  3850=>"000100000",
  3851=>"101000001",
  3852=>"000110100",
  3853=>"100111110",
  3854=>"010011000",
  3855=>"001010001",
  3856=>"111110100",
  3857=>"000100100",
  3858=>"100111100",
  3859=>"100000011",
  3860=>"100010011",
  3861=>"110100100",
  3862=>"000011100",
  3863=>"111110110",
  3864=>"101101111",
  3865=>"111001110",
  3866=>"111101010",
  3867=>"111010000",
  3868=>"111110011",
  3869=>"111001100",
  3870=>"000001000",
  3871=>"111010100",
  3872=>"101101001",
  3873=>"100000000",
  3874=>"001110011",
  3875=>"000000101",
  3876=>"000100100",
  3877=>"010101110",
  3878=>"000110101",
  3879=>"011010000",
  3880=>"010110010",
  3881=>"001100000",
  3882=>"011000000",
  3883=>"001010101",
  3884=>"101111110",
  3885=>"100000011",
  3886=>"010110000",
  3887=>"011101111",
  3888=>"111100111",
  3889=>"010000000",
  3890=>"011101100",
  3891=>"100011010",
  3892=>"011111111",
  3893=>"110111011",
  3894=>"000000010",
  3895=>"110110111",
  3896=>"100111011",
  3897=>"011010101",
  3898=>"010101100",
  3899=>"100100000",
  3900=>"001100000",
  3901=>"111011110",
  3902=>"000000101",
  3903=>"001000101",
  3904=>"010111001",
  3905=>"010011001",
  3906=>"110011010",
  3907=>"011101110",
  3908=>"100001100",
  3909=>"011010010",
  3910=>"110100000",
  3911=>"110110001",
  3912=>"010110111",
  3913=>"101111011",
  3914=>"001011010",
  3915=>"100001011",
  3916=>"001011111",
  3917=>"011111111",
  3918=>"001111110",
  3919=>"101000000",
  3920=>"100101101",
  3921=>"011001110",
  3922=>"110000011",
  3923=>"010110110",
  3924=>"001110011",
  3925=>"111010010",
  3926=>"111101100",
  3927=>"110001100",
  3928=>"110011111",
  3929=>"011111000",
  3930=>"110010001",
  3931=>"100101111",
  3932=>"110111010",
  3933=>"110110101",
  3934=>"011111000",
  3935=>"000100010",
  3936=>"111001010",
  3937=>"111011010",
  3938=>"001110010",
  3939=>"000000010",
  3940=>"000010001",
  3941=>"010000010",
  3942=>"001010101",
  3943=>"100001010",
  3944=>"001001111",
  3945=>"111111010",
  3946=>"000100101",
  3947=>"011101110",
  3948=>"001100000",
  3949=>"101000001",
  3950=>"100100111",
  3951=>"100110101",
  3952=>"010001010",
  3953=>"110011111",
  3954=>"100011011",
  3955=>"100101100",
  3956=>"000010001",
  3957=>"100110110",
  3958=>"101011100",
  3959=>"000101010",
  3960=>"111001111",
  3961=>"011001110",
  3962=>"101110001",
  3963=>"010110111",
  3964=>"110110111",
  3965=>"010110110",
  3966=>"011110001",
  3967=>"011100101",
  3968=>"101010111",
  3969=>"010011101",
  3970=>"111110101",
  3971=>"001100010",
  3972=>"100100001",
  3973=>"010111000",
  3974=>"100101001",
  3975=>"110001001",
  3976=>"110010111",
  3977=>"000100011",
  3978=>"010001010",
  3979=>"001010000",
  3980=>"010100110",
  3981=>"101001000",
  3982=>"010101110",
  3983=>"110010001",
  3984=>"101111100",
  3985=>"100010000",
  3986=>"011111100",
  3987=>"110110010",
  3988=>"110011101",
  3989=>"001111110",
  3990=>"000001110",
  3991=>"011111011",
  3992=>"111010001",
  3993=>"111101111",
  3994=>"001010110",
  3995=>"010111100",
  3996=>"101110111",
  3997=>"001110010",
  3998=>"101101000",
  3999=>"100011110",
  4000=>"010100101",
  4001=>"101001000",
  4002=>"101010100",
  4003=>"011111101",
  4004=>"001110101",
  4005=>"101000010",
  4006=>"000011101",
  4007=>"100000000",
  4008=>"100111111",
  4009=>"000100001",
  4010=>"010101001",
  4011=>"110010100",
  4012=>"010010100",
  4013=>"011010010",
  4014=>"101111001",
  4015=>"011101100",
  4016=>"001000000",
  4017=>"110010100",
  4018=>"100001011",
  4019=>"110000011",
  4020=>"000111000",
  4021=>"001010101",
  4022=>"001001111",
  4023=>"010001010",
  4024=>"000111111",
  4025=>"100001110",
  4026=>"110111001",
  4027=>"011111000",
  4028=>"010100111",
  4029=>"111100010",
  4030=>"010011111",
  4031=>"111010001",
  4032=>"101010111",
  4033=>"111011010",
  4034=>"010110110",
  4035=>"100111111",
  4036=>"101011010",
  4037=>"100111001",
  4038=>"001001001",
  4039=>"100100101",
  4040=>"001011111",
  4041=>"110100111",
  4042=>"111110111",
  4043=>"011000001",
  4044=>"100010110",
  4045=>"000000101",
  4046=>"110100010",
  4047=>"011010000",
  4048=>"101010111",
  4049=>"100000101",
  4050=>"000100000",
  4051=>"101111001",
  4052=>"110001101",
  4053=>"111101010",
  4054=>"001110010",
  4055=>"000011011",
  4056=>"101100111",
  4057=>"110101001",
  4058=>"111101010",
  4059=>"111010100",
  4060=>"011110001",
  4061=>"101110111",
  4062=>"111010011",
  4063=>"010100011",
  4064=>"100000010",
  4065=>"101010101",
  4066=>"001011001",
  4067=>"011001011",
  4068=>"110011001",
  4069=>"010001001",
  4070=>"001011100",
  4071=>"010001111",
  4072=>"110000110",
  4073=>"110110101",
  4074=>"010001001",
  4075=>"000110101",
  4076=>"000100010",
  4077=>"011010001",
  4078=>"010000000",
  4079=>"011111000",
  4080=>"001000100",
  4081=>"010011011",
  4082=>"111011110",
  4083=>"000110101",
  4084=>"110001001",
  4085=>"000001011",
  4086=>"000111101",
  4087=>"001111000",
  4088=>"001010110",
  4089=>"011001000",
  4090=>"011011011",
  4091=>"101100001",
  4092=>"010100000",
  4093=>"111100100",
  4094=>"100100100",
  4095=>"011100010",
  4096=>"001111011",
  4097=>"010111111",
  4098=>"100011101",
  4099=>"011110110",
  4100=>"011101011",
  4101=>"110101110",
  4102=>"001010110",
  4103=>"001000001",
  4104=>"111100111",
  4105=>"000011111",
  4106=>"000000011",
  4107=>"110010000",
  4108=>"010010001",
  4109=>"001100000",
  4110=>"110001000",
  4111=>"111010010",
  4112=>"100100001",
  4113=>"000111100",
  4114=>"111010110",
  4115=>"010011100",
  4116=>"000001011",
  4117=>"111101001",
  4118=>"000000110",
  4119=>"010010111",
  4120=>"001110100",
  4121=>"001000110",
  4122=>"010011110",
  4123=>"100011010",
  4124=>"101011000",
  4125=>"010101100",
  4126=>"010001101",
  4127=>"000111001",
  4128=>"001000010",
  4129=>"001110001",
  4130=>"101110001",
  4131=>"111110111",
  4132=>"011110011",
  4133=>"110010000",
  4134=>"001000010",
  4135=>"111111111",
  4136=>"010011100",
  4137=>"001010100",
  4138=>"010100000",
  4139=>"100110101",
  4140=>"001110110",
  4141=>"110010111",
  4142=>"111111101",
  4143=>"111000001",
  4144=>"101100000",
  4145=>"011011101",
  4146=>"111001010",
  4147=>"001011001",
  4148=>"110111011",
  4149=>"101111100",
  4150=>"000110000",
  4151=>"000100101",
  4152=>"100100101",
  4153=>"011100111",
  4154=>"001000010",
  4155=>"011110101",
  4156=>"011010000",
  4157=>"000010000",
  4158=>"100111111",
  4159=>"001010110",
  4160=>"011110001",
  4161=>"000010011",
  4162=>"010111010",
  4163=>"110101101",
  4164=>"101100101",
  4165=>"010000101",
  4166=>"111100001",
  4167=>"101110111",
  4168=>"111010000",
  4169=>"011000100",
  4170=>"001101101",
  4171=>"101000110",
  4172=>"010110000",
  4173=>"111100111",
  4174=>"111100011",
  4175=>"011100000",
  4176=>"100000110",
  4177=>"010111000",
  4178=>"101001011",
  4179=>"001110110",
  4180=>"010000001",
  4181=>"001001001",
  4182=>"000000100",
  4183=>"000101000",
  4184=>"000000011",
  4185=>"101011010",
  4186=>"100010011",
  4187=>"110100101",
  4188=>"111011111",
  4189=>"100101001",
  4190=>"000010010",
  4191=>"010001111",
  4192=>"111000001",
  4193=>"000111110",
  4194=>"101011110",
  4195=>"000110101",
  4196=>"101100100",
  4197=>"100100101",
  4198=>"110111101",
  4199=>"101001000",
  4200=>"101111101",
  4201=>"101111011",
  4202=>"101010100",
  4203=>"100001110",
  4204=>"101101101",
  4205=>"100000000",
  4206=>"001000110",
  4207=>"001010011",
  4208=>"111011111",
  4209=>"100001101",
  4210=>"101001011",
  4211=>"000010100",
  4212=>"101000110",
  4213=>"001000110",
  4214=>"110100010",
  4215=>"010100010",
  4216=>"000110101",
  4217=>"111011001",
  4218=>"111010110",
  4219=>"110010000",
  4220=>"101100000",
  4221=>"110110001",
  4222=>"111101101",
  4223=>"000010000",
  4224=>"000100000",
  4225=>"000010100",
  4226=>"101101111",
  4227=>"010110001",
  4228=>"111001111",
  4229=>"000100010",
  4230=>"011111000",
  4231=>"000100000",
  4232=>"011101111",
  4233=>"100000000",
  4234=>"101001000",
  4235=>"100101001",
  4236=>"001011100",
  4237=>"100010011",
  4238=>"000000111",
  4239=>"000010010",
  4240=>"010000100",
  4241=>"010001011",
  4242=>"001011011",
  4243=>"001101111",
  4244=>"101001000",
  4245=>"101010101",
  4246=>"001011001",
  4247=>"000100101",
  4248=>"101100100",
  4249=>"100011110",
  4250=>"011001101",
  4251=>"110111101",
  4252=>"110000011",
  4253=>"001010000",
  4254=>"010000001",
  4255=>"111001010",
  4256=>"001000010",
  4257=>"100001100",
  4258=>"101010001",
  4259=>"000010001",
  4260=>"010000111",
  4261=>"111010110",
  4262=>"100001101",
  4263=>"010100010",
  4264=>"111101000",
  4265=>"111111001",
  4266=>"010100100",
  4267=>"111010101",
  4268=>"011111011",
  4269=>"111111000",
  4270=>"110111111",
  4271=>"101111110",
  4272=>"011011101",
  4273=>"100111000",
  4274=>"100011010",
  4275=>"111101110",
  4276=>"010101001",
  4277=>"000110000",
  4278=>"101101111",
  4279=>"010001110",
  4280=>"110010010",
  4281=>"010011001",
  4282=>"101110001",
  4283=>"011011010",
  4284=>"001011101",
  4285=>"110101100",
  4286=>"100110111",
  4287=>"011011001",
  4288=>"111110001",
  4289=>"111110001",
  4290=>"000001011",
  4291=>"100010011",
  4292=>"111010011",
  4293=>"010010111",
  4294=>"100000100",
  4295=>"100011111",
  4296=>"000011101",
  4297=>"010011100",
  4298=>"010000111",
  4299=>"111010001",
  4300=>"110000101",
  4301=>"110111001",
  4302=>"010001011",
  4303=>"010011001",
  4304=>"001100000",
  4305=>"100010101",
  4306=>"101000000",
  4307=>"001010111",
  4308=>"111100011",
  4309=>"111101010",
  4310=>"101000001",
  4311=>"110001010",
  4312=>"000001111",
  4313=>"100001000",
  4314=>"111010110",
  4315=>"010100101",
  4316=>"010010010",
  4317=>"111001110",
  4318=>"110010000",
  4319=>"100011000",
  4320=>"100101100",
  4321=>"000101000",
  4322=>"000101000",
  4323=>"111000000",
  4324=>"011001111",
  4325=>"000001101",
  4326=>"001101001",
  4327=>"001101111",
  4328=>"101001110",
  4329=>"000100111",
  4330=>"001100101",
  4331=>"111000011",
  4332=>"101010101",
  4333=>"000101001",
  4334=>"100010110",
  4335=>"010110110",
  4336=>"101001101",
  4337=>"010001010",
  4338=>"000111000",
  4339=>"100101010",
  4340=>"100100110",
  4341=>"011100100",
  4342=>"101011111",
  4343=>"000101110",
  4344=>"011001010",
  4345=>"111101001",
  4346=>"000111001",
  4347=>"001000010",
  4348=>"010000100",
  4349=>"000010010",
  4350=>"110101011",
  4351=>"011010100",
  4352=>"110001110",
  4353=>"101110010",
  4354=>"111111000",
  4355=>"101101010",
  4356=>"101000101",
  4357=>"001100101",
  4358=>"000000100",
  4359=>"101100100",
  4360=>"100111001",
  4361=>"101010011",
  4362=>"101110110",
  4363=>"111100011",
  4364=>"110100001",
  4365=>"110001001",
  4366=>"010100100",
  4367=>"110110110",
  4368=>"111111111",
  4369=>"101011000",
  4370=>"100000010",
  4371=>"010111000",
  4372=>"110000011",
  4373=>"101100000",
  4374=>"011101010",
  4375=>"000110101",
  4376=>"101001011",
  4377=>"000011010",
  4378=>"011001001",
  4379=>"001110111",
  4380=>"000001010",
  4381=>"001111001",
  4382=>"010100101",
  4383=>"011101100",
  4384=>"010100101",
  4385=>"010011011",
  4386=>"001011000",
  4387=>"010000100",
  4388=>"011100100",
  4389=>"100111100",
  4390=>"010010101",
  4391=>"110011110",
  4392=>"010101001",
  4393=>"110001000",
  4394=>"101101101",
  4395=>"100111010",
  4396=>"100000000",
  4397=>"010011000",
  4398=>"101001001",
  4399=>"000101010",
  4400=>"001000010",
  4401=>"111111010",
  4402=>"010111101",
  4403=>"111111000",
  4404=>"101101000",
  4405=>"100111001",
  4406=>"100111001",
  4407=>"011000110",
  4408=>"010110111",
  4409=>"100000010",
  4410=>"000110100",
  4411=>"110000111",
  4412=>"111001001",
  4413=>"101100001",
  4414=>"110111011",
  4415=>"001001010",
  4416=>"001101000",
  4417=>"110101111",
  4418=>"100111010",
  4419=>"011110010",
  4420=>"101100110",
  4421=>"110100111",
  4422=>"110100110",
  4423=>"001110010",
  4424=>"000001011",
  4425=>"000000001",
  4426=>"101110101",
  4427=>"100001110",
  4428=>"110001100",
  4429=>"011100011",
  4430=>"001001100",
  4431=>"111011011",
  4432=>"000011000",
  4433=>"111000000",
  4434=>"001011010",
  4435=>"101100110",
  4436=>"101101101",
  4437=>"110010110",
  4438=>"001010001",
  4439=>"000001001",
  4440=>"110010101",
  4441=>"111101111",
  4442=>"101001111",
  4443=>"010011111",
  4444=>"001011100",
  4445=>"100110111",
  4446=>"111011010",
  4447=>"001010000",
  4448=>"110001000",
  4449=>"000011101",
  4450=>"000010001",
  4451=>"101101000",
  4452=>"101110010",
  4453=>"110000001",
  4454=>"110000110",
  4455=>"100111010",
  4456=>"010011111",
  4457=>"100110000",
  4458=>"000111010",
  4459=>"110000011",
  4460=>"111101001",
  4461=>"000011000",
  4462=>"111111001",
  4463=>"001000111",
  4464=>"010001010",
  4465=>"111001001",
  4466=>"111110010",
  4467=>"100010100",
  4468=>"101001010",
  4469=>"010101100",
  4470=>"101111001",
  4471=>"000001010",
  4472=>"100001000",
  4473=>"110011100",
  4474=>"100111110",
  4475=>"000100100",
  4476=>"000100100",
  4477=>"001110001",
  4478=>"110001010",
  4479=>"000101010",
  4480=>"000010100",
  4481=>"111011010",
  4482=>"100001001",
  4483=>"010011111",
  4484=>"011110100",
  4485=>"101101100",
  4486=>"101000111",
  4487=>"101111000",
  4488=>"000011011",
  4489=>"011111101",
  4490=>"110111111",
  4491=>"001100011",
  4492=>"100101001",
  4493=>"101001100",
  4494=>"100110101",
  4495=>"010000111",
  4496=>"101011000",
  4497=>"101011010",
  4498=>"111011110",
  4499=>"111010101",
  4500=>"100100010",
  4501=>"001010010",
  4502=>"110100100",
  4503=>"101111010",
  4504=>"111111101",
  4505=>"001001001",
  4506=>"101101100",
  4507=>"001111110",
  4508=>"101001100",
  4509=>"000101101",
  4510=>"010100110",
  4511=>"011101000",
  4512=>"101011100",
  4513=>"100101100",
  4514=>"001001011",
  4515=>"011010100",
  4516=>"111111100",
  4517=>"011111000",
  4518=>"111101101",
  4519=>"111101010",
  4520=>"011000010",
  4521=>"101101010",
  4522=>"000100001",
  4523=>"001000111",
  4524=>"010111001",
  4525=>"011100000",
  4526=>"111111100",
  4527=>"100010101",
  4528=>"010001110",
  4529=>"000101011",
  4530=>"001101111",
  4531=>"001101101",
  4532=>"101101010",
  4533=>"100101011",
  4534=>"011111111",
  4535=>"000000001",
  4536=>"001001011",
  4537=>"101111000",
  4538=>"001110010",
  4539=>"100001101",
  4540=>"101001001",
  4541=>"101010111",
  4542=>"011101001",
  4543=>"100111000",
  4544=>"000001000",
  4545=>"001001101",
  4546=>"100111110",
  4547=>"101110110",
  4548=>"111011010",
  4549=>"110100010",
  4550=>"111001110",
  4551=>"110001111",
  4552=>"010110100",
  4553=>"000101001",
  4554=>"000100011",
  4555=>"101011100",
  4556=>"101010000",
  4557=>"111110011",
  4558=>"001010001",
  4559=>"100101110",
  4560=>"110111111",
  4561=>"110010010",
  4562=>"011010001",
  4563=>"111110000",
  4564=>"110011111",
  4565=>"000100011",
  4566=>"110010111",
  4567=>"010010110",
  4568=>"000110001",
  4569=>"010010101",
  4570=>"011010001",
  4571=>"110100101",
  4572=>"100010101",
  4573=>"101100010",
  4574=>"111001000",
  4575=>"000010000",
  4576=>"001001110",
  4577=>"001111000",
  4578=>"011011011",
  4579=>"101110010",
  4580=>"000000010",
  4581=>"101010111",
  4582=>"101001010",
  4583=>"010000101",
  4584=>"111000011",
  4585=>"001000110",
  4586=>"000010100",
  4587=>"000000011",
  4588=>"000000010",
  4589=>"011101100",
  4590=>"000011100",
  4591=>"100110001",
  4592=>"011100110",
  4593=>"111110001",
  4594=>"110010110",
  4595=>"111110000",
  4596=>"010110000",
  4597=>"000000011",
  4598=>"000111000",
  4599=>"111110000",
  4600=>"011011000",
  4601=>"101011111",
  4602=>"111001010",
  4603=>"111101011",
  4604=>"111001110",
  4605=>"101001000",
  4606=>"101001011",
  4607=>"110010111",
  4608=>"010101100",
  4609=>"110001011",
  4610=>"111111010",
  4611=>"010101000",
  4612=>"111110011",
  4613=>"011010100",
  4614=>"000111110",
  4615=>"100100101",
  4616=>"000110001",
  4617=>"100110000",
  4618=>"110010010",
  4619=>"101000000",
  4620=>"001011011",
  4621=>"101100100",
  4622=>"001100010",
  4623=>"011101111",
  4624=>"011111011",
  4625=>"001010011",
  4626=>"100110111",
  4627=>"001110010",
  4628=>"001101110",
  4629=>"100010111",
  4630=>"000101000",
  4631=>"101010100",
  4632=>"111010001",
  4633=>"101101010",
  4634=>"100000001",
  4635=>"000101101",
  4636=>"111100000",
  4637=>"100100001",
  4638=>"111110100",
  4639=>"100110011",
  4640=>"011110010",
  4641=>"010101111",
  4642=>"100100000",
  4643=>"010001010",
  4644=>"000001100",
  4645=>"100001111",
  4646=>"000111100",
  4647=>"100000011",
  4648=>"011000010",
  4649=>"110110110",
  4650=>"110101101",
  4651=>"110010000",
  4652=>"010101101",
  4653=>"011010101",
  4654=>"111010000",
  4655=>"000011010",
  4656=>"000000101",
  4657=>"001111011",
  4658=>"101110100",
  4659=>"101111000",
  4660=>"011001011",
  4661=>"100111001",
  4662=>"101000110",
  4663=>"100010110",
  4664=>"111011101",
  4665=>"101010000",
  4666=>"100110100",
  4667=>"111001110",
  4668=>"101011001",
  4669=>"111001011",
  4670=>"111110111",
  4671=>"011101111",
  4672=>"000101100",
  4673=>"011000000",
  4674=>"111101010",
  4675=>"100110010",
  4676=>"011000001",
  4677=>"101011000",
  4678=>"100101000",
  4679=>"111010011",
  4680=>"001010100",
  4681=>"101110010",
  4682=>"011110110",
  4683=>"111000000",
  4684=>"000110010",
  4685=>"000110100",
  4686=>"010010100",
  4687=>"001011011",
  4688=>"100111100",
  4689=>"100000101",
  4690=>"001100100",
  4691=>"001011100",
  4692=>"001011000",
  4693=>"110001011",
  4694=>"001110000",
  4695=>"011111000",
  4696=>"011001101",
  4697=>"000111101",
  4698=>"001011101",
  4699=>"111011100",
  4700=>"010111010",
  4701=>"100101110",
  4702=>"000111111",
  4703=>"010111111",
  4704=>"010111101",
  4705=>"010001001",
  4706=>"011000010",
  4707=>"011000111",
  4708=>"000111010",
  4709=>"111100010",
  4710=>"011000101",
  4711=>"010111110",
  4712=>"111010101",
  4713=>"110111100",
  4714=>"001011101",
  4715=>"000000100",
  4716=>"000111111",
  4717=>"100101000",
  4718=>"011100101",
  4719=>"010000011",
  4720=>"011000101",
  4721=>"001111101",
  4722=>"000100100",
  4723=>"111101011",
  4724=>"101011010",
  4725=>"010110111",
  4726=>"100000100",
  4727=>"000001000",
  4728=>"100101001",
  4729=>"100001101",
  4730=>"101010111",
  4731=>"011110011",
  4732=>"010011101",
  4733=>"010010101",
  4734=>"010100000",
  4735=>"111110100",
  4736=>"110011011",
  4737=>"110000111",
  4738=>"000001111",
  4739=>"011000110",
  4740=>"011100011",
  4741=>"110010100",
  4742=>"110001001",
  4743=>"010010010",
  4744=>"100011000",
  4745=>"101010011",
  4746=>"111101111",
  4747=>"110000110",
  4748=>"101000101",
  4749=>"001111100",
  4750=>"011000001",
  4751=>"111011011",
  4752=>"010000001",
  4753=>"111101000",
  4754=>"011111110",
  4755=>"001111111",
  4756=>"011010011",
  4757=>"100001100",
  4758=>"010010011",
  4759=>"011111101",
  4760=>"010001011",
  4761=>"011111101",
  4762=>"010011011",
  4763=>"000101101",
  4764=>"011010000",
  4765=>"100010101",
  4766=>"110011101",
  4767=>"001010110",
  4768=>"011010101",
  4769=>"010011100",
  4770=>"010011100",
  4771=>"000000111",
  4772=>"110110101",
  4773=>"010100000",
  4774=>"101000001",
  4775=>"100111111",
  4776=>"001111000",
  4777=>"111011000",
  4778=>"100110100",
  4779=>"101111111",
  4780=>"000101101",
  4781=>"111110011",
  4782=>"001100010",
  4783=>"101010110",
  4784=>"101000000",
  4785=>"001010000",
  4786=>"000001011",
  4787=>"000101111",
  4788=>"011000101",
  4789=>"101010101",
  4790=>"000111010",
  4791=>"101100001",
  4792=>"101000011",
  4793=>"101010111",
  4794=>"011111001",
  4795=>"110001110",
  4796=>"101010011",
  4797=>"000010101",
  4798=>"000000011",
  4799=>"001011101",
  4800=>"100110101",
  4801=>"010001000",
  4802=>"010110110",
  4803=>"011010100",
  4804=>"100101001",
  4805=>"100011111",
  4806=>"000010001",
  4807=>"011011010",
  4808=>"011011011",
  4809=>"101101011",
  4810=>"011101101",
  4811=>"111110011",
  4812=>"011010101",
  4813=>"100010010",
  4814=>"001100000",
  4815=>"101011111",
  4816=>"001000110",
  4817=>"011000000",
  4818=>"100111010",
  4819=>"011111111",
  4820=>"000001110",
  4821=>"110011000",
  4822=>"100011001",
  4823=>"010101100",
  4824=>"100010011",
  4825=>"101101001",
  4826=>"100100100",
  4827=>"000001000",
  4828=>"100101111",
  4829=>"000110011",
  4830=>"110100111",
  4831=>"011100000",
  4832=>"010110110",
  4833=>"011001001",
  4834=>"111011000",
  4835=>"110111011",
  4836=>"110100101",
  4837=>"101001110",
  4838=>"111101001",
  4839=>"001101111",
  4840=>"011100000",
  4841=>"101010011",
  4842=>"010001110",
  4843=>"010010010",
  4844=>"111111001",
  4845=>"010110010",
  4846=>"110001001",
  4847=>"000110110",
  4848=>"011010010",
  4849=>"110010000",
  4850=>"001000100",
  4851=>"110000000",
  4852=>"011101000",
  4853=>"011111010",
  4854=>"000001100",
  4855=>"100011101",
  4856=>"110110011",
  4857=>"011000110",
  4858=>"101101101",
  4859=>"100101100",
  4860=>"010010000",
  4861=>"000010010",
  4862=>"101111100",
  4863=>"101001110",
  4864=>"101011101",
  4865=>"100101001",
  4866=>"000111001",
  4867=>"111110001",
  4868=>"010111011",
  4869=>"010010101",
  4870=>"111101110",
  4871=>"101000100",
  4872=>"000000000",
  4873=>"000000011",
  4874=>"111001111",
  4875=>"101010111",
  4876=>"101111011",
  4877=>"001010100",
  4878=>"010010010",
  4879=>"011001100",
  4880=>"010000100",
  4881=>"000100111",
  4882=>"011000100",
  4883=>"101010100",
  4884=>"010011100",
  4885=>"101001001",
  4886=>"000001011",
  4887=>"000000100",
  4888=>"001011000",
  4889=>"100101001",
  4890=>"100000011",
  4891=>"110110110",
  4892=>"101111010",
  4893=>"110110001",
  4894=>"000011000",
  4895=>"001111111",
  4896=>"110111010",
  4897=>"101001101",
  4898=>"101010000",
  4899=>"101011010",
  4900=>"001111001",
  4901=>"101010001",
  4902=>"000000100",
  4903=>"010100110",
  4904=>"011111101",
  4905=>"101111111",
  4906=>"010001100",
  4907=>"011001101",
  4908=>"011011000",
  4909=>"010001000",
  4910=>"000000000",
  4911=>"100010011",
  4912=>"010100100",
  4913=>"101001111",
  4914=>"101100011",
  4915=>"101100111",
  4916=>"111100010",
  4917=>"100110111",
  4918=>"101011000",
  4919=>"110011101",
  4920=>"110011000",
  4921=>"010010100",
  4922=>"100001000",
  4923=>"001101010",
  4924=>"001101100",
  4925=>"001001101",
  4926=>"111000100",
  4927=>"011100010",
  4928=>"110001001",
  4929=>"111010010",
  4930=>"001111101",
  4931=>"100100010",
  4932=>"010100110",
  4933=>"111110111",
  4934=>"000111011",
  4935=>"000000110",
  4936=>"001010110",
  4937=>"101101100",
  4938=>"100010110",
  4939=>"101010110",
  4940=>"011110000",
  4941=>"100001110",
  4942=>"100001100",
  4943=>"010000111",
  4944=>"111010101",
  4945=>"110011011",
  4946=>"111010111",
  4947=>"100000011",
  4948=>"000101101",
  4949=>"000101000",
  4950=>"100111101",
  4951=>"100111110",
  4952=>"010010010",
  4953=>"101000011",
  4954=>"100100010",
  4955=>"001001001",
  4956=>"100000100",
  4957=>"000100111",
  4958=>"001110011",
  4959=>"101010110",
  4960=>"110011110",
  4961=>"010010101",
  4962=>"011111101",
  4963=>"110100010",
  4964=>"001010010",
  4965=>"111000010",
  4966=>"110001100",
  4967=>"100101000",
  4968=>"110010100",
  4969=>"000111101",
  4970=>"111010110",
  4971=>"000000101",
  4972=>"111100100",
  4973=>"100100001",
  4974=>"010101000",
  4975=>"011011111",
  4976=>"111001011",
  4977=>"010001101",
  4978=>"100010010",
  4979=>"101101011",
  4980=>"011001000",
  4981=>"010011110",
  4982=>"111010101",
  4983=>"110000000",
  4984=>"110101000",
  4985=>"111011110",
  4986=>"011001011",
  4987=>"000110110",
  4988=>"011011000",
  4989=>"110000011",
  4990=>"100100000",
  4991=>"111101111",
  4992=>"101001110",
  4993=>"000101001",
  4994=>"100100111",
  4995=>"100101111",
  4996=>"000011100",
  4997=>"111111000",
  4998=>"001000010",
  4999=>"001101010",
  5000=>"010101101",
  5001=>"101110100",
  5002=>"100000101",
  5003=>"111000001",
  5004=>"000100100",
  5005=>"100111000",
  5006=>"001010001",
  5007=>"000010001",
  5008=>"110000001",
  5009=>"001011001",
  5010=>"100011000",
  5011=>"100000000",
  5012=>"011010000",
  5013=>"000010011",
  5014=>"001110011",
  5015=>"001101001",
  5016=>"111110110",
  5017=>"011101101",
  5018=>"100000111",
  5019=>"000101110",
  5020=>"010010011",
  5021=>"011110110",
  5022=>"000101101",
  5023=>"101000100",
  5024=>"100101010",
  5025=>"011110011",
  5026=>"110100000",
  5027=>"101010101",
  5028=>"011000000",
  5029=>"000001011",
  5030=>"111111110",
  5031=>"101000100",
  5032=>"000111111",
  5033=>"010000101",
  5034=>"011011101",
  5035=>"010000010",
  5036=>"101010100",
  5037=>"111111000",
  5038=>"110100110",
  5039=>"010000110",
  5040=>"000101111",
  5041=>"111111011",
  5042=>"000010010",
  5043=>"110011011",
  5044=>"000000110",
  5045=>"101000111",
  5046=>"011110110",
  5047=>"000000110",
  5048=>"100100111",
  5049=>"100010010",
  5050=>"111000001",
  5051=>"110101001",
  5052=>"100101111",
  5053=>"110101111",
  5054=>"111001100",
  5055=>"010101011",
  5056=>"000100001",
  5057=>"110110111",
  5058=>"001000101",
  5059=>"011010011",
  5060=>"000000100",
  5061=>"101001011",
  5062=>"110101000",
  5063=>"011100111",
  5064=>"100110100",
  5065=>"000011101",
  5066=>"011101101",
  5067=>"111111110",
  5068=>"111001111",
  5069=>"000010001",
  5070=>"110110001",
  5071=>"101001101",
  5072=>"100010111",
  5073=>"010111000",
  5074=>"000001100",
  5075=>"100010101",
  5076=>"000000001",
  5077=>"100001001",
  5078=>"100010001",
  5079=>"110000101",
  5080=>"101011010",
  5081=>"110101110",
  5082=>"100110001",
  5083=>"010101011",
  5084=>"011010101",
  5085=>"110011011",
  5086=>"111010011",
  5087=>"000100010",
  5088=>"000100000",
  5089=>"101000000",
  5090=>"110000111",
  5091=>"000010110",
  5092=>"101100011",
  5093=>"110111101",
  5094=>"011100000",
  5095=>"100011111",
  5096=>"000000000",
  5097=>"000000100",
  5098=>"001100001",
  5099=>"101000010",
  5100=>"110111011",
  5101=>"111000010",
  5102=>"011001111",
  5103=>"000010011",
  5104=>"011000000",
  5105=>"110110111",
  5106=>"111101111",
  5107=>"011001011",
  5108=>"110010001",
  5109=>"101011110",
  5110=>"000111100",
  5111=>"001011110",
  5112=>"100111010",
  5113=>"100111110",
  5114=>"100100001",
  5115=>"100111110",
  5116=>"011110111",
  5117=>"000100111",
  5118=>"000000100",
  5119=>"011001010",
  5120=>"011011100",
  5121=>"100111111",
  5122=>"100110010",
  5123=>"111000000",
  5124=>"111010001",
  5125=>"001011011",
  5126=>"000100000",
  5127=>"110000100",
  5128=>"011011110",
  5129=>"100011001",
  5130=>"110101000",
  5131=>"101110110",
  5132=>"001100001",
  5133=>"101110101",
  5134=>"111010101",
  5135=>"110101000",
  5136=>"111001010",
  5137=>"111011010",
  5138=>"001111011",
  5139=>"000000101",
  5140=>"111111011",
  5141=>"110010110",
  5142=>"100001001",
  5143=>"100011100",
  5144=>"100100000",
  5145=>"101111101",
  5146=>"010100000",
  5147=>"000010110",
  5148=>"011001110",
  5149=>"111111010",
  5150=>"101101111",
  5151=>"000110010",
  5152=>"010111000",
  5153=>"000010001",
  5154=>"100010111",
  5155=>"101100111",
  5156=>"000111001",
  5157=>"101110001",
  5158=>"000101001",
  5159=>"111000111",
  5160=>"001111111",
  5161=>"111110000",
  5162=>"110100011",
  5163=>"111011111",
  5164=>"100001010",
  5165=>"011110001",
  5166=>"100111011",
  5167=>"100000000",
  5168=>"010000111",
  5169=>"011101001",
  5170=>"100001000",
  5171=>"110011001",
  5172=>"011100101",
  5173=>"001100010",
  5174=>"001001100",
  5175=>"010010111",
  5176=>"001111100",
  5177=>"011010000",
  5178=>"000010010",
  5179=>"111010111",
  5180=>"100011001",
  5181=>"000010000",
  5182=>"001011010",
  5183=>"010111000",
  5184=>"101000011",
  5185=>"010000001",
  5186=>"111001001",
  5187=>"001100010",
  5188=>"100100100",
  5189=>"101101111",
  5190=>"011011101",
  5191=>"010001110",
  5192=>"101100010",
  5193=>"111111110",
  5194=>"111010101",
  5195=>"111110000",
  5196=>"011100010",
  5197=>"111101111",
  5198=>"011101010",
  5199=>"100110101",
  5200=>"000000001",
  5201=>"100100100",
  5202=>"000100011",
  5203=>"110011110",
  5204=>"011111001",
  5205=>"001000000",
  5206=>"111100011",
  5207=>"001111000",
  5208=>"110110111",
  5209=>"110001100",
  5210=>"100100011",
  5211=>"010110011",
  5212=>"011000000",
  5213=>"111011000",
  5214=>"110110101",
  5215=>"001000011",
  5216=>"011001110",
  5217=>"101111001",
  5218=>"000001111",
  5219=>"000110100",
  5220=>"000100000",
  5221=>"001001000",
  5222=>"100000100",
  5223=>"011101011",
  5224=>"001111111",
  5225=>"010100110",
  5226=>"010110111",
  5227=>"011100010",
  5228=>"000111100",
  5229=>"000011011",
  5230=>"100110000",
  5231=>"101100101",
  5232=>"101000111",
  5233=>"010011100",
  5234=>"100110000",
  5235=>"100000010",
  5236=>"101001010",
  5237=>"100001010",
  5238=>"101110001",
  5239=>"011101101",
  5240=>"000001110",
  5241=>"001010000",
  5242=>"101010110",
  5243=>"000011110",
  5244=>"111111111",
  5245=>"110011101",
  5246=>"011101111",
  5247=>"011000000",
  5248=>"011111111",
  5249=>"011111001",
  5250=>"110010101",
  5251=>"001111100",
  5252=>"100000011",
  5253=>"101100000",
  5254=>"001110111",
  5255=>"010110111",
  5256=>"101110010",
  5257=>"110001000",
  5258=>"011000110",
  5259=>"001001111",
  5260=>"100000011",
  5261=>"111001101",
  5262=>"100100001",
  5263=>"101000000",
  5264=>"111000000",
  5265=>"101010000",
  5266=>"111100010",
  5267=>"000100010",
  5268=>"111010010",
  5269=>"001101101",
  5270=>"100001110",
  5271=>"101001000",
  5272=>"110111000",
  5273=>"110111000",
  5274=>"001010000",
  5275=>"001010111",
  5276=>"100100010",
  5277=>"010001010",
  5278=>"011110000",
  5279=>"001001010",
  5280=>"001001101",
  5281=>"111010110",
  5282=>"011011000",
  5283=>"100010101",
  5284=>"110111011",
  5285=>"010111001",
  5286=>"001000001",
  5287=>"001011010",
  5288=>"000010000",
  5289=>"010010001",
  5290=>"001010011",
  5291=>"001001110",
  5292=>"101100010",
  5293=>"101011001",
  5294=>"010011010",
  5295=>"111001000",
  5296=>"000000011",
  5297=>"101000010",
  5298=>"110011100",
  5299=>"110010000",
  5300=>"110010001",
  5301=>"101101101",
  5302=>"000100101",
  5303=>"000011100",
  5304=>"100111001",
  5305=>"101010100",
  5306=>"101100010",
  5307=>"000000110",
  5308=>"001010011",
  5309=>"000111111",
  5310=>"011011001",
  5311=>"111001001",
  5312=>"000000110",
  5313=>"011011110",
  5314=>"101101001",
  5315=>"001111100",
  5316=>"011011000",
  5317=>"110011001",
  5318=>"111110001",
  5319=>"100001001",
  5320=>"101001111",
  5321=>"001111101",
  5322=>"001001011",
  5323=>"110111111",
  5324=>"011000101",
  5325=>"110111010",
  5326=>"010110101",
  5327=>"000010010",
  5328=>"010000010",
  5329=>"001001101",
  5330=>"110000111",
  5331=>"000101111",
  5332=>"101101110",
  5333=>"100000011",
  5334=>"110010101",
  5335=>"110111011",
  5336=>"000011001",
  5337=>"111100111",
  5338=>"011101010",
  5339=>"111110000",
  5340=>"110110001",
  5341=>"000000000",
  5342=>"100001001",
  5343=>"000101110",
  5344=>"001110010",
  5345=>"000001000",
  5346=>"111011000",
  5347=>"001100011",
  5348=>"111001110",
  5349=>"000111011",
  5350=>"001001010",
  5351=>"001001111",
  5352=>"010101010",
  5353=>"100000010",
  5354=>"000011000",
  5355=>"001011111",
  5356=>"111110101",
  5357=>"001000010",
  5358=>"101000110",
  5359=>"001001111",
  5360=>"100001000",
  5361=>"101101101",
  5362=>"011001010",
  5363=>"100011100",
  5364=>"110000010",
  5365=>"110010001",
  5366=>"100000110",
  5367=>"000000100",
  5368=>"010110010",
  5369=>"010111010",
  5370=>"111010100",
  5371=>"011001100",
  5372=>"000110011",
  5373=>"001011001",
  5374=>"111111111",
  5375=>"010101100",
  5376=>"001000101",
  5377=>"010101111",
  5378=>"011001011",
  5379=>"111010010",
  5380=>"011000000",
  5381=>"010100110",
  5382=>"010001010",
  5383=>"111110100",
  5384=>"001111101",
  5385=>"100010001",
  5386=>"111110110",
  5387=>"100000111",
  5388=>"011111011",
  5389=>"011111010",
  5390=>"101101011",
  5391=>"101000011",
  5392=>"111111111",
  5393=>"100001110",
  5394=>"101111010",
  5395=>"111010000",
  5396=>"111110110",
  5397=>"000000011",
  5398=>"100000101",
  5399=>"110101100",
  5400=>"010100111",
  5401=>"010110110",
  5402=>"000100001",
  5403=>"101011001",
  5404=>"101001100",
  5405=>"111111111",
  5406=>"111110011",
  5407=>"101110111",
  5408=>"000001111",
  5409=>"100101110",
  5410=>"101111010",
  5411=>"010001001",
  5412=>"011000000",
  5413=>"100100110",
  5414=>"100011110",
  5415=>"010000101",
  5416=>"001000100",
  5417=>"100010001",
  5418=>"100110000",
  5419=>"001000001",
  5420=>"000000000",
  5421=>"000001000",
  5422=>"001001000",
  5423=>"001001011",
  5424=>"000110100",
  5425=>"110001011",
  5426=>"011001100",
  5427=>"111110111",
  5428=>"000011110",
  5429=>"101101001",
  5430=>"000001011",
  5431=>"010010001",
  5432=>"111110100",
  5433=>"001010110",
  5434=>"000001110",
  5435=>"011011110",
  5436=>"100001000",
  5437=>"000111000",
  5438=>"011111010",
  5439=>"110011101",
  5440=>"100010111",
  5441=>"110110001",
  5442=>"011010000",
  5443=>"010011011",
  5444=>"110100110",
  5445=>"101100010",
  5446=>"000010011",
  5447=>"100110100",
  5448=>"110100000",
  5449=>"101000100",
  5450=>"101010101",
  5451=>"011110100",
  5452=>"110010010",
  5453=>"100110101",
  5454=>"100000011",
  5455=>"110001011",
  5456=>"110101111",
  5457=>"101111110",
  5458=>"110111110",
  5459=>"111110100",
  5460=>"100010010",
  5461=>"011010101",
  5462=>"010010001",
  5463=>"100110000",
  5464=>"000101000",
  5465=>"110000010",
  5466=>"010001100",
  5467=>"001111111",
  5468=>"100110000",
  5469=>"111101011",
  5470=>"101000101",
  5471=>"010101001",
  5472=>"000111111",
  5473=>"010011010",
  5474=>"110110111",
  5475=>"111001011",
  5476=>"100100100",
  5477=>"110001110",
  5478=>"110001100",
  5479=>"101001111",
  5480=>"010011010",
  5481=>"101000000",
  5482=>"011000110",
  5483=>"101001001",
  5484=>"000101111",
  5485=>"110101011",
  5486=>"001101110",
  5487=>"001100000",
  5488=>"001010010",
  5489=>"001011111",
  5490=>"100101000",
  5491=>"110001001",
  5492=>"001101000",
  5493=>"101110011",
  5494=>"101111000",
  5495=>"101011100",
  5496=>"001100110",
  5497=>"110010100",
  5498=>"111001011",
  5499=>"101010011",
  5500=>"010100100",
  5501=>"101000000",
  5502=>"101100100",
  5503=>"100011111",
  5504=>"111101100",
  5505=>"100000010",
  5506=>"001100111",
  5507=>"111000000",
  5508=>"001000000",
  5509=>"110001011",
  5510=>"010100110",
  5511=>"100001110",
  5512=>"001010100",
  5513=>"000100000",
  5514=>"011010110",
  5515=>"111111011",
  5516=>"100101000",
  5517=>"000010010",
  5518=>"001101111",
  5519=>"010101011",
  5520=>"000001010",
  5521=>"111101101",
  5522=>"111011111",
  5523=>"000000001",
  5524=>"110100101",
  5525=>"010100111",
  5526=>"000001011",
  5527=>"001001011",
  5528=>"011111010",
  5529=>"101000010",
  5530=>"101110110",
  5531=>"000011001",
  5532=>"101111101",
  5533=>"001001001",
  5534=>"010001100",
  5535=>"100100001",
  5536=>"110101110",
  5537=>"010000010",
  5538=>"000111101",
  5539=>"001001100",
  5540=>"011000000",
  5541=>"100000000",
  5542=>"111010011",
  5543=>"100000110",
  5544=>"010101110",
  5545=>"101010010",
  5546=>"101001100",
  5547=>"110111000",
  5548=>"101001100",
  5549=>"110111011",
  5550=>"001010010",
  5551=>"010110011",
  5552=>"011101010",
  5553=>"000000110",
  5554=>"001111110",
  5555=>"001101011",
  5556=>"011110111",
  5557=>"100011100",
  5558=>"110100110",
  5559=>"111010011",
  5560=>"001101001",
  5561=>"101111101",
  5562=>"011100011",
  5563=>"000011111",
  5564=>"110010000",
  5565=>"100100001",
  5566=>"000011100",
  5567=>"000101000",
  5568=>"001101111",
  5569=>"011100101",
  5570=>"110100100",
  5571=>"101100110",
  5572=>"111011111",
  5573=>"100110110",
  5574=>"000101000",
  5575=>"001000000",
  5576=>"111011111",
  5577=>"000111000",
  5578=>"110110100",
  5579=>"011001000",
  5580=>"011111010",
  5581=>"010010110",
  5582=>"100000110",
  5583=>"010111111",
  5584=>"101001110",
  5585=>"101101000",
  5586=>"010100011",
  5587=>"001001101",
  5588=>"111111101",
  5589=>"100111101",
  5590=>"111101000",
  5591=>"010100001",
  5592=>"110101110",
  5593=>"110010010",
  5594=>"100010101",
  5595=>"001001101",
  5596=>"110010000",
  5597=>"001110010",
  5598=>"111110000",
  5599=>"011100011",
  5600=>"001010011",
  5601=>"101000010",
  5602=>"100001110",
  5603=>"001011001",
  5604=>"010111011",
  5605=>"100101001",
  5606=>"011001100",
  5607=>"101100000",
  5608=>"111100000",
  5609=>"110110010",
  5610=>"110011100",
  5611=>"010000000",
  5612=>"001110101",
  5613=>"011101110",
  5614=>"011010101",
  5615=>"000100010",
  5616=>"011000101",
  5617=>"110111101",
  5618=>"101111000",
  5619=>"000110001",
  5620=>"101010110",
  5621=>"011111010",
  5622=>"011100000",
  5623=>"111001110",
  5624=>"011101001",
  5625=>"010100110",
  5626=>"000010100",
  5627=>"101011101",
  5628=>"110011011",
  5629=>"001101011",
  5630=>"010010011",
  5631=>"100101101",
  5632=>"110001100",
  5633=>"101001010",
  5634=>"111111111",
  5635=>"001111000",
  5636=>"110010111",
  5637=>"101010001",
  5638=>"010001001",
  5639=>"101101100",
  5640=>"001111000",
  5641=>"001011101",
  5642=>"101000000",
  5643=>"000000001",
  5644=>"101010110",
  5645=>"010001110",
  5646=>"100001100",
  5647=>"011101111",
  5648=>"100110011",
  5649=>"110110011",
  5650=>"100010110",
  5651=>"100001100",
  5652=>"010110001",
  5653=>"111001111",
  5654=>"110010001",
  5655=>"110011110",
  5656=>"010101010",
  5657=>"111000010",
  5658=>"100100010",
  5659=>"101100100",
  5660=>"111010011",
  5661=>"000000111",
  5662=>"010010101",
  5663=>"001001000",
  5664=>"100000100",
  5665=>"010110100",
  5666=>"000100111",
  5667=>"011100111",
  5668=>"101011100",
  5669=>"001001101",
  5670=>"001101101",
  5671=>"101011100",
  5672=>"001101010",
  5673=>"111001011",
  5674=>"101101011",
  5675=>"111011110",
  5676=>"011100110",
  5677=>"001001110",
  5678=>"001001101",
  5679=>"100010101",
  5680=>"000101010",
  5681=>"000011011",
  5682=>"110110111",
  5683=>"100000101",
  5684=>"000101011",
  5685=>"111000111",
  5686=>"101111010",
  5687=>"000000001",
  5688=>"000101011",
  5689=>"110111001",
  5690=>"011100001",
  5691=>"111000001",
  5692=>"110000100",
  5693=>"000000010",
  5694=>"001011101",
  5695=>"010101000",
  5696=>"111100010",
  5697=>"110000100",
  5698=>"000011001",
  5699=>"011111011",
  5700=>"100010111",
  5701=>"010001100",
  5702=>"111111001",
  5703=>"100110000",
  5704=>"100000110",
  5705=>"010101011",
  5706=>"010111001",
  5707=>"100010101",
  5708=>"110110000",
  5709=>"011101000",
  5710=>"011101010",
  5711=>"000101001",
  5712=>"000110100",
  5713=>"011110101",
  5714=>"000001001",
  5715=>"110001100",
  5716=>"011100111",
  5717=>"100111110",
  5718=>"111101110",
  5719=>"010111010",
  5720=>"101101111",
  5721=>"010001011",
  5722=>"011011010",
  5723=>"011000100",
  5724=>"111010001",
  5725=>"000001101",
  5726=>"010111011",
  5727=>"011001010",
  5728=>"010010001",
  5729=>"010100101",
  5730=>"111011001",
  5731=>"100100101",
  5732=>"111011111",
  5733=>"110001111",
  5734=>"110111101",
  5735=>"100111110",
  5736=>"001010101",
  5737=>"110110001",
  5738=>"111110111",
  5739=>"000001001",
  5740=>"000101000",
  5741=>"000100101",
  5742=>"100000000",
  5743=>"001100101",
  5744=>"100101001",
  5745=>"011010101",
  5746=>"110010110",
  5747=>"000001010",
  5748=>"100100111",
  5749=>"100011010",
  5750=>"011110010",
  5751=>"100110101",
  5752=>"010011011",
  5753=>"000111000",
  5754=>"000001010",
  5755=>"010000100",
  5756=>"100100011",
  5757=>"101000100",
  5758=>"110000100",
  5759=>"010111010",
  5760=>"110010000",
  5761=>"111010111",
  5762=>"111010101",
  5763=>"011001011",
  5764=>"101100100",
  5765=>"011110001",
  5766=>"010001110",
  5767=>"100010010",
  5768=>"111111001",
  5769=>"001001111",
  5770=>"001001111",
  5771=>"011110001",
  5772=>"110000100",
  5773=>"101110001",
  5774=>"110101111",
  5775=>"111111011",
  5776=>"011100111",
  5777=>"010110110",
  5778=>"101000000",
  5779=>"101111000",
  5780=>"001001011",
  5781=>"000011000",
  5782=>"101111110",
  5783=>"010000010",
  5784=>"100110000",
  5785=>"101001010",
  5786=>"011011110",
  5787=>"110011100",
  5788=>"010111010",
  5789=>"101000010",
  5790=>"011111101",
  5791=>"000100011",
  5792=>"000011000",
  5793=>"100100110",
  5794=>"011011000",
  5795=>"010000110",
  5796=>"010010101",
  5797=>"001001010",
  5798=>"011010110",
  5799=>"100011000",
  5800=>"110100111",
  5801=>"110010111",
  5802=>"100000010",
  5803=>"000010000",
  5804=>"111011110",
  5805=>"110001110",
  5806=>"000010110",
  5807=>"111011011",
  5808=>"100011000",
  5809=>"001100101",
  5810=>"110110101",
  5811=>"001101101",
  5812=>"110110100",
  5813=>"011110000",
  5814=>"100111001",
  5815=>"100111110",
  5816=>"111111010",
  5817=>"101010000",
  5818=>"011011010",
  5819=>"000011010",
  5820=>"111101101",
  5821=>"100000100",
  5822=>"000111100",
  5823=>"111101100",
  5824=>"111101001",
  5825=>"100111011",
  5826=>"011000000",
  5827=>"100001110",
  5828=>"101011101",
  5829=>"000111000",
  5830=>"000100101",
  5831=>"100111010",
  5832=>"011000011",
  5833=>"100101010",
  5834=>"110010101",
  5835=>"111010110",
  5836=>"100110110",
  5837=>"010101110",
  5838=>"001001001",
  5839=>"111001101",
  5840=>"110000000",
  5841=>"100000110",
  5842=>"000010101",
  5843=>"111111010",
  5844=>"010110111",
  5845=>"010011001",
  5846=>"001110010",
  5847=>"010010010",
  5848=>"110011101",
  5849=>"001111001",
  5850=>"111010000",
  5851=>"011001000",
  5852=>"101111111",
  5853=>"101101010",
  5854=>"011100011",
  5855=>"100000101",
  5856=>"000011100",
  5857=>"011001111",
  5858=>"011111100",
  5859=>"011011111",
  5860=>"000101001",
  5861=>"000001100",
  5862=>"100110111",
  5863=>"000111001",
  5864=>"111100000",
  5865=>"111001100",
  5866=>"111000110",
  5867=>"001001000",
  5868=>"000000010",
  5869=>"101100100",
  5870=>"100101001",
  5871=>"111010101",
  5872=>"100011011",
  5873=>"100000111",
  5874=>"000001100",
  5875=>"011111001",
  5876=>"100011011",
  5877=>"111110110",
  5878=>"010111001",
  5879=>"001000011",
  5880=>"111101010",
  5881=>"110111110",
  5882=>"000011010",
  5883=>"001101010",
  5884=>"000101111",
  5885=>"110011110",
  5886=>"110100010",
  5887=>"100100111",
  5888=>"011000000",
  5889=>"000110000",
  5890=>"010100101",
  5891=>"010100001",
  5892=>"111101000",
  5893=>"001100100",
  5894=>"010111000",
  5895=>"111000101",
  5896=>"111100111",
  5897=>"010000001",
  5898=>"001010001",
  5899=>"000011111",
  5900=>"011011100",
  5901=>"110110010",
  5902=>"011000000",
  5903=>"001001101",
  5904=>"111110100",
  5905=>"011110000",
  5906=>"101101100",
  5907=>"000100111",
  5908=>"010101001",
  5909=>"111001100",
  5910=>"101111101",
  5911=>"001101001",
  5912=>"100100110",
  5913=>"010100011",
  5914=>"010111110",
  5915=>"000001110",
  5916=>"011001011",
  5917=>"001001101",
  5918=>"011001111",
  5919=>"000010011",
  5920=>"101101111",
  5921=>"000000000",
  5922=>"111110101",
  5923=>"000101000",
  5924=>"111111111",
  5925=>"100000111",
  5926=>"010111111",
  5927=>"010001001",
  5928=>"110111011",
  5929=>"010011010",
  5930=>"110101010",
  5931=>"011100001",
  5932=>"100011010",
  5933=>"011001111",
  5934=>"100010110",
  5935=>"111010111",
  5936=>"100000011",
  5937=>"110110011",
  5938=>"000100110",
  5939=>"100000011",
  5940=>"011000101",
  5941=>"110001101",
  5942=>"010001000",
  5943=>"101010010",
  5944=>"000000110",
  5945=>"110000111",
  5946=>"110111100",
  5947=>"010001100",
  5948=>"111000010",
  5949=>"001101101",
  5950=>"010101001",
  5951=>"000000100",
  5952=>"011100111",
  5953=>"100110111",
  5954=>"100000001",
  5955=>"001010000",
  5956=>"100011111",
  5957=>"001001011",
  5958=>"110010011",
  5959=>"001110010",
  5960=>"111110010",
  5961=>"001110101",
  5962=>"101011010",
  5963=>"011010000",
  5964=>"011001101",
  5965=>"111000101",
  5966=>"010100110",
  5967=>"111111111",
  5968=>"101001011",
  5969=>"001011101",
  5970=>"010010011",
  5971=>"101110000",
  5972=>"101010010",
  5973=>"111111011",
  5974=>"010101100",
  5975=>"111011010",
  5976=>"011100001",
  5977=>"110110011",
  5978=>"101000001",
  5979=>"000001001",
  5980=>"000001110",
  5981=>"110101111",
  5982=>"110001010",
  5983=>"010111010",
  5984=>"100000111",
  5985=>"000100111",
  5986=>"111101100",
  5987=>"000100011",
  5988=>"011100000",
  5989=>"001001001",
  5990=>"000010000",
  5991=>"111101001",
  5992=>"001100010",
  5993=>"001011010",
  5994=>"101101111",
  5995=>"001010000",
  5996=>"011101011",
  5997=>"110001001",
  5998=>"111000011",
  5999=>"010100010",
  6000=>"011010100",
  6001=>"101101110",
  6002=>"001010111",
  6003=>"100000010",
  6004=>"110001011",
  6005=>"101111000",
  6006=>"011001010",
  6007=>"010011000",
  6008=>"001000001",
  6009=>"011101000",
  6010=>"100111010",
  6011=>"111000011",
  6012=>"010011111",
  6013=>"011110110",
  6014=>"110011010",
  6015=>"101101100",
  6016=>"101011011",
  6017=>"111111000",
  6018=>"100100100",
  6019=>"101110100",
  6020=>"111011111",
  6021=>"011000101",
  6022=>"101001001",
  6023=>"001001000",
  6024=>"001100100",
  6025=>"000100101",
  6026=>"100011001",
  6027=>"010000001",
  6028=>"111101010",
  6029=>"010001011",
  6030=>"100000010",
  6031=>"101101011",
  6032=>"100000110",
  6033=>"100010111",
  6034=>"100111101",
  6035=>"111011011",
  6036=>"000101000",
  6037=>"100011110",
  6038=>"100010111",
  6039=>"111010110",
  6040=>"010100010",
  6041=>"000010101",
  6042=>"111110010",
  6043=>"000111110",
  6044=>"110000010",
  6045=>"000000011",
  6046=>"000000001",
  6047=>"001101100",
  6048=>"000111001",
  6049=>"001011100",
  6050=>"111110000",
  6051=>"001011001",
  6052=>"011100101",
  6053=>"110110111",
  6054=>"101100001",
  6055=>"111010010",
  6056=>"110001110",
  6057=>"100001011",
  6058=>"001001111",
  6059=>"110011000",
  6060=>"010101011",
  6061=>"110001010",
  6062=>"111000110",
  6063=>"110100011",
  6064=>"111010110",
  6065=>"110111000",
  6066=>"011111010",
  6067=>"010101000",
  6068=>"000110010",
  6069=>"110110111",
  6070=>"110111110",
  6071=>"101010110",
  6072=>"111100000",
  6073=>"001010101",
  6074=>"000110101",
  6075=>"110101100",
  6076=>"100100100",
  6077=>"001101001",
  6078=>"011100101",
  6079=>"111111000",
  6080=>"101011100",
  6081=>"101010101",
  6082=>"001101110",
  6083=>"001100011",
  6084=>"110101101",
  6085=>"000111100",
  6086=>"111001011",
  6087=>"110011001",
  6088=>"100000111",
  6089=>"111011000",
  6090=>"101111000",
  6091=>"111111111",
  6092=>"100110000",
  6093=>"010101101",
  6094=>"000101111",
  6095=>"010101000",
  6096=>"111000010",
  6097=>"000111010",
  6098=>"001100100",
  6099=>"010100100",
  6100=>"000110001",
  6101=>"100110101",
  6102=>"000110111",
  6103=>"010001111",
  6104=>"110101101",
  6105=>"011010000",
  6106=>"000101011",
  6107=>"100111000",
  6108=>"011110111",
  6109=>"101000000",
  6110=>"010110001",
  6111=>"101000110",
  6112=>"100101110",
  6113=>"111011010",
  6114=>"010010010",
  6115=>"110011101",
  6116=>"000110100",
  6117=>"011010001",
  6118=>"001110000",
  6119=>"111101001",
  6120=>"010010000",
  6121=>"100100010",
  6122=>"110010100",
  6123=>"100010100",
  6124=>"010001001",
  6125=>"011011010",
  6126=>"011101000",
  6127=>"101100001",
  6128=>"000011110",
  6129=>"100111000",
  6130=>"010011101",
  6131=>"110010110",
  6132=>"111000100",
  6133=>"111111110",
  6134=>"000001001",
  6135=>"100110100",
  6136=>"011001011",
  6137=>"111100000",
  6138=>"011001001",
  6139=>"111010100",
  6140=>"101110111",
  6141=>"001100001",
  6142=>"001111010",
  6143=>"101011001",
  6144=>"110001000",
  6145=>"111111011",
  6146=>"100101101",
  6147=>"100011101",
  6148=>"001010100",
  6149=>"110011111",
  6150=>"011100110",
  6151=>"100000101",
  6152=>"001011101",
  6153=>"111010011",
  6154=>"111111100",
  6155=>"111110100",
  6156=>"000101001",
  6157=>"111110100",
  6158=>"110111111",
  6159=>"111110110",
  6160=>"000000111",
  6161=>"111101111",
  6162=>"111100010",
  6163=>"010110011",
  6164=>"100001011",
  6165=>"011011101",
  6166=>"100011010",
  6167=>"010001010",
  6168=>"000001000",
  6169=>"101000101",
  6170=>"101010101",
  6171=>"101111110",
  6172=>"100010110",
  6173=>"001101001",
  6174=>"101100010",
  6175=>"010110101",
  6176=>"001001100",
  6177=>"110101000",
  6178=>"100011011",
  6179=>"001001011",
  6180=>"011001101",
  6181=>"101000000",
  6182=>"011110101",
  6183=>"110011000",
  6184=>"100101100",
  6185=>"000001101",
  6186=>"110001111",
  6187=>"110111001",
  6188=>"011010110",
  6189=>"111111101",
  6190=>"110100011",
  6191=>"101011010",
  6192=>"010100001",
  6193=>"100101111",
  6194=>"001110111",
  6195=>"011100010",
  6196=>"001001001",
  6197=>"011101110",
  6198=>"100110010",
  6199=>"010101010",
  6200=>"000000100",
  6201=>"110011000",
  6202=>"000100000",
  6203=>"111100100",
  6204=>"100000001",
  6205=>"101000011",
  6206=>"101111111",
  6207=>"110001000",
  6208=>"011000010",
  6209=>"000100100",
  6210=>"111110011",
  6211=>"110000100",
  6212=>"000010111",
  6213=>"010001000",
  6214=>"001011101",
  6215=>"110000011",
  6216=>"001100010",
  6217=>"111001110",
  6218=>"000000010",
  6219=>"010100001",
  6220=>"000100101",
  6221=>"000011110",
  6222=>"101010010",
  6223=>"111101011",
  6224=>"110010101",
  6225=>"010110110",
  6226=>"110010100",
  6227=>"101011111",
  6228=>"101101110",
  6229=>"000100101",
  6230=>"111001011",
  6231=>"100000000",
  6232=>"101011011",
  6233=>"010000110",
  6234=>"100111100",
  6235=>"100011100",
  6236=>"001010001",
  6237=>"011111001",
  6238=>"111011001",
  6239=>"001000000",
  6240=>"100110001",
  6241=>"010000010",
  6242=>"111101111",
  6243=>"111001010",
  6244=>"111010101",
  6245=>"000001010",
  6246=>"010011011",
  6247=>"101010100",
  6248=>"010001001",
  6249=>"000000011",
  6250=>"001111111",
  6251=>"111001001",
  6252=>"000110011",
  6253=>"101111010",
  6254=>"000101100",
  6255=>"010011010",
  6256=>"111001000",
  6257=>"110011010",
  6258=>"000000111",
  6259=>"010000110",
  6260=>"110000001",
  6261=>"010010001",
  6262=>"110100010",
  6263=>"000010110",
  6264=>"100101011",
  6265=>"100111101",
  6266=>"110011000",
  6267=>"100000001",
  6268=>"100100110",
  6269=>"000001111",
  6270=>"000011110",
  6271=>"101001001",
  6272=>"001010101",
  6273=>"110010100",
  6274=>"110111011",
  6275=>"100100000",
  6276=>"000010000",
  6277=>"100010111",
  6278=>"110010001",
  6279=>"110001100",
  6280=>"001000111",
  6281=>"100001000",
  6282=>"001110000",
  6283=>"110000110",
  6284=>"110110000",
  6285=>"111011111",
  6286=>"011000000",
  6287=>"000001110",
  6288=>"110010101",
  6289=>"100001010",
  6290=>"000111001",
  6291=>"111011111",
  6292=>"111101111",
  6293=>"111100000",
  6294=>"010010110",
  6295=>"111010101",
  6296=>"000010001",
  6297=>"110100001",
  6298=>"000111111",
  6299=>"001101000",
  6300=>"101101011",
  6301=>"110110000",
  6302=>"011110011",
  6303=>"110011011",
  6304=>"011111011",
  6305=>"010011000",
  6306=>"101001010",
  6307=>"101101001",
  6308=>"100111010",
  6309=>"101010011",
  6310=>"100001011",
  6311=>"100100101",
  6312=>"101110101",
  6313=>"101111000",
  6314=>"101000100",
  6315=>"011100101",
  6316=>"110110110",
  6317=>"010011001",
  6318=>"101000001",
  6319=>"011111011",
  6320=>"000011100",
  6321=>"111001101",
  6322=>"011111011",
  6323=>"100010001",
  6324=>"000111101",
  6325=>"100000011",
  6326=>"000001101",
  6327=>"110100101",
  6328=>"000110101",
  6329=>"000100001",
  6330=>"011111000",
  6331=>"000011010",
  6332=>"010111101",
  6333=>"001101100",
  6334=>"101100111",
  6335=>"111110000",
  6336=>"101110110",
  6337=>"001111010",
  6338=>"111010110",
  6339=>"111110000",
  6340=>"111101111",
  6341=>"000100000",
  6342=>"111011001",
  6343=>"001111011",
  6344=>"001011001",
  6345=>"111111110",
  6346=>"101010010",
  6347=>"011100101",
  6348=>"010101100",
  6349=>"100010111",
  6350=>"010010010",
  6351=>"001000001",
  6352=>"100110100",
  6353=>"011100010",
  6354=>"111000111",
  6355=>"001001001",
  6356=>"001101001",
  6357=>"100010101",
  6358=>"010101000",
  6359=>"100110000",
  6360=>"011110010",
  6361=>"110001110",
  6362=>"100101110",
  6363=>"001101000",
  6364=>"111110111",
  6365=>"011101011",
  6366=>"101001001",
  6367=>"100101000",
  6368=>"010001111",
  6369=>"111011110",
  6370=>"110111100",
  6371=>"010100010",
  6372=>"110100001",
  6373=>"001101010",
  6374=>"011000101",
  6375=>"100001001",
  6376=>"011001110",
  6377=>"001100010",
  6378=>"111011111",
  6379=>"010001101",
  6380=>"110101110",
  6381=>"111000111",
  6382=>"101111101",
  6383=>"100000110",
  6384=>"111111000",
  6385=>"101010111",
  6386=>"000010100",
  6387=>"110101101",
  6388=>"001101001",
  6389=>"000011001",
  6390=>"001100111",
  6391=>"111001011",
  6392=>"111001101",
  6393=>"001111100",
  6394=>"101101101",
  6395=>"000001010",
  6396=>"000111110",
  6397=>"111111111",
  6398=>"000001010",
  6399=>"001000010",
  6400=>"011001111",
  6401=>"100111110",
  6402=>"101110110",
  6403=>"100011010",
  6404=>"010111000",
  6405=>"100111110",
  6406=>"100011010",
  6407=>"000001111",
  6408=>"011001101",
  6409=>"100101000",
  6410=>"010010100",
  6411=>"100011101",
  6412=>"101111011",
  6413=>"100101111",
  6414=>"011101011",
  6415=>"110110100",
  6416=>"100010010",
  6417=>"011110111",
  6418=>"110011010",
  6419=>"111101101",
  6420=>"000000000",
  6421=>"001111110",
  6422=>"110000101",
  6423=>"011000110",
  6424=>"110010010",
  6425=>"111011100",
  6426=>"000110100",
  6427=>"010011111",
  6428=>"011010001",
  6429=>"010011111",
  6430=>"011110100",
  6431=>"011011101",
  6432=>"011011101",
  6433=>"011100010",
  6434=>"110100110",
  6435=>"000000101",
  6436=>"110111010",
  6437=>"110101011",
  6438=>"000011101",
  6439=>"010100010",
  6440=>"101010010",
  6441=>"100110001",
  6442=>"000001100",
  6443=>"100000100",
  6444=>"010111100",
  6445=>"000111101",
  6446=>"100010000",
  6447=>"011100010",
  6448=>"110101001",
  6449=>"101110110",
  6450=>"000111001",
  6451=>"000000101",
  6452=>"001101101",
  6453=>"111101110",
  6454=>"101100001",
  6455=>"111001100",
  6456=>"000010010",
  6457=>"111010100",
  6458=>"001111100",
  6459=>"110100110",
  6460=>"110001010",
  6461=>"001110110",
  6462=>"100111100",
  6463=>"000000001",
  6464=>"110011110",
  6465=>"111100001",
  6466=>"010000100",
  6467=>"101010110",
  6468=>"010000000",
  6469=>"000000010",
  6470=>"010100111",
  6471=>"001110110",
  6472=>"101000101",
  6473=>"110011010",
  6474=>"101100011",
  6475=>"001101011",
  6476=>"000110000",
  6477=>"101011101",
  6478=>"100101010",
  6479=>"101111101",
  6480=>"001000101",
  6481=>"100000111",
  6482=>"111111100",
  6483=>"101000010",
  6484=>"011001010",
  6485=>"101001010",
  6486=>"110001011",
  6487=>"011100001",
  6488=>"010001101",
  6489=>"111010111",
  6490=>"010001010",
  6491=>"011010000",
  6492=>"001011000",
  6493=>"111001001",
  6494=>"000010111",
  6495=>"000110101",
  6496=>"001011011",
  6497=>"100100010",
  6498=>"010011001",
  6499=>"100111011",
  6500=>"010111011",
  6501=>"111010011",
  6502=>"010011000",
  6503=>"110010111",
  6504=>"011010111",
  6505=>"101001110",
  6506=>"100001001",
  6507=>"000010111",
  6508=>"000010101",
  6509=>"000111101",
  6510=>"100000111",
  6511=>"000101000",
  6512=>"000101001",
  6513=>"111100010",
  6514=>"100101000",
  6515=>"111011110",
  6516=>"010010001",
  6517=>"000000010",
  6518=>"010001111",
  6519=>"000110000",
  6520=>"100101000",
  6521=>"011011000",
  6522=>"010111011",
  6523=>"101110000",
  6524=>"011000110",
  6525=>"111010011",
  6526=>"110010100",
  6527=>"001001000",
  6528=>"101001101",
  6529=>"010000111",
  6530=>"010011000",
  6531=>"011000000",
  6532=>"001100001",
  6533=>"010011000",
  6534=>"100110000",
  6535=>"101011101",
  6536=>"100111110",
  6537=>"011110001",
  6538=>"011100000",
  6539=>"000101010",
  6540=>"100011000",
  6541=>"011010001",
  6542=>"110111011",
  6543=>"010001110",
  6544=>"011100010",
  6545=>"111000101",
  6546=>"001100111",
  6547=>"010110011",
  6548=>"110110001",
  6549=>"011010111",
  6550=>"100011101",
  6551=>"010111001",
  6552=>"011001101",
  6553=>"110110110",
  6554=>"111011101",
  6555=>"110001101",
  6556=>"011011100",
  6557=>"000001000",
  6558=>"001110110",
  6559=>"110000010",
  6560=>"000001011",
  6561=>"010100111",
  6562=>"111010000",
  6563=>"001110010",
  6564=>"001001111",
  6565=>"100101001",
  6566=>"110011110",
  6567=>"010001001",
  6568=>"110011010",
  6569=>"001011000",
  6570=>"001111101",
  6571=>"001011110",
  6572=>"101101011",
  6573=>"011000110",
  6574=>"010000100",
  6575=>"010011110",
  6576=>"101100111",
  6577=>"001010010",
  6578=>"111011000",
  6579=>"101011110",
  6580=>"001100100",
  6581=>"010101001",
  6582=>"111010111",
  6583=>"100011111",
  6584=>"001010101",
  6585=>"101111010",
  6586=>"001000110",
  6587=>"001100101",
  6588=>"001010100",
  6589=>"001010001",
  6590=>"010100100",
  6591=>"010110111",
  6592=>"111010010",
  6593=>"100110111",
  6594=>"101000010",
  6595=>"110001111",
  6596=>"000010110",
  6597=>"100011101",
  6598=>"001000101",
  6599=>"101000001",
  6600=>"101111010",
  6601=>"001010001",
  6602=>"111110111",
  6603=>"100100001",
  6604=>"111011001",
  6605=>"101001111",
  6606=>"001111111",
  6607=>"111100000",
  6608=>"010101001",
  6609=>"100101111",
  6610=>"011001100",
  6611=>"011010110",
  6612=>"000110010",
  6613=>"101111111",
  6614=>"101110000",
  6615=>"111101011",
  6616=>"011111101",
  6617=>"010111110",
  6618=>"001111111",
  6619=>"011000111",
  6620=>"101011001",
  6621=>"110000010",
  6622=>"100110010",
  6623=>"110101100",
  6624=>"000000010",
  6625=>"110011100",
  6626=>"111010101",
  6627=>"010001101",
  6628=>"110000111",
  6629=>"010001010",
  6630=>"101001111",
  6631=>"000000001",
  6632=>"100000000",
  6633=>"000100111",
  6634=>"000010100",
  6635=>"111011100",
  6636=>"010101100",
  6637=>"011110000",
  6638=>"110100110",
  6639=>"010110000",
  6640=>"101100100",
  6641=>"100011010",
  6642=>"101111000",
  6643=>"011111110",
  6644=>"100100101",
  6645=>"111101110",
  6646=>"000111110",
  6647=>"101110100",
  6648=>"100111001",
  6649=>"101111111",
  6650=>"111010111",
  6651=>"000000111",
  6652=>"000111110",
  6653=>"101101100",
  6654=>"101100100",
  6655=>"110100000",
  6656=>"010001001",
  6657=>"101000110",
  6658=>"000000000",
  6659=>"010010000",
  6660=>"111111110",
  6661=>"111111111",
  6662=>"110000111",
  6663=>"110010111",
  6664=>"101100110",
  6665=>"101110000",
  6666=>"000000001",
  6667=>"111011001",
  6668=>"011100000",
  6669=>"000111010",
  6670=>"000010101",
  6671=>"001011010",
  6672=>"000011111",
  6673=>"011011111",
  6674=>"001110110",
  6675=>"001000111",
  6676=>"100011001",
  6677=>"110001010",
  6678=>"110100101",
  6679=>"000101010",
  6680=>"111110011",
  6681=>"101000101",
  6682=>"001100010",
  6683=>"011011000",
  6684=>"110101011",
  6685=>"111011101",
  6686=>"001001010",
  6687=>"111011010",
  6688=>"111000000",
  6689=>"001001110",
  6690=>"000111100",
  6691=>"001100111",
  6692=>"110011101",
  6693=>"111101100",
  6694=>"011101110",
  6695=>"001101100",
  6696=>"000010111",
  6697=>"001101000",
  6698=>"111110010",
  6699=>"110010000",
  6700=>"111000111",
  6701=>"001011001",
  6702=>"010010100",
  6703=>"110101100",
  6704=>"101110000",
  6705=>"001111000",
  6706=>"011010000",
  6707=>"000001010",
  6708=>"010100110",
  6709=>"010110100",
  6710=>"011110110",
  6711=>"011001101",
  6712=>"001110010",
  6713=>"100101110",
  6714=>"110101100",
  6715=>"000001000",
  6716=>"001110011",
  6717=>"000010110",
  6718=>"001111000",
  6719=>"101011111",
  6720=>"101101110",
  6721=>"101001111",
  6722=>"100000100",
  6723=>"100000110",
  6724=>"011101100",
  6725=>"000010010",
  6726=>"111111001",
  6727=>"010001011",
  6728=>"100010000",
  6729=>"000110111",
  6730=>"010100001",
  6731=>"100101101",
  6732=>"111100100",
  6733=>"010010110",
  6734=>"010001100",
  6735=>"001010010",
  6736=>"101100110",
  6737=>"111001000",
  6738=>"111000111",
  6739=>"111000110",
  6740=>"100110111",
  6741=>"111001011",
  6742=>"000000100",
  6743=>"000100101",
  6744=>"011100011",
  6745=>"010101001",
  6746=>"100000010",
  6747=>"111000011",
  6748=>"110110100",
  6749=>"111011010",
  6750=>"100110000",
  6751=>"100011101",
  6752=>"100110111",
  6753=>"100110110",
  6754=>"110011010",
  6755=>"101101000",
  6756=>"010100000",
  6757=>"001111100",
  6758=>"100011111",
  6759=>"110111110",
  6760=>"011001111",
  6761=>"011001101",
  6762=>"001100010",
  6763=>"011110011",
  6764=>"000001100",
  6765=>"101101001",
  6766=>"000001010",
  6767=>"110010010",
  6768=>"111001001",
  6769=>"000110001",
  6770=>"011101000",
  6771=>"010011110",
  6772=>"000000000",
  6773=>"010011100",
  6774=>"000011110",
  6775=>"110010110",
  6776=>"011010011",
  6777=>"011011111",
  6778=>"110001000",
  6779=>"000100001",
  6780=>"010001000",
  6781=>"101101001",
  6782=>"101010100",
  6783=>"101001101",
  6784=>"011101101",
  6785=>"000001010",
  6786=>"001001000",
  6787=>"101111010",
  6788=>"001011000",
  6789=>"101000010",
  6790=>"101101111",
  6791=>"110111011",
  6792=>"001000010",
  6793=>"000110011",
  6794=>"011101011",
  6795=>"010111100",
  6796=>"110011110",
  6797=>"010001111",
  6798=>"111010100",
  6799=>"110001011",
  6800=>"110110110",
  6801=>"110001110",
  6802=>"111101010",
  6803=>"011101000",
  6804=>"010100100",
  6805=>"110111001",
  6806=>"110110100",
  6807=>"010000111",
  6808=>"110010001",
  6809=>"011100000",
  6810=>"010100100",
  6811=>"000100001",
  6812=>"000101110",
  6813=>"000000110",
  6814=>"111000100",
  6815=>"001101111",
  6816=>"101001110",
  6817=>"000010000",
  6818=>"010110011",
  6819=>"011000010",
  6820=>"010010100",
  6821=>"100110000",
  6822=>"111000000",
  6823=>"110010000",
  6824=>"101010011",
  6825=>"110100110",
  6826=>"001101000",
  6827=>"111011100",
  6828=>"000010011",
  6829=>"101101100",
  6830=>"000100001",
  6831=>"001101000",
  6832=>"001010100",
  6833=>"101100010",
  6834=>"000000100",
  6835=>"001011011",
  6836=>"000100010",
  6837=>"000000111",
  6838=>"001110011",
  6839=>"010101011",
  6840=>"001101010",
  6841=>"010001010",
  6842=>"010100010",
  6843=>"000000001",
  6844=>"111011101",
  6845=>"010010110",
  6846=>"000100001",
  6847=>"110011110",
  6848=>"111010101",
  6849=>"111011001",
  6850=>"100111111",
  6851=>"100101010",
  6852=>"001001100",
  6853=>"001000111",
  6854=>"101101010",
  6855=>"110010001",
  6856=>"101010100",
  6857=>"111101001",
  6858=>"000110101",
  6859=>"000000001",
  6860=>"001011110",
  6861=>"110101011",
  6862=>"001000010",
  6863=>"111111111",
  6864=>"010010010",
  6865=>"111100000",
  6866=>"010101011",
  6867=>"011111110",
  6868=>"000001011",
  6869=>"000101100",
  6870=>"110011101",
  6871=>"000101100",
  6872=>"111110100",
  6873=>"101110111",
  6874=>"111100000",
  6875=>"111100100",
  6876=>"010100110",
  6877=>"000001011",
  6878=>"001001010",
  6879=>"010110000",
  6880=>"111110100",
  6881=>"110010000",
  6882=>"010100000",
  6883=>"001001111",
  6884=>"000010100",
  6885=>"011101111",
  6886=>"010011011",
  6887=>"110100010",
  6888=>"010010100",
  6889=>"001000010",
  6890=>"010111000",
  6891=>"001000100",
  6892=>"011011011",
  6893=>"101110101",
  6894=>"111100010",
  6895=>"111110011",
  6896=>"101110001",
  6897=>"100110110",
  6898=>"100001000",
  6899=>"010000000",
  6900=>"011000000",
  6901=>"011101110",
  6902=>"010101011",
  6903=>"110101100",
  6904=>"100110101",
  6905=>"111100101",
  6906=>"001010011",
  6907=>"111011111",
  6908=>"101011101",
  6909=>"010100000",
  6910=>"000100001",
  6911=>"010100111",
  6912=>"010010010",
  6913=>"100101011",
  6914=>"010111110",
  6915=>"001101011",
  6916=>"010000100",
  6917=>"001001011",
  6918=>"110010011",
  6919=>"010011100",
  6920=>"110100100",
  6921=>"000100001",
  6922=>"000010000",
  6923=>"011110110",
  6924=>"101011110",
  6925=>"110100100",
  6926=>"010000111",
  6927=>"000101000",
  6928=>"001010100",
  6929=>"101000000",
  6930=>"100000100",
  6931=>"111000111",
  6932=>"000100111",
  6933=>"000110101",
  6934=>"100001000",
  6935=>"100111110",
  6936=>"101001011",
  6937=>"010011001",
  6938=>"001111100",
  6939=>"001001010",
  6940=>"000111010",
  6941=>"000101101",
  6942=>"110000110",
  6943=>"111010011",
  6944=>"101001110",
  6945=>"011101011",
  6946=>"001001001",
  6947=>"111011111",
  6948=>"101010101",
  6949=>"000000001",
  6950=>"101011100",
  6951=>"001010001",
  6952=>"011010110",
  6953=>"000111100",
  6954=>"000010000",
  6955=>"001111100",
  6956=>"010010010",
  6957=>"111011001",
  6958=>"000110000",
  6959=>"101100001",
  6960=>"010001011",
  6961=>"001101110",
  6962=>"011111110",
  6963=>"111101010",
  6964=>"011011011",
  6965=>"011000000",
  6966=>"001001001",
  6967=>"100100001",
  6968=>"001000011",
  6969=>"100101111",
  6970=>"100111110",
  6971=>"100111101",
  6972=>"011100101",
  6973=>"111111111",
  6974=>"000001000",
  6975=>"111111111",
  6976=>"101011101",
  6977=>"101011010",
  6978=>"100010001",
  6979=>"100011010",
  6980=>"110001100",
  6981=>"110010100",
  6982=>"101101010",
  6983=>"111001111",
  6984=>"010100011",
  6985=>"100011010",
  6986=>"111111011",
  6987=>"000011110",
  6988=>"101110000",
  6989=>"101100000",
  6990=>"110100110",
  6991=>"101101101",
  6992=>"101101110",
  6993=>"001100101",
  6994=>"000010110",
  6995=>"111100110",
  6996=>"000001001",
  6997=>"010110011",
  6998=>"011010101",
  6999=>"010011011",
  7000=>"100101111",
  7001=>"110100101",
  7002=>"100100110",
  7003=>"010110011",
  7004=>"010101101",
  7005=>"010110111",
  7006=>"101001111",
  7007=>"000101010",
  7008=>"010110111",
  7009=>"011111110",
  7010=>"000111111",
  7011=>"111110100",
  7012=>"001110011",
  7013=>"101001000",
  7014=>"101100001",
  7015=>"100101000",
  7016=>"110001101",
  7017=>"010000101",
  7018=>"001010110",
  7019=>"011110010",
  7020=>"101100101",
  7021=>"111000001",
  7022=>"000110001",
  7023=>"001100010",
  7024=>"100110000",
  7025=>"111011110",
  7026=>"011000110",
  7027=>"001000110",
  7028=>"010100111",
  7029=>"000110101",
  7030=>"011101111",
  7031=>"111100001",
  7032=>"011010111",
  7033=>"011111000",
  7034=>"011100011",
  7035=>"101000010",
  7036=>"000001001",
  7037=>"001000100",
  7038=>"111111000",
  7039=>"001101111",
  7040=>"111111111",
  7041=>"110110101",
  7042=>"111101010",
  7043=>"011111010",
  7044=>"010100011",
  7045=>"111001001",
  7046=>"100001001",
  7047=>"001010101",
  7048=>"111001000",
  7049=>"000101110",
  7050=>"100001110",
  7051=>"000100000",
  7052=>"001100110",
  7053=>"000010000",
  7054=>"111000110",
  7055=>"110011101",
  7056=>"110001101",
  7057=>"111011111",
  7058=>"101000111",
  7059=>"010001010",
  7060=>"000100000",
  7061=>"001101111",
  7062=>"100101100",
  7063=>"110101011",
  7064=>"111111110",
  7065=>"000000110",
  7066=>"111111011",
  7067=>"101110011",
  7068=>"011101000",
  7069=>"101011110",
  7070=>"011101101",
  7071=>"101111001",
  7072=>"100000000",
  7073=>"011001000",
  7074=>"010011011",
  7075=>"111111111",
  7076=>"000000010",
  7077=>"111110001",
  7078=>"100101010",
  7079=>"111110000",
  7080=>"001011111",
  7081=>"001000000",
  7082=>"001100100",
  7083=>"100100110",
  7084=>"111100101",
  7085=>"111100110",
  7086=>"100000001",
  7087=>"110001001",
  7088=>"011011001",
  7089=>"101101100",
  7090=>"010100111",
  7091=>"111001010",
  7092=>"111101001",
  7093=>"011010000",
  7094=>"101010101",
  7095=>"000100011",
  7096=>"111110100",
  7097=>"011000100",
  7098=>"000011001",
  7099=>"010010101",
  7100=>"010001000",
  7101=>"111111111",
  7102=>"011001111",
  7103=>"001001011",
  7104=>"010010101",
  7105=>"001001001",
  7106=>"110001111",
  7107=>"010001001",
  7108=>"010000101",
  7109=>"000001101",
  7110=>"011101000",
  7111=>"100110101",
  7112=>"100000001",
  7113=>"011001011",
  7114=>"100010100",
  7115=>"001111001",
  7116=>"011000101",
  7117=>"010010000",
  7118=>"001000000",
  7119=>"000000000",
  7120=>"101101010",
  7121=>"001001011",
  7122=>"111111001",
  7123=>"001101100",
  7124=>"001000000",
  7125=>"111101110",
  7126=>"011000000",
  7127=>"110111100",
  7128=>"110001101",
  7129=>"011011110",
  7130=>"011100110",
  7131=>"111111010",
  7132=>"110110001",
  7133=>"000001110",
  7134=>"001111010",
  7135=>"010011001",
  7136=>"111001111",
  7137=>"100111101",
  7138=>"010111100",
  7139=>"111001010",
  7140=>"111100000",
  7141=>"011101011",
  7142=>"011100011",
  7143=>"001010010",
  7144=>"101111100",
  7145=>"010111110",
  7146=>"010100110",
  7147=>"011000101",
  7148=>"010001011",
  7149=>"010110110",
  7150=>"100011011",
  7151=>"010101000",
  7152=>"111101010",
  7153=>"011110111",
  7154=>"010111110",
  7155=>"111111101",
  7156=>"001110111",
  7157=>"100011111",
  7158=>"100111010",
  7159=>"001010101",
  7160=>"011101001",
  7161=>"010101100",
  7162=>"101010101",
  7163=>"001100000",
  7164=>"000000011",
  7165=>"110010010",
  7166=>"010110010",
  7167=>"000111011",
  7168=>"101000000",
  7169=>"101101101",
  7170=>"000110011",
  7171=>"111111001",
  7172=>"111000001",
  7173=>"100011000",
  7174=>"101001110",
  7175=>"000000001",
  7176=>"101110001",
  7177=>"101010001",
  7178=>"001110010",
  7179=>"001110110",
  7180=>"100100110",
  7181=>"001101110",
  7182=>"110000110",
  7183=>"111101110",
  7184=>"000000101",
  7185=>"011101111",
  7186=>"101000100",
  7187=>"110001010",
  7188=>"111001110",
  7189=>"111001111",
  7190=>"000000101",
  7191=>"101011011",
  7192=>"111010010",
  7193=>"110010100",
  7194=>"000001000",
  7195=>"000000101",
  7196=>"011101101",
  7197=>"000000011",
  7198=>"110101010",
  7199=>"111110111",
  7200=>"011000001",
  7201=>"110000001",
  7202=>"111011101",
  7203=>"001110110",
  7204=>"101011101",
  7205=>"110010111",
  7206=>"110101000",
  7207=>"010100111",
  7208=>"001000110",
  7209=>"100000110",
  7210=>"010110101",
  7211=>"001011010",
  7212=>"000000000",
  7213=>"101101010",
  7214=>"010100011",
  7215=>"111000010",
  7216=>"001111011",
  7217=>"101101001",
  7218=>"110110000",
  7219=>"000100010",
  7220=>"111101010",
  7221=>"111000000",
  7222=>"010001010",
  7223=>"000000001",
  7224=>"000000100",
  7225=>"101001110",
  7226=>"101010010",
  7227=>"101100001",
  7228=>"101000000",
  7229=>"110101110",
  7230=>"000010000",
  7231=>"011010001",
  7232=>"001111110",
  7233=>"001001101",
  7234=>"110000001",
  7235=>"101000010",
  7236=>"011010000",
  7237=>"100100100",
  7238=>"011101100",
  7239=>"000000011",
  7240=>"110110100",
  7241=>"101011111",
  7242=>"000100000",
  7243=>"011001001",
  7244=>"110100000",
  7245=>"100101000",
  7246=>"101110101",
  7247=>"101001011",
  7248=>"100100101",
  7249=>"100111111",
  7250=>"000010110",
  7251=>"001010111",
  7252=>"001010000",
  7253=>"111011111",
  7254=>"110110100",
  7255=>"001100101",
  7256=>"110101111",
  7257=>"101000000",
  7258=>"100000001",
  7259=>"011000001",
  7260=>"110110011",
  7261=>"101101100",
  7262=>"010101100",
  7263=>"000100101",
  7264=>"010101011",
  7265=>"110100100",
  7266=>"110100011",
  7267=>"010011010",
  7268=>"000011101",
  7269=>"100100000",
  7270=>"001011010",
  7271=>"100000010",
  7272=>"001011011",
  7273=>"001010010",
  7274=>"110000111",
  7275=>"110100000",
  7276=>"101101110",
  7277=>"111011010",
  7278=>"001011111",
  7279=>"110110101",
  7280=>"110001000",
  7281=>"110000000",
  7282=>"111111110",
  7283=>"000101100",
  7284=>"010101000",
  7285=>"111100100",
  7286=>"001100001",
  7287=>"011100101",
  7288=>"101110001",
  7289=>"111111001",
  7290=>"001111001",
  7291=>"111000011",
  7292=>"010101110",
  7293=>"111101010",
  7294=>"100110100",
  7295=>"100000000",
  7296=>"010000100",
  7297=>"110110010",
  7298=>"001101010",
  7299=>"001001000",
  7300=>"011101100",
  7301=>"011100001",
  7302=>"000111111",
  7303=>"100111000",
  7304=>"011000010",
  7305=>"110011101",
  7306=>"101011000",
  7307=>"001000111",
  7308=>"100011101",
  7309=>"111001110",
  7310=>"100110010",
  7311=>"101001011",
  7312=>"001010101",
  7313=>"000111110",
  7314=>"111000110",
  7315=>"100000100",
  7316=>"000000100",
  7317=>"011001010",
  7318=>"101000000",
  7319=>"001011110",
  7320=>"000110101",
  7321=>"000001000",
  7322=>"010111000",
  7323=>"000111111",
  7324=>"011100000",
  7325=>"110100110",
  7326=>"000111000",
  7327=>"111011101",
  7328=>"100001101",
  7329=>"011010110",
  7330=>"010101000",
  7331=>"000001000",
  7332=>"000101111",
  7333=>"000010111",
  7334=>"110100000",
  7335=>"110110111",
  7336=>"101001100",
  7337=>"000111110",
  7338=>"101110101",
  7339=>"110001100",
  7340=>"101001010",
  7341=>"100010110",
  7342=>"100101100",
  7343=>"101100000",
  7344=>"000100101",
  7345=>"010011010",
  7346=>"011001110",
  7347=>"100001111",
  7348=>"111110001",
  7349=>"011011100",
  7350=>"101101001",
  7351=>"101001011",
  7352=>"011000001",
  7353=>"100110010",
  7354=>"111111111",
  7355=>"101011101",
  7356=>"101110100",
  7357=>"111001101",
  7358=>"001001100",
  7359=>"000101101",
  7360=>"100000101",
  7361=>"111101000",
  7362=>"111000010",
  7363=>"110111000",
  7364=>"001100110",
  7365=>"101111111",
  7366=>"000111010",
  7367=>"110101110",
  7368=>"110000110",
  7369=>"001011001",
  7370=>"011001101",
  7371=>"111000000",
  7372=>"011010000",
  7373=>"011000100",
  7374=>"000101000",
  7375=>"100111101",
  7376=>"011011111",
  7377=>"010001111",
  7378=>"101100010",
  7379=>"110011101",
  7380=>"011010000",
  7381=>"000111111",
  7382=>"101011010",
  7383=>"010100111",
  7384=>"100000100",
  7385=>"111011011",
  7386=>"001100011",
  7387=>"000000110",
  7388=>"100110101",
  7389=>"100010111",
  7390=>"001110110",
  7391=>"110001101",
  7392=>"101011101",
  7393=>"001101110",
  7394=>"110011000",
  7395=>"111001111",
  7396=>"111111011",
  7397=>"001101000",
  7398=>"111010110",
  7399=>"010010110",
  7400=>"100100101",
  7401=>"000101000",
  7402=>"010100100",
  7403=>"010101100",
  7404=>"010011001",
  7405=>"001111101",
  7406=>"001001100",
  7407=>"100110011",
  7408=>"000001010",
  7409=>"111011010",
  7410=>"011101001",
  7411=>"000011010",
  7412=>"000111001",
  7413=>"011100111",
  7414=>"011010100",
  7415=>"111000001",
  7416=>"010000110",
  7417=>"010111101",
  7418=>"111111111",
  7419=>"100101011",
  7420=>"101111101",
  7421=>"111011000",
  7422=>"000010010",
  7423=>"001011101",
  7424=>"101101110",
  7425=>"011011111",
  7426=>"010010110",
  7427=>"110011000",
  7428=>"101100010",
  7429=>"000110111",
  7430=>"101101000",
  7431=>"001001110",
  7432=>"001001010",
  7433=>"101110010",
  7434=>"101011111",
  7435=>"111110100",
  7436=>"101111101",
  7437=>"111011101",
  7438=>"100110110",
  7439=>"000001101",
  7440=>"110010010",
  7441=>"110001100",
  7442=>"010000100",
  7443=>"101010001",
  7444=>"101001010",
  7445=>"000010011",
  7446=>"111111111",
  7447=>"101100100",
  7448=>"111110001",
  7449=>"101001010",
  7450=>"101100000",
  7451=>"111110100",
  7452=>"010101010",
  7453=>"011000000",
  7454=>"011111000",
  7455=>"100100001",
  7456=>"000000001",
  7457=>"101001110",
  7458=>"111110000",
  7459=>"000100010",
  7460=>"001110100",
  7461=>"010000111",
  7462=>"110000111",
  7463=>"110001111",
  7464=>"011101001",
  7465=>"101101101",
  7466=>"101000100",
  7467=>"000010110",
  7468=>"011000110",
  7469=>"101001011",
  7470=>"100011100",
  7471=>"110001110",
  7472=>"100000100",
  7473=>"110111010",
  7474=>"101101101",
  7475=>"101010000",
  7476=>"000110111",
  7477=>"011000011",
  7478=>"111110001",
  7479=>"010010101",
  7480=>"001000000",
  7481=>"100011011",
  7482=>"011010000",
  7483=>"001000111",
  7484=>"111100000",
  7485=>"111101010",
  7486=>"011001111",
  7487=>"111100000",
  7488=>"100100100",
  7489=>"001111000",
  7490=>"111110011",
  7491=>"011101100",
  7492=>"101000001",
  7493=>"000011011",
  7494=>"000011000",
  7495=>"101001000",
  7496=>"011011101",
  7497=>"000011010",
  7498=>"001101000",
  7499=>"010000111",
  7500=>"100000110",
  7501=>"100011001",
  7502=>"010010001",
  7503=>"100110101",
  7504=>"001111110",
  7505=>"111101000",
  7506=>"110100010",
  7507=>"100010100",
  7508=>"000000110",
  7509=>"000101010",
  7510=>"111100010",
  7511=>"111001000",
  7512=>"001100100",
  7513=>"101011111",
  7514=>"000001101",
  7515=>"110100111",
  7516=>"111110110",
  7517=>"111010100",
  7518=>"110000010",
  7519=>"011101101",
  7520=>"111100110",
  7521=>"010011100",
  7522=>"110110111",
  7523=>"011001100",
  7524=>"101000000",
  7525=>"000001001",
  7526=>"111110011",
  7527=>"111100100",
  7528=>"010010111",
  7529=>"101011000",
  7530=>"010011010",
  7531=>"001000110",
  7532=>"000110100",
  7533=>"011111010",
  7534=>"111100111",
  7535=>"000001000",
  7536=>"101111101",
  7537=>"000000100",
  7538=>"010110001",
  7539=>"110100001",
  7540=>"000100010",
  7541=>"110110100",
  7542=>"110001001",
  7543=>"111101110",
  7544=>"101011000",
  7545=>"100100111",
  7546=>"101111111",
  7547=>"001001000",
  7548=>"111001010",
  7549=>"010000110",
  7550=>"101101001",
  7551=>"010101000",
  7552=>"110101110",
  7553=>"000001110",
  7554=>"101110101",
  7555=>"110000001",
  7556=>"010101101",
  7557=>"001100011",
  7558=>"110011111",
  7559=>"100101100",
  7560=>"110001011",
  7561=>"011010011",
  7562=>"001011000",
  7563=>"000010000",
  7564=>"000110001",
  7565=>"001000000",
  7566=>"100000100",
  7567=>"110011011",
  7568=>"111100011",
  7569=>"011000010",
  7570=>"110001011",
  7571=>"000010011",
  7572=>"000100101",
  7573=>"101000001",
  7574=>"010000000",
  7575=>"111111001",
  7576=>"100011001",
  7577=>"100001010",
  7578=>"100111101",
  7579=>"000010001",
  7580=>"100111101",
  7581=>"111110001",
  7582=>"110010000",
  7583=>"000011101",
  7584=>"111001100",
  7585=>"100000111",
  7586=>"000010011",
  7587=>"010000000",
  7588=>"001010010",
  7589=>"001000000",
  7590=>"011000110",
  7591=>"100001001",
  7592=>"001011000",
  7593=>"001010001",
  7594=>"010000111",
  7595=>"111110100",
  7596=>"110101011",
  7597=>"110110101",
  7598=>"000110010",
  7599=>"111110100",
  7600=>"111000100",
  7601=>"111000110",
  7602=>"101011110",
  7603=>"000100011",
  7604=>"010000000",
  7605=>"001000001",
  7606=>"110101000",
  7607=>"000001011",
  7608=>"110100101",
  7609=>"111001110",
  7610=>"110000101",
  7611=>"011100010",
  7612=>"111011101",
  7613=>"111111111",
  7614=>"101101011",
  7615=>"010101001",
  7616=>"000011111",
  7617=>"000100110",
  7618=>"011001101",
  7619=>"110101100",
  7620=>"101001000",
  7621=>"101011100",
  7622=>"000011001",
  7623=>"000000001",
  7624=>"010001111",
  7625=>"101111111",
  7626=>"100101001",
  7627=>"110011110",
  7628=>"000001010",
  7629=>"010110010",
  7630=>"111101110",
  7631=>"110011001",
  7632=>"111010011",
  7633=>"001110100",
  7634=>"001001011",
  7635=>"010111011",
  7636=>"101111000",
  7637=>"100000011",
  7638=>"100100001",
  7639=>"111110110",
  7640=>"001010010",
  7641=>"000011010",
  7642=>"111111011",
  7643=>"100110100",
  7644=>"101010110",
  7645=>"001100010",
  7646=>"101010110",
  7647=>"110011010",
  7648=>"001010100",
  7649=>"111100110",
  7650=>"111001000",
  7651=>"100110110",
  7652=>"110100110",
  7653=>"100100100",
  7654=>"110101100",
  7655=>"000001011",
  7656=>"011100000",
  7657=>"001110011",
  7658=>"111010100",
  7659=>"100001000",
  7660=>"001101101",
  7661=>"000100010",
  7662=>"011111100",
  7663=>"100101011",
  7664=>"010000101",
  7665=>"100011001",
  7666=>"000111110",
  7667=>"010011000",
  7668=>"110110100",
  7669=>"100110100",
  7670=>"101111111",
  7671=>"100010000",
  7672=>"100101011",
  7673=>"111110001",
  7674=>"001111010",
  7675=>"000001001",
  7676=>"100001010",
  7677=>"000000100",
  7678=>"100011011",
  7679=>"111011100",
  7680=>"011110101",
  7681=>"001110101",
  7682=>"011100110",
  7683=>"000000010",
  7684=>"000111100",
  7685=>"001100000",
  7686=>"110011101",
  7687=>"111101011",
  7688=>"111011110",
  7689=>"000111101",
  7690=>"110111011",
  7691=>"010010010",
  7692=>"010010001",
  7693=>"101111100",
  7694=>"000011101",
  7695=>"011010100",
  7696=>"100100110",
  7697=>"011110111",
  7698=>"100011000",
  7699=>"101111100",
  7700=>"000001000",
  7701=>"000001011",
  7702=>"110000110",
  7703=>"111011010",
  7704=>"100010000",
  7705=>"001101111",
  7706=>"011010111",
  7707=>"011011111",
  7708=>"101000000",
  7709=>"111110110",
  7710=>"001111000",
  7711=>"010010011",
  7712=>"000100011",
  7713=>"110111001",
  7714=>"011010101",
  7715=>"111111111",
  7716=>"001011110",
  7717=>"101001011",
  7718=>"100001001",
  7719=>"110100000",
  7720=>"011011001",
  7721=>"001110101",
  7722=>"000100011",
  7723=>"001101010",
  7724=>"001001110",
  7725=>"001001001",
  7726=>"001101110",
  7727=>"100100100",
  7728=>"010111001",
  7729=>"010111111",
  7730=>"011011110",
  7731=>"101011001",
  7732=>"001100110",
  7733=>"110101010",
  7734=>"110010111",
  7735=>"001000001",
  7736=>"100110001",
  7737=>"110000101",
  7738=>"000110111",
  7739=>"110101100",
  7740=>"000110100",
  7741=>"100011100",
  7742=>"100010100",
  7743=>"000111000",
  7744=>"111110011",
  7745=>"100000100",
  7746=>"100001111",
  7747=>"000111001",
  7748=>"011000010",
  7749=>"010111000",
  7750=>"000100000",
  7751=>"100110111",
  7752=>"101110100",
  7753=>"000010011",
  7754=>"110011111",
  7755=>"100000011",
  7756=>"110111000",
  7757=>"100001111",
  7758=>"000001011",
  7759=>"101010011",
  7760=>"001111100",
  7761=>"111000100",
  7762=>"010100001",
  7763=>"001001011",
  7764=>"001011001",
  7765=>"010000011",
  7766=>"001000010",
  7767=>"101001010",
  7768=>"111111111",
  7769=>"100010100",
  7770=>"001011100",
  7771=>"100001100",
  7772=>"000110000",
  7773=>"100100010",
  7774=>"001000111",
  7775=>"010110010",
  7776=>"100111000",
  7777=>"110011011",
  7778=>"000101111",
  7779=>"111001001",
  7780=>"011000010",
  7781=>"001001111",
  7782=>"100100001",
  7783=>"110001110",
  7784=>"011010000",
  7785=>"111111111",
  7786=>"001000010",
  7787=>"001000000",
  7788=>"100001110",
  7789=>"101111010",
  7790=>"011000110",
  7791=>"100001101",
  7792=>"011010001",
  7793=>"011010000",
  7794=>"110111011",
  7795=>"101000010",
  7796=>"001000010",
  7797=>"000000011",
  7798=>"011111100",
  7799=>"000010111",
  7800=>"000011111",
  7801=>"101100000",
  7802=>"011111100",
  7803=>"110000110",
  7804=>"101000100",
  7805=>"010010101",
  7806=>"111111101",
  7807=>"010101001",
  7808=>"100101010",
  7809=>"111001011",
  7810=>"011101010",
  7811=>"001001000",
  7812=>"110011011",
  7813=>"100100000",
  7814=>"000000110",
  7815=>"011001010",
  7816=>"011101000",
  7817=>"100001010",
  7818=>"101111101",
  7819=>"011000011",
  7820=>"000001000",
  7821=>"000000010",
  7822=>"100100010",
  7823=>"110111101",
  7824=>"011110110",
  7825=>"011100111",
  7826=>"100010000",
  7827=>"100011101",
  7828=>"100110100",
  7829=>"011111001",
  7830=>"001010101",
  7831=>"100010011",
  7832=>"111011111",
  7833=>"111010000",
  7834=>"000010010",
  7835=>"101111100",
  7836=>"000011111",
  7837=>"111101001",
  7838=>"010111111",
  7839=>"001101000",
  7840=>"000000000",
  7841=>"111000111",
  7842=>"100011010",
  7843=>"101010011",
  7844=>"111111101",
  7845=>"001110010",
  7846=>"001011000",
  7847=>"101000010",
  7848=>"010010010",
  7849=>"010100010",
  7850=>"010000001",
  7851=>"011010000",
  7852=>"011110101",
  7853=>"110110000",
  7854=>"111011110",
  7855=>"000011110",
  7856=>"000001101",
  7857=>"000010101",
  7858=>"100101110",
  7859=>"010001111",
  7860=>"100011110",
  7861=>"111100010",
  7862=>"111010001",
  7863=>"010010010",
  7864=>"111011001",
  7865=>"111101110",
  7866=>"001101000",
  7867=>"000110110",
  7868=>"001010001",
  7869=>"100110011",
  7870=>"101000111",
  7871=>"101011110",
  7872=>"101010000",
  7873=>"100011001",
  7874=>"011010111",
  7875=>"111001010",
  7876=>"101001011",
  7877=>"000001110",
  7878=>"010001010",
  7879=>"101011010",
  7880=>"110010001",
  7881=>"110001100",
  7882=>"001101110",
  7883=>"100100010",
  7884=>"010010000",
  7885=>"011001011",
  7886=>"001111101",
  7887=>"010000100",
  7888=>"100001110",
  7889=>"011000110",
  7890=>"111010100",
  7891=>"010011011",
  7892=>"000010010",
  7893=>"110000011",
  7894=>"010101001",
  7895=>"011111001",
  7896=>"100000101",
  7897=>"111101111",
  7898=>"111011100",
  7899=>"111110000",
  7900=>"101101101",
  7901=>"010100010",
  7902=>"011111100",
  7903=>"000000111",
  7904=>"001100011",
  7905=>"101110110",
  7906=>"111011111",
  7907=>"111010111",
  7908=>"100101001",
  7909=>"111100001",
  7910=>"000110100",
  7911=>"010101011",
  7912=>"101111011",
  7913=>"000100000",
  7914=>"000100101",
  7915=>"001001011",
  7916=>"101001011",
  7917=>"001111101",
  7918=>"001110010",
  7919=>"001011111",
  7920=>"010000111",
  7921=>"010110111",
  7922=>"001111111",
  7923=>"000110110",
  7924=>"100001101",
  7925=>"101101010",
  7926=>"100000111",
  7927=>"100001000",
  7928=>"011011100",
  7929=>"101010000",
  7930=>"110011100",
  7931=>"010110101",
  7932=>"100111100",
  7933=>"000000100",
  7934=>"001110100",
  7935=>"100010010",
  7936=>"010101011",
  7937=>"001111011",
  7938=>"101101000",
  7939=>"111110100",
  7940=>"101110010",
  7941=>"100011111",
  7942=>"111001110",
  7943=>"000001000",
  7944=>"110100010",
  7945=>"010011110",
  7946=>"111000110",
  7947=>"001111011",
  7948=>"111001000",
  7949=>"000011010",
  7950=>"100010110",
  7951=>"111011011",
  7952=>"010000000",
  7953=>"010001000",
  7954=>"110110000",
  7955=>"100011101",
  7956=>"010010100",
  7957=>"110011000",
  7958=>"011000011",
  7959=>"011101011",
  7960=>"111101101",
  7961=>"010101000",
  7962=>"001000001",
  7963=>"111010111",
  7964=>"011010110",
  7965=>"111101111",
  7966=>"010001101",
  7967=>"010101111",
  7968=>"000100011",
  7969=>"111100101",
  7970=>"111101101",
  7971=>"111011001",
  7972=>"111011001",
  7973=>"100101111",
  7974=>"101101000",
  7975=>"011110111",
  7976=>"011101010",
  7977=>"000001100",
  7978=>"000110001",
  7979=>"010100110",
  7980=>"000110111",
  7981=>"101100011",
  7982=>"100000010",
  7983=>"100100100",
  7984=>"001010110",
  7985=>"010110101",
  7986=>"000001011",
  7987=>"111100101",
  7988=>"001001000",
  7989=>"100101001",
  7990=>"111011001",
  7991=>"100000001",
  7992=>"101111110",
  7993=>"000000111",
  7994=>"001011100",
  7995=>"101011001",
  7996=>"110111000",
  7997=>"001100111",
  7998=>"100110100",
  7999=>"001100000",
  8000=>"111010111",
  8001=>"011111011",
  8002=>"000100010",
  8003=>"110001111",
  8004=>"101101110",
  8005=>"011000011",
  8006=>"100100001",
  8007=>"010001101",
  8008=>"110101111",
  8009=>"011000100",
  8010=>"100111010",
  8011=>"000110110",
  8012=>"101001011",
  8013=>"001000110",
  8014=>"100001101",
  8015=>"100010001",
  8016=>"110000011",
  8017=>"111101000",
  8018=>"111110000",
  8019=>"001110101",
  8020=>"000111011",
  8021=>"010111111",
  8022=>"001101001",
  8023=>"001010010",
  8024=>"111101111",
  8025=>"100111011",
  8026=>"011110111",
  8027=>"011111101",
  8028=>"001000100",
  8029=>"101000001",
  8030=>"000110110",
  8031=>"101110000",
  8032=>"001011100",
  8033=>"000011001",
  8034=>"101000110",
  8035=>"111010100",
  8036=>"100001100",
  8037=>"011010010",
  8038=>"110101001",
  8039=>"101101110",
  8040=>"001101000",
  8041=>"011110101",
  8042=>"001110100",
  8043=>"100010111",
  8044=>"001110001",
  8045=>"010100100",
  8046=>"001110110",
  8047=>"111111010",
  8048=>"000110111",
  8049=>"011001101",
  8050=>"110011101",
  8051=>"001001000",
  8052=>"000001010",
  8053=>"100001111",
  8054=>"101110010",
  8055=>"111100100",
  8056=>"001000111",
  8057=>"010101011",
  8058=>"110011101",
  8059=>"110000101",
  8060=>"011100000",
  8061=>"100101101",
  8062=>"101010100",
  8063=>"001101101",
  8064=>"111010001",
  8065=>"010100010",
  8066=>"100100101",
  8067=>"010111010",
  8068=>"010110100",
  8069=>"010000101",
  8070=>"001111100",
  8071=>"111111011",
  8072=>"010111000",
  8073=>"011111110",
  8074=>"101101111",
  8075=>"010000001",
  8076=>"000001001",
  8077=>"100001101",
  8078=>"111001111",
  8079=>"111001110",
  8080=>"111000000",
  8081=>"000010101",
  8082=>"011110110",
  8083=>"011000010",
  8084=>"001001111",
  8085=>"000111001",
  8086=>"010110011",
  8087=>"000100011",
  8088=>"000001000",
  8089=>"111101111",
  8090=>"100110001",
  8091=>"000000100",
  8092=>"110000000",
  8093=>"111010000",
  8094=>"001001001",
  8095=>"100110000",
  8096=>"000000001",
  8097=>"110011000",
  8098=>"111100100",
  8099=>"100001000",
  8100=>"111000000",
  8101=>"001101111",
  8102=>"100100000",
  8103=>"110000111",
  8104=>"001100010",
  8105=>"110100111",
  8106=>"000111100",
  8107=>"000110000",
  8108=>"110010001",
  8109=>"100011001",
  8110=>"001101010",
  8111=>"000110101",
  8112=>"000111000",
  8113=>"110001010",
  8114=>"011000111",
  8115=>"100000001",
  8116=>"000001011",
  8117=>"111111101",
  8118=>"111110100",
  8119=>"110101011",
  8120=>"101101001",
  8121=>"111111001",
  8122=>"011111011",
  8123=>"011010100",
  8124=>"101001100",
  8125=>"010000000",
  8126=>"011011100",
  8127=>"110001000",
  8128=>"100011000",
  8129=>"000111011",
  8130=>"101011000",
  8131=>"001011011",
  8132=>"010100111",
  8133=>"110011110",
  8134=>"100101011",
  8135=>"000110100",
  8136=>"000010001",
  8137=>"111010100",
  8138=>"100101001",
  8139=>"100000010",
  8140=>"000000111",
  8141=>"101000111",
  8142=>"111000000",
  8143=>"110001101",
  8144=>"100011001",
  8145=>"100000010",
  8146=>"000101001",
  8147=>"110000100",
  8148=>"011110010",
  8149=>"010101101",
  8150=>"010011011",
  8151=>"110110111",
  8152=>"110110111",
  8153=>"001011010",
  8154=>"101111110",
  8155=>"000001111",
  8156=>"000110101",
  8157=>"011011001",
  8158=>"000000110",
  8159=>"011010111",
  8160=>"100110001",
  8161=>"010010101",
  8162=>"001011011",
  8163=>"101001111",
  8164=>"100100100",
  8165=>"001001011",
  8166=>"110000100",
  8167=>"110100100",
  8168=>"001000010",
  8169=>"111111001",
  8170=>"010011100",
  8171=>"101011010",
  8172=>"011111100",
  8173=>"000000011",
  8174=>"100000111",
  8175=>"011010010",
  8176=>"100001110",
  8177=>"101100111",
  8178=>"101111100",
  8179=>"101000111",
  8180=>"001011011",
  8181=>"001100101",
  8182=>"101000000",
  8183=>"011111111",
  8184=>"000001100",
  8185=>"110110011",
  8186=>"000101111",
  8187=>"100110011",
  8188=>"010011000",
  8189=>"010000001",
  8190=>"011110000",
  8191=>"100111111",
  8192=>"101001100",
  8193=>"011010101",
  8194=>"010001000",
  8195=>"000100101",
  8196=>"101111010",
  8197=>"110100111",
  8198=>"111100100",
  8199=>"000110010",
  8200=>"001000111",
  8201=>"101001000",
  8202=>"110000110",
  8203=>"001010010",
  8204=>"111101011",
  8205=>"110110000",
  8206=>"011010000",
  8207=>"111111100",
  8208=>"001001001",
  8209=>"101111101",
  8210=>"111100010",
  8211=>"010000000",
  8212=>"001111100",
  8213=>"100000010",
  8214=>"000001110",
  8215=>"101101001",
  8216=>"110000100",
  8217=>"100010000",
  8218=>"010010100",
  8219=>"000000001",
  8220=>"100001001",
  8221=>"101010011",
  8222=>"110110011",
  8223=>"011000001",
  8224=>"011111110",
  8225=>"100111100",
  8226=>"001111010",
  8227=>"101001000",
  8228=>"111011000",
  8229=>"001001000",
  8230=>"010110011",
  8231=>"100111110",
  8232=>"111011101",
  8233=>"010111100",
  8234=>"110110100",
  8235=>"101001101",
  8236=>"110101111",
  8237=>"000101001",
  8238=>"000010100",
  8239=>"001010110",
  8240=>"100010111",
  8241=>"111001011",
  8242=>"101011100",
  8243=>"010001011",
  8244=>"100010011",
  8245=>"101011011",
  8246=>"011000101",
  8247=>"000010000",
  8248=>"100100011",
  8249=>"011100100",
  8250=>"000100100",
  8251=>"011111110",
  8252=>"111111011",
  8253=>"000000111",
  8254=>"011001000",
  8255=>"101110110",
  8256=>"111011001",
  8257=>"001100110",
  8258=>"110010110",
  8259=>"001010110",
  8260=>"101011110",
  8261=>"010100101",
  8262=>"101111011",
  8263=>"111001101",
  8264=>"100000010",
  8265=>"001000101",
  8266=>"111001101",
  8267=>"101011111",
  8268=>"100001010",
  8269=>"110001001",
  8270=>"000010000",
  8271=>"100100000",
  8272=>"000010000",
  8273=>"111111011",
  8274=>"000100110",
  8275=>"101001011",
  8276=>"111000100",
  8277=>"100010001",
  8278=>"000010001",
  8279=>"101001001",
  8280=>"100101100",
  8281=>"101001011",
  8282=>"000101010",
  8283=>"111000100",
  8284=>"101100110",
  8285=>"100100101",
  8286=>"100101100",
  8287=>"000000001",
  8288=>"000011001",
  8289=>"111001101",
  8290=>"000100111",
  8291=>"010010111",
  8292=>"011111111",
  8293=>"000010110",
  8294=>"000001000",
  8295=>"010011110",
  8296=>"100011111",
  8297=>"000010001",
  8298=>"110110000",
  8299=>"011110011",
  8300=>"100001100",
  8301=>"011100000",
  8302=>"000000011",
  8303=>"011010000",
  8304=>"110011110",
  8305=>"110000001",
  8306=>"001100100",
  8307=>"110110010",
  8308=>"000001000",
  8309=>"100010110",
  8310=>"001000110",
  8311=>"001101111",
  8312=>"110100010",
  8313=>"111011101",
  8314=>"001100000",
  8315=>"101101100",
  8316=>"011000000",
  8317=>"110111110",
  8318=>"111011101",
  8319=>"100101111",
  8320=>"110110010",
  8321=>"111100111",
  8322=>"000000011",
  8323=>"000110010",
  8324=>"011000001",
  8325=>"111100110",
  8326=>"110110110",
  8327=>"011000011",
  8328=>"100100010",
  8329=>"111011011",
  8330=>"011000001",
  8331=>"111011111",
  8332=>"101010010",
  8333=>"100100000",
  8334=>"111101010",
  8335=>"011010110",
  8336=>"110010101",
  8337=>"100100101",
  8338=>"010001000",
  8339=>"111111110",
  8340=>"000111110",
  8341=>"001000010",
  8342=>"001110101",
  8343=>"000100000",
  8344=>"100111010",
  8345=>"101011110",
  8346=>"101110001",
  8347=>"100011011",
  8348=>"010011110",
  8349=>"000101110",
  8350=>"111101101",
  8351=>"010010100",
  8352=>"101111100",
  8353=>"011010101",
  8354=>"101011100",
  8355=>"001011111",
  8356=>"101111100",
  8357=>"111111111",
  8358=>"011110011",
  8359=>"011101101",
  8360=>"010010100",
  8361=>"110011011",
  8362=>"111101011",
  8363=>"100000111",
  8364=>"010111111",
  8365=>"100010000",
  8366=>"101100110",
  8367=>"100011100",
  8368=>"000100010",
  8369=>"000111111",
  8370=>"111010010",
  8371=>"011001110",
  8372=>"001011000",
  8373=>"101011000",
  8374=>"010111001",
  8375=>"101000001",
  8376=>"010000100",
  8377=>"001010010",
  8378=>"011011000",
  8379=>"000101110",
  8380=>"001011011",
  8381=>"100100010",
  8382=>"010010010",
  8383=>"000110010",
  8384=>"000010101",
  8385=>"111010110",
  8386=>"101110101",
  8387=>"001011111",
  8388=>"000001101",
  8389=>"111111100",
  8390=>"110101010",
  8391=>"101001001",
  8392=>"010111011",
  8393=>"101101111",
  8394=>"000110111",
  8395=>"010000111",
  8396=>"100011111",
  8397=>"001000101",
  8398=>"011011001",
  8399=>"111001100",
  8400=>"100111110",
  8401=>"100111011",
  8402=>"100010101",
  8403=>"000100010",
  8404=>"101110000",
  8405=>"000110010",
  8406=>"011100110",
  8407=>"001010011",
  8408=>"101101101",
  8409=>"001100000",
  8410=>"111101101",
  8411=>"111001011",
  8412=>"010110101",
  8413=>"101011101",
  8414=>"001110001",
  8415=>"100100101",
  8416=>"011100100",
  8417=>"111101111",
  8418=>"001010110",
  8419=>"101100100",
  8420=>"000010001",
  8421=>"000000000",
  8422=>"001100000",
  8423=>"111111001",
  8424=>"111011011",
  8425=>"110101100",
  8426=>"110100110",
  8427=>"001110101",
  8428=>"111001100",
  8429=>"100111100",
  8430=>"100110010",
  8431=>"010011001",
  8432=>"010000111",
  8433=>"011110110",
  8434=>"011001111",
  8435=>"011011000",
  8436=>"111011110",
  8437=>"001101110",
  8438=>"101101011",
  8439=>"111100110",
  8440=>"011111100",
  8441=>"111111110",
  8442=>"001011110",
  8443=>"001000100",
  8444=>"111110101",
  8445=>"111101111",
  8446=>"000000110",
  8447=>"100000101",
  8448=>"011011000",
  8449=>"011100110",
  8450=>"100001011",
  8451=>"101011000",
  8452=>"001000001",
  8453=>"011110110",
  8454=>"011101110",
  8455=>"111001111",
  8456=>"010100010",
  8457=>"110110111",
  8458=>"010000110",
  8459=>"110000100",
  8460=>"110000000",
  8461=>"111011100",
  8462=>"101000011",
  8463=>"000000111",
  8464=>"011001011",
  8465=>"001001000",
  8466=>"010011100",
  8467=>"111010001",
  8468=>"110011011",
  8469=>"101111010",
  8470=>"100110100",
  8471=>"001100011",
  8472=>"101110000",
  8473=>"100000101",
  8474=>"011000101",
  8475=>"000001010",
  8476=>"001100000",
  8477=>"100100000",
  8478=>"110011110",
  8479=>"010011001",
  8480=>"010000110",
  8481=>"001100001",
  8482=>"101000010",
  8483=>"111101100",
  8484=>"001000010",
  8485=>"111011010",
  8486=>"001111111",
  8487=>"000010010",
  8488=>"000111100",
  8489=>"010111111",
  8490=>"101100011",
  8491=>"010111100",
  8492=>"101110001",
  8493=>"111101101",
  8494=>"110011110",
  8495=>"110101000",
  8496=>"101110001",
  8497=>"010000010",
  8498=>"001100110",
  8499=>"000010000",
  8500=>"100000010",
  8501=>"100001111",
  8502=>"011100111",
  8503=>"100111010",
  8504=>"011111110",
  8505=>"000101111",
  8506=>"111101101",
  8507=>"000001010",
  8508=>"001110111",
  8509=>"001001110",
  8510=>"000010001",
  8511=>"101000010",
  8512=>"111111011",
  8513=>"100111011",
  8514=>"011011100",
  8515=>"100011001",
  8516=>"111011001",
  8517=>"100010110",
  8518=>"000100000",
  8519=>"010100100",
  8520=>"101000000",
  8521=>"101111011",
  8522=>"101000111",
  8523=>"111000101",
  8524=>"001010011",
  8525=>"111111010",
  8526=>"001011010",
  8527=>"111000000",
  8528=>"011001010",
  8529=>"100010000",
  8530=>"100011000",
  8531=>"000000000",
  8532=>"100000110",
  8533=>"111001010",
  8534=>"000001110",
  8535=>"111010111",
  8536=>"000110011",
  8537=>"111001110",
  8538=>"001000001",
  8539=>"011000011",
  8540=>"101111001",
  8541=>"010001100",
  8542=>"111110010",
  8543=>"100010110",
  8544=>"011011111",
  8545=>"000001011",
  8546=>"000011101",
  8547=>"000000111",
  8548=>"001010000",
  8549=>"110100101",
  8550=>"101000111",
  8551=>"110110000",
  8552=>"000101110",
  8553=>"111101010",
  8554=>"101010000",
  8555=>"100011101",
  8556=>"101110001",
  8557=>"000011111",
  8558=>"001000110",
  8559=>"000010110",
  8560=>"001100001",
  8561=>"001100111",
  8562=>"100111011",
  8563=>"100000001",
  8564=>"100001000",
  8565=>"011100001",
  8566=>"111011110",
  8567=>"000001111",
  8568=>"011110011",
  8569=>"100101010",
  8570=>"010010101",
  8571=>"010011001",
  8572=>"111100010",
  8573=>"011000000",
  8574=>"111010010",
  8575=>"011000011",
  8576=>"100100110",
  8577=>"000011111",
  8578=>"101010011",
  8579=>"001101100",
  8580=>"111111000",
  8581=>"010110110",
  8582=>"101110011",
  8583=>"011000101",
  8584=>"100001011",
  8585=>"111110110",
  8586=>"111001101",
  8587=>"100111111",
  8588=>"100110110",
  8589=>"111001000",
  8590=>"110010000",
  8591=>"100100010",
  8592=>"101000000",
  8593=>"011000000",
  8594=>"101110010",
  8595=>"010111011",
  8596=>"111010100",
  8597=>"001001011",
  8598=>"001000000",
  8599=>"011001101",
  8600=>"001000010",
  8601=>"000100111",
  8602=>"101011011",
  8603=>"101101100",
  8604=>"100100001",
  8605=>"111011111",
  8606=>"011011111",
  8607=>"110100011",
  8608=>"101101000",
  8609=>"000001111",
  8610=>"000001101",
  8611=>"001111100",
  8612=>"101111110",
  8613=>"111100011",
  8614=>"110011010",
  8615=>"000001100",
  8616=>"110110100",
  8617=>"001100111",
  8618=>"010110011",
  8619=>"011101000",
  8620=>"000101001",
  8621=>"000110010",
  8622=>"001000000",
  8623=>"111001111",
  8624=>"110001110",
  8625=>"100110111",
  8626=>"000101101",
  8627=>"101011101",
  8628=>"010111110",
  8629=>"010100010",
  8630=>"101101010",
  8631=>"111001101",
  8632=>"010100000",
  8633=>"000000011",
  8634=>"001110101",
  8635=>"000110011",
  8636=>"010101111",
  8637=>"001001101",
  8638=>"100000110",
  8639=>"001110000",
  8640=>"010100000",
  8641=>"011110100",
  8642=>"110110110",
  8643=>"100000000",
  8644=>"001111001",
  8645=>"111111111",
  8646=>"000100000",
  8647=>"111101101",
  8648=>"001110000",
  8649=>"011100010",
  8650=>"110000100",
  8651=>"110001101",
  8652=>"010000010",
  8653=>"000001110",
  8654=>"100111011",
  8655=>"100101011",
  8656=>"011101100",
  8657=>"011011010",
  8658=>"100011010",
  8659=>"011101111",
  8660=>"000110001",
  8661=>"001111011",
  8662=>"100100100",
  8663=>"101000111",
  8664=>"100001000",
  8665=>"101100011",
  8666=>"010000010",
  8667=>"111001111",
  8668=>"010010010",
  8669=>"111110001",
  8670=>"000111111",
  8671=>"001011111",
  8672=>"110011111",
  8673=>"011100011",
  8674=>"111100001",
  8675=>"010011101",
  8676=>"010100111",
  8677=>"110100000",
  8678=>"011111000",
  8679=>"111101001",
  8680=>"110010101",
  8681=>"101011110",
  8682=>"110010100",
  8683=>"011001110",
  8684=>"101000001",
  8685=>"101100010",
  8686=>"010100011",
  8687=>"000000110",
  8688=>"110110110",
  8689=>"011001001",
  8690=>"010111101",
  8691=>"011011010",
  8692=>"011011110",
  8693=>"000000110",
  8694=>"010110100",
  8695=>"010111001",
  8696=>"011101001",
  8697=>"111111011",
  8698=>"101001110",
  8699=>"101001111",
  8700=>"011001100",
  8701=>"110010111",
  8702=>"001111000",
  8703=>"011011010",
  8704=>"110001010",
  8705=>"100010010",
  8706=>"110101101",
  8707=>"001000110",
  8708=>"001010011",
  8709=>"111110000",
  8710=>"000110100",
  8711=>"010000001",
  8712=>"011001110",
  8713=>"101000000",
  8714=>"010000111",
  8715=>"011101101",
  8716=>"000100001",
  8717=>"111110001",
  8718=>"000101000",
  8719=>"000110100",
  8720=>"111111101",
  8721=>"010110111",
  8722=>"100000101",
  8723=>"111000001",
  8724=>"010011011",
  8725=>"110011010",
  8726=>"000101000",
  8727=>"000100101",
  8728=>"001010101",
  8729=>"001011000",
  8730=>"001000110",
  8731=>"110101111",
  8732=>"101100011",
  8733=>"001001111",
  8734=>"101100011",
  8735=>"100100111",
  8736=>"010010111",
  8737=>"000001011",
  8738=>"101001000",
  8739=>"000000000",
  8740=>"101011111",
  8741=>"110011111",
  8742=>"111101111",
  8743=>"000000001",
  8744=>"100000111",
  8745=>"111010101",
  8746=>"100101101",
  8747=>"110000111",
  8748=>"011001110",
  8749=>"000000011",
  8750=>"000100000",
  8751=>"110110100",
  8752=>"001110000",
  8753=>"110011111",
  8754=>"110001111",
  8755=>"000100110",
  8756=>"010101111",
  8757=>"011101001",
  8758=>"011001001",
  8759=>"010000111",
  8760=>"100111101",
  8761=>"010011110",
  8762=>"101110010",
  8763=>"010010011",
  8764=>"100110111",
  8765=>"100011101",
  8766=>"011100110",
  8767=>"011011001",
  8768=>"100001001",
  8769=>"110111010",
  8770=>"111101000",
  8771=>"010101001",
  8772=>"000101101",
  8773=>"100101110",
  8774=>"111000100",
  8775=>"101010001",
  8776=>"101010110",
  8777=>"000001100",
  8778=>"000011100",
  8779=>"111001111",
  8780=>"010101110",
  8781=>"101101010",
  8782=>"110100000",
  8783=>"110001011",
  8784=>"110101000",
  8785=>"111101011",
  8786=>"101101111",
  8787=>"011100000",
  8788=>"100110110",
  8789=>"101011101",
  8790=>"101110010",
  8791=>"111011001",
  8792=>"101100111",
  8793=>"110101011",
  8794=>"011110011",
  8795=>"100001010",
  8796=>"001101011",
  8797=>"010110001",
  8798=>"101000000",
  8799=>"100001101",
  8800=>"010010001",
  8801=>"111101011",
  8802=>"001101100",
  8803=>"000111111",
  8804=>"101111001",
  8805=>"010110001",
  8806=>"001001001",
  8807=>"000101111",
  8808=>"011111001",
  8809=>"110010110",
  8810=>"101110111",
  8811=>"101001000",
  8812=>"101010001",
  8813=>"011110101",
  8814=>"010110000",
  8815=>"001011101",
  8816=>"001111101",
  8817=>"100101010",
  8818=>"000100100",
  8819=>"100001000",
  8820=>"101011111",
  8821=>"010000100",
  8822=>"111101000",
  8823=>"101100110",
  8824=>"000100010",
  8825=>"110101100",
  8826=>"101001000",
  8827=>"110010111",
  8828=>"001101000",
  8829=>"000001101",
  8830=>"110000010",
  8831=>"011000011",
  8832=>"110011001",
  8833=>"110011110",
  8834=>"110001111",
  8835=>"110010010",
  8836=>"110110110",
  8837=>"111110111",
  8838=>"110011100",
  8839=>"110000111",
  8840=>"011101000",
  8841=>"010101000",
  8842=>"100000111",
  8843=>"101110101",
  8844=>"011111100",
  8845=>"101100110",
  8846=>"101100011",
  8847=>"000001100",
  8848=>"000001001",
  8849=>"001111111",
  8850=>"111111110",
  8851=>"000011101",
  8852=>"010010100",
  8853=>"101011100",
  8854=>"101001111",
  8855=>"000101011",
  8856=>"010100100",
  8857=>"000111011",
  8858=>"101111110",
  8859=>"000000101",
  8860=>"001011000",
  8861=>"100101010",
  8862=>"111101111",
  8863=>"100000011",
  8864=>"111111101",
  8865=>"011110111",
  8866=>"101110101",
  8867=>"101101010",
  8868=>"111010001",
  8869=>"011011011",
  8870=>"100001011",
  8871=>"111100101",
  8872=>"001110000",
  8873=>"011000111",
  8874=>"001011100",
  8875=>"101101000",
  8876=>"110100011",
  8877=>"101111010",
  8878=>"111000100",
  8879=>"000111010",
  8880=>"101100110",
  8881=>"000111100",
  8882=>"110101011",
  8883=>"001001001",
  8884=>"011101110",
  8885=>"101110000",
  8886=>"111100011",
  8887=>"110101010",
  8888=>"111000111",
  8889=>"000111000",
  8890=>"011011001",
  8891=>"011000011",
  8892=>"011011000",
  8893=>"010001000",
  8894=>"001101011",
  8895=>"101000100",
  8896=>"111011011",
  8897=>"000101100",
  8898=>"000001111",
  8899=>"010001000",
  8900=>"100111101",
  8901=>"111011100",
  8902=>"101001110",
  8903=>"100000110",
  8904=>"011010110",
  8905=>"000101001",
  8906=>"000001100",
  8907=>"100000111",
  8908=>"000101111",
  8909=>"011001100",
  8910=>"011101000",
  8911=>"111110010",
  8912=>"111111001",
  8913=>"011001100",
  8914=>"101100101",
  8915=>"001000000",
  8916=>"000110100",
  8917=>"100111010",
  8918=>"011011000",
  8919=>"000111000",
  8920=>"111001011",
  8921=>"001010111",
  8922=>"101100000",
  8923=>"100001011",
  8924=>"001110011",
  8925=>"001001010",
  8926=>"011111000",
  8927=>"110011000",
  8928=>"011000100",
  8929=>"111011110",
  8930=>"111010001",
  8931=>"000111010",
  8932=>"011010011",
  8933=>"111000101",
  8934=>"010010001",
  8935=>"011010100",
  8936=>"101110010",
  8937=>"111100100",
  8938=>"010011101",
  8939=>"001011011",
  8940=>"101001001",
  8941=>"001100111",
  8942=>"101001001",
  8943=>"111100000",
  8944=>"111111000",
  8945=>"001000011",
  8946=>"000001110",
  8947=>"100011001",
  8948=>"011000010",
  8949=>"111000000",
  8950=>"000000100",
  8951=>"111111100",
  8952=>"001111101",
  8953=>"101011101",
  8954=>"100000111",
  8955=>"011010001",
  8956=>"101100100",
  8957=>"010011111",
  8958=>"110010001",
  8959=>"000001111",
  8960=>"110111001",
  8961=>"100001111",
  8962=>"011110010",
  8963=>"010001111",
  8964=>"000110000",
  8965=>"100001000",
  8966=>"001010101",
  8967=>"011011010",
  8968=>"100000001",
  8969=>"110110000",
  8970=>"110001001",
  8971=>"001000000",
  8972=>"111110100",
  8973=>"100100010",
  8974=>"011100111",
  8975=>"100111100",
  8976=>"010001111",
  8977=>"110110011",
  8978=>"111101100",
  8979=>"001001110",
  8980=>"000011111",
  8981=>"011110001",
  8982=>"011110100",
  8983=>"010000110",
  8984=>"000001000",
  8985=>"100001001",
  8986=>"111110100",
  8987=>"110111110",
  8988=>"001010000",
  8989=>"001010101",
  8990=>"111011000",
  8991=>"110110100",
  8992=>"110111101",
  8993=>"111101101",
  8994=>"110111111",
  8995=>"101100001",
  8996=>"000101110",
  8997=>"111010001",
  8998=>"010111011",
  8999=>"100000010",
  9000=>"000010010",
  9001=>"001111111",
  9002=>"100100111",
  9003=>"010101100",
  9004=>"000111000",
  9005=>"000011111",
  9006=>"101110000",
  9007=>"101101110",
  9008=>"101100110",
  9009=>"111110111",
  9010=>"010110101",
  9011=>"011101000",
  9012=>"101111001",
  9013=>"000010101",
  9014=>"100111001",
  9015=>"110101110",
  9016=>"101011111",
  9017=>"101100110",
  9018=>"010110110",
  9019=>"001101010",
  9020=>"100000000",
  9021=>"000110001",
  9022=>"100001111",
  9023=>"010010000",
  9024=>"001111000",
  9025=>"011001111",
  9026=>"001001010",
  9027=>"100001100",
  9028=>"000111010",
  9029=>"100101110",
  9030=>"001010111",
  9031=>"010000111",
  9032=>"101110010",
  9033=>"010010001",
  9034=>"101001011",
  9035=>"110110110",
  9036=>"100001001",
  9037=>"011000001",
  9038=>"111110101",
  9039=>"001010111",
  9040=>"100000011",
  9041=>"100111000",
  9042=>"101101011",
  9043=>"111101000",
  9044=>"111100101",
  9045=>"100100110",
  9046=>"111000100",
  9047=>"011001010",
  9048=>"000011011",
  9049=>"100000101",
  9050=>"110100100",
  9051=>"111101001",
  9052=>"111000110",
  9053=>"100110110",
  9054=>"001101011",
  9055=>"010001100",
  9056=>"111111010",
  9057=>"001100000",
  9058=>"000000001",
  9059=>"001101001",
  9060=>"100010011",
  9061=>"000110111",
  9062=>"100011001",
  9063=>"111000010",
  9064=>"111111111",
  9065=>"000111110",
  9066=>"011110110",
  9067=>"100101111",
  9068=>"010100001",
  9069=>"101001100",
  9070=>"000111111",
  9071=>"110010011",
  9072=>"101100000",
  9073=>"101001011",
  9074=>"111000101",
  9075=>"011101101",
  9076=>"100000001",
  9077=>"011111101",
  9078=>"110111110",
  9079=>"010011101",
  9080=>"111110110",
  9081=>"000110110",
  9082=>"101011010",
  9083=>"001000101",
  9084=>"011001001",
  9085=>"010011010",
  9086=>"101100000",
  9087=>"010010100",
  9088=>"110010100",
  9089=>"111110110",
  9090=>"100000000",
  9091=>"100010000",
  9092=>"100110001",
  9093=>"001111001",
  9094=>"010000000",
  9095=>"110101110",
  9096=>"101001001",
  9097=>"101100111",
  9098=>"010100000",
  9099=>"101110001",
  9100=>"001011110",
  9101=>"011011110",
  9102=>"111100111",
  9103=>"101101011",
  9104=>"000111000",
  9105=>"011100100",
  9106=>"110010000",
  9107=>"011101111",
  9108=>"011011011",
  9109=>"110100101",
  9110=>"000100110",
  9111=>"000100111",
  9112=>"011001000",
  9113=>"100111101",
  9114=>"001100001",
  9115=>"010000101",
  9116=>"001011101",
  9117=>"011111000",
  9118=>"111010101",
  9119=>"101110110",
  9120=>"000110010",
  9121=>"011111011",
  9122=>"111001000",
  9123=>"100101000",
  9124=>"101101101",
  9125=>"010001100",
  9126=>"101110001",
  9127=>"111000010",
  9128=>"011000100",
  9129=>"111001101",
  9130=>"100001010",
  9131=>"100001011",
  9132=>"001101110",
  9133=>"011011010",
  9134=>"001000000",
  9135=>"000101110",
  9136=>"101010011",
  9137=>"101100100",
  9138=>"111011011",
  9139=>"101101101",
  9140=>"100100011",
  9141=>"000111111",
  9142=>"010010111",
  9143=>"100110011",
  9144=>"100100100",
  9145=>"010100001",
  9146=>"110000000",
  9147=>"111001010",
  9148=>"100011011",
  9149=>"010001010",
  9150=>"101110101",
  9151=>"100000101",
  9152=>"011101100",
  9153=>"111000101",
  9154=>"000101101",
  9155=>"100101101",
  9156=>"100001000",
  9157=>"001100100",
  9158=>"000011001",
  9159=>"010010010",
  9160=>"011111010",
  9161=>"111101110",
  9162=>"001011010",
  9163=>"000000110",
  9164=>"100110010",
  9165=>"100000001",
  9166=>"100000111",
  9167=>"110000000",
  9168=>"000100111",
  9169=>"101110001",
  9170=>"110010100",
  9171=>"010011110",
  9172=>"000000011",
  9173=>"000110010",
  9174=>"100101011",
  9175=>"000010111",
  9176=>"111101111",
  9177=>"000011111",
  9178=>"000001111",
  9179=>"111100010",
  9180=>"000001110",
  9181=>"001111000",
  9182=>"001100000",
  9183=>"000111100",
  9184=>"001000100",
  9185=>"111011010",
  9186=>"101010001",
  9187=>"110000000",
  9188=>"010101001",
  9189=>"000101100",
  9190=>"111111010",
  9191=>"110101000",
  9192=>"000101001",
  9193=>"000001000",
  9194=>"100011110",
  9195=>"010111010",
  9196=>"000111111",
  9197=>"000011011",
  9198=>"110000010",
  9199=>"101001100",
  9200=>"010110011",
  9201=>"111011011",
  9202=>"000100001",
  9203=>"011111110",
  9204=>"111110111",
  9205=>"001101111",
  9206=>"100001111",
  9207=>"010001001",
  9208=>"011010000",
  9209=>"100110100",
  9210=>"100111111",
  9211=>"110000000",
  9212=>"011001101",
  9213=>"101001110",
  9214=>"100111000",
  9215=>"011010010",
  9216=>"011101110",
  9217=>"001110110",
  9218=>"101101011",
  9219=>"000001110",
  9220=>"111111100",
  9221=>"110111001",
  9222=>"011011100",
  9223=>"000111000",
  9224=>"100010110",
  9225=>"110000001",
  9226=>"010000001",
  9227=>"101001101",
  9228=>"000000010",
  9229=>"100000011",
  9230=>"101111001",
  9231=>"110011101",
  9232=>"011001100",
  9233=>"101010000",
  9234=>"100111101",
  9235=>"011000010",
  9236=>"000000001",
  9237=>"000000010",
  9238=>"011000010",
  9239=>"111010000",
  9240=>"111001011",
  9241=>"110111010",
  9242=>"011011011",
  9243=>"110001000",
  9244=>"111000101",
  9245=>"101101100",
  9246=>"011011010",
  9247=>"001001000",
  9248=>"100100001",
  9249=>"111001110",
  9250=>"111100000",
  9251=>"011100110",
  9252=>"110011000",
  9253=>"101011011",
  9254=>"011010000",
  9255=>"001000011",
  9256=>"010110111",
  9257=>"010010000",
  9258=>"101000110",
  9259=>"001111011",
  9260=>"110101111",
  9261=>"000101100",
  9262=>"100000000",
  9263=>"101010101",
  9264=>"000011010",
  9265=>"000000101",
  9266=>"000000000",
  9267=>"101111110",
  9268=>"100100011",
  9269=>"000011000",
  9270=>"101110101",
  9271=>"100011010",
  9272=>"010001010",
  9273=>"100101100",
  9274=>"010000100",
  9275=>"110100101",
  9276=>"001110110",
  9277=>"111101110",
  9278=>"001110110",
  9279=>"100000000",
  9280=>"000101000",
  9281=>"000010101",
  9282=>"000000010",
  9283=>"100100001",
  9284=>"110000111",
  9285=>"110111111",
  9286=>"011001101",
  9287=>"110001100",
  9288=>"001100011",
  9289=>"100010100",
  9290=>"010001000",
  9291=>"101100000",
  9292=>"001000111",
  9293=>"110011100",
  9294=>"111101111",
  9295=>"000111011",
  9296=>"011000010",
  9297=>"111101101",
  9298=>"011001000",
  9299=>"100011001",
  9300=>"101010100",
  9301=>"000100000",
  9302=>"011010010",
  9303=>"110000000",
  9304=>"000100000",
  9305=>"001010111",
  9306=>"001010001",
  9307=>"101101101",
  9308=>"010101101",
  9309=>"000110010",
  9310=>"100110111",
  9311=>"001000010",
  9312=>"001111100",
  9313=>"010010000",
  9314=>"100001000",
  9315=>"111010101",
  9316=>"100001110",
  9317=>"101111000",
  9318=>"001110010",
  9319=>"100000101",
  9320=>"100010010",
  9321=>"101101111",
  9322=>"101011000",
  9323=>"100000110",
  9324=>"111011100",
  9325=>"101001101",
  9326=>"110000011",
  9327=>"000011000",
  9328=>"001011001",
  9329=>"111000110",
  9330=>"110100111",
  9331=>"000000010",
  9332=>"000100110",
  9333=>"001001101",
  9334=>"110001101",
  9335=>"101000101",
  9336=>"001000011",
  9337=>"111111010",
  9338=>"101101110",
  9339=>"100110011",
  9340=>"110001000",
  9341=>"001001000",
  9342=>"111101110",
  9343=>"001010111",
  9344=>"011110001",
  9345=>"001010101",
  9346=>"101110010",
  9347=>"000000000",
  9348=>"011000001",
  9349=>"011000111",
  9350=>"000111111",
  9351=>"001001011",
  9352=>"010110110",
  9353=>"110110100",
  9354=>"001101101",
  9355=>"111000101",
  9356=>"111010100",
  9357=>"000010010",
  9358=>"110111000",
  9359=>"100101001",
  9360=>"011001100",
  9361=>"010101101",
  9362=>"100100110",
  9363=>"101111001",
  9364=>"110111100",
  9365=>"100111111",
  9366=>"100010001",
  9367=>"100001011",
  9368=>"010011000",
  9369=>"110010100",
  9370=>"000000000",
  9371=>"110111011",
  9372=>"110010010",
  9373=>"000101001",
  9374=>"110010001",
  9375=>"001010010",
  9376=>"100010000",
  9377=>"011100010",
  9378=>"001011111",
  9379=>"000111100",
  9380=>"011010111",
  9381=>"100011110",
  9382=>"101010101",
  9383=>"010010000",
  9384=>"010010011",
  9385=>"000000001",
  9386=>"100011101",
  9387=>"000111000",
  9388=>"000101101",
  9389=>"111101110",
  9390=>"101111111",
  9391=>"010110110",
  9392=>"111011101",
  9393=>"111001001",
  9394=>"000100001",
  9395=>"000100110",
  9396=>"010001110",
  9397=>"000000000",
  9398=>"010101011",
  9399=>"011101011",
  9400=>"000001110",
  9401=>"001011001",
  9402=>"011100101",
  9403=>"000001111",
  9404=>"000110111",
  9405=>"000110011",
  9406=>"011110101",
  9407=>"010101010",
  9408=>"000011100",
  9409=>"101101010",
  9410=>"000010000",
  9411=>"111111011",
  9412=>"111101100",
  9413=>"010101101",
  9414=>"100001111",
  9415=>"111000001",
  9416=>"011100110",
  9417=>"000101001",
  9418=>"000100010",
  9419=>"110010100",
  9420=>"111000011",
  9421=>"010111011",
  9422=>"100110011",
  9423=>"000110110",
  9424=>"001001011",
  9425=>"111101000",
  9426=>"000011010",
  9427=>"011011001",
  9428=>"001011100",
  9429=>"100011111",
  9430=>"010001011",
  9431=>"001010111",
  9432=>"011001010",
  9433=>"011011100",
  9434=>"111010011",
  9435=>"011001100",
  9436=>"000101111",
  9437=>"111001010",
  9438=>"100111010",
  9439=>"101011010",
  9440=>"001111100",
  9441=>"101111111",
  9442=>"010011111",
  9443=>"101101100",
  9444=>"110101101",
  9445=>"101000000",
  9446=>"001101110",
  9447=>"110100000",
  9448=>"101110100",
  9449=>"011011110",
  9450=>"111101010",
  9451=>"001101100",
  9452=>"101001000",
  9453=>"011110000",
  9454=>"100010110",
  9455=>"000100000",
  9456=>"011011000",
  9457=>"000100010",
  9458=>"000110100",
  9459=>"001000111",
  9460=>"000010101",
  9461=>"111111010",
  9462=>"011011000",
  9463=>"000010001",
  9464=>"110001110",
  9465=>"010010001",
  9466=>"001010111",
  9467=>"101111000",
  9468=>"101000110",
  9469=>"100100011",
  9470=>"101001011",
  9471=>"011010111",
  9472=>"011011111",
  9473=>"100101101",
  9474=>"011111110",
  9475=>"100001110",
  9476=>"100001101",
  9477=>"110011000",
  9478=>"101110101",
  9479=>"000110101",
  9480=>"011010001",
  9481=>"100111111",
  9482=>"000100010",
  9483=>"010000100",
  9484=>"101101001",
  9485=>"110001110",
  9486=>"111100001",
  9487=>"000110010",
  9488=>"101101111",
  9489=>"100100100",
  9490=>"001001001",
  9491=>"101011101",
  9492=>"011111000",
  9493=>"110110111",
  9494=>"110110011",
  9495=>"011001111",
  9496=>"000011000",
  9497=>"011101010",
  9498=>"000101001",
  9499=>"011000000",
  9500=>"111000111",
  9501=>"100000000",
  9502=>"011011011",
  9503=>"101011001",
  9504=>"001011010",
  9505=>"100110111",
  9506=>"010000010",
  9507=>"100110110",
  9508=>"101110111",
  9509=>"001101100",
  9510=>"001000011",
  9511=>"101101110",
  9512=>"011011100",
  9513=>"100100111",
  9514=>"101110110",
  9515=>"000111000",
  9516=>"011001111",
  9517=>"000001011",
  9518=>"111101110",
  9519=>"100110110",
  9520=>"010000100",
  9521=>"110011111",
  9522=>"111000001",
  9523=>"010100000",
  9524=>"000011001",
  9525=>"000000110",
  9526=>"110000001",
  9527=>"000101101",
  9528=>"011010101",
  9529=>"100110001",
  9530=>"101111010",
  9531=>"110100111",
  9532=>"100110010",
  9533=>"100100100",
  9534=>"101001010",
  9535=>"001001001",
  9536=>"111100001",
  9537=>"011011011",
  9538=>"111100111",
  9539=>"001000000",
  9540=>"001011010",
  9541=>"011011100",
  9542=>"001001010",
  9543=>"100111100",
  9544=>"000000001",
  9545=>"100000111",
  9546=>"101000110",
  9547=>"000010001",
  9548=>"100100101",
  9549=>"000010010",
  9550=>"000001100",
  9551=>"010001011",
  9552=>"010110101",
  9553=>"001110000",
  9554=>"001001100",
  9555=>"110101111",
  9556=>"100110000",
  9557=>"010111101",
  9558=>"000100110",
  9559=>"111111101",
  9560=>"011001001",
  9561=>"100111001",
  9562=>"001000011",
  9563=>"100010001",
  9564=>"000010011",
  9565=>"000111011",
  9566=>"101110001",
  9567=>"111000000",
  9568=>"001010111",
  9569=>"101101011",
  9570=>"000000000",
  9571=>"010010001",
  9572=>"010000111",
  9573=>"111111010",
  9574=>"001100010",
  9575=>"010010000",
  9576=>"011101000",
  9577=>"001011011",
  9578=>"000101010",
  9579=>"001100100",
  9580=>"010111010",
  9581=>"111101100",
  9582=>"001010010",
  9583=>"011100000",
  9584=>"101101110",
  9585=>"110001010",
  9586=>"110001111",
  9587=>"101100000",
  9588=>"010011001",
  9589=>"100010010",
  9590=>"010000001",
  9591=>"001101101",
  9592=>"111000111",
  9593=>"101001101",
  9594=>"011011101",
  9595=>"110101000",
  9596=>"000001110",
  9597=>"000001010",
  9598=>"110111101",
  9599=>"101010110",
  9600=>"010100110",
  9601=>"000000010",
  9602=>"110011010",
  9603=>"010101010",
  9604=>"010100101",
  9605=>"010000001",
  9606=>"111000010",
  9607=>"010001001",
  9608=>"000011011",
  9609=>"111101011",
  9610=>"110011110",
  9611=>"000001011",
  9612=>"111101010",
  9613=>"101000000",
  9614=>"010011001",
  9615=>"000101011",
  9616=>"001111111",
  9617=>"000001001",
  9618=>"001000010",
  9619=>"000010100",
  9620=>"100000100",
  9621=>"100100000",
  9622=>"111101111",
  9623=>"101001010",
  9624=>"101001110",
  9625=>"101000101",
  9626=>"010011011",
  9627=>"001001101",
  9628=>"111111101",
  9629=>"111111111",
  9630=>"010011010",
  9631=>"011111000",
  9632=>"011101110",
  9633=>"101111110",
  9634=>"011101100",
  9635=>"011011101",
  9636=>"101101000",
  9637=>"101100101",
  9638=>"000111010",
  9639=>"011101010",
  9640=>"001011100",
  9641=>"010101110",
  9642=>"011101000",
  9643=>"000111010",
  9644=>"000010010",
  9645=>"010001111",
  9646=>"110011010",
  9647=>"000001111",
  9648=>"100000100",
  9649=>"001010011",
  9650=>"011111111",
  9651=>"111000110",
  9652=>"101111110",
  9653=>"100101010",
  9654=>"111110111",
  9655=>"000101010",
  9656=>"010110001",
  9657=>"001111100",
  9658=>"111101101",
  9659=>"101110001",
  9660=>"010101010",
  9661=>"111011101",
  9662=>"001110111",
  9663=>"010101010",
  9664=>"000010011",
  9665=>"001101100",
  9666=>"110010110",
  9667=>"011100011",
  9668=>"000000001",
  9669=>"101011111",
  9670=>"100010010",
  9671=>"000100001",
  9672=>"010110100",
  9673=>"010110010",
  9674=>"011001010",
  9675=>"000111110",
  9676=>"100110010",
  9677=>"111101001",
  9678=>"011111111",
  9679=>"000111001",
  9680=>"000100111",
  9681=>"111011010",
  9682=>"001011111",
  9683=>"010100110",
  9684=>"000111011",
  9685=>"000100011",
  9686=>"010010000",
  9687=>"101000111",
  9688=>"001111011",
  9689=>"000001111",
  9690=>"010111011",
  9691=>"101110010",
  9692=>"111001001",
  9693=>"100010101",
  9694=>"001000011",
  9695=>"001001101",
  9696=>"010010101",
  9697=>"000010110",
  9698=>"110111101",
  9699=>"010100101",
  9700=>"000001000",
  9701=>"111111011",
  9702=>"110110010",
  9703=>"010010111",
  9704=>"001011010",
  9705=>"111011111",
  9706=>"000101001",
  9707=>"110101010",
  9708=>"110011111",
  9709=>"000111101",
  9710=>"000100001",
  9711=>"110000001",
  9712=>"011001010",
  9713=>"010111001",
  9714=>"110111101",
  9715=>"001111111",
  9716=>"000000001",
  9717=>"100100110",
  9718=>"010011001",
  9719=>"111101001",
  9720=>"010000000",
  9721=>"010001100",
  9722=>"111111010",
  9723=>"111000000",
  9724=>"111111100",
  9725=>"111011100",
  9726=>"111101011",
  9727=>"000001111",
  9728=>"010010010",
  9729=>"110001111",
  9730=>"000011010",
  9731=>"000010100",
  9732=>"010010110",
  9733=>"100111110",
  9734=>"100100010",
  9735=>"000100011",
  9736=>"011001100",
  9737=>"000100100",
  9738=>"000101000",
  9739=>"000011100",
  9740=>"101010111",
  9741=>"001001100",
  9742=>"000111010",
  9743=>"011000001",
  9744=>"100101010",
  9745=>"010000100",
  9746=>"000111010",
  9747=>"101001011",
  9748=>"001000111",
  9749=>"101010001",
  9750=>"110101011",
  9751=>"001101011",
  9752=>"101001000",
  9753=>"001000101",
  9754=>"111011010",
  9755=>"100000110",
  9756=>"111111111",
  9757=>"111101110",
  9758=>"010100111",
  9759=>"010100101",
  9760=>"010010010",
  9761=>"101101100",
  9762=>"001100100",
  9763=>"110100011",
  9764=>"010011011",
  9765=>"110110111",
  9766=>"101101010",
  9767=>"010010001",
  9768=>"011110101",
  9769=>"001110100",
  9770=>"100010010",
  9771=>"011000000",
  9772=>"101100001",
  9773=>"000011110",
  9774=>"001000100",
  9775=>"001111001",
  9776=>"111011000",
  9777=>"010011100",
  9778=>"101101111",
  9779=>"001100110",
  9780=>"001000011",
  9781=>"010100001",
  9782=>"110010011",
  9783=>"100111111",
  9784=>"101101110",
  9785=>"010111101",
  9786=>"100010110",
  9787=>"001000111",
  9788=>"111101011",
  9789=>"000111101",
  9790=>"011001011",
  9791=>"001001101",
  9792=>"000111000",
  9793=>"001001111",
  9794=>"000011011",
  9795=>"101010001",
  9796=>"111011101",
  9797=>"111010001",
  9798=>"000111101",
  9799=>"000101001",
  9800=>"101000000",
  9801=>"110001010",
  9802=>"010110110",
  9803=>"111101100",
  9804=>"011101011",
  9805=>"101100100",
  9806=>"000011011",
  9807=>"010010001",
  9808=>"100001000",
  9809=>"100000010",
  9810=>"000101110",
  9811=>"000011000",
  9812=>"010110101",
  9813=>"000110101",
  9814=>"001101111",
  9815=>"100110001",
  9816=>"011101010",
  9817=>"111000101",
  9818=>"110000111",
  9819=>"100101101",
  9820=>"000011011",
  9821=>"011000000",
  9822=>"001111101",
  9823=>"101101100",
  9824=>"111110111",
  9825=>"000111110",
  9826=>"001111111",
  9827=>"110001101",
  9828=>"011101001",
  9829=>"110111111",
  9830=>"101000111",
  9831=>"000010110",
  9832=>"000000000",
  9833=>"011010100",
  9834=>"111100000",
  9835=>"001111001",
  9836=>"111101001",
  9837=>"110100101",
  9838=>"100110100",
  9839=>"110001111",
  9840=>"111100111",
  9841=>"000101100",
  9842=>"000011000",
  9843=>"001001100",
  9844=>"100001011",
  9845=>"000110100",
  9846=>"011000001",
  9847=>"000010011",
  9848=>"101000010",
  9849=>"101110000",
  9850=>"101111010",
  9851=>"111101010",
  9852=>"001000010",
  9853=>"111000111",
  9854=>"000100000",
  9855=>"110111101",
  9856=>"001010100",
  9857=>"010101101",
  9858=>"111000110",
  9859=>"000000000",
  9860=>"000100111",
  9861=>"101010001",
  9862=>"101010000",
  9863=>"100101001",
  9864=>"011000100",
  9865=>"000100010",
  9866=>"110100001",
  9867=>"000010000",
  9868=>"010111011",
  9869=>"011001000",
  9870=>"100011001",
  9871=>"111100010",
  9872=>"111001010",
  9873=>"101101000",
  9874=>"011100100",
  9875=>"000100000",
  9876=>"010000000",
  9877=>"101111011",
  9878=>"101010100",
  9879=>"111001000",
  9880=>"110001010",
  9881=>"101000011",
  9882=>"101101010",
  9883=>"010111111",
  9884=>"010101001",
  9885=>"111100101",
  9886=>"111110100",
  9887=>"001011110",
  9888=>"011010000",
  9889=>"010001011",
  9890=>"110100100",
  9891=>"110100011",
  9892=>"111100100",
  9893=>"111010010",
  9894=>"000010011",
  9895=>"000000100",
  9896=>"110111010",
  9897=>"010100000",
  9898=>"101011110",
  9899=>"110010011",
  9900=>"111000011",
  9901=>"000011100",
  9902=>"101100000",
  9903=>"110011110",
  9904=>"100000110",
  9905=>"000111011",
  9906=>"100011000",
  9907=>"010100111",
  9908=>"110101011",
  9909=>"001100010",
  9910=>"010011100",
  9911=>"010011110",
  9912=>"111011110",
  9913=>"001000110",
  9914=>"111111111",
  9915=>"100110001",
  9916=>"001100010",
  9917=>"110101010",
  9918=>"001101101",
  9919=>"100111100",
  9920=>"110111111",
  9921=>"101100000",
  9922=>"000001101",
  9923=>"010011000",
  9924=>"110110111",
  9925=>"000010010",
  9926=>"000100010",
  9927=>"110011001",
  9928=>"100111100",
  9929=>"001010101",
  9930=>"100110000",
  9931=>"110000001",
  9932=>"101100110",
  9933=>"000101001",
  9934=>"001000111",
  9935=>"011000000",
  9936=>"000100011",
  9937=>"011001110",
  9938=>"001010010",
  9939=>"011000110",
  9940=>"101000000",
  9941=>"000001110",
  9942=>"110110100",
  9943=>"111010001",
  9944=>"000010111",
  9945=>"011100111",
  9946=>"000110100",
  9947=>"000111100",
  9948=>"010000110",
  9949=>"111101011",
  9950=>"011101101",
  9951=>"000000000",
  9952=>"000010000",
  9953=>"010111001",
  9954=>"000010000",
  9955=>"001111111",
  9956=>"111111101",
  9957=>"110110000",
  9958=>"110001100",
  9959=>"100001100",
  9960=>"101011010",
  9961=>"010010110",
  9962=>"111010101",
  9963=>"011010101",
  9964=>"110000001",
  9965=>"000010011",
  9966=>"101111101",
  9967=>"001001000",
  9968=>"110010000",
  9969=>"010011000",
  9970=>"111101111",
  9971=>"010010011",
  9972=>"110101101",
  9973=>"000101010",
  9974=>"001111001",
  9975=>"101111111",
  9976=>"001010001",
  9977=>"011010110",
  9978=>"010001010",
  9979=>"101000111",
  9980=>"110011001",
  9981=>"001001000",
  9982=>"101001010",
  9983=>"101001101",
  9984=>"011111111",
  9985=>"110111011",
  9986=>"011001010",
  9987=>"000001001",
  9988=>"000100001",
  9989=>"000100111",
  9990=>"000001100",
  9991=>"110110011",
  9992=>"110011111",
  9993=>"001111000",
  9994=>"100111011",
  9995=>"110100110",
  9996=>"000101111",
  9997=>"110100000",
  9998=>"011100001",
  9999=>"000000010",
  10000=>"010101110",
  10001=>"001000111",
  10002=>"001111100",
  10003=>"010011011",
  10004=>"010111101",
  10005=>"011000010",
  10006=>"110111001",
  10007=>"111010110",
  10008=>"110110010",
  10009=>"110101000",
  10010=>"001000100",
  10011=>"100001010",
  10012=>"010000001",
  10013=>"000010111",
  10014=>"000101101",
  10015=>"001010101",
  10016=>"101010010",
  10017=>"111100111",
  10018=>"011010100",
  10019=>"110011101",
  10020=>"011011001",
  10021=>"101000111",
  10022=>"000011001",
  10023=>"001100110",
  10024=>"000010111",
  10025=>"000110010",
  10026=>"100010111",
  10027=>"001011010",
  10028=>"010011010",
  10029=>"001000101",
  10030=>"111111101",
  10031=>"111110011",
  10032=>"101110011",
  10033=>"101101101",
  10034=>"110000001",
  10035=>"101111001",
  10036=>"010011011",
  10037=>"100011111",
  10038=>"111101100",
  10039=>"111000110",
  10040=>"111111111",
  10041=>"011010010",
  10042=>"100110000",
  10043=>"111100111",
  10044=>"001100110",
  10045=>"011110110",
  10046=>"110011100",
  10047=>"010010011",
  10048=>"111100100",
  10049=>"011011010",
  10050=>"010111111",
  10051=>"111100000",
  10052=>"000100000",
  10053=>"110100010",
  10054=>"010000001",
  10055=>"101110101",
  10056=>"000001000",
  10057=>"111110110",
  10058=>"101111111",
  10059=>"111000000",
  10060=>"111100101",
  10061=>"101000001",
  10062=>"100001001",
  10063=>"000011000",
  10064=>"011011001",
  10065=>"000100100",
  10066=>"000110001",
  10067=>"000110101",
  10068=>"011110011",
  10069=>"101110110",
  10070=>"010010101",
  10071=>"000001000",
  10072=>"001100101",
  10073=>"100010010",
  10074=>"010000011",
  10075=>"001100110",
  10076=>"110100100",
  10077=>"111101001",
  10078=>"110010010",
  10079=>"101110001",
  10080=>"100101001",
  10081=>"100101001",
  10082=>"010000000",
  10083=>"001010010",
  10084=>"010111100",
  10085=>"111000010",
  10086=>"001101111",
  10087=>"010110111",
  10088=>"010001101",
  10089=>"101001010",
  10090=>"101111111",
  10091=>"100111101",
  10092=>"110100001",
  10093=>"000101010",
  10094=>"100001110",
  10095=>"111111100",
  10096=>"000100011",
  10097=>"000110000",
  10098=>"100010101",
  10099=>"110100100",
  10100=>"000011100",
  10101=>"101001000",
  10102=>"000010000",
  10103=>"101110110",
  10104=>"011000000",
  10105=>"011100110",
  10106=>"011110001",
  10107=>"011111100",
  10108=>"101000000",
  10109=>"111101110",
  10110=>"101010111",
  10111=>"100100001",
  10112=>"111101101",
  10113=>"111110011",
  10114=>"100001010",
  10115=>"111101100",
  10116=>"010000001",
  10117=>"001000100",
  10118=>"110000000",
  10119=>"110000111",
  10120=>"101110001",
  10121=>"001110101",
  10122=>"001100001",
  10123=>"111111010",
  10124=>"110001010",
  10125=>"001011110",
  10126=>"110000101",
  10127=>"011111001",
  10128=>"100000110",
  10129=>"111111010",
  10130=>"000001000",
  10131=>"010100010",
  10132=>"100110011",
  10133=>"000010110",
  10134=>"000010101",
  10135=>"000001111",
  10136=>"110101101",
  10137=>"000111000",
  10138=>"101111110",
  10139=>"001101101",
  10140=>"000111011",
  10141=>"100100111",
  10142=>"000001010",
  10143=>"010001001",
  10144=>"011100000",
  10145=>"110111011",
  10146=>"001000001",
  10147=>"001000010",
  10148=>"010001111",
  10149=>"110011011",
  10150=>"010111110",
  10151=>"110010000",
  10152=>"000110001",
  10153=>"000010000",
  10154=>"010010110",
  10155=>"001101101",
  10156=>"100110100",
  10157=>"100110001",
  10158=>"011101010",
  10159=>"000011001",
  10160=>"010110000",
  10161=>"111111101",
  10162=>"101010110",
  10163=>"100010101",
  10164=>"010110000",
  10165=>"000001011",
  10166=>"110100010",
  10167=>"111100000",
  10168=>"001001011",
  10169=>"000111010",
  10170=>"001011111",
  10171=>"011010100",
  10172=>"000001000",
  10173=>"010010010",
  10174=>"110111101",
  10175=>"101001101",
  10176=>"000111000",
  10177=>"100001011",
  10178=>"010110010",
  10179=>"001011011",
  10180=>"101000000",
  10181=>"000001001",
  10182=>"010101000",
  10183=>"001100000",
  10184=>"101100011",
  10185=>"111110111",
  10186=>"001111101",
  10187=>"011001101",
  10188=>"110010000",
  10189=>"011001000",
  10190=>"001011011",
  10191=>"111110000",
  10192=>"000010110",
  10193=>"111000011",
  10194=>"101010000",
  10195=>"110100000",
  10196=>"111101111",
  10197=>"000101110",
  10198=>"011000001",
  10199=>"000111110",
  10200=>"101110010",
  10201=>"000001100",
  10202=>"011110000",
  10203=>"001001011",
  10204=>"011100111",
  10205=>"101001000",
  10206=>"101010110",
  10207=>"110100101",
  10208=>"111010101",
  10209=>"110101100",
  10210=>"010100100",
  10211=>"010110110",
  10212=>"111100101",
  10213=>"000000010",
  10214=>"011001110",
  10215=>"101100010",
  10216=>"111011001",
  10217=>"101111010",
  10218=>"101111100",
  10219=>"010110010",
  10220=>"101101111",
  10221=>"101111011",
  10222=>"001010000",
  10223=>"110010001",
  10224=>"101111111",
  10225=>"100011001",
  10226=>"110101111",
  10227=>"010110110",
  10228=>"011000111",
  10229=>"111101101",
  10230=>"100110101",
  10231=>"110110100",
  10232=>"000110100",
  10233=>"001000110",
  10234=>"101111110",
  10235=>"111011011",
  10236=>"101111100",
  10237=>"101111001",
  10238=>"001010100",
  10239=>"001010110",
  10240=>"110101111",
  10241=>"001000101",
  10242=>"010101110",
  10243=>"010011111",
  10244=>"100110101",
  10245=>"001011000",
  10246=>"111100001",
  10247=>"000011110",
  10248=>"111101101",
  10249=>"101111111",
  10250=>"000001101",
  10251=>"101101111",
  10252=>"011101111",
  10253=>"011011001",
  10254=>"010100111",
  10255=>"001111111",
  10256=>"101000000",
  10257=>"110110111",
  10258=>"000110101",
  10259=>"110110011",
  10260=>"101110100",
  10261=>"100001010",
  10262=>"111011000",
  10263=>"100000010",
  10264=>"100001111",
  10265=>"000110000",
  10266=>"011001101",
  10267=>"000111000",
  10268=>"011100000",
  10269=>"110001001",
  10270=>"110011011",
  10271=>"110100110",
  10272=>"110001011",
  10273=>"000010001",
  10274=>"100000100",
  10275=>"000000000",
  10276=>"000000101",
  10277=>"101110101",
  10278=>"110110100",
  10279=>"011100111",
  10280=>"001001011",
  10281=>"001001011",
  10282=>"111001100",
  10283=>"001001101",
  10284=>"100111011",
  10285=>"001111101",
  10286=>"001101110",
  10287=>"000101010",
  10288=>"000000100",
  10289=>"010001011",
  10290=>"000001010",
  10291=>"000111011",
  10292=>"101110000",
  10293=>"100010010",
  10294=>"000001010",
  10295=>"101111111",
  10296=>"111010111",
  10297=>"011110001",
  10298=>"011111011",
  10299=>"010111100",
  10300=>"010011011",
  10301=>"000000011",
  10302=>"100101101",
  10303=>"101001001",
  10304=>"001010101",
  10305=>"101000111",
  10306=>"011001000",
  10307=>"011100000",
  10308=>"110101011",
  10309=>"111101001",
  10310=>"010111001",
  10311=>"100111010",
  10312=>"111110010",
  10313=>"101010010",
  10314=>"110010000",
  10315=>"001110001",
  10316=>"011010010",
  10317=>"101001010",
  10318=>"001001001",
  10319=>"100100111",
  10320=>"010011010",
  10321=>"110000111",
  10322=>"111111000",
  10323=>"010101000",
  10324=>"000001110",
  10325=>"001001110",
  10326=>"101001001",
  10327=>"000101100",
  10328=>"111001101",
  10329=>"111011110",
  10330=>"000011000",
  10331=>"000000100",
  10332=>"100001000",
  10333=>"011011111",
  10334=>"000101010",
  10335=>"101011000",
  10336=>"111011010",
  10337=>"000011010",
  10338=>"001011011",
  10339=>"011110010",
  10340=>"111010010",
  10341=>"100000101",
  10342=>"110100110",
  10343=>"100110111",
  10344=>"001101100",
  10345=>"100110000",
  10346=>"011011110",
  10347=>"010000111",
  10348=>"000000000",
  10349=>"000110001",
  10350=>"101001001",
  10351=>"010010000",
  10352=>"001001110",
  10353=>"011011111",
  10354=>"010110011",
  10355=>"001111111",
  10356=>"010010010",
  10357=>"110011111",
  10358=>"100000001",
  10359=>"001011000",
  10360=>"100110101",
  10361=>"101011100",
  10362=>"000001010",
  10363=>"100010110",
  10364=>"011001000",
  10365=>"101101011",
  10366=>"100000100",
  10367=>"111110000",
  10368=>"011101000",
  10369=>"001000100",
  10370=>"111100100",
  10371=>"111011101",
  10372=>"110000110",
  10373=>"010111010",
  10374=>"010110111",
  10375=>"110110110",
  10376=>"110001110",
  10377=>"111101010",
  10378=>"000011100",
  10379=>"000100111",
  10380=>"000011101",
  10381=>"110101111",
  10382=>"001111100",
  10383=>"110101010",
  10384=>"111101011",
  10385=>"100001001",
  10386=>"001001110",
  10387=>"010010110",
  10388=>"010011101",
  10389=>"001000000",
  10390=>"100100000",
  10391=>"101101111",
  10392=>"010001000",
  10393=>"100001101",
  10394=>"111000100",
  10395=>"101001000",
  10396=>"000111101",
  10397=>"111111010",
  10398=>"001100000",
  10399=>"010100110",
  10400=>"100011001",
  10401=>"100011101",
  10402=>"011111101",
  10403=>"000001111",
  10404=>"011100000",
  10405=>"101010000",
  10406=>"101101111",
  10407=>"010101100",
  10408=>"101010101",
  10409=>"000000001",
  10410=>"010000101",
  10411=>"111100010",
  10412=>"110011001",
  10413=>"110101110",
  10414=>"100011111",
  10415=>"100011011",
  10416=>"101001010",
  10417=>"001110101",
  10418=>"110010010",
  10419=>"100100110",
  10420=>"101111101",
  10421=>"100001100",
  10422=>"011001011",
  10423=>"100011110",
  10424=>"100000001",
  10425=>"101011001",
  10426=>"111100000",
  10427=>"001110100",
  10428=>"011110001",
  10429=>"101100010",
  10430=>"101101111",
  10431=>"100010101",
  10432=>"111010000",
  10433=>"110010100",
  10434=>"100011110",
  10435=>"010000001",
  10436=>"000010011",
  10437=>"110000010",
  10438=>"000101010",
  10439=>"010001111",
  10440=>"101110001",
  10441=>"100111000",
  10442=>"001101111",
  10443=>"100000000",
  10444=>"100011110",
  10445=>"010111000",
  10446=>"000000011",
  10447=>"111000001",
  10448=>"100010100",
  10449=>"100010101",
  10450=>"011111010",
  10451=>"010010100",
  10452=>"000010000",
  10453=>"111110010",
  10454=>"011001110",
  10455=>"111111111",
  10456=>"101001110",
  10457=>"000000111",
  10458=>"010111001",
  10459=>"110011011",
  10460=>"111011000",
  10461=>"111001001",
  10462=>"011101001",
  10463=>"111110110",
  10464=>"000110110",
  10465=>"001110100",
  10466=>"101001100",
  10467=>"011000110",
  10468=>"111010110",
  10469=>"010000001",
  10470=>"101100111",
  10471=>"001010100",
  10472=>"010111011",
  10473=>"111010010",
  10474=>"100010011",
  10475=>"101111001",
  10476=>"100110001",
  10477=>"010101110",
  10478=>"111100101",
  10479=>"100100000",
  10480=>"011100101",
  10481=>"110110011",
  10482=>"110011001",
  10483=>"101001001",
  10484=>"111011101",
  10485=>"010001010",
  10486=>"100011000",
  10487=>"100110111",
  10488=>"111001001",
  10489=>"000100000",
  10490=>"100100100",
  10491=>"100011011",
  10492=>"100010100",
  10493=>"101010001",
  10494=>"100000010",
  10495=>"010110101",
  10496=>"010110011",
  10497=>"100011101",
  10498=>"100010001",
  10499=>"111111100",
  10500=>"111101011",
  10501=>"101000101",
  10502=>"001100111",
  10503=>"101111100",
  10504=>"111100100",
  10505=>"111110010",
  10506=>"011101101",
  10507=>"000011010",
  10508=>"000100010",
  10509=>"000000000",
  10510=>"101001101",
  10511=>"110011111",
  10512=>"001111110",
  10513=>"110010101",
  10514=>"101010000",
  10515=>"001101110",
  10516=>"010000111",
  10517=>"010100100",
  10518=>"010010011",
  10519=>"000110111",
  10520=>"101100000",
  10521=>"001000100",
  10522=>"010111000",
  10523=>"111011111",
  10524=>"010110000",
  10525=>"101100101",
  10526=>"110101001",
  10527=>"000101011",
  10528=>"000010111",
  10529=>"011000010",
  10530=>"101000111",
  10531=>"100101110",
  10532=>"010110010",
  10533=>"110011001",
  10534=>"000111110",
  10535=>"011111100",
  10536=>"110101011",
  10537=>"111101001",
  10538=>"100010101",
  10539=>"110101000",
  10540=>"110101010",
  10541=>"011011010",
  10542=>"111000001",
  10543=>"010101111",
  10544=>"001101010",
  10545=>"000110001",
  10546=>"111110101",
  10547=>"111001010",
  10548=>"011000011",
  10549=>"111011100",
  10550=>"000111011",
  10551=>"001001001",
  10552=>"010000011",
  10553=>"000010000",
  10554=>"111010111",
  10555=>"000000101",
  10556=>"100101011",
  10557=>"101001010",
  10558=>"111101001",
  10559=>"111011110",
  10560=>"000101100",
  10561=>"001110111",
  10562=>"011101110",
  10563=>"101011001",
  10564=>"010010000",
  10565=>"111101011",
  10566=>"111111000",
  10567=>"001000000",
  10568=>"111110000",
  10569=>"100101111",
  10570=>"001100001",
  10571=>"101110011",
  10572=>"110010011",
  10573=>"000100001",
  10574=>"011110100",
  10575=>"111111110",
  10576=>"001101011",
  10577=>"101110001",
  10578=>"010111011",
  10579=>"110011011",
  10580=>"001011000",
  10581=>"001111000",
  10582=>"100001101",
  10583=>"010010100",
  10584=>"100011110",
  10585=>"011000010",
  10586=>"011100000",
  10587=>"100101000",
  10588=>"111010101",
  10589=>"101001101",
  10590=>"000010111",
  10591=>"111110111",
  10592=>"100000000",
  10593=>"100000110",
  10594=>"011110011",
  10595=>"001001011",
  10596=>"100110001",
  10597=>"100100010",
  10598=>"100000111",
  10599=>"101100100",
  10600=>"001011010",
  10601=>"001110000",
  10602=>"000010000",
  10603=>"100000100",
  10604=>"011101101",
  10605=>"111010000",
  10606=>"001001100",
  10607=>"000110000",
  10608=>"011010010",
  10609=>"010101111",
  10610=>"100111000",
  10611=>"011101100",
  10612=>"111111101",
  10613=>"000011011",
  10614=>"111000111",
  10615=>"000001000",
  10616=>"101111101",
  10617=>"100010100",
  10618=>"110101111",
  10619=>"001001010",
  10620=>"011101011",
  10621=>"001001011",
  10622=>"101000010",
  10623=>"100000001",
  10624=>"000101111",
  10625=>"100111001",
  10626=>"000101010",
  10627=>"010111110",
  10628=>"110100101",
  10629=>"100010111",
  10630=>"111010110",
  10631=>"110100111",
  10632=>"011100111",
  10633=>"110000111",
  10634=>"001110111",
  10635=>"101111000",
  10636=>"111010110",
  10637=>"010110001",
  10638=>"010011100",
  10639=>"111110000",
  10640=>"000111100",
  10641=>"100110011",
  10642=>"110001010",
  10643=>"111100111",
  10644=>"111111101",
  10645=>"000100111",
  10646=>"011001111",
  10647=>"111011100",
  10648=>"101001101",
  10649=>"011100111",
  10650=>"011000110",
  10651=>"110011111",
  10652=>"001011110",
  10653=>"000110101",
  10654=>"111111010",
  10655=>"101101100",
  10656=>"100101011",
  10657=>"110000000",
  10658=>"101101111",
  10659=>"010000000",
  10660=>"110101000",
  10661=>"110101001",
  10662=>"100011011",
  10663=>"111001001",
  10664=>"110100101",
  10665=>"111011001",
  10666=>"000101111",
  10667=>"010011110",
  10668=>"100001011",
  10669=>"011100111",
  10670=>"110111101",
  10671=>"111100111",
  10672=>"101101001",
  10673=>"100110011",
  10674=>"101111001",
  10675=>"001011100",
  10676=>"010111000",
  10677=>"001001000",
  10678=>"111001101",
  10679=>"100100001",
  10680=>"100000100",
  10681=>"111000101",
  10682=>"000000111",
  10683=>"100011000",
  10684=>"110001011",
  10685=>"110001001",
  10686=>"001011101",
  10687=>"011010111",
  10688=>"111100110",
  10689=>"101011000",
  10690=>"111101010",
  10691=>"100100011",
  10692=>"010100010",
  10693=>"101111001",
  10694=>"110001000",
  10695=>"010110011",
  10696=>"111011101",
  10697=>"001101001",
  10698=>"000010010",
  10699=>"101011100",
  10700=>"011111110",
  10701=>"010011011",
  10702=>"101011011",
  10703=>"111011110",
  10704=>"011011100",
  10705=>"000000010",
  10706=>"010101100",
  10707=>"011100110",
  10708=>"100111001",
  10709=>"100101100",
  10710=>"011001011",
  10711=>"100101100",
  10712=>"101111101",
  10713=>"101001101",
  10714=>"111010101",
  10715=>"001010101",
  10716=>"000110011",
  10717=>"000010001",
  10718=>"110011001",
  10719=>"001001101",
  10720=>"111000000",
  10721=>"110010011",
  10722=>"100000101",
  10723=>"110001011",
  10724=>"000010010",
  10725=>"010000101",
  10726=>"001001010",
  10727=>"010111010",
  10728=>"110110001",
  10729=>"000100100",
  10730=>"101000000",
  10731=>"010000010",
  10732=>"111001000",
  10733=>"100010010",
  10734=>"100001001",
  10735=>"111011111",
  10736=>"100100001",
  10737=>"111010011",
  10738=>"111100011",
  10739=>"011110100",
  10740=>"011100101",
  10741=>"100100001",
  10742=>"110011010",
  10743=>"011111000",
  10744=>"000010101",
  10745=>"101011110",
  10746=>"111000111",
  10747=>"110110001",
  10748=>"010111101",
  10749=>"000011111",
  10750=>"010101111",
  10751=>"110110011",
  10752=>"100000000",
  10753=>"000001000",
  10754=>"010011011",
  10755=>"010011111",
  10756=>"000001101",
  10757=>"100101101",
  10758=>"100110111",
  10759=>"011111000",
  10760=>"011011001",
  10761=>"001000101",
  10762=>"011111110",
  10763=>"010000011",
  10764=>"100111011",
  10765=>"010011000",
  10766=>"000001110",
  10767=>"101111111",
  10768=>"011000110",
  10769=>"001001010",
  10770=>"000010110",
  10771=>"100000111",
  10772=>"101010101",
  10773=>"100010010",
  10774=>"111101111",
  10775=>"001000100",
  10776=>"100001101",
  10777=>"011100000",
  10778=>"001110100",
  10779=>"101011000",
  10780=>"111000010",
  10781=>"001101001",
  10782=>"010110011",
  10783=>"000010100",
  10784=>"000100001",
  10785=>"011001010",
  10786=>"000011110",
  10787=>"110011000",
  10788=>"000010110",
  10789=>"011100001",
  10790=>"011110010",
  10791=>"101010111",
  10792=>"101110100",
  10793=>"101011110",
  10794=>"011010111",
  10795=>"011110111",
  10796=>"101000101",
  10797=>"000000011",
  10798=>"110110011",
  10799=>"000101111",
  10800=>"000011100",
  10801=>"110001101",
  10802=>"101110010",
  10803=>"110111110",
  10804=>"111101100",
  10805=>"110111110",
  10806=>"011110100",
  10807=>"001011011",
  10808=>"111111011",
  10809=>"100101110",
  10810=>"101101100",
  10811=>"001110011",
  10812=>"111111001",
  10813=>"010111111",
  10814=>"100010010",
  10815=>"100100000",
  10816=>"111011111",
  10817=>"110101110",
  10818=>"001001011",
  10819=>"000011011",
  10820=>"011010110",
  10821=>"001000010",
  10822=>"000100111",
  10823=>"001100110",
  10824=>"001101110",
  10825=>"000111000",
  10826=>"000000100",
  10827=>"100110101",
  10828=>"011010100",
  10829=>"000110111",
  10830=>"110000110",
  10831=>"110100011",
  10832=>"101100010",
  10833=>"110111110",
  10834=>"000001101",
  10835=>"100000010",
  10836=>"011100111",
  10837=>"011101110",
  10838=>"110111011",
  10839=>"010100011",
  10840=>"101011101",
  10841=>"111110001",
  10842=>"110100010",
  10843=>"110111110",
  10844=>"010000001",
  10845=>"101000110",
  10846=>"110101100",
  10847=>"010010101",
  10848=>"110111011",
  10849=>"001111110",
  10850=>"110010100",
  10851=>"100111100",
  10852=>"000000000",
  10853=>"110111011",
  10854=>"010000001",
  10855=>"000110101",
  10856=>"000110011",
  10857=>"000101010",
  10858=>"000100000",
  10859=>"010001101",
  10860=>"100011110",
  10861=>"011111111",
  10862=>"011111011",
  10863=>"111010111",
  10864=>"000011000",
  10865=>"001111000",
  10866=>"100011000",
  10867=>"000000010",
  10868=>"001001010",
  10869=>"010100110",
  10870=>"111000001",
  10871=>"101111011",
  10872=>"011001100",
  10873=>"001011111",
  10874=>"011000101",
  10875=>"111111001",
  10876=>"100110111",
  10877=>"011111000",
  10878=>"101011000",
  10879=>"111100101",
  10880=>"000000110",
  10881=>"110101110",
  10882=>"010110010",
  10883=>"111011110",
  10884=>"100011011",
  10885=>"100010110",
  10886=>"101010011",
  10887=>"001000110",
  10888=>"001000100",
  10889=>"110110011",
  10890=>"001100111",
  10891=>"000011101",
  10892=>"001111110",
  10893=>"100101101",
  10894=>"101101001",
  10895=>"100100111",
  10896=>"101001110",
  10897=>"001001100",
  10898=>"101001110",
  10899=>"100111111",
  10900=>"101111010",
  10901=>"010011101",
  10902=>"111111111",
  10903=>"000011100",
  10904=>"110000011",
  10905=>"111101010",
  10906=>"111000100",
  10907=>"101111010",
  10908=>"000000110",
  10909=>"111110001",
  10910=>"000010010",
  10911=>"110100000",
  10912=>"100110100",
  10913=>"011011001",
  10914=>"100110101",
  10915=>"011111111",
  10916=>"001010100",
  10917=>"100100010",
  10918=>"111111010",
  10919=>"001001111",
  10920=>"011110000",
  10921=>"010111001",
  10922=>"110101000",
  10923=>"000110111",
  10924=>"010100110",
  10925=>"010000001",
  10926=>"010111000",
  10927=>"011011011",
  10928=>"110111010",
  10929=>"000010000",
  10930=>"110011010",
  10931=>"100011101",
  10932=>"001010101",
  10933=>"000100001",
  10934=>"111011101",
  10935=>"110111001",
  10936=>"011100101",
  10937=>"100101111",
  10938=>"011010000",
  10939=>"000100101",
  10940=>"101000110",
  10941=>"100010111",
  10942=>"010010101",
  10943=>"100100111",
  10944=>"111001110",
  10945=>"101111111",
  10946=>"000000011",
  10947=>"101100000",
  10948=>"101100110",
  10949=>"011110100",
  10950=>"011010100",
  10951=>"101010110",
  10952=>"100011011",
  10953=>"011111001",
  10954=>"010110100",
  10955=>"101000001",
  10956=>"110111001",
  10957=>"011010000",
  10958=>"000001001",
  10959=>"100101111",
  10960=>"011101000",
  10961=>"000011001",
  10962=>"101100001",
  10963=>"100110110",
  10964=>"100101000",
  10965=>"011100100",
  10966=>"011110001",
  10967=>"010110110",
  10968=>"000111100",
  10969=>"101101100",
  10970=>"010000001",
  10971=>"111010011",
  10972=>"000110001",
  10973=>"101011001",
  10974=>"100001011",
  10975=>"011011001",
  10976=>"010011110",
  10977=>"100000110",
  10978=>"100111011",
  10979=>"110001100",
  10980=>"000110000",
  10981=>"011111110",
  10982=>"110011000",
  10983=>"000011011",
  10984=>"001001000",
  10985=>"101111101",
  10986=>"110101100",
  10987=>"110110111",
  10988=>"100100110",
  10989=>"101010000",
  10990=>"111000000",
  10991=>"110100110",
  10992=>"001011000",
  10993=>"111011111",
  10994=>"001011100",
  10995=>"100001101",
  10996=>"011110101",
  10997=>"001001000",
  10998=>"010000100",
  10999=>"110001010",
  11000=>"101100001",
  11001=>"011100110",
  11002=>"111000010",
  11003=>"010100001",
  11004=>"001011101",
  11005=>"001001000",
  11006=>"101100011",
  11007=>"111110011",
  11008=>"110111011",
  11009=>"100010110",
  11010=>"010011010",
  11011=>"001010001",
  11012=>"101000100",
  11013=>"101011110",
  11014=>"000010111",
  11015=>"000101111",
  11016=>"100001010",
  11017=>"101000000",
  11018=>"001000000",
  11019=>"110111000",
  11020=>"001001101",
  11021=>"010011001",
  11022=>"011111011",
  11023=>"001000100",
  11024=>"101100001",
  11025=>"100011010",
  11026=>"010101101",
  11027=>"100100011",
  11028=>"011010111",
  11029=>"101001101",
  11030=>"001100010",
  11031=>"100010101",
  11032=>"011001010",
  11033=>"000111111",
  11034=>"111111101",
  11035=>"101100001",
  11036=>"010000010",
  11037=>"111000110",
  11038=>"100001100",
  11039=>"001011111",
  11040=>"000100011",
  11041=>"100001000",
  11042=>"000001010",
  11043=>"110111001",
  11044=>"111000111",
  11045=>"010110100",
  11046=>"000110011",
  11047=>"110101010",
  11048=>"011000010",
  11049=>"010101000",
  11050=>"000001010",
  11051=>"001011111",
  11052=>"011000100",
  11053=>"000111101",
  11054=>"111011110",
  11055=>"010110000",
  11056=>"001101000",
  11057=>"101100001",
  11058=>"111000010",
  11059=>"101000111",
  11060=>"000000100",
  11061=>"111111111",
  11062=>"011110110",
  11063=>"000010010",
  11064=>"110011010",
  11065=>"100100110",
  11066=>"111010011",
  11067=>"101010001",
  11068=>"101001110",
  11069=>"000100100",
  11070=>"000000100",
  11071=>"000000111",
  11072=>"100111110",
  11073=>"010000100",
  11074=>"011011100",
  11075=>"001110010",
  11076=>"011011100",
  11077=>"111000100",
  11078=>"100101010",
  11079=>"000100110",
  11080=>"000010110",
  11081=>"111001100",
  11082=>"100010011",
  11083=>"100100010",
  11084=>"110010111",
  11085=>"110111101",
  11086=>"111100101",
  11087=>"010000000",
  11088=>"000010101",
  11089=>"100111100",
  11090=>"101000101",
  11091=>"100010100",
  11092=>"101001011",
  11093=>"011100010",
  11094=>"111001101",
  11095=>"011011110",
  11096=>"101010001",
  11097=>"011100011",
  11098=>"011011000",
  11099=>"110111010",
  11100=>"110000110",
  11101=>"110111011",
  11102=>"111011101",
  11103=>"000010100",
  11104=>"111011001",
  11105=>"011010010",
  11106=>"110101010",
  11107=>"110100110",
  11108=>"100101110",
  11109=>"110001100",
  11110=>"001100000",
  11111=>"001011111",
  11112=>"111011001",
  11113=>"100101111",
  11114=>"011000000",
  11115=>"100110110",
  11116=>"101111111",
  11117=>"011111101",
  11118=>"100000110",
  11119=>"000010000",
  11120=>"100101100",
  11121=>"001100110",
  11122=>"000110110",
  11123=>"101000010",
  11124=>"001110110",
  11125=>"010111100",
  11126=>"110010010",
  11127=>"000101011",
  11128=>"000101000",
  11129=>"111111000",
  11130=>"001101110",
  11131=>"101011100",
  11132=>"000000100",
  11133=>"000010000",
  11134=>"000010000",
  11135=>"110000110",
  11136=>"101110101",
  11137=>"000010001",
  11138=>"001001000",
  11139=>"111110101",
  11140=>"101100111",
  11141=>"100110111",
  11142=>"001101000",
  11143=>"010111100",
  11144=>"111110100",
  11145=>"111010000",
  11146=>"010110011",
  11147=>"011001010",
  11148=>"110111101",
  11149=>"000111101",
  11150=>"011110010",
  11151=>"001010101",
  11152=>"101101111",
  11153=>"110111111",
  11154=>"100000010",
  11155=>"001001110",
  11156=>"100001011",
  11157=>"001101010",
  11158=>"110100100",
  11159=>"100111111",
  11160=>"110101011",
  11161=>"010110100",
  11162=>"110110110",
  11163=>"000110000",
  11164=>"000011100",
  11165=>"111110100",
  11166=>"101001001",
  11167=>"100010001",
  11168=>"010100001",
  11169=>"010010111",
  11170=>"101101101",
  11171=>"111111000",
  11172=>"000111010",
  11173=>"011111001",
  11174=>"010110110",
  11175=>"110011010",
  11176=>"010001100",
  11177=>"000010000",
  11178=>"101011110",
  11179=>"100010000",
  11180=>"111000011",
  11181=>"000100001",
  11182=>"101010010",
  11183=>"011110011",
  11184=>"001010000",
  11185=>"011011111",
  11186=>"010100000",
  11187=>"100110100",
  11188=>"111011110",
  11189=>"010101010",
  11190=>"100111110",
  11191=>"100010111",
  11192=>"111110110",
  11193=>"101011000",
  11194=>"110010011",
  11195=>"111000100",
  11196=>"000101000",
  11197=>"110010011",
  11198=>"001011000",
  11199=>"111101011",
  11200=>"100111100",
  11201=>"000010100",
  11202=>"110000100",
  11203=>"000010100",
  11204=>"000001101",
  11205=>"110111111",
  11206=>"010000101",
  11207=>"101101001",
  11208=>"010100001",
  11209=>"101100110",
  11210=>"001101111",
  11211=>"000100101",
  11212=>"101001001",
  11213=>"001111001",
  11214=>"101110001",
  11215=>"001110001",
  11216=>"000101001",
  11217=>"000000110",
  11218=>"111011000",
  11219=>"100101110",
  11220=>"110111110",
  11221=>"000000110",
  11222=>"001001111",
  11223=>"011100010",
  11224=>"100000111",
  11225=>"101100010",
  11226=>"011111011",
  11227=>"111011011",
  11228=>"100110101",
  11229=>"100100100",
  11230=>"110000001",
  11231=>"100001000",
  11232=>"111001000",
  11233=>"000110010",
  11234=>"001010110",
  11235=>"000100111",
  11236=>"110000110",
  11237=>"111000101",
  11238=>"101110000",
  11239=>"001100100",
  11240=>"010111110",
  11241=>"011100101",
  11242=>"000010111",
  11243=>"011101110",
  11244=>"101011111",
  11245=>"011101011",
  11246=>"110010011",
  11247=>"110001000",
  11248=>"000100101",
  11249=>"000010100",
  11250=>"001100101",
  11251=>"101011010",
  11252=>"100111110",
  11253=>"000000000",
  11254=>"010011110",
  11255=>"111101010",
  11256=>"110111110",
  11257=>"100000111",
  11258=>"000100001",
  11259=>"001010001",
  11260=>"011010111",
  11261=>"100011001",
  11262=>"110011000",
  11263=>"000001011",
  11264=>"000100010",
  11265=>"101100110",
  11266=>"011000111",
  11267=>"100010011",
  11268=>"111010100",
  11269=>"101101110",
  11270=>"011100010",
  11271=>"101111000",
  11272=>"011011010",
  11273=>"001001101",
  11274=>"001011011",
  11275=>"011101001",
  11276=>"010010000",
  11277=>"110111000",
  11278=>"100100110",
  11279=>"001010010",
  11280=>"100010110",
  11281=>"011111110",
  11282=>"110111000",
  11283=>"111101011",
  11284=>"100010100",
  11285=>"010100100",
  11286=>"001001010",
  11287=>"000011111",
  11288=>"111110001",
  11289=>"101110000",
  11290=>"010111111",
  11291=>"101010110",
  11292=>"011011000",
  11293=>"101000001",
  11294=>"011101111",
  11295=>"100110011",
  11296=>"000111010",
  11297=>"100001000",
  11298=>"101010111",
  11299=>"001001011",
  11300=>"000010001",
  11301=>"000010001",
  11302=>"011101110",
  11303=>"100000000",
  11304=>"111001000",
  11305=>"001011110",
  11306=>"110011101",
  11307=>"001010100",
  11308=>"011010011",
  11309=>"100001011",
  11310=>"101100001",
  11311=>"110010111",
  11312=>"111110000",
  11313=>"010101100",
  11314=>"100100101",
  11315=>"100100111",
  11316=>"000100101",
  11317=>"001000011",
  11318=>"111011111",
  11319=>"101110101",
  11320=>"001110100",
  11321=>"011000101",
  11322=>"110111100",
  11323=>"110011010",
  11324=>"010111011",
  11325=>"110111000",
  11326=>"100110001",
  11327=>"101010001",
  11328=>"001000010",
  11329=>"001111111",
  11330=>"111111010",
  11331=>"100101000",
  11332=>"111010111",
  11333=>"100000001",
  11334=>"001111100",
  11335=>"110101110",
  11336=>"100001100",
  11337=>"010011101",
  11338=>"110111100",
  11339=>"111111001",
  11340=>"010111000",
  11341=>"010000011",
  11342=>"110000001",
  11343=>"000010000",
  11344=>"000100011",
  11345=>"111111101",
  11346=>"101000111",
  11347=>"010000111",
  11348=>"110101010",
  11349=>"011000001",
  11350=>"100000110",
  11351=>"101100110",
  11352=>"110001011",
  11353=>"010110100",
  11354=>"011110100",
  11355=>"100110001",
  11356=>"000011001",
  11357=>"101101010",
  11358=>"101101001",
  11359=>"101001000",
  11360=>"110001000",
  11361=>"000111001",
  11362=>"110000101",
  11363=>"100000110",
  11364=>"101001011",
  11365=>"010011011",
  11366=>"011000110",
  11367=>"101010000",
  11368=>"100110111",
  11369=>"001111101",
  11370=>"111011111",
  11371=>"111010010",
  11372=>"110011110",
  11373=>"111100000",
  11374=>"001011001",
  11375=>"110101001",
  11376=>"110110111",
  11377=>"111101111",
  11378=>"110111011",
  11379=>"010111011",
  11380=>"101011010",
  11381=>"011101000",
  11382=>"100101100",
  11383=>"101101111",
  11384=>"110001000",
  11385=>"100011011",
  11386=>"000111011",
  11387=>"010000100",
  11388=>"110100000",
  11389=>"110110100",
  11390=>"010001010",
  11391=>"100101000",
  11392=>"001101110",
  11393=>"011101110",
  11394=>"000010010",
  11395=>"110010001",
  11396=>"000110110",
  11397=>"110110100",
  11398=>"101001010",
  11399=>"101000111",
  11400=>"000011010",
  11401=>"110011110",
  11402=>"101000110",
  11403=>"101100000",
  11404=>"011111111",
  11405=>"010111111",
  11406=>"000000001",
  11407=>"101111111",
  11408=>"000010101",
  11409=>"110001100",
  11410=>"100101010",
  11411=>"100010101",
  11412=>"111001110",
  11413=>"100001111",
  11414=>"000101110",
  11415=>"000011000",
  11416=>"001000010",
  11417=>"100100101",
  11418=>"000100100",
  11419=>"101101100",
  11420=>"110011110",
  11421=>"000001111",
  11422=>"110101101",
  11423=>"010110000",
  11424=>"011000000",
  11425=>"100111011",
  11426=>"001111101",
  11427=>"111111101",
  11428=>"101001011",
  11429=>"100000011",
  11430=>"011110110",
  11431=>"000101101",
  11432=>"001111100",
  11433=>"110001011",
  11434=>"111111001",
  11435=>"100110000",
  11436=>"101110001",
  11437=>"001111010",
  11438=>"101101011",
  11439=>"110100101",
  11440=>"101100110",
  11441=>"100110000",
  11442=>"010101001",
  11443=>"010010001",
  11444=>"010110100",
  11445=>"111010001",
  11446=>"100111110",
  11447=>"000110000",
  11448=>"111110111",
  11449=>"110111010",
  11450=>"100110001",
  11451=>"110101000",
  11452=>"010011010",
  11453=>"111010000",
  11454=>"111110111",
  11455=>"100000001",
  11456=>"011101111",
  11457=>"001000100",
  11458=>"101010111",
  11459=>"100111000",
  11460=>"010101001",
  11461=>"101111101",
  11462=>"101001000",
  11463=>"011111001",
  11464=>"000100011",
  11465=>"011101010",
  11466=>"101011101",
  11467=>"000001011",
  11468=>"001010111",
  11469=>"010011010",
  11470=>"111001110",
  11471=>"010001110",
  11472=>"001000000",
  11473=>"110010010",
  11474=>"000001000",
  11475=>"000101011",
  11476=>"000000111",
  11477=>"110100001",
  11478=>"100100000",
  11479=>"100110011",
  11480=>"000101001",
  11481=>"100111111",
  11482=>"101000110",
  11483=>"000101101",
  11484=>"111101001",
  11485=>"010010000",
  11486=>"010100110",
  11487=>"111011100",
  11488=>"110011101",
  11489=>"101011101",
  11490=>"001110110",
  11491=>"001010011",
  11492=>"000000010",
  11493=>"110111000",
  11494=>"100111010",
  11495=>"101111110",
  11496=>"111110001",
  11497=>"001110111",
  11498=>"000011110",
  11499=>"101101000",
  11500=>"110111110",
  11501=>"110011010",
  11502=>"101100110",
  11503=>"100011110",
  11504=>"010101111",
  11505=>"001100100",
  11506=>"110011010",
  11507=>"001000111",
  11508=>"111011110",
  11509=>"100000000",
  11510=>"110111110",
  11511=>"100101001",
  11512=>"000001101",
  11513=>"110001101",
  11514=>"110110111",
  11515=>"000001111",
  11516=>"001000011",
  11517=>"101111100",
  11518=>"000110010",
  11519=>"101011011",
  11520=>"110011000",
  11521=>"001001100",
  11522=>"110000101",
  11523=>"111011100",
  11524=>"001110101",
  11525=>"100001010",
  11526=>"100101001",
  11527=>"100001001",
  11528=>"111010010",
  11529=>"011000100",
  11530=>"001001010",
  11531=>"000110111",
  11532=>"100011110",
  11533=>"000011110",
  11534=>"111100110",
  11535=>"100111010",
  11536=>"101100011",
  11537=>"111111101",
  11538=>"010110011",
  11539=>"110111100",
  11540=>"010101100",
  11541=>"100000110",
  11542=>"110001100",
  11543=>"001010001",
  11544=>"011110010",
  11545=>"110010000",
  11546=>"111010001",
  11547=>"100010001",
  11548=>"010010000",
  11549=>"010110111",
  11550=>"110100110",
  11551=>"011111001",
  11552=>"111101010",
  11553=>"011011001",
  11554=>"100000011",
  11555=>"010101100",
  11556=>"111011000",
  11557=>"100101011",
  11558=>"111110110",
  11559=>"100110111",
  11560=>"011010100",
  11561=>"111001111",
  11562=>"000001011",
  11563=>"011011100",
  11564=>"010101000",
  11565=>"001100010",
  11566=>"110111111",
  11567=>"010000110",
  11568=>"010111111",
  11569=>"100000011",
  11570=>"000010000",
  11571=>"110010100",
  11572=>"011000110",
  11573=>"111100001",
  11574=>"011100010",
  11575=>"010011000",
  11576=>"011111001",
  11577=>"010000111",
  11578=>"110101111",
  11579=>"111001001",
  11580=>"111011111",
  11581=>"011001111",
  11582=>"010010111",
  11583=>"111001011",
  11584=>"110100001",
  11585=>"110100101",
  11586=>"001111110",
  11587=>"110011001",
  11588=>"100011110",
  11589=>"000011101",
  11590=>"011101100",
  11591=>"110101110",
  11592=>"011010111",
  11593=>"011011011",
  11594=>"111100011",
  11595=>"100111100",
  11596=>"100111011",
  11597=>"100010010",
  11598=>"110001101",
  11599=>"101000011",
  11600=>"111010101",
  11601=>"101011101",
  11602=>"000110110",
  11603=>"101101100",
  11604=>"101010000",
  11605=>"010010001",
  11606=>"001110110",
  11607=>"011111001",
  11608=>"001111111",
  11609=>"001011111",
  11610=>"001001101",
  11611=>"001001010",
  11612=>"100000000",
  11613=>"011111110",
  11614=>"100011001",
  11615=>"110000010",
  11616=>"001000101",
  11617=>"000101011",
  11618=>"111110010",
  11619=>"101110010",
  11620=>"001000100",
  11621=>"001001010",
  11622=>"111110111",
  11623=>"111000010",
  11624=>"100011000",
  11625=>"001101110",
  11626=>"001001110",
  11627=>"001110011",
  11628=>"100010100",
  11629=>"110001101",
  11630=>"100100010",
  11631=>"110010011",
  11632=>"110110110",
  11633=>"111001011",
  11634=>"100001011",
  11635=>"111100111",
  11636=>"110001011",
  11637=>"001111000",
  11638=>"001100011",
  11639=>"001100111",
  11640=>"101001001",
  11641=>"101110100",
  11642=>"010011110",
  11643=>"111001000",
  11644=>"101100001",
  11645=>"110101000",
  11646=>"110111000",
  11647=>"000101011",
  11648=>"000110101",
  11649=>"010000011",
  11650=>"000001110",
  11651=>"011101010",
  11652=>"110111011",
  11653=>"011011010",
  11654=>"010011011",
  11655=>"101100111",
  11656=>"110001000",
  11657=>"011100101",
  11658=>"000001011",
  11659=>"101110001",
  11660=>"000101011",
  11661=>"000001111",
  11662=>"100011111",
  11663=>"111001010",
  11664=>"001001010",
  11665=>"110110110",
  11666=>"011001101",
  11667=>"111111010",
  11668=>"100000000",
  11669=>"100011011",
  11670=>"100111111",
  11671=>"010111111",
  11672=>"110000111",
  11673=>"100101001",
  11674=>"010101110",
  11675=>"010010011",
  11676=>"110010101",
  11677=>"010010010",
  11678=>"000111010",
  11679=>"101111111",
  11680=>"111111101",
  11681=>"100011010",
  11682=>"010010101",
  11683=>"101100111",
  11684=>"011100111",
  11685=>"011010000",
  11686=>"001001111",
  11687=>"101100111",
  11688=>"110111000",
  11689=>"111001101",
  11690=>"100100010",
  11691=>"000000000",
  11692=>"111001110",
  11693=>"000001011",
  11694=>"101010010",
  11695=>"101100001",
  11696=>"110101011",
  11697=>"001011111",
  11698=>"000100111",
  11699=>"111111111",
  11700=>"000000000",
  11701=>"100000010",
  11702=>"110101111",
  11703=>"000010111",
  11704=>"001011000",
  11705=>"000011001",
  11706=>"000100010",
  11707=>"010010100",
  11708=>"100100001",
  11709=>"111110011",
  11710=>"111000001",
  11711=>"101110000",
  11712=>"011110101",
  11713=>"000000000",
  11714=>"101111111",
  11715=>"100010111",
  11716=>"000111011",
  11717=>"101111110",
  11718=>"100100000",
  11719=>"111010001",
  11720=>"100101101",
  11721=>"010100100",
  11722=>"001010001",
  11723=>"000001100",
  11724=>"110010000",
  11725=>"100001110",
  11726=>"001111000",
  11727=>"000010101",
  11728=>"010100110",
  11729=>"111010111",
  11730=>"010110000",
  11731=>"010001010",
  11732=>"011000001",
  11733=>"010001001",
  11734=>"001000010",
  11735=>"000100111",
  11736=>"101011010",
  11737=>"010100101",
  11738=>"010100010",
  11739=>"001110101",
  11740=>"110111011",
  11741=>"110010010",
  11742=>"010001111",
  11743=>"110101101",
  11744=>"111111111",
  11745=>"000110110",
  11746=>"110100110",
  11747=>"001101011",
  11748=>"010110000",
  11749=>"001110111",
  11750=>"100011111",
  11751=>"110010100",
  11752=>"111111101",
  11753=>"000111111",
  11754=>"110010010",
  11755=>"010101101",
  11756=>"010010011",
  11757=>"001100000",
  11758=>"111111100",
  11759=>"110000000",
  11760=>"111100110",
  11761=>"000011011",
  11762=>"010001110",
  11763=>"100000110",
  11764=>"110010000",
  11765=>"000111110",
  11766=>"110101001",
  11767=>"111000011",
  11768=>"111110000",
  11769=>"101010010",
  11770=>"101110110",
  11771=>"001011010",
  11772=>"111010101",
  11773=>"100001001",
  11774=>"010011101",
  11775=>"101111111",
  11776=>"110011100",
  11777=>"100001111",
  11778=>"011100011",
  11779=>"101101011",
  11780=>"011001100",
  11781=>"011100110",
  11782=>"101110110",
  11783=>"000001100",
  11784=>"111100011",
  11785=>"001001001",
  11786=>"111001000",
  11787=>"011001001",
  11788=>"101010101",
  11789=>"110100010",
  11790=>"000011011",
  11791=>"100000000",
  11792=>"001100011",
  11793=>"011110000",
  11794=>"101110101",
  11795=>"001010000",
  11796=>"011001000",
  11797=>"000101111",
  11798=>"110001010",
  11799=>"111111111",
  11800=>"111000100",
  11801=>"100111110",
  11802=>"101111100",
  11803=>"000000100",
  11804=>"000000010",
  11805=>"000001111",
  11806=>"111001000",
  11807=>"001100001",
  11808=>"110011111",
  11809=>"111001111",
  11810=>"111111111",
  11811=>"000111010",
  11812=>"000011000",
  11813=>"101011011",
  11814=>"000000000",
  11815=>"110010110",
  11816=>"010001010",
  11817=>"110011010",
  11818=>"100001000",
  11819=>"111110001",
  11820=>"100100001",
  11821=>"111001001",
  11822=>"010001001",
  11823=>"111000000",
  11824=>"001000000",
  11825=>"111111101",
  11826=>"110111100",
  11827=>"110011000",
  11828=>"001100010",
  11829=>"111111001",
  11830=>"100100011",
  11831=>"011000110",
  11832=>"000100011",
  11833=>"010011110",
  11834=>"110101111",
  11835=>"101111001",
  11836=>"011001111",
  11837=>"000110100",
  11838=>"111111011",
  11839=>"001111101",
  11840=>"000110010",
  11841=>"011011000",
  11842=>"000111111",
  11843=>"011110010",
  11844=>"110100000",
  11845=>"011010101",
  11846=>"000101111",
  11847=>"011001011",
  11848=>"111011110",
  11849=>"000001100",
  11850=>"111110000",
  11851=>"010011000",
  11852=>"101110011",
  11853=>"011111001",
  11854=>"110010101",
  11855=>"000110100",
  11856=>"110010000",
  11857=>"010011011",
  11858=>"111001011",
  11859=>"110111101",
  11860=>"110111110",
  11861=>"101111110",
  11862=>"101111111",
  11863=>"111101111",
  11864=>"000110000",
  11865=>"001011010",
  11866=>"110111001",
  11867=>"011000100",
  11868=>"100000010",
  11869=>"111100100",
  11870=>"000110111",
  11871=>"100101010",
  11872=>"010100000",
  11873=>"111110011",
  11874=>"000011011",
  11875=>"011100110",
  11876=>"100001101",
  11877=>"110011111",
  11878=>"001000110",
  11879=>"000000000",
  11880=>"000101010",
  11881=>"111110000",
  11882=>"100101011",
  11883=>"000101011",
  11884=>"100001011",
  11885=>"101111011",
  11886=>"111101111",
  11887=>"101011100",
  11888=>"110011111",
  11889=>"010110000",
  11890=>"110000011",
  11891=>"000000100",
  11892=>"000010101",
  11893=>"111111110",
  11894=>"001000011",
  11895=>"110110100",
  11896=>"011100100",
  11897=>"100100101",
  11898=>"000111110",
  11899=>"011010110",
  11900=>"001111110",
  11901=>"000101101",
  11902=>"100000010",
  11903=>"111011100",
  11904=>"100000111",
  11905=>"111100000",
  11906=>"100010001",
  11907=>"110100101",
  11908=>"000110111",
  11909=>"100000100",
  11910=>"000000001",
  11911=>"101001100",
  11912=>"000001001",
  11913=>"100101010",
  11914=>"011011100",
  11915=>"000001100",
  11916=>"111001110",
  11917=>"111111000",
  11918=>"011001110",
  11919=>"101111011",
  11920=>"000111011",
  11921=>"001111010",
  11922=>"011001000",
  11923=>"101100011",
  11924=>"101101010",
  11925=>"000001110",
  11926=>"111111100",
  11927=>"100100001",
  11928=>"111011000",
  11929=>"101011001",
  11930=>"010000011",
  11931=>"101111110",
  11932=>"110111100",
  11933=>"000000010",
  11934=>"000100000",
  11935=>"111001111",
  11936=>"011101010",
  11937=>"010011001",
  11938=>"001011001",
  11939=>"011100101",
  11940=>"110110110",
  11941=>"101110110",
  11942=>"100001100",
  11943=>"010101000",
  11944=>"000000100",
  11945=>"100100101",
  11946=>"101001000",
  11947=>"101000001",
  11948=>"000000101",
  11949=>"101100000",
  11950=>"000000110",
  11951=>"101010101",
  11952=>"111010000",
  11953=>"110110001",
  11954=>"110101011",
  11955=>"111011010",
  11956=>"000011011",
  11957=>"111101011",
  11958=>"101010001",
  11959=>"101001111",
  11960=>"110011101",
  11961=>"001101111",
  11962=>"101100001",
  11963=>"010110011",
  11964=>"100111011",
  11965=>"100100010",
  11966=>"011111111",
  11967=>"110111100",
  11968=>"100100011",
  11969=>"110100010",
  11970=>"111011001",
  11971=>"010110101",
  11972=>"010100000",
  11973=>"110001000",
  11974=>"110100110",
  11975=>"010111110",
  11976=>"111100011",
  11977=>"011011111",
  11978=>"001000010",
  11979=>"001110011",
  11980=>"010010100",
  11981=>"010101001",
  11982=>"000111111",
  11983=>"010000100",
  11984=>"001111011",
  11985=>"111000110",
  11986=>"101011010",
  11987=>"100011100",
  11988=>"011101011",
  11989=>"000101011",
  11990=>"011010110",
  11991=>"001111111",
  11992=>"000000110",
  11993=>"001011000",
  11994=>"110000101",
  11995=>"010000101",
  11996=>"111010010",
  11997=>"100000101",
  11998=>"000000111",
  11999=>"000101100",
  12000=>"000001001",
  12001=>"001101010",
  12002=>"101000111",
  12003=>"101100111",
  12004=>"111000101",
  12005=>"101001011",
  12006=>"000110101",
  12007=>"101011111",
  12008=>"011001001",
  12009=>"111001011",
  12010=>"001001100",
  12011=>"000011000",
  12012=>"001111011",
  12013=>"010100110",
  12014=>"111100101",
  12015=>"110101110",
  12016=>"010110011",
  12017=>"000111101",
  12018=>"100111110",
  12019=>"011111011",
  12020=>"011011010",
  12021=>"001001001",
  12022=>"100011111",
  12023=>"110001101",
  12024=>"010110010",
  12025=>"010101011",
  12026=>"011101111",
  12027=>"101010011",
  12028=>"110111011",
  12029=>"010100000",
  12030=>"010111011",
  12031=>"100011101",
  12032=>"000000000",
  12033=>"000101100",
  12034=>"111101110",
  12035=>"100111110",
  12036=>"011100110",
  12037=>"010011110",
  12038=>"111001000",
  12039=>"111111110",
  12040=>"101001010",
  12041=>"000000000",
  12042=>"011001100",
  12043=>"111101110",
  12044=>"011000010",
  12045=>"100010010",
  12046=>"110010011",
  12047=>"100011100",
  12048=>"110010110",
  12049=>"100111010",
  12050=>"010110100",
  12051=>"111011010",
  12052=>"100110110",
  12053=>"110001001",
  12054=>"010110110",
  12055=>"001010111",
  12056=>"000000100",
  12057=>"001000110",
  12058=>"011011011",
  12059=>"011111000",
  12060=>"011101111",
  12061=>"111100101",
  12062=>"101001110",
  12063=>"000100001",
  12064=>"011011101",
  12065=>"101010000",
  12066=>"110100011",
  12067=>"110000101",
  12068=>"100101111",
  12069=>"111011001",
  12070=>"011000001",
  12071=>"101100011",
  12072=>"100100101",
  12073=>"010001010",
  12074=>"101010010",
  12075=>"110011001",
  12076=>"000001011",
  12077=>"010111111",
  12078=>"110101101",
  12079=>"110100111",
  12080=>"010001110",
  12081=>"011110100",
  12082=>"111000110",
  12083=>"111101000",
  12084=>"100101000",
  12085=>"111110001",
  12086=>"101010110",
  12087=>"111101000",
  12088=>"000010110",
  12089=>"011101011",
  12090=>"101011101",
  12091=>"111010101",
  12092=>"011000111",
  12093=>"101110111",
  12094=>"111010100",
  12095=>"010100100",
  12096=>"000110010",
  12097=>"010001001",
  12098=>"101101001",
  12099=>"100001011",
  12100=>"100010010",
  12101=>"011000101",
  12102=>"111100110",
  12103=>"110000111",
  12104=>"110010101",
  12105=>"110011001",
  12106=>"000011000",
  12107=>"111110110",
  12108=>"010100010",
  12109=>"011101011",
  12110=>"011010001",
  12111=>"011100010",
  12112=>"010100010",
  12113=>"111011101",
  12114=>"000010100",
  12115=>"110011101",
  12116=>"100000000",
  12117=>"100001100",
  12118=>"111010001",
  12119=>"110011111",
  12120=>"111111101",
  12121=>"000010011",
  12122=>"100111101",
  12123=>"110000010",
  12124=>"110101000",
  12125=>"111000011",
  12126=>"000101000",
  12127=>"110011011",
  12128=>"010001001",
  12129=>"000011111",
  12130=>"010111110",
  12131=>"100101011",
  12132=>"110110000",
  12133=>"101111111",
  12134=>"000100111",
  12135=>"110111111",
  12136=>"001000110",
  12137=>"001011101",
  12138=>"001101110",
  12139=>"100110001",
  12140=>"111011100",
  12141=>"111010011",
  12142=>"110011111",
  12143=>"001101000",
  12144=>"110001111",
  12145=>"010111110",
  12146=>"100001011",
  12147=>"110110111",
  12148=>"100110010",
  12149=>"111000000",
  12150=>"010100010",
  12151=>"011110000",
  12152=>"100101110",
  12153=>"011111011",
  12154=>"101101100",
  12155=>"010101101",
  12156=>"000100010",
  12157=>"111000111",
  12158=>"011110101",
  12159=>"011111101",
  12160=>"010000000",
  12161=>"010001101",
  12162=>"101101011",
  12163=>"010111001",
  12164=>"001101111",
  12165=>"010000010",
  12166=>"101001000",
  12167=>"110111011",
  12168=>"100011110",
  12169=>"000011001",
  12170=>"011100010",
  12171=>"110111100",
  12172=>"100100010",
  12173=>"110000000",
  12174=>"010100110",
  12175=>"000110111",
  12176=>"010000111",
  12177=>"110000110",
  12178=>"000111101",
  12179=>"101111110",
  12180=>"011010001",
  12181=>"101100100",
  12182=>"001000111",
  12183=>"011011000",
  12184=>"101101011",
  12185=>"111100111",
  12186=>"110101001",
  12187=>"111100011",
  12188=>"110100101",
  12189=>"010001011",
  12190=>"100101110",
  12191=>"100100110",
  12192=>"010100100",
  12193=>"110100101",
  12194=>"110111000",
  12195=>"001001111",
  12196=>"110111100",
  12197=>"001111011",
  12198=>"011011001",
  12199=>"101101010",
  12200=>"101001000",
  12201=>"111110111",
  12202=>"100101101",
  12203=>"000100101",
  12204=>"000111001",
  12205=>"001001001",
  12206=>"111000100",
  12207=>"001100001",
  12208=>"000101001",
  12209=>"010101110",
  12210=>"001011010",
  12211=>"010010011",
  12212=>"110111110",
  12213=>"101010100",
  12214=>"101111000",
  12215=>"101101110",
  12216=>"111100100",
  12217=>"110011101",
  12218=>"001100101",
  12219=>"010101010",
  12220=>"110100001",
  12221=>"100111100",
  12222=>"000100011",
  12223=>"000011010",
  12224=>"111001101",
  12225=>"110000111",
  12226=>"111011110",
  12227=>"110011110",
  12228=>"100000000",
  12229=>"110011111",
  12230=>"101011001",
  12231=>"100001111",
  12232=>"101011111",
  12233=>"001110001",
  12234=>"000001111",
  12235=>"001101100",
  12236=>"111011111",
  12237=>"100111010",
  12238=>"101001011",
  12239=>"110101100",
  12240=>"101011000",
  12241=>"111101010",
  12242=>"110001010",
  12243=>"000001010",
  12244=>"000010001",
  12245=>"000010111",
  12246=>"100100111",
  12247=>"101100100",
  12248=>"110000111",
  12249=>"001000101",
  12250=>"111101010",
  12251=>"110001001",
  12252=>"101110000",
  12253=>"010100100",
  12254=>"100101000",
  12255=>"011000111",
  12256=>"111000110",
  12257=>"100001011",
  12258=>"000001111",
  12259=>"000000110",
  12260=>"111110110",
  12261=>"010000000",
  12262=>"111110011",
  12263=>"010101011",
  12264=>"111100010",
  12265=>"111110101",
  12266=>"010100010",
  12267=>"001111011",
  12268=>"001110010",
  12269=>"110010011",
  12270=>"000001001",
  12271=>"100100000",
  12272=>"010111001",
  12273=>"000010011",
  12274=>"111111100",
  12275=>"011010111",
  12276=>"000000010",
  12277=>"001111000",
  12278=>"101010100",
  12279=>"010000001",
  12280=>"101100110",
  12281=>"010001100",
  12282=>"101111011",
  12283=>"010010010",
  12284=>"110101000",
  12285=>"000111010",
  12286=>"111101111",
  12287=>"000110110",
  12288=>"111111111",
  12289=>"000010101",
  12290=>"010001011",
  12291=>"110100110",
  12292=>"011111011",
  12293=>"011100001",
  12294=>"110100011",
  12295=>"000101101",
  12296=>"001000000",
  12297=>"001001100",
  12298=>"000110001",
  12299=>"010101101",
  12300=>"000100101",
  12301=>"011011110",
  12302=>"011000010",
  12303=>"111110000",
  12304=>"001000110",
  12305=>"110010100",
  12306=>"100011110",
  12307=>"111001100",
  12308=>"001111110",
  12309=>"101001011",
  12310=>"101010010",
  12311=>"011011010",
  12312=>"100000001",
  12313=>"000000111",
  12314=>"011110000",
  12315=>"011000010",
  12316=>"111001000",
  12317=>"110011001",
  12318=>"111110101",
  12319=>"110100010",
  12320=>"001110101",
  12321=>"000010011",
  12322=>"100100101",
  12323=>"110011100",
  12324=>"100010101",
  12325=>"110101011",
  12326=>"011110011",
  12327=>"111001101",
  12328=>"001100111",
  12329=>"101001001",
  12330=>"000000001",
  12331=>"011111101",
  12332=>"011111100",
  12333=>"000101001",
  12334=>"110000010",
  12335=>"000010111",
  12336=>"100011010",
  12337=>"000110010",
  12338=>"000001101",
  12339=>"100101000",
  12340=>"111110011",
  12341=>"011001000",
  12342=>"001000000",
  12343=>"101000000",
  12344=>"001111111",
  12345=>"001111010",
  12346=>"000101110",
  12347=>"010101110",
  12348=>"000011101",
  12349=>"111111000",
  12350=>"001011001",
  12351=>"110000100",
  12352=>"001011110",
  12353=>"010111000",
  12354=>"101001101",
  12355=>"101011111",
  12356=>"111101001",
  12357=>"111011010",
  12358=>"011111010",
  12359=>"110011110",
  12360=>"011110001",
  12361=>"001000000",
  12362=>"110101101",
  12363=>"110011111",
  12364=>"111011100",
  12365=>"000110010",
  12366=>"010100000",
  12367=>"111101111",
  12368=>"011000100",
  12369=>"000011001",
  12370=>"110001110",
  12371=>"000001010",
  12372=>"010101101",
  12373=>"011010111",
  12374=>"010111110",
  12375=>"001010001",
  12376=>"000001111",
  12377=>"101010100",
  12378=>"001010000",
  12379=>"100001010",
  12380=>"001000111",
  12381=>"100010000",
  12382=>"111101010",
  12383=>"011000100",
  12384=>"111010010",
  12385=>"111100101",
  12386=>"010010001",
  12387=>"110110110",
  12388=>"001110010",
  12389=>"101100110",
  12390=>"000010110",
  12391=>"001001000",
  12392=>"010011110",
  12393=>"101011011",
  12394=>"000111001",
  12395=>"010100000",
  12396=>"111110110",
  12397=>"001010110",
  12398=>"100000110",
  12399=>"110100100",
  12400=>"110011010",
  12401=>"000010100",
  12402=>"010111000",
  12403=>"100101100",
  12404=>"001101011",
  12405=>"101011000",
  12406=>"001011011",
  12407=>"111101001",
  12408=>"001100100",
  12409=>"001000011",
  12410=>"111011101",
  12411=>"011001111",
  12412=>"100001001",
  12413=>"001011111",
  12414=>"010110100",
  12415=>"011011100",
  12416=>"000000000",
  12417=>"001110110",
  12418=>"100000010",
  12419=>"110101110",
  12420=>"000000001",
  12421=>"010111110",
  12422=>"010000011",
  12423=>"011111100",
  12424=>"000011111",
  12425=>"000101101",
  12426=>"110001111",
  12427=>"011111111",
  12428=>"001100110",
  12429=>"011101010",
  12430=>"010101011",
  12431=>"101010110",
  12432=>"001000011",
  12433=>"011010011",
  12434=>"011111011",
  12435=>"011110001",
  12436=>"100101111",
  12437=>"010000111",
  12438=>"010100110",
  12439=>"000100101",
  12440=>"111101111",
  12441=>"111110100",
  12442=>"100101001",
  12443=>"111011100",
  12444=>"101011000",
  12445=>"010111111",
  12446=>"010001011",
  12447=>"000010110",
  12448=>"000110101",
  12449=>"101110111",
  12450=>"101000100",
  12451=>"000110000",
  12452=>"001000111",
  12453=>"001101111",
  12454=>"110111001",
  12455=>"100111011",
  12456=>"001001111",
  12457=>"100100011",
  12458=>"100100000",
  12459=>"101111011",
  12460=>"011011111",
  12461=>"101110001",
  12462=>"101100011",
  12463=>"001001111",
  12464=>"010111010",
  12465=>"000010110",
  12466=>"010100100",
  12467=>"111001001",
  12468=>"110011110",
  12469=>"110010010",
  12470=>"000101111",
  12471=>"011110011",
  12472=>"111010011",
  12473=>"110101111",
  12474=>"000101101",
  12475=>"110101000",
  12476=>"100010100",
  12477=>"111001100",
  12478=>"010110011",
  12479=>"000110001",
  12480=>"011001011",
  12481=>"010000011",
  12482=>"000001110",
  12483=>"101000010",
  12484=>"011001000",
  12485=>"011010100",
  12486=>"010000110",
  12487=>"000000000",
  12488=>"111010111",
  12489=>"001001110",
  12490=>"111110100",
  12491=>"111011111",
  12492=>"100110001",
  12493=>"110010100",
  12494=>"100011100",
  12495=>"110011100",
  12496=>"010100011",
  12497=>"010010110",
  12498=>"100001000",
  12499=>"011011100",
  12500=>"111010001",
  12501=>"101100101",
  12502=>"010011001",
  12503=>"111100010",
  12504=>"101111000",
  12505=>"000110010",
  12506=>"010110101",
  12507=>"011011000",
  12508=>"011001010",
  12509=>"100010100",
  12510=>"011110010",
  12511=>"100010010",
  12512=>"100110100",
  12513=>"010010100",
  12514=>"011000111",
  12515=>"110110000",
  12516=>"100110001",
  12517=>"010110001",
  12518=>"010110110",
  12519=>"011000111",
  12520=>"111101101",
  12521=>"111011110",
  12522=>"010001010",
  12523=>"000010001",
  12524=>"001110101",
  12525=>"000100011",
  12526=>"110011111",
  12527=>"110010010",
  12528=>"011011011",
  12529=>"010010001",
  12530=>"111011001",
  12531=>"100101011",
  12532=>"001011011",
  12533=>"101100000",
  12534=>"111011100",
  12535=>"001011101",
  12536=>"110010100",
  12537=>"001101001",
  12538=>"100000110",
  12539=>"101100001",
  12540=>"001000100",
  12541=>"001000010",
  12542=>"111111111",
  12543=>"101001011",
  12544=>"110001001",
  12545=>"010101111",
  12546=>"011110101",
  12547=>"010110000",
  12548=>"000001011",
  12549=>"011111100",
  12550=>"111000100",
  12551=>"100101011",
  12552=>"001010111",
  12553=>"111100100",
  12554=>"000011010",
  12555=>"001000100",
  12556=>"111110010",
  12557=>"101111111",
  12558=>"000001000",
  12559=>"111110010",
  12560=>"101110011",
  12561=>"100010101",
  12562=>"001101001",
  12563=>"011001101",
  12564=>"011111110",
  12565=>"010000110",
  12566=>"101101011",
  12567=>"010010101",
  12568=>"001111011",
  12569=>"011111111",
  12570=>"111100000",
  12571=>"010101011",
  12572=>"111110001",
  12573=>"101101011",
  12574=>"110011100",
  12575=>"001001001",
  12576=>"100000010",
  12577=>"110110111",
  12578=>"110001001",
  12579=>"111100110",
  12580=>"011111111",
  12581=>"000111010",
  12582=>"111000001",
  12583=>"000100000",
  12584=>"001100000",
  12585=>"001000111",
  12586=>"111011110",
  12587=>"100000101",
  12588=>"001011000",
  12589=>"001000010",
  12590=>"000000101",
  12591=>"100011101",
  12592=>"101100101",
  12593=>"000011001",
  12594=>"100110011",
  12595=>"001100100",
  12596=>"010101110",
  12597=>"000000001",
  12598=>"111010010",
  12599=>"101101000",
  12600=>"111111110",
  12601=>"100111001",
  12602=>"000101111",
  12603=>"010001011",
  12604=>"010011000",
  12605=>"110001010",
  12606=>"111111101",
  12607=>"110010011",
  12608=>"000011101",
  12609=>"101100110",
  12610=>"011001000",
  12611=>"011000010",
  12612=>"010011111",
  12613=>"000100100",
  12614=>"101011010",
  12615=>"001001011",
  12616=>"011111111",
  12617=>"100000000",
  12618=>"000011100",
  12619=>"111010110",
  12620=>"001110001",
  12621=>"100001100",
  12622=>"000111001",
  12623=>"110001001",
  12624=>"101100110",
  12625=>"111011111",
  12626=>"010010000",
  12627=>"000111001",
  12628=>"110101010",
  12629=>"001001111",
  12630=>"100001101",
  12631=>"001110101",
  12632=>"010010001",
  12633=>"000001000",
  12634=>"011111111",
  12635=>"111111000",
  12636=>"101001001",
  12637=>"100001101",
  12638=>"111010011",
  12639=>"111000011",
  12640=>"111110100",
  12641=>"111000011",
  12642=>"000110100",
  12643=>"000000011",
  12644=>"011111101",
  12645=>"000000100",
  12646=>"001000110",
  12647=>"111110111",
  12648=>"011101010",
  12649=>"010100110",
  12650=>"111001111",
  12651=>"110110011",
  12652=>"001111111",
  12653=>"100111010",
  12654=>"011110000",
  12655=>"100110000",
  12656=>"000101010",
  12657=>"001110011",
  12658=>"000101010",
  12659=>"100100001",
  12660=>"111010001",
  12661=>"111011111",
  12662=>"101011101",
  12663=>"100101101",
  12664=>"110010010",
  12665=>"100000001",
  12666=>"111110110",
  12667=>"100110111",
  12668=>"010001110",
  12669=>"110010100",
  12670=>"111001100",
  12671=>"110111100",
  12672=>"011011000",
  12673=>"000001110",
  12674=>"110001011",
  12675=>"001001001",
  12676=>"011110001",
  12677=>"110011011",
  12678=>"001100110",
  12679=>"110110110",
  12680=>"011001000",
  12681=>"011001010",
  12682=>"011010101",
  12683=>"010001101",
  12684=>"101010111",
  12685=>"110011001",
  12686=>"001001011",
  12687=>"100100001",
  12688=>"101101101",
  12689=>"100000000",
  12690=>"100101101",
  12691=>"100010010",
  12692=>"110010110",
  12693=>"000001110",
  12694=>"100101111",
  12695=>"010000100",
  12696=>"100100001",
  12697=>"111100001",
  12698=>"010110000",
  12699=>"001001010",
  12700=>"101001000",
  12701=>"000100000",
  12702=>"000110100",
  12703=>"100010100",
  12704=>"001101100",
  12705=>"100111001",
  12706=>"000100001",
  12707=>"110010011",
  12708=>"101000001",
  12709=>"100110111",
  12710=>"000101000",
  12711=>"001000001",
  12712=>"010010110",
  12713=>"010011111",
  12714=>"010110101",
  12715=>"101000010",
  12716=>"111001000",
  12717=>"011101101",
  12718=>"010001000",
  12719=>"100101111",
  12720=>"010000011",
  12721=>"111111001",
  12722=>"101100000",
  12723=>"111110100",
  12724=>"010110000",
  12725=>"000111111",
  12726=>"111011111",
  12727=>"000111001",
  12728=>"010010010",
  12729=>"100100100",
  12730=>"001000001",
  12731=>"111011110",
  12732=>"101010110",
  12733=>"010000001",
  12734=>"110001010",
  12735=>"101001001",
  12736=>"001100101",
  12737=>"000010001",
  12738=>"100001001",
  12739=>"000010011",
  12740=>"001000001",
  12741=>"100001000",
  12742=>"010001000",
  12743=>"100010001",
  12744=>"100001100",
  12745=>"001101110",
  12746=>"100101001",
  12747=>"111100100",
  12748=>"100111000",
  12749=>"101010010",
  12750=>"000101100",
  12751=>"010000010",
  12752=>"100111111",
  12753=>"011010111",
  12754=>"101111000",
  12755=>"100110110",
  12756=>"011110110",
  12757=>"100101100",
  12758=>"111101011",
  12759=>"010100001",
  12760=>"011010000",
  12761=>"100010110",
  12762=>"010010111",
  12763=>"111101111",
  12764=>"011010101",
  12765=>"110100010",
  12766=>"011111101",
  12767=>"010110111",
  12768=>"101111011",
  12769=>"110101000",
  12770=>"111100111",
  12771=>"111100101",
  12772=>"001011111",
  12773=>"101011111",
  12774=>"001110101",
  12775=>"101110100",
  12776=>"011111101",
  12777=>"011110001",
  12778=>"100000001",
  12779=>"001011011",
  12780=>"111110110",
  12781=>"001110001",
  12782=>"011001110",
  12783=>"100011100",
  12784=>"000010000",
  12785=>"111010011",
  12786=>"011101011",
  12787=>"100000001",
  12788=>"110001000",
  12789=>"000001111",
  12790=>"000011001",
  12791=>"111010001",
  12792=>"000111011",
  12793=>"111101001",
  12794=>"110101011",
  12795=>"101101110",
  12796=>"010011110",
  12797=>"111010111",
  12798=>"010111101",
  12799=>"000110101",
  12800=>"001100010",
  12801=>"001100000",
  12802=>"110100101",
  12803=>"101111101",
  12804=>"111101011",
  12805=>"000000100",
  12806=>"011111100",
  12807=>"111001101",
  12808=>"000011001",
  12809=>"100100111",
  12810=>"011101010",
  12811=>"110011100",
  12812=>"011000000",
  12813=>"010101111",
  12814=>"000001101",
  12815=>"000101110",
  12816=>"110000010",
  12817=>"111100010",
  12818=>"001100100",
  12819=>"110111111",
  12820=>"001001101",
  12821=>"000001000",
  12822=>"001110101",
  12823=>"100101111",
  12824=>"010011011",
  12825=>"000011010",
  12826=>"000001110",
  12827=>"111011100",
  12828=>"010110001",
  12829=>"011001110",
  12830=>"110111001",
  12831=>"011110110",
  12832=>"110100010",
  12833=>"010001001",
  12834=>"101111001",
  12835=>"110010011",
  12836=>"111110101",
  12837=>"000001110",
  12838=>"101011111",
  12839=>"100110010",
  12840=>"110101101",
  12841=>"000110010",
  12842=>"100000110",
  12843=>"110101001",
  12844=>"111011110",
  12845=>"100001001",
  12846=>"100000010",
  12847=>"000011111",
  12848=>"100000011",
  12849=>"110010000",
  12850=>"110101100",
  12851=>"100010111",
  12852=>"000101001",
  12853=>"011101001",
  12854=>"100110101",
  12855=>"001110010",
  12856=>"111011010",
  12857=>"010011000",
  12858=>"001010011",
  12859=>"010011001",
  12860=>"111111000",
  12861=>"100001010",
  12862=>"010001010",
  12863=>"001010110",
  12864=>"110110010",
  12865=>"011111110",
  12866=>"100000111",
  12867=>"111111000",
  12868=>"101110100",
  12869=>"111100101",
  12870=>"100100001",
  12871=>"010001101",
  12872=>"010001000",
  12873=>"000010110",
  12874=>"000101000",
  12875=>"100000001",
  12876=>"101111011",
  12877=>"100001000",
  12878=>"100001001",
  12879=>"110001000",
  12880=>"010011110",
  12881=>"111110010",
  12882=>"101111111",
  12883=>"100101000",
  12884=>"101110100",
  12885=>"101001111",
  12886=>"011001000",
  12887=>"001001000",
  12888=>"111111110",
  12889=>"000011110",
  12890=>"001100010",
  12891=>"111000111",
  12892=>"100001000",
  12893=>"000010100",
  12894=>"110000010",
  12895=>"100010111",
  12896=>"001001001",
  12897=>"101000001",
  12898=>"010101110",
  12899=>"000000111",
  12900=>"110110111",
  12901=>"111101111",
  12902=>"000100100",
  12903=>"001111000",
  12904=>"001000000",
  12905=>"100111000",
  12906=>"101011001",
  12907=>"101010110",
  12908=>"000001010",
  12909=>"111010111",
  12910=>"111011010",
  12911=>"011001100",
  12912=>"111011010",
  12913=>"010101101",
  12914=>"010000001",
  12915=>"100101111",
  12916=>"111011010",
  12917=>"000110010",
  12918=>"111010010",
  12919=>"011000000",
  12920=>"011010000",
  12921=>"010110111",
  12922=>"111010111",
  12923=>"000000001",
  12924=>"100000000",
  12925=>"010001100",
  12926=>"110111110",
  12927=>"100100001",
  12928=>"111111011",
  12929=>"100000010",
  12930=>"111010011",
  12931=>"011100110",
  12932=>"111110111",
  12933=>"000000000",
  12934=>"111011111",
  12935=>"010000000",
  12936=>"001110000",
  12937=>"111000110",
  12938=>"010101000",
  12939=>"110011010",
  12940=>"001000000",
  12941=>"001000100",
  12942=>"011011110",
  12943=>"000000011",
  12944=>"101110011",
  12945=>"100000011",
  12946=>"101001010",
  12947=>"110100110",
  12948=>"101011000",
  12949=>"011001011",
  12950=>"101011011",
  12951=>"100110000",
  12952=>"001000111",
  12953=>"110110010",
  12954=>"111000100",
  12955=>"010111000",
  12956=>"100010111",
  12957=>"111000011",
  12958=>"001010110",
  12959=>"010111100",
  12960=>"011111000",
  12961=>"100011100",
  12962=>"011001101",
  12963=>"001101111",
  12964=>"101110110",
  12965=>"111100101",
  12966=>"101011000",
  12967=>"100100100",
  12968=>"000001001",
  12969=>"111001111",
  12970=>"111010011",
  12971=>"000111111",
  12972=>"101111110",
  12973=>"011111111",
  12974=>"110011100",
  12975=>"000011110",
  12976=>"010001001",
  12977=>"010111010",
  12978=>"100011010",
  12979=>"111101010",
  12980=>"011111011",
  12981=>"111111000",
  12982=>"111011110",
  12983=>"000111100",
  12984=>"010000100",
  12985=>"110011111",
  12986=>"110101110",
  12987=>"011110101",
  12988=>"101000001",
  12989=>"000111101",
  12990=>"001100100",
  12991=>"001001101",
  12992=>"001000001",
  12993=>"101010110",
  12994=>"011011101",
  12995=>"110101110",
  12996=>"111010011",
  12997=>"111001100",
  12998=>"100110111",
  12999=>"000101001",
  13000=>"010000000",
  13001=>"100011110",
  13002=>"101010001",
  13003=>"001110001",
  13004=>"000110000",
  13005=>"000000010",
  13006=>"101111000",
  13007=>"011011011",
  13008=>"111010001",
  13009=>"001101010",
  13010=>"101010110",
  13011=>"011011111",
  13012=>"000001100",
  13013=>"110011010",
  13014=>"111001101",
  13015=>"100100111",
  13016=>"001010111",
  13017=>"000110010",
  13018=>"011101011",
  13019=>"000110100",
  13020=>"101010001",
  13021=>"000010011",
  13022=>"101101101",
  13023=>"000010000",
  13024=>"001001101",
  13025=>"001111100",
  13026=>"111011010",
  13027=>"001010011",
  13028=>"101011111",
  13029=>"100111010",
  13030=>"100000111",
  13031=>"000101010",
  13032=>"001101110",
  13033=>"010000010",
  13034=>"001010001",
  13035=>"110110011",
  13036=>"010111000",
  13037=>"111100001",
  13038=>"101001001",
  13039=>"111000100",
  13040=>"100101100",
  13041=>"110101110",
  13042=>"000001010",
  13043=>"100111001",
  13044=>"110111010",
  13045=>"011001010",
  13046=>"001011010",
  13047=>"011010010",
  13048=>"010011101",
  13049=>"101111100",
  13050=>"110001110",
  13051=>"000101101",
  13052=>"001010111",
  13053=>"000001100",
  13054=>"001001010",
  13055=>"011110110",
  13056=>"111100111",
  13057=>"110101101",
  13058=>"001101100",
  13059=>"110111011",
  13060=>"100000100",
  13061=>"010111100",
  13062=>"011100110",
  13063=>"000001010",
  13064=>"001110011",
  13065=>"001010100",
  13066=>"010100110",
  13067=>"110100001",
  13068=>"111011100",
  13069=>"110000001",
  13070=>"101011010",
  13071=>"100110011",
  13072=>"100011100",
  13073=>"011011010",
  13074=>"110110111",
  13075=>"000000000",
  13076=>"011100001",
  13077=>"100000111",
  13078=>"011111000",
  13079=>"000000010",
  13080=>"101011100",
  13081=>"101001000",
  13082=>"111011110",
  13083=>"001101011",
  13084=>"011010000",
  13085=>"100001110",
  13086=>"000011000",
  13087=>"010101111",
  13088=>"111011010",
  13089=>"101010001",
  13090=>"010110111",
  13091=>"110010111",
  13092=>"111111100",
  13093=>"100110000",
  13094=>"010011111",
  13095=>"111111001",
  13096=>"101101000",
  13097=>"101111010",
  13098=>"100101010",
  13099=>"001010011",
  13100=>"010111011",
  13101=>"000001101",
  13102=>"101001010",
  13103=>"011100000",
  13104=>"101011101",
  13105=>"000011010",
  13106=>"110000010",
  13107=>"101101111",
  13108=>"000010001",
  13109=>"001101101",
  13110=>"100001001",
  13111=>"011101100",
  13112=>"010110000",
  13113=>"100000011",
  13114=>"111100001",
  13115=>"100001001",
  13116=>"101101111",
  13117=>"111000001",
  13118=>"111000000",
  13119=>"010011100",
  13120=>"011011100",
  13121=>"011000000",
  13122=>"011110000",
  13123=>"111101110",
  13124=>"000111011",
  13125=>"100101111",
  13126=>"110010111",
  13127=>"100010010",
  13128=>"010000010",
  13129=>"000100001",
  13130=>"010001001",
  13131=>"000110000",
  13132=>"110110000",
  13133=>"011000100",
  13134=>"001010101",
  13135=>"010111110",
  13136=>"011100000",
  13137=>"111111111",
  13138=>"011111110",
  13139=>"101111101",
  13140=>"010000011",
  13141=>"101000010",
  13142=>"011100100",
  13143=>"010010101",
  13144=>"000000100",
  13145=>"010101111",
  13146=>"000011111",
  13147=>"101011000",
  13148=>"111001011",
  13149=>"000001110",
  13150=>"010100110",
  13151=>"100110000",
  13152=>"000000001",
  13153=>"100111010",
  13154=>"001110100",
  13155=>"011000000",
  13156=>"100101000",
  13157=>"000000000",
  13158=>"100000010",
  13159=>"000001111",
  13160=>"000100011",
  13161=>"110001111",
  13162=>"111100100",
  13163=>"110110111",
  13164=>"101011000",
  13165=>"010100101",
  13166=>"101010000",
  13167=>"111101111",
  13168=>"101100101",
  13169=>"101111010",
  13170=>"001110011",
  13171=>"010100000",
  13172=>"101001011",
  13173=>"111101011",
  13174=>"001000111",
  13175=>"100000000",
  13176=>"001111011",
  13177=>"001010100",
  13178=>"000101001",
  13179=>"010111001",
  13180=>"011101111",
  13181=>"101001101",
  13182=>"000001010",
  13183=>"001110111",
  13184=>"101011100",
  13185=>"110100101",
  13186=>"001100001",
  13187=>"111000110",
  13188=>"010100100",
  13189=>"000011111",
  13190=>"001111110",
  13191=>"100111000",
  13192=>"001011100",
  13193=>"011000110",
  13194=>"100010010",
  13195=>"011000000",
  13196=>"100100100",
  13197=>"001011001",
  13198=>"100010100",
  13199=>"001011010",
  13200=>"000010110",
  13201=>"000101010",
  13202=>"100001111",
  13203=>"100111101",
  13204=>"011010111",
  13205=>"100111001",
  13206=>"011111111",
  13207=>"001001110",
  13208=>"010101011",
  13209=>"101111100",
  13210=>"111111100",
  13211=>"010001100",
  13212=>"001110001",
  13213=>"101101000",
  13214=>"000000111",
  13215=>"101111100",
  13216=>"001101101",
  13217=>"001101110",
  13218=>"010111000",
  13219=>"100001110",
  13220=>"100110001",
  13221=>"101110101",
  13222=>"011001111",
  13223=>"111101110",
  13224=>"101011000",
  13225=>"001111110",
  13226=>"001010000",
  13227=>"111111001",
  13228=>"000111000",
  13229=>"010011010",
  13230=>"011001000",
  13231=>"011000111",
  13232=>"010010100",
  13233=>"100110011",
  13234=>"101000110",
  13235=>"100100111",
  13236=>"000010001",
  13237=>"001111010",
  13238=>"111011100",
  13239=>"111001001",
  13240=>"111110000",
  13241=>"111101010",
  13242=>"000111000",
  13243=>"010101101",
  13244=>"010011010",
  13245=>"100110000",
  13246=>"111000111",
  13247=>"010000000",
  13248=>"010001110",
  13249=>"011010101",
  13250=>"101010100",
  13251=>"011010000",
  13252=>"101001100",
  13253=>"111101010",
  13254=>"101010100",
  13255=>"111101011",
  13256=>"100001101",
  13257=>"111000001",
  13258=>"000011100",
  13259=>"000001110",
  13260=>"000101000",
  13261=>"111010000",
  13262=>"011001101",
  13263=>"110100100",
  13264=>"111101111",
  13265=>"100110100",
  13266=>"101101110",
  13267=>"010001101",
  13268=>"000100000",
  13269=>"101011000",
  13270=>"010001100",
  13271=>"000110011",
  13272=>"001001101",
  13273=>"111100101",
  13274=>"100001010",
  13275=>"100000010",
  13276=>"111100001",
  13277=>"100100001",
  13278=>"111011010",
  13279=>"111111100",
  13280=>"011110100",
  13281=>"100010000",
  13282=>"100110110",
  13283=>"000111010",
  13284=>"000100000",
  13285=>"111111101",
  13286=>"001010100",
  13287=>"111111001",
  13288=>"110000001",
  13289=>"101000101",
  13290=>"000010011",
  13291=>"011010011",
  13292=>"100110101",
  13293=>"100101000",
  13294=>"000010101",
  13295=>"010010000",
  13296=>"010110000",
  13297=>"101110110",
  13298=>"110100101",
  13299=>"100110011",
  13300=>"110101111",
  13301=>"110010010",
  13302=>"010010001",
  13303=>"111110110",
  13304=>"010110011",
  13305=>"000010010",
  13306=>"101111001",
  13307=>"011100011",
  13308=>"011011100",
  13309=>"011010101",
  13310=>"110001000",
  13311=>"111100000",
  13312=>"101000010",
  13313=>"011001000",
  13314=>"000000010",
  13315=>"001101000",
  13316=>"100011010",
  13317=>"111010000",
  13318=>"100111101",
  13319=>"010101100",
  13320=>"110011101",
  13321=>"110000110",
  13322=>"000001000",
  13323=>"011110111",
  13324=>"111111100",
  13325=>"111110011",
  13326=>"001001010",
  13327=>"010110111",
  13328=>"000101101",
  13329=>"001000000",
  13330=>"100001110",
  13331=>"101110010",
  13332=>"110010000",
  13333=>"010111100",
  13334=>"111110110",
  13335=>"111111000",
  13336=>"111001010",
  13337=>"110100101",
  13338=>"111101100",
  13339=>"001010111",
  13340=>"100110011",
  13341=>"101010011",
  13342=>"101011011",
  13343=>"111011111",
  13344=>"111000110",
  13345=>"101010101",
  13346=>"101111010",
  13347=>"001000001",
  13348=>"001011110",
  13349=>"011111100",
  13350=>"010111001",
  13351=>"000000100",
  13352=>"000001100",
  13353=>"000101011",
  13354=>"101010000",
  13355=>"100101110",
  13356=>"110101000",
  13357=>"101100101",
  13358=>"110000001",
  13359=>"001000101",
  13360=>"000001011",
  13361=>"001101110",
  13362=>"001000110",
  13363=>"000001101",
  13364=>"011110011",
  13365=>"001010011",
  13366=>"010101011",
  13367=>"000000111",
  13368=>"000010110",
  13369=>"111001100",
  13370=>"001010111",
  13371=>"111011000",
  13372=>"100000000",
  13373=>"111000001",
  13374=>"011010100",
  13375=>"110111010",
  13376=>"010100000",
  13377=>"001001100",
  13378=>"010000101",
  13379=>"100110001",
  13380=>"010100110",
  13381=>"111110001",
  13382=>"001010101",
  13383=>"100110011",
  13384=>"100100001",
  13385=>"100010110",
  13386=>"101110001",
  13387=>"001011110",
  13388=>"010001110",
  13389=>"010000101",
  13390=>"100111111",
  13391=>"000110011",
  13392=>"010111110",
  13393=>"111111011",
  13394=>"100110111",
  13395=>"011100111",
  13396=>"011111000",
  13397=>"001100001",
  13398=>"010100111",
  13399=>"101110110",
  13400=>"001010001",
  13401=>"111111111",
  13402=>"000000101",
  13403=>"001011100",
  13404=>"101011100",
  13405=>"101010111",
  13406=>"111110111",
  13407=>"101100100",
  13408=>"000111111",
  13409=>"100001000",
  13410=>"000011011",
  13411=>"010010001",
  13412=>"011111001",
  13413=>"110010100",
  13414=>"001000010",
  13415=>"000000100",
  13416=>"001000100",
  13417=>"000011001",
  13418=>"001011100",
  13419=>"000100111",
  13420=>"100000100",
  13421=>"000001110",
  13422=>"111111000",
  13423=>"110000010",
  13424=>"011011100",
  13425=>"000111010",
  13426=>"111001000",
  13427=>"100011011",
  13428=>"101000011",
  13429=>"110010010",
  13430=>"111101110",
  13431=>"110011111",
  13432=>"001111001",
  13433=>"001111110",
  13434=>"001011110",
  13435=>"010010111",
  13436=>"100010000",
  13437=>"100011000",
  13438=>"110010010",
  13439=>"000000010",
  13440=>"110110011",
  13441=>"110111100",
  13442=>"000011001",
  13443=>"110000111",
  13444=>"001011000",
  13445=>"100001011",
  13446=>"111100010",
  13447=>"010000100",
  13448=>"001100110",
  13449=>"001011111",
  13450=>"111001101",
  13451=>"011110001",
  13452=>"001111111",
  13453=>"011010000",
  13454=>"111001011",
  13455=>"101011000",
  13456=>"000101001",
  13457=>"000100111",
  13458=>"101011100",
  13459=>"111011000",
  13460=>"000000110",
  13461=>"000100000",
  13462=>"001100000",
  13463=>"011000000",
  13464=>"011101101",
  13465=>"010011001",
  13466=>"111101001",
  13467=>"110010100",
  13468=>"101111100",
  13469=>"000010011",
  13470=>"100101101",
  13471=>"011000101",
  13472=>"101010000",
  13473=>"100110010",
  13474=>"011110011",
  13475=>"111111111",
  13476=>"101000010",
  13477=>"001100111",
  13478=>"001000110",
  13479=>"100000011",
  13480=>"111101001",
  13481=>"011001000",
  13482=>"100011110",
  13483=>"111001000",
  13484=>"100100010",
  13485=>"100000000",
  13486=>"111010101",
  13487=>"101100111",
  13488=>"011111011",
  13489=>"010110011",
  13490=>"111100110",
  13491=>"000101001",
  13492=>"010000000",
  13493=>"001001011",
  13494=>"101000001",
  13495=>"001110011",
  13496=>"101110101",
  13497=>"101001100",
  13498=>"110011010",
  13499=>"101110011",
  13500=>"100101001",
  13501=>"000001011",
  13502=>"010000011",
  13503=>"101000010",
  13504=>"001101100",
  13505=>"000100111",
  13506=>"001011101",
  13507=>"001011001",
  13508=>"100111110",
  13509=>"111011000",
  13510=>"110101000",
  13511=>"001000000",
  13512=>"011010100",
  13513=>"000010101",
  13514=>"001110100",
  13515=>"101001110",
  13516=>"011010100",
  13517=>"110000101",
  13518=>"110011010",
  13519=>"100010100",
  13520=>"010110000",
  13521=>"010010001",
  13522=>"101100001",
  13523=>"100000101",
  13524=>"100011001",
  13525=>"101000000",
  13526=>"001010101",
  13527=>"111000011",
  13528=>"001010000",
  13529=>"001110110",
  13530=>"110011110",
  13531=>"011110111",
  13532=>"011101000",
  13533=>"111101101",
  13534=>"101000001",
  13535=>"000100011",
  13536=>"001110001",
  13537=>"010011111",
  13538=>"110110000",
  13539=>"110000010",
  13540=>"101000111",
  13541=>"000001111",
  13542=>"111111111",
  13543=>"001001010",
  13544=>"001011101",
  13545=>"011001100",
  13546=>"101001010",
  13547=>"111010010",
  13548=>"011000101",
  13549=>"101111100",
  13550=>"001001001",
  13551=>"001100000",
  13552=>"101111011",
  13553=>"101101001",
  13554=>"110101000",
  13555=>"111010001",
  13556=>"110000011",
  13557=>"110110100",
  13558=>"111110110",
  13559=>"100111000",
  13560=>"001001010",
  13561=>"011111000",
  13562=>"000000010",
  13563=>"011000000",
  13564=>"110000011",
  13565=>"110111011",
  13566=>"001111011",
  13567=>"010010100",
  13568=>"100011100",
  13569=>"001111000",
  13570=>"000100011",
  13571=>"001111100",
  13572=>"011000011",
  13573=>"100010001",
  13574=>"010001011",
  13575=>"101001001",
  13576=>"001010011",
  13577=>"101010110",
  13578=>"111111111",
  13579=>"000111110",
  13580=>"100010101",
  13581=>"101100100",
  13582=>"000000101",
  13583=>"000111101",
  13584=>"001110111",
  13585=>"100110111",
  13586=>"000110010",
  13587=>"111011001",
  13588=>"010111010",
  13589=>"110011101",
  13590=>"010101111",
  13591=>"010011111",
  13592=>"001010101",
  13593=>"010000110",
  13594=>"101011001",
  13595=>"011111000",
  13596=>"100010110",
  13597=>"110001001",
  13598=>"101010010",
  13599=>"101101001",
  13600=>"010111011",
  13601=>"110110000",
  13602=>"101111111",
  13603=>"100010010",
  13604=>"011011000",
  13605=>"111101101",
  13606=>"010001000",
  13607=>"110100101",
  13608=>"100001110",
  13609=>"110000001",
  13610=>"110110110",
  13611=>"011100000",
  13612=>"100111001",
  13613=>"110001000",
  13614=>"110001111",
  13615=>"110010010",
  13616=>"110101000",
  13617=>"000111011",
  13618=>"111111010",
  13619=>"111111100",
  13620=>"000000100",
  13621=>"000000110",
  13622=>"000111010",
  13623=>"001000110",
  13624=>"001111001",
  13625=>"001101001",
  13626=>"100010001",
  13627=>"010100000",
  13628=>"010000101",
  13629=>"100101111",
  13630=>"110010111",
  13631=>"000111011",
  13632=>"011011000",
  13633=>"011110000",
  13634=>"000000010",
  13635=>"010101111",
  13636=>"101101011",
  13637=>"111101100",
  13638=>"010010110",
  13639=>"110001001",
  13640=>"111000001",
  13641=>"001100100",
  13642=>"111000111",
  13643=>"011010010",
  13644=>"101001010",
  13645=>"110001110",
  13646=>"110011010",
  13647=>"110001110",
  13648=>"000011100",
  13649=>"100001001",
  13650=>"111000111",
  13651=>"001101111",
  13652=>"011100100",
  13653=>"101001011",
  13654=>"000010101",
  13655=>"111101101",
  13656=>"000111000",
  13657=>"101110111",
  13658=>"010011000",
  13659=>"010000011",
  13660=>"000010010",
  13661=>"111001001",
  13662=>"011011011",
  13663=>"001000010",
  13664=>"101110101",
  13665=>"011011001",
  13666=>"111110010",
  13667=>"101111100",
  13668=>"110001001",
  13669=>"100110110",
  13670=>"000010011",
  13671=>"000001111",
  13672=>"110010000",
  13673=>"000001110",
  13674=>"100101101",
  13675=>"111110100",
  13676=>"001101110",
  13677=>"011101110",
  13678=>"010010100",
  13679=>"001001101",
  13680=>"010001011",
  13681=>"001101000",
  13682=>"101100101",
  13683=>"001011001",
  13684=>"010001100",
  13685=>"101010010",
  13686=>"001101101",
  13687=>"010010000",
  13688=>"101011011",
  13689=>"010000010",
  13690=>"100110100",
  13691=>"100000001",
  13692=>"011111001",
  13693=>"001101001",
  13694=>"010010100",
  13695=>"101101101",
  13696=>"000000111",
  13697=>"100000111",
  13698=>"100000011",
  13699=>"101011010",
  13700=>"110100111",
  13701=>"100101101",
  13702=>"011100010",
  13703=>"011000100",
  13704=>"001011101",
  13705=>"100101111",
  13706=>"000010001",
  13707=>"111110111",
  13708=>"010101101",
  13709=>"111010111",
  13710=>"111011111",
  13711=>"000001011",
  13712=>"110111100",
  13713=>"100000111",
  13714=>"000100010",
  13715=>"100101111",
  13716=>"111101111",
  13717=>"101101100",
  13718=>"100100010",
  13719=>"110001000",
  13720=>"000000010",
  13721=>"001000100",
  13722=>"100010000",
  13723=>"000111101",
  13724=>"001101000",
  13725=>"010110000",
  13726=>"010000101",
  13727=>"100001010",
  13728=>"100100011",
  13729=>"111010001",
  13730=>"101001100",
  13731=>"000110111",
  13732=>"000110100",
  13733=>"010101111",
  13734=>"010001010",
  13735=>"111010110",
  13736=>"100101001",
  13737=>"011001011",
  13738=>"000100000",
  13739=>"101111110",
  13740=>"100001001",
  13741=>"010100001",
  13742=>"101100111",
  13743=>"011000010",
  13744=>"011011110",
  13745=>"100011010",
  13746=>"001000010",
  13747=>"000111111",
  13748=>"111111001",
  13749=>"011011000",
  13750=>"011110111",
  13751=>"100110010",
  13752=>"010100000",
  13753=>"100110111",
  13754=>"111101100",
  13755=>"011011010",
  13756=>"010011111",
  13757=>"100101010",
  13758=>"110001010",
  13759=>"010011101",
  13760=>"101011111",
  13761=>"011010110",
  13762=>"010111101",
  13763=>"111101101",
  13764=>"010000110",
  13765=>"011101110",
  13766=>"010010000",
  13767=>"001101110",
  13768=>"100101011",
  13769=>"011101011",
  13770=>"110011111",
  13771=>"100000001",
  13772=>"000010011",
  13773=>"110100110",
  13774=>"101000110",
  13775=>"111100001",
  13776=>"111010101",
  13777=>"110111111",
  13778=>"100001111",
  13779=>"000111000",
  13780=>"110010101",
  13781=>"011010101",
  13782=>"001101001",
  13783=>"111001010",
  13784=>"101101000",
  13785=>"101001000",
  13786=>"100100001",
  13787=>"011101000",
  13788=>"111011101",
  13789=>"100100011",
  13790=>"101011101",
  13791=>"000001100",
  13792=>"100111111",
  13793=>"001111010",
  13794=>"010110111",
  13795=>"111110101",
  13796=>"001100101",
  13797=>"011110011",
  13798=>"001101100",
  13799=>"101101010",
  13800=>"111011110",
  13801=>"001000100",
  13802=>"110000100",
  13803=>"110110000",
  13804=>"001100000",
  13805=>"100010100",
  13806=>"111001011",
  13807=>"111111100",
  13808=>"110011111",
  13809=>"000010001",
  13810=>"110000001",
  13811=>"100100000",
  13812=>"111010111",
  13813=>"101100011",
  13814=>"010010110",
  13815=>"110011010",
  13816=>"000000001",
  13817=>"111111101",
  13818=>"100000001",
  13819=>"001010011",
  13820=>"110111001",
  13821=>"010110001",
  13822=>"001010011",
  13823=>"101100110",
  13824=>"110101111",
  13825=>"001100011",
  13826=>"001000000",
  13827=>"001111101",
  13828=>"101111000",
  13829=>"100000001",
  13830=>"010000000",
  13831=>"111111100",
  13832=>"111110100",
  13833=>"011111011",
  13834=>"011111001",
  13835=>"011101010",
  13836=>"110001111",
  13837=>"101110101",
  13838=>"000000000",
  13839=>"111011011",
  13840=>"011001110",
  13841=>"100100000",
  13842=>"001001100",
  13843=>"011101101",
  13844=>"011000010",
  13845=>"100001110",
  13846=>"110010110",
  13847=>"101000000",
  13848=>"100100011",
  13849=>"011000101",
  13850=>"101011001",
  13851=>"110001110",
  13852=>"001010111",
  13853=>"101101101",
  13854=>"011000001",
  13855=>"000001000",
  13856=>"001010010",
  13857=>"100101000",
  13858=>"111111001",
  13859=>"110010010",
  13860=>"011011000",
  13861=>"111110000",
  13862=>"001010001",
  13863=>"100100110",
  13864=>"111110011",
  13865=>"101101001",
  13866=>"111000001",
  13867=>"110101001",
  13868=>"110001011",
  13869=>"101110101",
  13870=>"100011100",
  13871=>"010001010",
  13872=>"110010000",
  13873=>"101111101",
  13874=>"010100001",
  13875=>"010000010",
  13876=>"111001111",
  13877=>"001011011",
  13878=>"110110001",
  13879=>"000101100",
  13880=>"000010010",
  13881=>"100101011",
  13882=>"001110101",
  13883=>"110100101",
  13884=>"001100111",
  13885=>"110001010",
  13886=>"001011010",
  13887=>"110001001",
  13888=>"001111101",
  13889=>"000111001",
  13890=>"000000101",
  13891=>"011011011",
  13892=>"011011101",
  13893=>"011001101",
  13894=>"000101111",
  13895=>"001100001",
  13896=>"110101101",
  13897=>"010110011",
  13898=>"000101110",
  13899=>"100100110",
  13900=>"101010010",
  13901=>"110010110",
  13902=>"010010100",
  13903=>"110011100",
  13904=>"001011001",
  13905=>"111100000",
  13906=>"100010100",
  13907=>"010111101",
  13908=>"111000010",
  13909=>"110100010",
  13910=>"111101110",
  13911=>"011101010",
  13912=>"101111010",
  13913=>"110001111",
  13914=>"111000001",
  13915=>"001110001",
  13916=>"100001000",
  13917=>"100101000",
  13918=>"100100010",
  13919=>"001000101",
  13920=>"100001001",
  13921=>"011000011",
  13922=>"111001111",
  13923=>"101000010",
  13924=>"101100011",
  13925=>"110011010",
  13926=>"001101110",
  13927=>"101000111",
  13928=>"000110011",
  13929=>"100010100",
  13930=>"100111100",
  13931=>"101000100",
  13932=>"100101010",
  13933=>"001101011",
  13934=>"111101110",
  13935=>"000001010",
  13936=>"111001110",
  13937=>"010101000",
  13938=>"011000000",
  13939=>"000000110",
  13940=>"101101100",
  13941=>"000110110",
  13942=>"001010111",
  13943=>"001111100",
  13944=>"000010000",
  13945=>"101000110",
  13946=>"111001010",
  13947=>"000101011",
  13948=>"001001000",
  13949=>"100101011",
  13950=>"010000111",
  13951=>"111011100",
  13952=>"101010010",
  13953=>"100000100",
  13954=>"000001101",
  13955=>"111010100",
  13956=>"101000110",
  13957=>"101100110",
  13958=>"110010010",
  13959=>"110001011",
  13960=>"000011111",
  13961=>"000000101",
  13962=>"110111110",
  13963=>"010010101",
  13964=>"110101000",
  13965=>"001001000",
  13966=>"100000001",
  13967=>"000000100",
  13968=>"110111001",
  13969=>"001100100",
  13970=>"110100111",
  13971=>"000111101",
  13972=>"000111101",
  13973=>"100011011",
  13974=>"100001010",
  13975=>"001101001",
  13976=>"001101111",
  13977=>"111111010",
  13978=>"100100101",
  13979=>"011111110",
  13980=>"001011001",
  13981=>"001011010",
  13982=>"111110011",
  13983=>"100110110",
  13984=>"100011011",
  13985=>"001010010",
  13986=>"011010000",
  13987=>"101111101",
  13988=>"101001011",
  13989=>"010001100",
  13990=>"110101110",
  13991=>"000001110",
  13992=>"110000100",
  13993=>"001100000",
  13994=>"111101001",
  13995=>"001000110",
  13996=>"010100010",
  13997=>"101110110",
  13998=>"101100000",
  13999=>"101101101",
  14000=>"011101000",
  14001=>"100111110",
  14002=>"110101100",
  14003=>"100000100",
  14004=>"101010010",
  14005=>"111011101",
  14006=>"101010001",
  14007=>"001110110",
  14008=>"101101100",
  14009=>"011111111",
  14010=>"111001100",
  14011=>"010010100",
  14012=>"101110001",
  14013=>"110011011",
  14014=>"110011011",
  14015=>"110110101",
  14016=>"001001110",
  14017=>"010010000",
  14018=>"010100111",
  14019=>"111110001",
  14020=>"010001111",
  14021=>"010001110",
  14022=>"101100110",
  14023=>"100001100",
  14024=>"001001000",
  14025=>"000001111",
  14026=>"000010010",
  14027=>"001010100",
  14028=>"111010100",
  14029=>"110110000",
  14030=>"000001111",
  14031=>"101000100",
  14032=>"010000000",
  14033=>"100101101",
  14034=>"111110100",
  14035=>"000000101",
  14036=>"010000100",
  14037=>"101111111",
  14038=>"000011111",
  14039=>"100101111",
  14040=>"010000000",
  14041=>"101000011",
  14042=>"001100101",
  14043=>"011010111",
  14044=>"010000100",
  14045=>"101101000",
  14046=>"000111101",
  14047=>"010110111",
  14048=>"010101000",
  14049=>"011010011",
  14050=>"000011001",
  14051=>"101011111",
  14052=>"100101110",
  14053=>"110010010",
  14054=>"101100001",
  14055=>"111101100",
  14056=>"111000010",
  14057=>"110100110",
  14058=>"011011011",
  14059=>"111000111",
  14060=>"011010010",
  14061=>"001011101",
  14062=>"100100001",
  14063=>"101001010",
  14064=>"011111010",
  14065=>"000101011",
  14066=>"111000110",
  14067=>"010101010",
  14068=>"001101011",
  14069=>"101011000",
  14070=>"001101111",
  14071=>"101101111",
  14072=>"111100010",
  14073=>"100110101",
  14074=>"101111001",
  14075=>"101110011",
  14076=>"110010110",
  14077=>"000001011",
  14078=>"110110000",
  14079=>"111001110",
  14080=>"101010000",
  14081=>"000001101",
  14082=>"110001011",
  14083=>"110111111",
  14084=>"101010010",
  14085=>"000100110",
  14086=>"111101101",
  14087=>"111110101",
  14088=>"101000100",
  14089=>"001110101",
  14090=>"001000100",
  14091=>"100101010",
  14092=>"111111101",
  14093=>"011100001",
  14094=>"111000101",
  14095=>"011000100",
  14096=>"010000001",
  14097=>"000100111",
  14098=>"101000010",
  14099=>"110100101",
  14100=>"001010111",
  14101=>"001100111",
  14102=>"101011010",
  14103=>"101000111",
  14104=>"011010001",
  14105=>"000010100",
  14106=>"111110011",
  14107=>"111000000",
  14108=>"011101011",
  14109=>"100111111",
  14110=>"000100110",
  14111=>"011000001",
  14112=>"010000010",
  14113=>"001111010",
  14114=>"001101010",
  14115=>"010111100",
  14116=>"011011001",
  14117=>"000010001",
  14118=>"001000000",
  14119=>"001011001",
  14120=>"101010100",
  14121=>"011011111",
  14122=>"001110011",
  14123=>"000101110",
  14124=>"101100101",
  14125=>"101000011",
  14126=>"111110110",
  14127=>"001100000",
  14128=>"011011001",
  14129=>"001011001",
  14130=>"000111101",
  14131=>"001111111",
  14132=>"001001111",
  14133=>"100000111",
  14134=>"001110111",
  14135=>"011101000",
  14136=>"000111001",
  14137=>"000000001",
  14138=>"010010101",
  14139=>"110010100",
  14140=>"010100111",
  14141=>"101100000",
  14142=>"101010001",
  14143=>"110010111",
  14144=>"110000001",
  14145=>"010000000",
  14146=>"110010110",
  14147=>"010101010",
  14148=>"101000110",
  14149=>"001011111",
  14150=>"010011010",
  14151=>"110000011",
  14152=>"100101110",
  14153=>"001100010",
  14154=>"111011011",
  14155=>"101001100",
  14156=>"111100101",
  14157=>"000000000",
  14158=>"000110001",
  14159=>"011111101",
  14160=>"110110000",
  14161=>"110111011",
  14162=>"000000001",
  14163=>"000101111",
  14164=>"000110110",
  14165=>"111100011",
  14166=>"110111100",
  14167=>"100000010",
  14168=>"000111010",
  14169=>"110110001",
  14170=>"110000010",
  14171=>"100111100",
  14172=>"110010101",
  14173=>"110101000",
  14174=>"011000001",
  14175=>"000000111",
  14176=>"100101110",
  14177=>"000000001",
  14178=>"010000110",
  14179=>"111011111",
  14180=>"101111000",
  14181=>"111001000",
  14182=>"111110100",
  14183=>"010011010",
  14184=>"100010000",
  14185=>"111101000",
  14186=>"000011000",
  14187=>"100000110",
  14188=>"010011001",
  14189=>"101101101",
  14190=>"111001000",
  14191=>"111100001",
  14192=>"100111111",
  14193=>"011101001",
  14194=>"010000110",
  14195=>"000111011",
  14196=>"000110101",
  14197=>"010011001",
  14198=>"111111011",
  14199=>"100001000",
  14200=>"001101110",
  14201=>"000000000",
  14202=>"010111000",
  14203=>"001101000",
  14204=>"010100111",
  14205=>"100011110",
  14206=>"101101110",
  14207=>"000110110",
  14208=>"101100110",
  14209=>"101011110",
  14210=>"101111001",
  14211=>"000100010",
  14212=>"101100101",
  14213=>"101111010",
  14214=>"011100010",
  14215=>"001100111",
  14216=>"011001110",
  14217=>"110011100",
  14218=>"011011011",
  14219=>"000001110",
  14220=>"100011011",
  14221=>"110011000",
  14222=>"000111111",
  14223=>"110001100",
  14224=>"000100100",
  14225=>"100110100",
  14226=>"000010111",
  14227=>"001110001",
  14228=>"011000001",
  14229=>"101111110",
  14230=>"000101101",
  14231=>"011110001",
  14232=>"110010111",
  14233=>"100000101",
  14234=>"100000100",
  14235=>"000000000",
  14236=>"001111100",
  14237=>"101110101",
  14238=>"011000100",
  14239=>"101101101",
  14240=>"010010000",
  14241=>"000100100",
  14242=>"110010101",
  14243=>"000001110",
  14244=>"111111111",
  14245=>"001000001",
  14246=>"110000011",
  14247=>"001110010",
  14248=>"110011011",
  14249=>"100010111",
  14250=>"100011101",
  14251=>"000000011",
  14252=>"000111100",
  14253=>"100001110",
  14254=>"111010101",
  14255=>"110110000",
  14256=>"101001100",
  14257=>"011000110",
  14258=>"010001111",
  14259=>"100101000",
  14260=>"100100111",
  14261=>"111010000",
  14262=>"001111011",
  14263=>"111001001",
  14264=>"010010110",
  14265=>"111001101",
  14266=>"000101100",
  14267=>"111010000",
  14268=>"111111101",
  14269=>"010000001",
  14270=>"101110011",
  14271=>"101101000",
  14272=>"011001011",
  14273=>"100010001",
  14274=>"111000100",
  14275=>"010110010",
  14276=>"110000011",
  14277=>"100111000",
  14278=>"111000111",
  14279=>"111011100",
  14280=>"110000110",
  14281=>"101110111",
  14282=>"110110001",
  14283=>"111001100",
  14284=>"110000000",
  14285=>"110001100",
  14286=>"100000011",
  14287=>"001001000",
  14288=>"110100111",
  14289=>"000110001",
  14290=>"111011001",
  14291=>"100111010",
  14292=>"110000000",
  14293=>"101100000",
  14294=>"010001001",
  14295=>"011011001",
  14296=>"111111101",
  14297=>"110110011",
  14298=>"001100000",
  14299=>"111110111",
  14300=>"000001000",
  14301=>"100000001",
  14302=>"101111011",
  14303=>"100010010",
  14304=>"001111100",
  14305=>"000110110",
  14306=>"101010101",
  14307=>"101110000",
  14308=>"100011111",
  14309=>"100100101",
  14310=>"010111100",
  14311=>"100100000",
  14312=>"010011101",
  14313=>"100100101",
  14314=>"110110111",
  14315=>"000001110",
  14316=>"101100000",
  14317=>"001111100",
  14318=>"001111100",
  14319=>"100011010",
  14320=>"010111000",
  14321=>"101110101",
  14322=>"101101001",
  14323=>"101110001",
  14324=>"101111111",
  14325=>"110110000",
  14326=>"111000101",
  14327=>"000001111",
  14328=>"000010001",
  14329=>"000000011",
  14330=>"010010011",
  14331=>"100000000",
  14332=>"101101000",
  14333=>"100110110",
  14334=>"100001101",
  14335=>"010011001",
  14336=>"110000110",
  14337=>"101100100",
  14338=>"010010000",
  14339=>"001110101",
  14340=>"011010011",
  14341=>"000010100",
  14342=>"100010010",
  14343=>"001111011",
  14344=>"000101010",
  14345=>"111100100",
  14346=>"001000101",
  14347=>"011001100",
  14348=>"000101011",
  14349=>"000101110",
  14350=>"011000100",
  14351=>"110001011",
  14352=>"001100001",
  14353=>"001001101",
  14354=>"001011111",
  14355=>"011000101",
  14356=>"001111100",
  14357=>"010110100",
  14358=>"111101110",
  14359=>"110011010",
  14360=>"100010110",
  14361=>"110000111",
  14362=>"100100001",
  14363=>"101100000",
  14364=>"111111111",
  14365=>"011110010",
  14366=>"011001000",
  14367=>"011001010",
  14368=>"110110011",
  14369=>"010101000",
  14370=>"010001011",
  14371=>"111010001",
  14372=>"110001111",
  14373=>"111100100",
  14374=>"111001100",
  14375=>"111000110",
  14376=>"000010000",
  14377=>"001010101",
  14378=>"011111101",
  14379=>"010101010",
  14380=>"011110100",
  14381=>"110100101",
  14382=>"101100001",
  14383=>"101000010",
  14384=>"000000101",
  14385=>"110010001",
  14386=>"100100001",
  14387=>"100010100",
  14388=>"010011100",
  14389=>"001100110",
  14390=>"010111110",
  14391=>"110000001",
  14392=>"011010010",
  14393=>"011011001",
  14394=>"000000000",
  14395=>"111010000",
  14396=>"000100101",
  14397=>"010011101",
  14398=>"110011000",
  14399=>"010001111",
  14400=>"100100000",
  14401=>"110111011",
  14402=>"100011111",
  14403=>"011000110",
  14404=>"110110011",
  14405=>"010011000",
  14406=>"100100010",
  14407=>"100010100",
  14408=>"110110011",
  14409=>"000100011",
  14410=>"001101111",
  14411=>"000110111",
  14412=>"111111100",
  14413=>"001000111",
  14414=>"110000110",
  14415=>"101110001",
  14416=>"101111010",
  14417=>"100001101",
  14418=>"100110000",
  14419=>"011001010",
  14420=>"100000010",
  14421=>"001101001",
  14422=>"110000100",
  14423=>"100001001",
  14424=>"111010010",
  14425=>"000110110",
  14426=>"111001100",
  14427=>"011000010",
  14428=>"010111100",
  14429=>"100001110",
  14430=>"101010101",
  14431=>"000110001",
  14432=>"100001101",
  14433=>"000101000",
  14434=>"010001100",
  14435=>"111100010",
  14436=>"000010000",
  14437=>"001110111",
  14438=>"011100101",
  14439=>"000100011",
  14440=>"110000100",
  14441=>"000111110",
  14442=>"000100011",
  14443=>"110101111",
  14444=>"010011111",
  14445=>"011010110",
  14446=>"010001010",
  14447=>"010111010",
  14448=>"010011000",
  14449=>"000000000",
  14450=>"000101100",
  14451=>"110101101",
  14452=>"101010000",
  14453=>"011111010",
  14454=>"011100110",
  14455=>"111000010",
  14456=>"001111011",
  14457=>"111010100",
  14458=>"000011000",
  14459=>"101010101",
  14460=>"000001011",
  14461=>"000100000",
  14462=>"010101110",
  14463=>"101010000",
  14464=>"000011000",
  14465=>"100011100",
  14466=>"011100111",
  14467=>"100011110",
  14468=>"011100101",
  14469=>"101101100",
  14470=>"110111100",
  14471=>"110001011",
  14472=>"000100111",
  14473=>"111001000",
  14474=>"100011010",
  14475=>"101100000",
  14476=>"111111011",
  14477=>"100000110",
  14478=>"011110000",
  14479=>"010000010",
  14480=>"111000111",
  14481=>"100110111",
  14482=>"110001001",
  14483=>"110101101",
  14484=>"010101001",
  14485=>"010010110",
  14486=>"001000011",
  14487=>"111011001",
  14488=>"010011001",
  14489=>"110111001",
  14490=>"111100101",
  14491=>"010001101",
  14492=>"011000010",
  14493=>"001110011",
  14494=>"000111110",
  14495=>"100011011",
  14496=>"101001001",
  14497=>"100001001",
  14498=>"101101111",
  14499=>"110111100",
  14500=>"100001110",
  14501=>"101111010",
  14502=>"001100010",
  14503=>"000001000",
  14504=>"001000110",
  14505=>"100101000",
  14506=>"110111001",
  14507=>"010011111",
  14508=>"111001111",
  14509=>"000111111",
  14510=>"111010001",
  14511=>"111110010",
  14512=>"110100110",
  14513=>"111101011",
  14514=>"001001011",
  14515=>"010111100",
  14516=>"001000001",
  14517=>"010000110",
  14518=>"110001110",
  14519=>"110100111",
  14520=>"100111011",
  14521=>"010100110",
  14522=>"100010010",
  14523=>"100000011",
  14524=>"110100000",
  14525=>"010000110",
  14526=>"011110111",
  14527=>"000100111",
  14528=>"111010011",
  14529=>"000100110",
  14530=>"000010110",
  14531=>"001111001",
  14532=>"100010111",
  14533=>"011000001",
  14534=>"110111111",
  14535=>"011101011",
  14536=>"101010001",
  14537=>"011001111",
  14538=>"100011110",
  14539=>"111100010",
  14540=>"000001011",
  14541=>"111000010",
  14542=>"010010101",
  14543=>"010001000",
  14544=>"011001000",
  14545=>"111110001",
  14546=>"000001100",
  14547=>"011010000",
  14548=>"001011011",
  14549=>"101101111",
  14550=>"110111001",
  14551=>"011010001",
  14552=>"101101010",
  14553=>"011010011",
  14554=>"010101111",
  14555=>"100111001",
  14556=>"010101001",
  14557=>"000110100",
  14558=>"110110100",
  14559=>"111001111",
  14560=>"100010101",
  14561=>"010110100",
  14562=>"100110101",
  14563=>"010000010",
  14564=>"110110101",
  14565=>"010010110",
  14566=>"000111010",
  14567=>"101110011",
  14568=>"011011100",
  14569=>"011010011",
  14570=>"111010110",
  14571=>"011000110",
  14572=>"110111111",
  14573=>"011110110",
  14574=>"111111110",
  14575=>"110011011",
  14576=>"000000101",
  14577=>"001110110",
  14578=>"000111101",
  14579=>"100011010",
  14580=>"000010100",
  14581=>"111011001",
  14582=>"001110101",
  14583=>"010001101",
  14584=>"000100001",
  14585=>"001111001",
  14586=>"100001100",
  14587=>"110000111",
  14588=>"101000111",
  14589=>"100100101",
  14590=>"101111001",
  14591=>"111111011",
  14592=>"111010010",
  14593=>"000001101",
  14594=>"011011000",
  14595=>"111101000",
  14596=>"000011100",
  14597=>"010101111",
  14598=>"011000100",
  14599=>"000000110",
  14600=>"000110110",
  14601=>"100001000",
  14602=>"000000011",
  14603=>"011000111",
  14604=>"010110100",
  14605=>"101110101",
  14606=>"001010111",
  14607=>"101110110",
  14608=>"011100001",
  14609=>"110100011",
  14610=>"101100010",
  14611=>"011100011",
  14612=>"001011000",
  14613=>"011010000",
  14614=>"010101010",
  14615=>"101101011",
  14616=>"110101000",
  14617=>"111101001",
  14618=>"011001001",
  14619=>"000101101",
  14620=>"110000001",
  14621=>"101100000",
  14622=>"000011101",
  14623=>"101110001",
  14624=>"101011101",
  14625=>"110001110",
  14626=>"110011011",
  14627=>"101000011",
  14628=>"001000000",
  14629=>"100011111",
  14630=>"000110101",
  14631=>"111111010",
  14632=>"000101100",
  14633=>"010110010",
  14634=>"001100011",
  14635=>"001001101",
  14636=>"111100000",
  14637=>"100111001",
  14638=>"111001110",
  14639=>"000000100",
  14640=>"000110100",
  14641=>"011001101",
  14642=>"101010110",
  14643=>"010101110",
  14644=>"011110000",
  14645=>"101011111",
  14646=>"111000111",
  14647=>"010110000",
  14648=>"110110101",
  14649=>"101001101",
  14650=>"001110000",
  14651=>"011001010",
  14652=>"111100000",
  14653=>"011100111",
  14654=>"010101011",
  14655=>"001110010",
  14656=>"000100000",
  14657=>"010010000",
  14658=>"011010101",
  14659=>"000010101",
  14660=>"001110110",
  14661=>"001000000",
  14662=>"001000011",
  14663=>"111010000",
  14664=>"101000111",
  14665=>"000000010",
  14666=>"000011001",
  14667=>"000100100",
  14668=>"101111101",
  14669=>"100010100",
  14670=>"001010000",
  14671=>"111111101",
  14672=>"111100111",
  14673=>"001110000",
  14674=>"000000001",
  14675=>"100011110",
  14676=>"011110100",
  14677=>"000001110",
  14678=>"111111101",
  14679=>"000001001",
  14680=>"101100001",
  14681=>"010110100",
  14682=>"010101011",
  14683=>"111111000",
  14684=>"110100001",
  14685=>"110101000",
  14686=>"101101110",
  14687=>"101101001",
  14688=>"100011011",
  14689=>"001000000",
  14690=>"110011100",
  14691=>"100011101",
  14692=>"011011000",
  14693=>"100001000",
  14694=>"000011101",
  14695=>"011100010",
  14696=>"000111111",
  14697=>"110100010",
  14698=>"000100100",
  14699=>"000010100",
  14700=>"001011001",
  14701=>"110110111",
  14702=>"001110110",
  14703=>"001011110",
  14704=>"011000010",
  14705=>"111011100",
  14706=>"001000111",
  14707=>"000100000",
  14708=>"110011111",
  14709=>"100100111",
  14710=>"100010110",
  14711=>"101001000",
  14712=>"011000001",
  14713=>"010101111",
  14714=>"010101110",
  14715=>"001110111",
  14716=>"111010111",
  14717=>"111010111",
  14718=>"101110001",
  14719=>"110010000",
  14720=>"011000010",
  14721=>"010110000",
  14722=>"011010010",
  14723=>"010101010",
  14724=>"101011010",
  14725=>"111001110",
  14726=>"011001010",
  14727=>"000100000",
  14728=>"000000001",
  14729=>"110100100",
  14730=>"100111001",
  14731=>"111111111",
  14732=>"000011110",
  14733=>"000100010",
  14734=>"111000010",
  14735=>"110000000",
  14736=>"010000101",
  14737=>"000010001",
  14738=>"001100000",
  14739=>"111101110",
  14740=>"000101111",
  14741=>"011100110",
  14742=>"100010000",
  14743=>"101111010",
  14744=>"101001101",
  14745=>"001001000",
  14746=>"101001100",
  14747=>"001111101",
  14748=>"010111001",
  14749=>"010101101",
  14750=>"100010100",
  14751=>"100100100",
  14752=>"010001010",
  14753=>"011010010",
  14754=>"001001011",
  14755=>"101110111",
  14756=>"101111010",
  14757=>"111100011",
  14758=>"000111111",
  14759=>"011000001",
  14760=>"100110100",
  14761=>"011110010",
  14762=>"010100101",
  14763=>"000011011",
  14764=>"111110110",
  14765=>"110011111",
  14766=>"001110010",
  14767=>"001000000",
  14768=>"100110111",
  14769=>"111011001",
  14770=>"111111100",
  14771=>"000110110",
  14772=>"110100011",
  14773=>"000010101",
  14774=>"010111000",
  14775=>"100111011",
  14776=>"101111110",
  14777=>"100100101",
  14778=>"000110110",
  14779=>"101111110",
  14780=>"110110011",
  14781=>"001011001",
  14782=>"100010011",
  14783=>"111000001",
  14784=>"100001011",
  14785=>"010000011",
  14786=>"111011100",
  14787=>"010001010",
  14788=>"001111010",
  14789=>"001011111",
  14790=>"010111100",
  14791=>"110010010",
  14792=>"111101100",
  14793=>"100111101",
  14794=>"101111110",
  14795=>"100110111",
  14796=>"111101000",
  14797=>"010101110",
  14798=>"100000100",
  14799=>"010100000",
  14800=>"001100000",
  14801=>"110001101",
  14802=>"011011110",
  14803=>"101000101",
  14804=>"000001111",
  14805=>"001101111",
  14806=>"110000111",
  14807=>"111010000",
  14808=>"111010011",
  14809=>"111000001",
  14810=>"100011001",
  14811=>"101000100",
  14812=>"010111110",
  14813=>"011101011",
  14814=>"011110010",
  14815=>"111110111",
  14816=>"101100001",
  14817=>"000111101",
  14818=>"010100001",
  14819=>"100111110",
  14820=>"110000111",
  14821=>"100011110",
  14822=>"100010100",
  14823=>"111011101",
  14824=>"111000010",
  14825=>"001111111",
  14826=>"110100101",
  14827=>"010000111",
  14828=>"101001111",
  14829=>"100011111",
  14830=>"110111010",
  14831=>"000001100",
  14832=>"101101111",
  14833=>"110101101",
  14834=>"100011001",
  14835=>"110111110",
  14836=>"001001011",
  14837=>"001110011",
  14838=>"101101100",
  14839=>"110100101",
  14840=>"010001100",
  14841=>"000110111",
  14842=>"001101110",
  14843=>"010110010",
  14844=>"110100010",
  14845=>"111010011",
  14846=>"010000001",
  14847=>"101011011",
  14848=>"111010010",
  14849=>"100001101",
  14850=>"110100100",
  14851=>"010010001",
  14852=>"000110101",
  14853=>"111111101",
  14854=>"110001011",
  14855=>"011101011",
  14856=>"111000111",
  14857=>"001010011",
  14858=>"010100011",
  14859=>"101110010",
  14860=>"011000101",
  14861=>"011011101",
  14862=>"101001110",
  14863=>"110000000",
  14864=>"001011010",
  14865=>"100111000",
  14866=>"001011100",
  14867=>"111010001",
  14868=>"100111011",
  14869=>"001101011",
  14870=>"010111011",
  14871=>"110000100",
  14872=>"111011000",
  14873=>"011010100",
  14874=>"110001000",
  14875=>"101010100",
  14876=>"100010110",
  14877=>"111100101",
  14878=>"110110010",
  14879=>"110011110",
  14880=>"110011101",
  14881=>"010100101",
  14882=>"001010000",
  14883=>"010111110",
  14884=>"100010111",
  14885=>"111111101",
  14886=>"011001110",
  14887=>"001100001",
  14888=>"000100101",
  14889=>"111111101",
  14890=>"010001011",
  14891=>"110101001",
  14892=>"010111101",
  14893=>"101011111",
  14894=>"101111001",
  14895=>"101101100",
  14896=>"111010111",
  14897=>"111000001",
  14898=>"101100100",
  14899=>"000110010",
  14900=>"110001000",
  14901=>"001000111",
  14902=>"011100000",
  14903=>"110001011",
  14904=>"101000100",
  14905=>"000100000",
  14906=>"110111110",
  14907=>"111001010",
  14908=>"011111101",
  14909=>"011010001",
  14910=>"000001010",
  14911=>"111110001",
  14912=>"010110011",
  14913=>"100011111",
  14914=>"010110110",
  14915=>"011000011",
  14916=>"011101010",
  14917=>"000010010",
  14918=>"001000000",
  14919=>"010000111",
  14920=>"100011011",
  14921=>"101111000",
  14922=>"100011101",
  14923=>"111001110",
  14924=>"010010100",
  14925=>"110011011",
  14926=>"011000101",
  14927=>"100010101",
  14928=>"100110001",
  14929=>"001110010",
  14930=>"011110001",
  14931=>"110100000",
  14932=>"000010110",
  14933=>"001101101",
  14934=>"101010111",
  14935=>"110011100",
  14936=>"111101111",
  14937=>"101110100",
  14938=>"011110010",
  14939=>"000100100",
  14940=>"111010001",
  14941=>"010010011",
  14942=>"111110011",
  14943=>"001111110",
  14944=>"110100101",
  14945=>"100110111",
  14946=>"010100011",
  14947=>"011000110",
  14948=>"111000010",
  14949=>"001001000",
  14950=>"110011101",
  14951=>"011010111",
  14952=>"010000000",
  14953=>"111101111",
  14954=>"001101011",
  14955=>"111001111",
  14956=>"110010000",
  14957=>"000111011",
  14958=>"111100101",
  14959=>"001011100",
  14960=>"111011001",
  14961=>"100101000",
  14962=>"111111011",
  14963=>"101100100",
  14964=>"000001110",
  14965=>"000111101",
  14966=>"001010010",
  14967=>"100110000",
  14968=>"010000101",
  14969=>"111100010",
  14970=>"010000000",
  14971=>"000000010",
  14972=>"111111110",
  14973=>"101010001",
  14974=>"000001101",
  14975=>"001111010",
  14976=>"101000100",
  14977=>"101111111",
  14978=>"100100010",
  14979=>"001100000",
  14980=>"111010101",
  14981=>"000010001",
  14982=>"111111101",
  14983=>"110111011",
  14984=>"001001100",
  14985=>"000100011",
  14986=>"010010000",
  14987=>"000111101",
  14988=>"010000111",
  14989=>"010010011",
  14990=>"001100001",
  14991=>"001000111",
  14992=>"010111011",
  14993=>"001010100",
  14994=>"100111100",
  14995=>"010101110",
  14996=>"110110111",
  14997=>"101001011",
  14998=>"010110100",
  14999=>"001101100",
  15000=>"010101011",
  15001=>"011000011",
  15002=>"000111010",
  15003=>"010010101",
  15004=>"001011111",
  15005=>"001110001",
  15006=>"011100110",
  15007=>"001110010",
  15008=>"010110011",
  15009=>"100101011",
  15010=>"111111000",
  15011=>"110110011",
  15012=>"001111111",
  15013=>"111110001",
  15014=>"110000111",
  15015=>"011111010",
  15016=>"010110001",
  15017=>"000101110",
  15018=>"000111111",
  15019=>"101100001",
  15020=>"010100010",
  15021=>"110011110",
  15022=>"101110010",
  15023=>"010011010",
  15024=>"111011000",
  15025=>"101010000",
  15026=>"001100010",
  15027=>"000011001",
  15028=>"101000011",
  15029=>"010101010",
  15030=>"111001000",
  15031=>"000001001",
  15032=>"010110000",
  15033=>"010010100",
  15034=>"000011110",
  15035=>"010011111",
  15036=>"100010110",
  15037=>"000001100",
  15038=>"110110000",
  15039=>"010010011",
  15040=>"101110000",
  15041=>"100011111",
  15042=>"001001100",
  15043=>"010101000",
  15044=>"001101111",
  15045=>"100000110",
  15046=>"101001100",
  15047=>"010101110",
  15048=>"000001100",
  15049=>"001110100",
  15050=>"011101111",
  15051=>"100100010",
  15052=>"010011011",
  15053=>"101101110",
  15054=>"010100000",
  15055=>"010000111",
  15056=>"010000101",
  15057=>"000001000",
  15058=>"001111001",
  15059=>"000010001",
  15060=>"110010100",
  15061=>"010111010",
  15062=>"011100000",
  15063=>"110011101",
  15064=>"111100010",
  15065=>"100000100",
  15066=>"111100111",
  15067=>"101100101",
  15068=>"001011010",
  15069=>"011110001",
  15070=>"011011101",
  15071=>"011011101",
  15072=>"110010111",
  15073=>"000011010",
  15074=>"010000101",
  15075=>"000111010",
  15076=>"111010100",
  15077=>"000010110",
  15078=>"100111110",
  15079=>"100001110",
  15080=>"001101111",
  15081=>"101000110",
  15082=>"011101100",
  15083=>"001110000",
  15084=>"001101101",
  15085=>"101101101",
  15086=>"110001010",
  15087=>"000011011",
  15088=>"000010111",
  15089=>"111001001",
  15090=>"111000111",
  15091=>"010010111",
  15092=>"111100100",
  15093=>"100001000",
  15094=>"010111111",
  15095=>"111110001",
  15096=>"010000010",
  15097=>"110000111",
  15098=>"011100011",
  15099=>"101001010",
  15100=>"010010100",
  15101=>"110111010",
  15102=>"000010000",
  15103=>"010100111",
  15104=>"111010000",
  15105=>"001011011",
  15106=>"011111001",
  15107=>"011011110",
  15108=>"001001011",
  15109=>"000110101",
  15110=>"010110011",
  15111=>"011100011",
  15112=>"000100011",
  15113=>"000001001",
  15114=>"111000011",
  15115=>"001101101",
  15116=>"000100001",
  15117=>"110000010",
  15118=>"010010100",
  15119=>"000101001",
  15120=>"110100010",
  15121=>"001011010",
  15122=>"011011110",
  15123=>"011010001",
  15124=>"101001010",
  15125=>"100111111",
  15126=>"100100101",
  15127=>"110110011",
  15128=>"111001001",
  15129=>"010100001",
  15130=>"010010001",
  15131=>"110110010",
  15132=>"001000111",
  15133=>"001111011",
  15134=>"000101000",
  15135=>"001111001",
  15136=>"111110111",
  15137=>"010111110",
  15138=>"100111100",
  15139=>"110101011",
  15140=>"000001101",
  15141=>"000111010",
  15142=>"111111100",
  15143=>"110010011",
  15144=>"011101011",
  15145=>"111101001",
  15146=>"001010000",
  15147=>"100001101",
  15148=>"101101000",
  15149=>"000101111",
  15150=>"001011010",
  15151=>"010011101",
  15152=>"010010110",
  15153=>"000100011",
  15154=>"001010101",
  15155=>"100111111",
  15156=>"100010011",
  15157=>"001001111",
  15158=>"000010010",
  15159=>"001110000",
  15160=>"110111011",
  15161=>"010111111",
  15162=>"000000001",
  15163=>"111100011",
  15164=>"111000110",
  15165=>"001000001",
  15166=>"100101000",
  15167=>"000110100",
  15168=>"111101100",
  15169=>"011110000",
  15170=>"000001000",
  15171=>"010000001",
  15172=>"100000101",
  15173=>"100001101",
  15174=>"101001100",
  15175=>"000001001",
  15176=>"001001100",
  15177=>"010110110",
  15178=>"010100111",
  15179=>"111110010",
  15180=>"110010011",
  15181=>"101111001",
  15182=>"000100001",
  15183=>"101100000",
  15184=>"011000110",
  15185=>"101100110",
  15186=>"001110101",
  15187=>"011011000",
  15188=>"000010001",
  15189=>"100111111",
  15190=>"100001011",
  15191=>"101011001",
  15192=>"111000101",
  15193=>"100010111",
  15194=>"010111100",
  15195=>"101000101",
  15196=>"101010111",
  15197=>"001111111",
  15198=>"001110010",
  15199=>"110011001",
  15200=>"010001110",
  15201=>"110000010",
  15202=>"010110011",
  15203=>"100001100",
  15204=>"101011101",
  15205=>"010110011",
  15206=>"011011001",
  15207=>"010010000",
  15208=>"111110110",
  15209=>"111100011",
  15210=>"000011011",
  15211=>"101100000",
  15212=>"001001110",
  15213=>"000110000",
  15214=>"111100010",
  15215=>"110001000",
  15216=>"010111110",
  15217=>"011010000",
  15218=>"010110010",
  15219=>"111010000",
  15220=>"100000110",
  15221=>"100010100",
  15222=>"101001101",
  15223=>"001001100",
  15224=>"110111000",
  15225=>"111010011",
  15226=>"101010011",
  15227=>"101000010",
  15228=>"000001000",
  15229=>"001100001",
  15230=>"111000110",
  15231=>"010100101",
  15232=>"011110110",
  15233=>"101110101",
  15234=>"100010000",
  15235=>"111000001",
  15236=>"010010000",
  15237=>"011100100",
  15238=>"110110111",
  15239=>"111100101",
  15240=>"000111100",
  15241=>"000010011",
  15242=>"101011001",
  15243=>"100010010",
  15244=>"010010110",
  15245=>"100100010",
  15246=>"100011101",
  15247=>"001000110",
  15248=>"000100111",
  15249=>"001001111",
  15250=>"100110001",
  15251=>"111101110",
  15252=>"010011101",
  15253=>"111110001",
  15254=>"011101000",
  15255=>"001001110",
  15256=>"100110000",
  15257=>"001010001",
  15258=>"010010011",
  15259=>"101100011",
  15260=>"100111101",
  15261=>"110111111",
  15262=>"110011001",
  15263=>"011010001",
  15264=>"011110000",
  15265=>"111011110",
  15266=>"011001000",
  15267=>"011110100",
  15268=>"011000010",
  15269=>"101011011",
  15270=>"111100111",
  15271=>"010101000",
  15272=>"001000001",
  15273=>"111001001",
  15274=>"011001111",
  15275=>"111100111",
  15276=>"011100111",
  15277=>"001001001",
  15278=>"110010010",
  15279=>"011110111",
  15280=>"000011100",
  15281=>"101110010",
  15282=>"011000101",
  15283=>"111101001",
  15284=>"001101011",
  15285=>"111001101",
  15286=>"001001111",
  15287=>"000010011",
  15288=>"000100001",
  15289=>"101000010",
  15290=>"000001010",
  15291=>"110010110",
  15292=>"100001010",
  15293=>"001000001",
  15294=>"010000110",
  15295=>"000000000",
  15296=>"110110100",
  15297=>"011000111",
  15298=>"111011000",
  15299=>"001111111",
  15300=>"010010010",
  15301=>"011001101",
  15302=>"111110111",
  15303=>"110010001",
  15304=>"001010011",
  15305=>"100011011",
  15306=>"111000111",
  15307=>"110100101",
  15308=>"111101101",
  15309=>"111000101",
  15310=>"100100100",
  15311=>"011011110",
  15312=>"100111011",
  15313=>"100101100",
  15314=>"100000111",
  15315=>"000000011",
  15316=>"001001110",
  15317=>"010011111",
  15318=>"101110110",
  15319=>"000101111",
  15320=>"111101010",
  15321=>"100101010",
  15322=>"011110110",
  15323=>"001001100",
  15324=>"001110110",
  15325=>"010110101",
  15326=>"100001000",
  15327=>"100111101",
  15328=>"100011101",
  15329=>"110100001",
  15330=>"101101100",
  15331=>"010110000",
  15332=>"110011001",
  15333=>"100011101",
  15334=>"101011110",
  15335=>"010000011",
  15336=>"101110010",
  15337=>"110101110",
  15338=>"001100011",
  15339=>"001010010",
  15340=>"010011100",
  15341=>"011110011",
  15342=>"110001001",
  15343=>"000010011",
  15344=>"110001011",
  15345=>"001010100",
  15346=>"000000100",
  15347=>"000101001",
  15348=>"101111010",
  15349=>"001101111",
  15350=>"011110110",
  15351=>"010011010",
  15352=>"110000111",
  15353=>"001010100",
  15354=>"101110010",
  15355=>"101011000",
  15356=>"100001100",
  15357=>"000000001",
  15358=>"111001111",
  15359=>"010000011",
  15360=>"100000010",
  15361=>"110010011",
  15362=>"010111110",
  15363=>"001110100",
  15364=>"110101010",
  15365=>"011110110",
  15366=>"110110100",
  15367=>"100000010",
  15368=>"010111111",
  15369=>"001100000",
  15370=>"111110010",
  15371=>"100001001",
  15372=>"010111000",
  15373=>"111111010",
  15374=>"101111101",
  15375=>"111110101",
  15376=>"110011101",
  15377=>"111101111",
  15378=>"111000000",
  15379=>"011011110",
  15380=>"111000110",
  15381=>"110011010",
  15382=>"000110101",
  15383=>"101111101",
  15384=>"011110110",
  15385=>"101110010",
  15386=>"010000110",
  15387=>"010010100",
  15388=>"000011001",
  15389=>"000010000",
  15390=>"000010111",
  15391=>"110010111",
  15392=>"010000001",
  15393=>"111011101",
  15394=>"011100001",
  15395=>"011000000",
  15396=>"011101000",
  15397=>"010001010",
  15398=>"100010011",
  15399=>"111001010",
  15400=>"001011110",
  15401=>"101110101",
  15402=>"100110100",
  15403=>"011010001",
  15404=>"100100110",
  15405=>"110111000",
  15406=>"111101111",
  15407=>"011101111",
  15408=>"001000001",
  15409=>"110011111",
  15410=>"110011100",
  15411=>"110101100",
  15412=>"011001000",
  15413=>"001110001",
  15414=>"001001001",
  15415=>"110001101",
  15416=>"110010011",
  15417=>"110011000",
  15418=>"000000000",
  15419=>"101110110",
  15420=>"011101010",
  15421=>"010011011",
  15422=>"100100000",
  15423=>"111111110",
  15424=>"011110010",
  15425=>"101101111",
  15426=>"011000001",
  15427=>"110000111",
  15428=>"011010010",
  15429=>"000111010",
  15430=>"111110010",
  15431=>"010111101",
  15432=>"011101101",
  15433=>"110010100",
  15434=>"000001001",
  15435=>"000000011",
  15436=>"010111001",
  15437=>"011111000",
  15438=>"001111010",
  15439=>"000011001",
  15440=>"011101100",
  15441=>"000111000",
  15442=>"000010001",
  15443=>"000011000",
  15444=>"010101000",
  15445=>"000111111",
  15446=>"001001111",
  15447=>"010001100",
  15448=>"000001100",
  15449=>"110000001",
  15450=>"000100111",
  15451=>"111101010",
  15452=>"110000011",
  15453=>"110010110",
  15454=>"001110110",
  15455=>"011010001",
  15456=>"100010001",
  15457=>"010110010",
  15458=>"001111111",
  15459=>"111000111",
  15460=>"110001101",
  15461=>"000011010",
  15462=>"100111010",
  15463=>"001011001",
  15464=>"001100001",
  15465=>"000000111",
  15466=>"111100100",
  15467=>"011111111",
  15468=>"100100000",
  15469=>"100010000",
  15470=>"011010010",
  15471=>"111000000",
  15472=>"111101100",
  15473=>"110110101",
  15474=>"111000011",
  15475=>"000011101",
  15476=>"000011010",
  15477=>"101000000",
  15478=>"111011011",
  15479=>"010010111",
  15480=>"111111110",
  15481=>"011100011",
  15482=>"011010100",
  15483=>"110111000",
  15484=>"011001010",
  15485=>"000010010",
  15486=>"000001010",
  15487=>"001001001",
  15488=>"001001010",
  15489=>"100010010",
  15490=>"100010001",
  15491=>"111011101",
  15492=>"111101100",
  15493=>"000000100",
  15494=>"110001111",
  15495=>"100000110",
  15496=>"111011000",
  15497=>"111001011",
  15498=>"110011111",
  15499=>"110000000",
  15500=>"100110110",
  15501=>"000101101",
  15502=>"111000111",
  15503=>"000000000",
  15504=>"010100111",
  15505=>"110000000",
  15506=>"111110010",
  15507=>"001001101",
  15508=>"000100101",
  15509=>"010010001",
  15510=>"111111001",
  15511=>"010111111",
  15512=>"110010001",
  15513=>"110100010",
  15514=>"101010100",
  15515=>"000011001",
  15516=>"001001111",
  15517=>"001111101",
  15518=>"010000000",
  15519=>"010101011",
  15520=>"001011101",
  15521=>"011001011",
  15522=>"101100010",
  15523=>"110110111",
  15524=>"100011101",
  15525=>"011100001",
  15526=>"000111111",
  15527=>"111001001",
  15528=>"011000110",
  15529=>"000111001",
  15530=>"100000111",
  15531=>"111001001",
  15532=>"011111100",
  15533=>"000101010",
  15534=>"110110010",
  15535=>"010111111",
  15536=>"100110010",
  15537=>"011011101",
  15538=>"100111011",
  15539=>"100011010",
  15540=>"001111011",
  15541=>"100000101",
  15542=>"101001001",
  15543=>"111011010",
  15544=>"000111001",
  15545=>"100000110",
  15546=>"001000101",
  15547=>"101010000",
  15548=>"000011001",
  15549=>"010101011",
  15550=>"011001101",
  15551=>"110111010",
  15552=>"000000110",
  15553=>"010100100",
  15554=>"101100000",
  15555=>"000110010",
  15556=>"100111101",
  15557=>"110010110",
  15558=>"011101101",
  15559=>"101100111",
  15560=>"101101100",
  15561=>"000010101",
  15562=>"110001101",
  15563=>"001100010",
  15564=>"011110100",
  15565=>"111111110",
  15566=>"010011111",
  15567=>"001110101",
  15568=>"010111011",
  15569=>"110101000",
  15570=>"001001110",
  15571=>"100101111",
  15572=>"111000110",
  15573=>"100011111",
  15574=>"110101101",
  15575=>"111010010",
  15576=>"010101000",
  15577=>"000001100",
  15578=>"111111000",
  15579=>"010101001",
  15580=>"100010001",
  15581=>"011000011",
  15582=>"110100101",
  15583=>"111000001",
  15584=>"110111100",
  15585=>"010001010",
  15586=>"110000011",
  15587=>"001000000",
  15588=>"111110010",
  15589=>"000011000",
  15590=>"110111111",
  15591=>"101110010",
  15592=>"100100100",
  15593=>"111010001",
  15594=>"110001001",
  15595=>"111001011",
  15596=>"000101101",
  15597=>"000101010",
  15598=>"000000101",
  15599=>"000000000",
  15600=>"011011011",
  15601=>"001101000",
  15602=>"111010100",
  15603=>"011000000",
  15604=>"110110011",
  15605=>"011001111",
  15606=>"010110100",
  15607=>"111101111",
  15608=>"010101000",
  15609=>"100011001",
  15610=>"110011101",
  15611=>"111011011",
  15612=>"110001000",
  15613=>"010111111",
  15614=>"001000110",
  15615=>"011100000",
  15616=>"011010110",
  15617=>"111001110",
  15618=>"001010111",
  15619=>"110100011",
  15620=>"101100001",
  15621=>"000001011",
  15622=>"110111101",
  15623=>"101110110",
  15624=>"011101000",
  15625=>"011000100",
  15626=>"101101011",
  15627=>"001111111",
  15628=>"001001110",
  15629=>"010010100",
  15630=>"110111011",
  15631=>"000000011",
  15632=>"110110000",
  15633=>"111110000",
  15634=>"011101000",
  15635=>"000111110",
  15636=>"010000000",
  15637=>"011010110",
  15638=>"110111111",
  15639=>"100100111",
  15640=>"110011110",
  15641=>"111000000",
  15642=>"111001101",
  15643=>"100001010",
  15644=>"000000000",
  15645=>"111100010",
  15646=>"110101110",
  15647=>"000101111",
  15648=>"101010011",
  15649=>"101010110",
  15650=>"111111100",
  15651=>"001001101",
  15652=>"110110010",
  15653=>"001000001",
  15654=>"010000110",
  15655=>"111010100",
  15656=>"000100010",
  15657=>"101101111",
  15658=>"101101011",
  15659=>"111010000",
  15660=>"110100010",
  15661=>"111110100",
  15662=>"111010010",
  15663=>"010110110",
  15664=>"011101000",
  15665=>"001111010",
  15666=>"110101011",
  15667=>"010011001",
  15668=>"110000111",
  15669=>"101111101",
  15670=>"110011111",
  15671=>"000111010",
  15672=>"111111111",
  15673=>"101100010",
  15674=>"101100111",
  15675=>"001101000",
  15676=>"011110001",
  15677=>"100100001",
  15678=>"111110100",
  15679=>"001100010",
  15680=>"101010001",
  15681=>"111010001",
  15682=>"001110001",
  15683=>"111011110",
  15684=>"001111100",
  15685=>"010111101",
  15686=>"010110111",
  15687=>"111011011",
  15688=>"101000100",
  15689=>"011000011",
  15690=>"100001101",
  15691=>"001001000",
  15692=>"010000110",
  15693=>"110100000",
  15694=>"001011100",
  15695=>"101110011",
  15696=>"110100110",
  15697=>"001001101",
  15698=>"111100000",
  15699=>"000000110",
  15700=>"110011101",
  15701=>"000000111",
  15702=>"101100100",
  15703=>"000100101",
  15704=>"110101111",
  15705=>"101001011",
  15706=>"111101011",
  15707=>"011000011",
  15708=>"101011010",
  15709=>"001010101",
  15710=>"010111111",
  15711=>"000010010",
  15712=>"000000100",
  15713=>"000101000",
  15714=>"110010101",
  15715=>"101000001",
  15716=>"101011001",
  15717=>"001001110",
  15718=>"101000101",
  15719=>"110100111",
  15720=>"000001010",
  15721=>"101011100",
  15722=>"000100100",
  15723=>"010000010",
  15724=>"001001001",
  15725=>"001001100",
  15726=>"100100001",
  15727=>"010111100",
  15728=>"011101110",
  15729=>"101001101",
  15730=>"010101011",
  15731=>"000011100",
  15732=>"101010100",
  15733=>"111010111",
  15734=>"111011100",
  15735=>"011000011",
  15736=>"010001011",
  15737=>"110100010",
  15738=>"010110111",
  15739=>"001000001",
  15740=>"000000111",
  15741=>"000101111",
  15742=>"101010000",
  15743=>"110001101",
  15744=>"100011101",
  15745=>"011010100",
  15746=>"000000101",
  15747=>"001110001",
  15748=>"111100100",
  15749=>"101101111",
  15750=>"000110100",
  15751=>"110010110",
  15752=>"100000101",
  15753=>"110111110",
  15754=>"001001101",
  15755=>"100111000",
  15756=>"010001101",
  15757=>"111101111",
  15758=>"000111001",
  15759=>"011010011",
  15760=>"001011111",
  15761=>"001000111",
  15762=>"111001001",
  15763=>"010000100",
  15764=>"110110001",
  15765=>"000001111",
  15766=>"111000001",
  15767=>"001000000",
  15768=>"111101000",
  15769=>"100000110",
  15770=>"100101010",
  15771=>"101000110",
  15772=>"111000000",
  15773=>"001110000",
  15774=>"100100010",
  15775=>"000101110",
  15776=>"101001001",
  15777=>"000111110",
  15778=>"001111100",
  15779=>"111011110",
  15780=>"111011000",
  15781=>"000000010",
  15782=>"111111000",
  15783=>"000010000",
  15784=>"111001000",
  15785=>"111100100",
  15786=>"011100100",
  15787=>"011000110",
  15788=>"111110111",
  15789=>"001011000",
  15790=>"010010110",
  15791=>"010101000",
  15792=>"101000011",
  15793=>"100001111",
  15794=>"111010101",
  15795=>"001000000",
  15796=>"000100011",
  15797=>"000011011",
  15798=>"100011011",
  15799=>"010100101",
  15800=>"100000110",
  15801=>"001110001",
  15802=>"110000110",
  15803=>"110010111",
  15804=>"001010111",
  15805=>"110111101",
  15806=>"001000111",
  15807=>"111010010",
  15808=>"011001010",
  15809=>"111111011",
  15810=>"000001110",
  15811=>"011010001",
  15812=>"101011100",
  15813=>"111011000",
  15814=>"111001001",
  15815=>"111101111",
  15816=>"011101101",
  15817=>"111001111",
  15818=>"100110111",
  15819=>"100111010",
  15820=>"011100101",
  15821=>"110110000",
  15822=>"000100110",
  15823=>"100101101",
  15824=>"110101011",
  15825=>"111110100",
  15826=>"001110110",
  15827=>"000000010",
  15828=>"010111101",
  15829=>"110110101",
  15830=>"111011010",
  15831=>"001001100",
  15832=>"001110010",
  15833=>"010000000",
  15834=>"111010100",
  15835=>"100011101",
  15836=>"010000111",
  15837=>"110101101",
  15838=>"000111110",
  15839=>"000011111",
  15840=>"111011010",
  15841=>"111100111",
  15842=>"001111011",
  15843=>"100110011",
  15844=>"000110000",
  15845=>"000001011",
  15846=>"110011011",
  15847=>"101001101",
  15848=>"101101010",
  15849=>"010011111",
  15850=>"100111010",
  15851=>"000100111",
  15852=>"101110110",
  15853=>"101001110",
  15854=>"111010110",
  15855=>"000010110",
  15856=>"011000110",
  15857=>"110100110",
  15858=>"011111111",
  15859=>"000011111",
  15860=>"000101111",
  15861=>"111110101",
  15862=>"111010101",
  15863=>"001010000",
  15864=>"000011111",
  15865=>"010101001",
  15866=>"101100010",
  15867=>"010001101",
  15868=>"001000000",
  15869=>"011010000",
  15870=>"011111000",
  15871=>"010001110",
  15872=>"110000001",
  15873=>"000001001",
  15874=>"001011111",
  15875=>"111110010",
  15876=>"010011000",
  15877=>"010111100",
  15878=>"101011110",
  15879=>"111111010",
  15880=>"001000100",
  15881=>"011011000",
  15882=>"101110110",
  15883=>"000100011",
  15884=>"110011101",
  15885=>"000100100",
  15886=>"001100010",
  15887=>"101010010",
  15888=>"010001100",
  15889=>"101011100",
  15890=>"100010000",
  15891=>"110101001",
  15892=>"010110000",
  15893=>"011110110",
  15894=>"011010111",
  15895=>"011001110",
  15896=>"000011011",
  15897=>"000111000",
  15898=>"110000100",
  15899=>"010101001",
  15900=>"110111001",
  15901=>"101111001",
  15902=>"111101100",
  15903=>"100000111",
  15904=>"110111101",
  15905=>"111111011",
  15906=>"110101011",
  15907=>"011100011",
  15908=>"111100010",
  15909=>"110100011",
  15910=>"111000100",
  15911=>"001000010",
  15912=>"010001100",
  15913=>"111101001",
  15914=>"110010111",
  15915=>"001111100",
  15916=>"101110010",
  15917=>"001000010",
  15918=>"000111111",
  15919=>"100110100",
  15920=>"111000000",
  15921=>"001010110",
  15922=>"101000110",
  15923=>"111111110",
  15924=>"011011001",
  15925=>"110011011",
  15926=>"111101001",
  15927=>"000000100",
  15928=>"111100001",
  15929=>"011000010",
  15930=>"101101101",
  15931=>"100111000",
  15932=>"111110011",
  15933=>"010101111",
  15934=>"101101101",
  15935=>"110101001",
  15936=>"111010101",
  15937=>"110011110",
  15938=>"111100101",
  15939=>"100111001",
  15940=>"100100010",
  15941=>"010111000",
  15942=>"101001011",
  15943=>"011011100",
  15944=>"011010001",
  15945=>"011110010",
  15946=>"001111110",
  15947=>"101110100",
  15948=>"011100111",
  15949=>"001001011",
  15950=>"100001000",
  15951=>"011010110",
  15952=>"111110110",
  15953=>"110011110",
  15954=>"100001111",
  15955=>"001100000",
  15956=>"110100101",
  15957=>"111111011",
  15958=>"111100110",
  15959=>"110011011",
  15960=>"000000100",
  15961=>"110000001",
  15962=>"011110110",
  15963=>"101111100",
  15964=>"110001010",
  15965=>"110110101",
  15966=>"011011011",
  15967=>"111101000",
  15968=>"111000001",
  15969=>"110010110",
  15970=>"101000010",
  15971=>"100111100",
  15972=>"110111111",
  15973=>"111101111",
  15974=>"001001111",
  15975=>"001000111",
  15976=>"001110011",
  15977=>"001101011",
  15978=>"101000010",
  15979=>"001001101",
  15980=>"010110000",
  15981=>"011110001",
  15982=>"001110011",
  15983=>"111010001",
  15984=>"110111111",
  15985=>"111100110",
  15986=>"111010110",
  15987=>"001110101",
  15988=>"100010011",
  15989=>"000010000",
  15990=>"111010101",
  15991=>"011011111",
  15992=>"100011011",
  15993=>"100100100",
  15994=>"101100000",
  15995=>"111010010",
  15996=>"111011110",
  15997=>"000001011",
  15998=>"000111000",
  15999=>"111010100",
  16000=>"110111001",
  16001=>"101101100",
  16002=>"110110110",
  16003=>"100101011",
  16004=>"011001000",
  16005=>"001110111",
  16006=>"000001001",
  16007=>"010110101",
  16008=>"001100010",
  16009=>"010011001",
  16010=>"101011000",
  16011=>"011100101",
  16012=>"010000001",
  16013=>"110000001",
  16014=>"000100101",
  16015=>"100001000",
  16016=>"110101110",
  16017=>"010010011",
  16018=>"100000100",
  16019=>"011000110",
  16020=>"101101001",
  16021=>"111101111",
  16022=>"111011101",
  16023=>"100011110",
  16024=>"111001111",
  16025=>"001000000",
  16026=>"100111101",
  16027=>"110101010",
  16028=>"111111001",
  16029=>"100010100",
  16030=>"010110101",
  16031=>"111101101",
  16032=>"111011101",
  16033=>"111001010",
  16034=>"100101001",
  16035=>"000101100",
  16036=>"101001101",
  16037=>"011000100",
  16038=>"000001011",
  16039=>"111101111",
  16040=>"001001110",
  16041=>"110010100",
  16042=>"100101010",
  16043=>"101000010",
  16044=>"100001010",
  16045=>"000101110",
  16046=>"111110101",
  16047=>"100000001",
  16048=>"100011100",
  16049=>"100110100",
  16050=>"110011111",
  16051=>"000101011",
  16052=>"000010010",
  16053=>"000010110",
  16054=>"101000001",
  16055=>"001100100",
  16056=>"111111101",
  16057=>"110100111",
  16058=>"011101111",
  16059=>"110001100",
  16060=>"111011111",
  16061=>"010110101",
  16062=>"110111110",
  16063=>"111001111",
  16064=>"010011101",
  16065=>"000110111",
  16066=>"101010001",
  16067=>"000100011",
  16068=>"010110100",
  16069=>"000101111",
  16070=>"111111010",
  16071=>"010000011",
  16072=>"110111000",
  16073=>"000001011",
  16074=>"010100000",
  16075=>"010010111",
  16076=>"111001110",
  16077=>"011011111",
  16078=>"110010101",
  16079=>"100101010",
  16080=>"001111011",
  16081=>"110101011",
  16082=>"001110101",
  16083=>"100010000",
  16084=>"100100111",
  16085=>"111101111",
  16086=>"110111111",
  16087=>"101110110",
  16088=>"001011101",
  16089=>"001001110",
  16090=>"111000000",
  16091=>"011001001",
  16092=>"000000001",
  16093=>"100000001",
  16094=>"101011101",
  16095=>"110110000",
  16096=>"100101001",
  16097=>"011110100",
  16098=>"010011000",
  16099=>"110100101",
  16100=>"101001101",
  16101=>"011001000",
  16102=>"101000111",
  16103=>"011111110",
  16104=>"110000110",
  16105=>"011010100",
  16106=>"010001001",
  16107=>"011011011",
  16108=>"100101100",
  16109=>"101011001",
  16110=>"100100011",
  16111=>"000000000",
  16112=>"011100000",
  16113=>"110110101",
  16114=>"010100110",
  16115=>"010111000",
  16116=>"101101100",
  16117=>"001100000",
  16118=>"011010101",
  16119=>"000111010",
  16120=>"011010010",
  16121=>"010010010",
  16122=>"111101111",
  16123=>"000111001",
  16124=>"100000111",
  16125=>"011000100",
  16126=>"110001101",
  16127=>"001000100",
  16128=>"100100000",
  16129=>"101111100",
  16130=>"110001010",
  16131=>"111001001",
  16132=>"100110110",
  16133=>"011000111",
  16134=>"101110010",
  16135=>"101111100",
  16136=>"000111000",
  16137=>"101011100",
  16138=>"101001111",
  16139=>"010011000",
  16140=>"100010100",
  16141=>"010111111",
  16142=>"111000100",
  16143=>"010011101",
  16144=>"001010110",
  16145=>"001011101",
  16146=>"011010101",
  16147=>"010111100",
  16148=>"011010000",
  16149=>"010001001",
  16150=>"101001100",
  16151=>"101101111",
  16152=>"111000101",
  16153=>"111100000",
  16154=>"101011001",
  16155=>"011110000",
  16156=>"110000000",
  16157=>"011111111",
  16158=>"011011101",
  16159=>"110101100",
  16160=>"100011110",
  16161=>"100000001",
  16162=>"001100100",
  16163=>"111111010",
  16164=>"011011010",
  16165=>"100000100",
  16166=>"000111010",
  16167=>"100001010",
  16168=>"000010111",
  16169=>"110000110",
  16170=>"000110100",
  16171=>"101101101",
  16172=>"001011001",
  16173=>"110100000",
  16174=>"010101001",
  16175=>"000010110",
  16176=>"110000100",
  16177=>"000000111",
  16178=>"000010010",
  16179=>"111010110",
  16180=>"110010101",
  16181=>"001000011",
  16182=>"111111110",
  16183=>"010101000",
  16184=>"101101010",
  16185=>"011011010",
  16186=>"110001000",
  16187=>"001010001",
  16188=>"110011101",
  16189=>"110001110",
  16190=>"000000000",
  16191=>"000100110",
  16192=>"100001100",
  16193=>"001011000",
  16194=>"000000101",
  16195=>"100110000",
  16196=>"011000001",
  16197=>"000000101",
  16198=>"100000010",
  16199=>"101000111",
  16200=>"010110000",
  16201=>"011011101",
  16202=>"111010100",
  16203=>"101001100",
  16204=>"101010011",
  16205=>"100111111",
  16206=>"111101110",
  16207=>"000100011",
  16208=>"011000111",
  16209=>"100010010",
  16210=>"110010001",
  16211=>"111000101",
  16212=>"110000000",
  16213=>"110110011",
  16214=>"110000100",
  16215=>"101111001",
  16216=>"101000110",
  16217=>"101111000",
  16218=>"001001111",
  16219=>"010011101",
  16220=>"000000010",
  16221=>"010001011",
  16222=>"101100100",
  16223=>"111011001",
  16224=>"100000010",
  16225=>"011111000",
  16226=>"000110010",
  16227=>"100101101",
  16228=>"011011010",
  16229=>"011000111",
  16230=>"001010000",
  16231=>"110111101",
  16232=>"010111001",
  16233=>"111100000",
  16234=>"110100000",
  16235=>"011110110",
  16236=>"100110000",
  16237=>"110100000",
  16238=>"001001011",
  16239=>"010000101",
  16240=>"110001100",
  16241=>"100000110",
  16242=>"010100000",
  16243=>"000100101",
  16244=>"101101110",
  16245=>"010010110",
  16246=>"111000100",
  16247=>"001110010",
  16248=>"111110110",
  16249=>"000000000",
  16250=>"000101000",
  16251=>"100111101",
  16252=>"010100110",
  16253=>"111000000",
  16254=>"101001001",
  16255=>"000110110",
  16256=>"010101001",
  16257=>"111011000",
  16258=>"111010011",
  16259=>"111010001",
  16260=>"011001101",
  16261=>"011100010",
  16262=>"110001001",
  16263=>"110011110",
  16264=>"111011000",
  16265=>"111101010",
  16266=>"100110111",
  16267=>"111010111",
  16268=>"110111010",
  16269=>"110110111",
  16270=>"101101000",
  16271=>"001001100",
  16272=>"101100101",
  16273=>"010100101",
  16274=>"011000011",
  16275=>"100001110",
  16276=>"010110011",
  16277=>"110111111",
  16278=>"010011011",
  16279=>"011010110",
  16280=>"000001000",
  16281=>"100100101",
  16282=>"111111111",
  16283=>"010010111",
  16284=>"110010001",
  16285=>"101111010",
  16286=>"100001011",
  16287=>"101001100",
  16288=>"110000010",
  16289=>"111110110",
  16290=>"110001111",
  16291=>"101111101",
  16292=>"011101001",
  16293=>"010110101",
  16294=>"111101111",
  16295=>"111110110",
  16296=>"110010100",
  16297=>"100010100",
  16298=>"000111111",
  16299=>"110000111",
  16300=>"110001010",
  16301=>"001111111",
  16302=>"000010010",
  16303=>"110011001",
  16304=>"000111000",
  16305=>"111001000",
  16306=>"111001110",
  16307=>"011010010",
  16308=>"000000100",
  16309=>"101011111",
  16310=>"100011111",
  16311=>"000000011",
  16312=>"110000111",
  16313=>"111100100",
  16314=>"000100000",
  16315=>"011001010",
  16316=>"100111111",
  16317=>"101011011",
  16318=>"111100101",
  16319=>"111101111",
  16320=>"001010001",
  16321=>"100011111",
  16322=>"100110111",
  16323=>"000100100",
  16324=>"010011011",
  16325=>"110101111",
  16326=>"110010100",
  16327=>"001001111",
  16328=>"010001011",
  16329=>"011010010",
  16330=>"001111101",
  16331=>"100011110",
  16332=>"001011110",
  16333=>"010011011",
  16334=>"001101100",
  16335=>"110100001",
  16336=>"100000010",
  16337=>"001100000",
  16338=>"001110100",
  16339=>"101100000",
  16340=>"010101010",
  16341=>"001001110",
  16342=>"010111000",
  16343=>"111001111",
  16344=>"111100000",
  16345=>"001100110",
  16346=>"111111111",
  16347=>"011010101",
  16348=>"110110110",
  16349=>"110100100",
  16350=>"011000000",
  16351=>"000000010",
  16352=>"111100100",
  16353=>"100100110",
  16354=>"011010010",
  16355=>"110101010",
  16356=>"100101001",
  16357=>"111001000",
  16358=>"011101000",
  16359=>"111100000",
  16360=>"001111001",
  16361=>"111101100",
  16362=>"101110011",
  16363=>"111001011",
  16364=>"100101001",
  16365=>"101111001",
  16366=>"011111011",
  16367=>"011111100",
  16368=>"110000011",
  16369=>"011101011",
  16370=>"101001111",
  16371=>"111111011",
  16372=>"001001011",
  16373=>"101111101",
  16374=>"001110001",
  16375=>"111111101",
  16376=>"001110010",
  16377=>"111011101",
  16378=>"010011001",
  16379=>"101110101",
  16380=>"110011001",
  16381=>"010001111",
  16382=>"010010000",
  16383=>"001100001",
  16384=>"010111111",
  16385=>"101011010",
  16386=>"111101010",
  16387=>"101100110",
  16388=>"111011100",
  16389=>"010110000",
  16390=>"010000000",
  16391=>"000111000",
  16392=>"011100111",
  16393=>"011011000",
  16394=>"100110100",
  16395=>"111001101",
  16396=>"110000001",
  16397=>"110100011",
  16398=>"000100001",
  16399=>"101111101",
  16400=>"101110100",
  16401=>"000111000",
  16402=>"110000100",
  16403=>"111111111",
  16404=>"101100100",
  16405=>"100101000",
  16406=>"101000010",
  16407=>"000101110",
  16408=>"100100000",
  16409=>"000010010",
  16410=>"101011001",
  16411=>"111100000",
  16412=>"010011001",
  16413=>"000001000",
  16414=>"001001100",
  16415=>"100000011",
  16416=>"100000111",
  16417=>"011100100",
  16418=>"100011110",
  16419=>"101101100",
  16420=>"011101001",
  16421=>"000010111",
  16422=>"001000000",
  16423=>"010010011",
  16424=>"111101111",
  16425=>"111100110",
  16426=>"110100000",
  16427=>"111011101",
  16428=>"111010100",
  16429=>"001001101",
  16430=>"000000000",
  16431=>"100000110",
  16432=>"101111011",
  16433=>"111110001",
  16434=>"101110100",
  16435=>"000011010",
  16436=>"100100111",
  16437=>"000100010",
  16438=>"100011000",
  16439=>"101010010",
  16440=>"011010001",
  16441=>"100001111",
  16442=>"001001001",
  16443=>"111100011",
  16444=>"101110101",
  16445=>"110011001",
  16446=>"111100011",
  16447=>"000010100",
  16448=>"000011101",
  16449=>"000100010",
  16450=>"000110010",
  16451=>"010111101",
  16452=>"111011010",
  16453=>"000111010",
  16454=>"111100010",
  16455=>"110001101",
  16456=>"110111000",
  16457=>"000101011",
  16458=>"111110111",
  16459=>"111011111",
  16460=>"110100100",
  16461=>"110101011",
  16462=>"011010010",
  16463=>"111100111",
  16464=>"111010001",
  16465=>"011111000",
  16466=>"100101011",
  16467=>"111011010",
  16468=>"111001111",
  16469=>"001010001",
  16470=>"010100101",
  16471=>"101101000",
  16472=>"000100110",
  16473=>"111011111",
  16474=>"100000000",
  16475=>"101001100",
  16476=>"001000110",
  16477=>"001101010",
  16478=>"000111001",
  16479=>"101101110",
  16480=>"101000000",
  16481=>"110001010",
  16482=>"000100100",
  16483=>"110110011",
  16484=>"111110011",
  16485=>"111011101",
  16486=>"101010010",
  16487=>"110000101",
  16488=>"001100011",
  16489=>"000111011",
  16490=>"000011011",
  16491=>"010011010",
  16492=>"000101010",
  16493=>"100000011",
  16494=>"001011011",
  16495=>"010001101",
  16496=>"001001111",
  16497=>"111011101",
  16498=>"111010101",
  16499=>"011010000",
  16500=>"110001111",
  16501=>"110000111",
  16502=>"011101101",
  16503=>"111011111",
  16504=>"111010111",
  16505=>"011110110",
  16506=>"111000110",
  16507=>"010001100",
  16508=>"000001100",
  16509=>"011010010",
  16510=>"100100111",
  16511=>"101011011",
  16512=>"101001110",
  16513=>"001111110",
  16514=>"110100111",
  16515=>"011011010",
  16516=>"001010001",
  16517=>"101110111",
  16518=>"110101010",
  16519=>"011010000",
  16520=>"011000100",
  16521=>"010111110",
  16522=>"101101101",
  16523=>"011010011",
  16524=>"111111110",
  16525=>"101111010",
  16526=>"011110000",
  16527=>"100111000",
  16528=>"001000010",
  16529=>"001010110",
  16530=>"000001011",
  16531=>"100011011",
  16532=>"100111011",
  16533=>"010010110",
  16534=>"100100111",
  16535=>"011110001",
  16536=>"010110100",
  16537=>"000010000",
  16538=>"111100000",
  16539=>"100000100",
  16540=>"010010010",
  16541=>"000100110",
  16542=>"000001100",
  16543=>"001010111",
  16544=>"111000010",
  16545=>"010100011",
  16546=>"111010011",
  16547=>"010101000",
  16548=>"011100100",
  16549=>"001100101",
  16550=>"101000001",
  16551=>"011100111",
  16552=>"110011111",
  16553=>"101100101",
  16554=>"110101010",
  16555=>"000101001",
  16556=>"111011010",
  16557=>"101001011",
  16558=>"100011001",
  16559=>"000110001",
  16560=>"000011011",
  16561=>"001001000",
  16562=>"100000000",
  16563=>"000001001",
  16564=>"011001100",
  16565=>"100111000",
  16566=>"111110001",
  16567=>"010001101",
  16568=>"100111010",
  16569=>"101001111",
  16570=>"101011111",
  16571=>"011000001",
  16572=>"010010110",
  16573=>"110110000",
  16574=>"111011000",
  16575=>"011110000",
  16576=>"001001010",
  16577=>"010011011",
  16578=>"110110010",
  16579=>"100111100",
  16580=>"011111110",
  16581=>"010111101",
  16582=>"111100001",
  16583=>"001000010",
  16584=>"110011001",
  16585=>"011010011",
  16586=>"000001111",
  16587=>"011111110",
  16588=>"110011011",
  16589=>"110100101",
  16590=>"001010100",
  16591=>"000001111",
  16592=>"000000111",
  16593=>"011101001",
  16594=>"001000000",
  16595=>"011000000",
  16596=>"100000000",
  16597=>"000110100",
  16598=>"100001110",
  16599=>"001010110",
  16600=>"000001111",
  16601=>"011111110",
  16602=>"100010001",
  16603=>"011001101",
  16604=>"001110110",
  16605=>"001110101",
  16606=>"101101001",
  16607=>"000001000",
  16608=>"111100110",
  16609=>"110110000",
  16610=>"000010010",
  16611=>"011111001",
  16612=>"101110111",
  16613=>"111000001",
  16614=>"011011100",
  16615=>"011001111",
  16616=>"110010000",
  16617=>"110000000",
  16618=>"000011111",
  16619=>"111010001",
  16620=>"010101111",
  16621=>"000001100",
  16622=>"000011101",
  16623=>"001000010",
  16624=>"110110100",
  16625=>"000101100",
  16626=>"100001100",
  16627=>"101000010",
  16628=>"011001110",
  16629=>"011101000",
  16630=>"010001011",
  16631=>"111110100",
  16632=>"010100000",
  16633=>"010010011",
  16634=>"110010000",
  16635=>"100000001",
  16636=>"011110111",
  16637=>"000000101",
  16638=>"110010101",
  16639=>"101000111",
  16640=>"001000110",
  16641=>"001000000",
  16642=>"110010101",
  16643=>"000110111",
  16644=>"100000001",
  16645=>"110101101",
  16646=>"001100100",
  16647=>"011001011",
  16648=>"110001001",
  16649=>"100100111",
  16650=>"111010101",
  16651=>"101101100",
  16652=>"010010010",
  16653=>"100001110",
  16654=>"000010101",
  16655=>"011001111",
  16656=>"000111100",
  16657=>"111000000",
  16658=>"000010101",
  16659=>"010011001",
  16660=>"101101101",
  16661=>"010001100",
  16662=>"100011111",
  16663=>"000101000",
  16664=>"110110100",
  16665=>"011001100",
  16666=>"001001100",
  16667=>"111110000",
  16668=>"000101010",
  16669=>"001110001",
  16670=>"110101010",
  16671=>"111101110",
  16672=>"101110001",
  16673=>"111101101",
  16674=>"101011011",
  16675=>"101010010",
  16676=>"010100000",
  16677=>"010101111",
  16678=>"010110010",
  16679=>"011111010",
  16680=>"000000000",
  16681=>"010101110",
  16682=>"111001111",
  16683=>"001101110",
  16684=>"101001001",
  16685=>"011011011",
  16686=>"101101010",
  16687=>"011110011",
  16688=>"001000111",
  16689=>"011010100",
  16690=>"111101110",
  16691=>"101110110",
  16692=>"100101010",
  16693=>"101110001",
  16694=>"001000011",
  16695=>"000100101",
  16696=>"110100000",
  16697=>"011101101",
  16698=>"111010011",
  16699=>"111100101",
  16700=>"110111110",
  16701=>"000011010",
  16702=>"000001011",
  16703=>"111001011",
  16704=>"000011100",
  16705=>"100010000",
  16706=>"111111101",
  16707=>"100010100",
  16708=>"011011010",
  16709=>"011111111",
  16710=>"011100000",
  16711=>"011000101",
  16712=>"111010110",
  16713=>"100101001",
  16714=>"100010000",
  16715=>"110111111",
  16716=>"101011000",
  16717=>"010111010",
  16718=>"000110010",
  16719=>"001000110",
  16720=>"110110011",
  16721=>"011101110",
  16722=>"001000000",
  16723=>"011011101",
  16724=>"110110010",
  16725=>"110100100",
  16726=>"100000001",
  16727=>"111000000",
  16728=>"001111011",
  16729=>"000011000",
  16730=>"001001000",
  16731=>"010000000",
  16732=>"000010100",
  16733=>"001001001",
  16734=>"100001010",
  16735=>"001100111",
  16736=>"001101010",
  16737=>"011110010",
  16738=>"001001000",
  16739=>"010100011",
  16740=>"000000000",
  16741=>"011000010",
  16742=>"000100111",
  16743=>"011111000",
  16744=>"101000111",
  16745=>"101011101",
  16746=>"001000001",
  16747=>"101010010",
  16748=>"000100111",
  16749=>"100000011",
  16750=>"001010000",
  16751=>"001100000",
  16752=>"100001000",
  16753=>"111100011",
  16754=>"000010001",
  16755=>"010100011",
  16756=>"111100101",
  16757=>"011110001",
  16758=>"100000111",
  16759=>"011010111",
  16760=>"011110010",
  16761=>"100011000",
  16762=>"010000100",
  16763=>"011101011",
  16764=>"010101110",
  16765=>"000110010",
  16766=>"011011011",
  16767=>"011100011",
  16768=>"000000100",
  16769=>"001111011",
  16770=>"100101001",
  16771=>"010111010",
  16772=>"100110101",
  16773=>"000101111",
  16774=>"101101101",
  16775=>"111100111",
  16776=>"010111010",
  16777=>"101100000",
  16778=>"000001010",
  16779=>"110111111",
  16780=>"010001000",
  16781=>"010111001",
  16782=>"011000001",
  16783=>"001100001",
  16784=>"010001110",
  16785=>"001000110",
  16786=>"100111011",
  16787=>"010000100",
  16788=>"001110010",
  16789=>"100111010",
  16790=>"111100111",
  16791=>"101100001",
  16792=>"000001101",
  16793=>"010001110",
  16794=>"001100101",
  16795=>"011100101",
  16796=>"101100100",
  16797=>"111110110",
  16798=>"111111011",
  16799=>"111011110",
  16800=>"111001001",
  16801=>"000110000",
  16802=>"101010110",
  16803=>"011111010",
  16804=>"010100110",
  16805=>"001000111",
  16806=>"101111100",
  16807=>"001111111",
  16808=>"000101110",
  16809=>"110111000",
  16810=>"010001000",
  16811=>"000100011",
  16812=>"010000001",
  16813=>"101110001",
  16814=>"010111010",
  16815=>"110111111",
  16816=>"011000000",
  16817=>"011111011",
  16818=>"110000010",
  16819=>"101100111",
  16820=>"101000100",
  16821=>"110011110",
  16822=>"101111010",
  16823=>"001000000",
  16824=>"000100111",
  16825=>"111001111",
  16826=>"100110101",
  16827=>"101011010",
  16828=>"011001111",
  16829=>"001100000",
  16830=>"010110011",
  16831=>"010100000",
  16832=>"001000001",
  16833=>"001110100",
  16834=>"000001100",
  16835=>"110011001",
  16836=>"100010000",
  16837=>"101101110",
  16838=>"111101011",
  16839=>"100111100",
  16840=>"001001101",
  16841=>"110111100",
  16842=>"010000101",
  16843=>"011101011",
  16844=>"001101010",
  16845=>"011110111",
  16846=>"111101111",
  16847=>"110001011",
  16848=>"101100111",
  16849=>"001000100",
  16850=>"110011010",
  16851=>"110010110",
  16852=>"101110000",
  16853=>"000010011",
  16854=>"011001010",
  16855=>"000001011",
  16856=>"011101000",
  16857=>"001001010",
  16858=>"011110100",
  16859=>"000011000",
  16860=>"111001110",
  16861=>"111111101",
  16862=>"001101110",
  16863=>"000111101",
  16864=>"111110110",
  16865=>"010011010",
  16866=>"110110100",
  16867=>"100110011",
  16868=>"110100000",
  16869=>"001010011",
  16870=>"110100110",
  16871=>"100011000",
  16872=>"100100101",
  16873=>"010110000",
  16874=>"000000000",
  16875=>"000100110",
  16876=>"001001010",
  16877=>"001010110",
  16878=>"000101111",
  16879=>"100011101",
  16880=>"101001110",
  16881=>"110010001",
  16882=>"100110010",
  16883=>"110101110",
  16884=>"100001110",
  16885=>"111010101",
  16886=>"011010111",
  16887=>"000110011",
  16888=>"011101110",
  16889=>"111100011",
  16890=>"000000010",
  16891=>"101110011",
  16892=>"111001111",
  16893=>"000010111",
  16894=>"111011001",
  16895=>"110011010",
  16896=>"101110001",
  16897=>"110010101",
  16898=>"101110111",
  16899=>"001010011",
  16900=>"000010000",
  16901=>"100110001",
  16902=>"001011101",
  16903=>"111101000",
  16904=>"010000110",
  16905=>"001100111",
  16906=>"010011100",
  16907=>"010010111",
  16908=>"001001000",
  16909=>"000111000",
  16910=>"011010101",
  16911=>"001110010",
  16912=>"100000000",
  16913=>"100001010",
  16914=>"000101101",
  16915=>"100001101",
  16916=>"101100101",
  16917=>"000110010",
  16918=>"010100010",
  16919=>"011111110",
  16920=>"100011011",
  16921=>"101100101",
  16922=>"011010111",
  16923=>"101111001",
  16924=>"001101111",
  16925=>"110101110",
  16926=>"001011100",
  16927=>"010001111",
  16928=>"011011001",
  16929=>"100100001",
  16930=>"011100000",
  16931=>"000101111",
  16932=>"011010010",
  16933=>"000000101",
  16934=>"101001100",
  16935=>"101101100",
  16936=>"110001100",
  16937=>"010111000",
  16938=>"011001000",
  16939=>"001101000",
  16940=>"111101011",
  16941=>"001010001",
  16942=>"011101001",
  16943=>"100100000",
  16944=>"001110001",
  16945=>"100111000",
  16946=>"010011101",
  16947=>"111110001",
  16948=>"111010001",
  16949=>"010001100",
  16950=>"010000101",
  16951=>"100010101",
  16952=>"000101110",
  16953=>"000100001",
  16954=>"111110110",
  16955=>"010110010",
  16956=>"010001101",
  16957=>"111111100",
  16958=>"000000100",
  16959=>"011001011",
  16960=>"111001110",
  16961=>"110111100",
  16962=>"010001010",
  16963=>"111000000",
  16964=>"000011111",
  16965=>"111111001",
  16966=>"100010000",
  16967=>"001000010",
  16968=>"111001000",
  16969=>"000100000",
  16970=>"000101010",
  16971=>"001101110",
  16972=>"000101001",
  16973=>"100000010",
  16974=>"001010011",
  16975=>"100001101",
  16976=>"011010010",
  16977=>"010010100",
  16978=>"001001000",
  16979=>"011100101",
  16980=>"100000000",
  16981=>"100100000",
  16982=>"001100001",
  16983=>"101011000",
  16984=>"000010101",
  16985=>"101000011",
  16986=>"101011011",
  16987=>"011001111",
  16988=>"100010101",
  16989=>"001101000",
  16990=>"000000100",
  16991=>"100110001",
  16992=>"000001100",
  16993=>"100010111",
  16994=>"111010001",
  16995=>"000010011",
  16996=>"101000001",
  16997=>"001110111",
  16998=>"100001010",
  16999=>"110011010",
  17000=>"000011101",
  17001=>"100010000",
  17002=>"110010111",
  17003=>"111111111",
  17004=>"000001001",
  17005=>"111011001",
  17006=>"010001100",
  17007=>"110010101",
  17008=>"000010110",
  17009=>"100110110",
  17010=>"100001000",
  17011=>"011001100",
  17012=>"010001110",
  17013=>"111010101",
  17014=>"011101110",
  17015=>"011100110",
  17016=>"100110100",
  17017=>"110101010",
  17018=>"001101011",
  17019=>"010101101",
  17020=>"111110000",
  17021=>"010010000",
  17022=>"011111011",
  17023=>"110000010",
  17024=>"000010010",
  17025=>"101000100",
  17026=>"011000011",
  17027=>"101010011",
  17028=>"001111010",
  17029=>"000101100",
  17030=>"010110110",
  17031=>"000110101",
  17032=>"010100111",
  17033=>"110000101",
  17034=>"101111111",
  17035=>"101010000",
  17036=>"100111100",
  17037=>"011001100",
  17038=>"101010001",
  17039=>"110010101",
  17040=>"000100001",
  17041=>"100010010",
  17042=>"001010011",
  17043=>"011010000",
  17044=>"000000010",
  17045=>"001001101",
  17046=>"001110101",
  17047=>"110001100",
  17048=>"011011000",
  17049=>"000101001",
  17050=>"100100101",
  17051=>"111110100",
  17052=>"100111010",
  17053=>"010010001",
  17054=>"111010100",
  17055=>"010001100",
  17056=>"101100000",
  17057=>"010000101",
  17058=>"001101111",
  17059=>"101100101",
  17060=>"000110110",
  17061=>"001011000",
  17062=>"101110110",
  17063=>"000111001",
  17064=>"110110100",
  17065=>"100101011",
  17066=>"010111000",
  17067=>"010110011",
  17068=>"101100010",
  17069=>"101011011",
  17070=>"001000111",
  17071=>"000111101",
  17072=>"111001111",
  17073=>"100010000",
  17074=>"100001100",
  17075=>"110010000",
  17076=>"110011110",
  17077=>"001111000",
  17078=>"100110001",
  17079=>"001101011",
  17080=>"110011111",
  17081=>"001100011",
  17082=>"011111111",
  17083=>"010010110",
  17084=>"010100111",
  17085=>"110011010",
  17086=>"101101001",
  17087=>"111110111",
  17088=>"000111010",
  17089=>"110010010",
  17090=>"000111011",
  17091=>"110010111",
  17092=>"011111111",
  17093=>"010011000",
  17094=>"100101111",
  17095=>"000010101",
  17096=>"100011110",
  17097=>"010101001",
  17098=>"010101001",
  17099=>"011110011",
  17100=>"000011110",
  17101=>"110110010",
  17102=>"000100100",
  17103=>"111110110",
  17104=>"111011001",
  17105=>"100100001",
  17106=>"110111100",
  17107=>"000000001",
  17108=>"111010101",
  17109=>"010001101",
  17110=>"100001100",
  17111=>"010100111",
  17112=>"010100111",
  17113=>"100100110",
  17114=>"111110001",
  17115=>"101001101",
  17116=>"000001000",
  17117=>"001100011",
  17118=>"000010001",
  17119=>"110000101",
  17120=>"010101011",
  17121=>"011001000",
  17122=>"010010100",
  17123=>"111101011",
  17124=>"100000100",
  17125=>"011100011",
  17126=>"001001101",
  17127=>"110000010",
  17128=>"001111010",
  17129=>"101111010",
  17130=>"011101110",
  17131=>"111110110",
  17132=>"011000101",
  17133=>"111110001",
  17134=>"011000000",
  17135=>"000100000",
  17136=>"001000100",
  17137=>"010011001",
  17138=>"000000010",
  17139=>"001000010",
  17140=>"110101100",
  17141=>"001110100",
  17142=>"011111010",
  17143=>"010000111",
  17144=>"001111011",
  17145=>"011110100",
  17146=>"000111100",
  17147=>"010011100",
  17148=>"110111000",
  17149=>"010011011",
  17150=>"001010000",
  17151=>"001110110",
  17152=>"010101001",
  17153=>"000001111",
  17154=>"101001111",
  17155=>"000010110",
  17156=>"101001100",
  17157=>"101011001",
  17158=>"011100010",
  17159=>"001111010",
  17160=>"001000100",
  17161=>"110110010",
  17162=>"010000011",
  17163=>"111000100",
  17164=>"001010000",
  17165=>"101110111",
  17166=>"010110000",
  17167=>"010001100",
  17168=>"011000001",
  17169=>"001001000",
  17170=>"010010110",
  17171=>"001110111",
  17172=>"101011110",
  17173=>"010111100",
  17174=>"000110000",
  17175=>"100010101",
  17176=>"111100010",
  17177=>"010111100",
  17178=>"001000001",
  17179=>"101001101",
  17180=>"001000111",
  17181=>"000101110",
  17182=>"001010010",
  17183=>"011100011",
  17184=>"000010101",
  17185=>"100101111",
  17186=>"000101010",
  17187=>"001010011",
  17188=>"110100010",
  17189=>"000010001",
  17190=>"000111010",
  17191=>"000010011",
  17192=>"010101100",
  17193=>"001110100",
  17194=>"000010010",
  17195=>"101111001",
  17196=>"101010000",
  17197=>"000001011",
  17198=>"100001010",
  17199=>"001100111",
  17200=>"010110011",
  17201=>"110011111",
  17202=>"001101111",
  17203=>"110000101",
  17204=>"110010111",
  17205=>"011011111",
  17206=>"001111001",
  17207=>"010111010",
  17208=>"101010010",
  17209=>"001011111",
  17210=>"000001000",
  17211=>"100011001",
  17212=>"010111111",
  17213=>"111001000",
  17214=>"000101100",
  17215=>"011110110",
  17216=>"110101000",
  17217=>"010011100",
  17218=>"011000010",
  17219=>"111111101",
  17220=>"010100010",
  17221=>"001001001",
  17222=>"101111000",
  17223=>"011101101",
  17224=>"100100110",
  17225=>"011100100",
  17226=>"100010101",
  17227=>"010001010",
  17228=>"101000001",
  17229=>"011000110",
  17230=>"001111011",
  17231=>"100100001",
  17232=>"001000101",
  17233=>"101110001",
  17234=>"011100110",
  17235=>"011100111",
  17236=>"110110000",
  17237=>"001010001",
  17238=>"001101000",
  17239=>"011000000",
  17240=>"010000110",
  17241=>"101000010",
  17242=>"111001100",
  17243=>"000000111",
  17244=>"011101010",
  17245=>"111111011",
  17246=>"010000101",
  17247=>"001000110",
  17248=>"101101100",
  17249=>"100001011",
  17250=>"100100001",
  17251=>"011101100",
  17252=>"111100011",
  17253=>"100100010",
  17254=>"110000001",
  17255=>"011100001",
  17256=>"100011111",
  17257=>"010100011",
  17258=>"011101111",
  17259=>"101001101",
  17260=>"011111101",
  17261=>"100010010",
  17262=>"000000111",
  17263=>"100110111",
  17264=>"111010100",
  17265=>"011100100",
  17266=>"001100111",
  17267=>"010100111",
  17268=>"100100100",
  17269=>"100111101",
  17270=>"001100000",
  17271=>"011010011",
  17272=>"100001100",
  17273=>"011111010",
  17274=>"010100011",
  17275=>"001000110",
  17276=>"000000100",
  17277=>"100110001",
  17278=>"010101010",
  17279=>"111100111",
  17280=>"111000101",
  17281=>"000000000",
  17282=>"010110110",
  17283=>"111011100",
  17284=>"110111011",
  17285=>"000110101",
  17286=>"011000000",
  17287=>"100010011",
  17288=>"111111011",
  17289=>"001000111",
  17290=>"000000000",
  17291=>"000001000",
  17292=>"000111100",
  17293=>"110110100",
  17294=>"010111111",
  17295=>"000011011",
  17296=>"101010001",
  17297=>"010011110",
  17298=>"001000111",
  17299=>"000111100",
  17300=>"101100110",
  17301=>"011111000",
  17302=>"010010110",
  17303=>"100101111",
  17304=>"011100010",
  17305=>"100010001",
  17306=>"011001101",
  17307=>"101110000",
  17308=>"000000111",
  17309=>"000011101",
  17310=>"010011101",
  17311=>"010001110",
  17312=>"110110110",
  17313=>"110010100",
  17314=>"111000111",
  17315=>"011110000",
  17316=>"101111001",
  17317=>"011011100",
  17318=>"010001100",
  17319=>"001111011",
  17320=>"010001111",
  17321=>"111010001",
  17322=>"111000001",
  17323=>"011110011",
  17324=>"110011111",
  17325=>"011111000",
  17326=>"000011001",
  17327=>"001100011",
  17328=>"101111101",
  17329=>"111011110",
  17330=>"000111011",
  17331=>"010011001",
  17332=>"101000110",
  17333=>"001001101",
  17334=>"000010100",
  17335=>"101001001",
  17336=>"011111001",
  17337=>"010100010",
  17338=>"100101011",
  17339=>"011100110",
  17340=>"000101000",
  17341=>"001110111",
  17342=>"000000111",
  17343=>"011011011",
  17344=>"011100010",
  17345=>"001110111",
  17346=>"011100010",
  17347=>"100110000",
  17348=>"101000100",
  17349=>"000100110",
  17350=>"101000111",
  17351=>"100001000",
  17352=>"001101111",
  17353=>"101001001",
  17354=>"001000000",
  17355=>"100010101",
  17356=>"000000011",
  17357=>"110111001",
  17358=>"111100011",
  17359=>"000001001",
  17360=>"100100101",
  17361=>"010101011",
  17362=>"101010110",
  17363=>"101111100",
  17364=>"101100110",
  17365=>"000010010",
  17366=>"001011101",
  17367=>"100000111",
  17368=>"010011111",
  17369=>"010100010",
  17370=>"000001011",
  17371=>"101000111",
  17372=>"010010000",
  17373=>"110110011",
  17374=>"000001010",
  17375=>"100001001",
  17376=>"110011011",
  17377=>"111101011",
  17378=>"001111100",
  17379=>"110101010",
  17380=>"011111100",
  17381=>"001010001",
  17382=>"001000100",
  17383=>"111111100",
  17384=>"101011011",
  17385=>"010011101",
  17386=>"100011111",
  17387=>"111101010",
  17388=>"001111100",
  17389=>"110000010",
  17390=>"111100111",
  17391=>"110101111",
  17392=>"001101100",
  17393=>"011010010",
  17394=>"110110110",
  17395=>"001011011",
  17396=>"100111101",
  17397=>"110000000",
  17398=>"011100110",
  17399=>"001010010",
  17400=>"111110010",
  17401=>"111110011",
  17402=>"011101001",
  17403=>"111110011",
  17404=>"000111001",
  17405=>"111000000",
  17406=>"001110010",
  17407=>"011000111",
  17408=>"110011000",
  17409=>"000111001",
  17410=>"010100011",
  17411=>"001010000",
  17412=>"100011000",
  17413=>"111111101",
  17414=>"010101000",
  17415=>"111000110",
  17416=>"010110100",
  17417=>"100000110",
  17418=>"010111010",
  17419=>"110110010",
  17420=>"000011101",
  17421=>"101001100",
  17422=>"001000011",
  17423=>"100100010",
  17424=>"100111010",
  17425=>"000010001",
  17426=>"101011101",
  17427=>"100100100",
  17428=>"010011000",
  17429=>"111101011",
  17430=>"101100001",
  17431=>"111010001",
  17432=>"010111000",
  17433=>"001000000",
  17434=>"111010111",
  17435=>"100101100",
  17436=>"001100101",
  17437=>"101000100",
  17438=>"110100101",
  17439=>"011100111",
  17440=>"101100010",
  17441=>"010000101",
  17442=>"011100100",
  17443=>"110000011",
  17444=>"000000101",
  17445=>"011000001",
  17446=>"001101010",
  17447=>"101101100",
  17448=>"111100011",
  17449=>"110101100",
  17450=>"001001100",
  17451=>"110010100",
  17452=>"111110011",
  17453=>"111110111",
  17454=>"111010010",
  17455=>"111011101",
  17456=>"101011111",
  17457=>"000100101",
  17458=>"011110001",
  17459=>"010100110",
  17460=>"000101000",
  17461=>"110010000",
  17462=>"011011011",
  17463=>"010100111",
  17464=>"100101111",
  17465=>"000110011",
  17466=>"110000110",
  17467=>"001000110",
  17468=>"110011100",
  17469=>"111101011",
  17470=>"011000010",
  17471=>"101110000",
  17472=>"111110100",
  17473=>"000000110",
  17474=>"010001001",
  17475=>"001001110",
  17476=>"111000101",
  17477=>"000100001",
  17478=>"011110110",
  17479=>"000001001",
  17480=>"010000000",
  17481=>"111011000",
  17482=>"010010101",
  17483=>"001011011",
  17484=>"001010101",
  17485=>"100011011",
  17486=>"000011110",
  17487=>"010000100",
  17488=>"000010011",
  17489=>"101000001",
  17490=>"111110100",
  17491=>"011001001",
  17492=>"110110011",
  17493=>"011000100",
  17494=>"000111110",
  17495=>"111001111",
  17496=>"001011111",
  17497=>"100100100",
  17498=>"111000010",
  17499=>"001000010",
  17500=>"100100000",
  17501=>"100011010",
  17502=>"110110110",
  17503=>"101000100",
  17504=>"101101001",
  17505=>"110001000",
  17506=>"110010101",
  17507=>"011001000",
  17508=>"111000110",
  17509=>"101101000",
  17510=>"010100011",
  17511=>"010001010",
  17512=>"111001111",
  17513=>"011001101",
  17514=>"010110101",
  17515=>"110101001",
  17516=>"101101110",
  17517=>"010010011",
  17518=>"000010101",
  17519=>"110010001",
  17520=>"000001101",
  17521=>"110110010",
  17522=>"101010000",
  17523=>"100010100",
  17524=>"010011011",
  17525=>"110001100",
  17526=>"010110011",
  17527=>"111011101",
  17528=>"101011100",
  17529=>"001111010",
  17530=>"011110010",
  17531=>"000010010",
  17532=>"000000011",
  17533=>"111111110",
  17534=>"111100110",
  17535=>"010000101",
  17536=>"011001110",
  17537=>"011101001",
  17538=>"010000110",
  17539=>"001110011",
  17540=>"111111100",
  17541=>"110000110",
  17542=>"101000100",
  17543=>"000100010",
  17544=>"010001101",
  17545=>"011011010",
  17546=>"000111111",
  17547=>"001100000",
  17548=>"111111110",
  17549=>"001100100",
  17550=>"001001100",
  17551=>"000100010",
  17552=>"101111100",
  17553=>"100100111",
  17554=>"001100010",
  17555=>"101110011",
  17556=>"001010010",
  17557=>"100110101",
  17558=>"111101011",
  17559=>"100101101",
  17560=>"000011000",
  17561=>"011000001",
  17562=>"011001111",
  17563=>"011101100",
  17564=>"001110111",
  17565=>"111101010",
  17566=>"100101001",
  17567=>"001010100",
  17568=>"011011000",
  17569=>"101101100",
  17570=>"110110011",
  17571=>"001101010",
  17572=>"010001111",
  17573=>"110111101",
  17574=>"100110001",
  17575=>"000001111",
  17576=>"001110110",
  17577=>"100100011",
  17578=>"000000101",
  17579=>"000000101",
  17580=>"011110110",
  17581=>"010000000",
  17582=>"111101101",
  17583=>"000000111",
  17584=>"011100111",
  17585=>"110110101",
  17586=>"000001000",
  17587=>"001011001",
  17588=>"010001001",
  17589=>"011101110",
  17590=>"010100011",
  17591=>"011101111",
  17592=>"100011010",
  17593=>"101001100",
  17594=>"101001000",
  17595=>"111110111",
  17596=>"000101000",
  17597=>"000011010",
  17598=>"111000000",
  17599=>"011001111",
  17600=>"110110010",
  17601=>"011111011",
  17602=>"101101011",
  17603=>"100001110",
  17604=>"101100000",
  17605=>"000010001",
  17606=>"110111011",
  17607=>"101010001",
  17608=>"100000000",
  17609=>"100100100",
  17610=>"111100101",
  17611=>"011011000",
  17612=>"011110100",
  17613=>"001000011",
  17614=>"110000100",
  17615=>"101011100",
  17616=>"000100010",
  17617=>"100110010",
  17618=>"000001001",
  17619=>"000000101",
  17620=>"011111001",
  17621=>"000101010",
  17622=>"001101110",
  17623=>"000010101",
  17624=>"101000010",
  17625=>"000000110",
  17626=>"111111000",
  17627=>"011110110",
  17628=>"101011000",
  17629=>"101110011",
  17630=>"011111010",
  17631=>"000001010",
  17632=>"010000011",
  17633=>"101000110",
  17634=>"001010001",
  17635=>"101010101",
  17636=>"101111001",
  17637=>"010111101",
  17638=>"101100011",
  17639=>"101010110",
  17640=>"000010100",
  17641=>"010011110",
  17642=>"011010010",
  17643=>"001100101",
  17644=>"000010111",
  17645=>"110110101",
  17646=>"100101101",
  17647=>"011101000",
  17648=>"011001101",
  17649=>"010011010",
  17650=>"000010110",
  17651=>"011001001",
  17652=>"101001100",
  17653=>"110111001",
  17654=>"010011101",
  17655=>"000011011",
  17656=>"111001101",
  17657=>"111001000",
  17658=>"011001000",
  17659=>"110011000",
  17660=>"011110010",
  17661=>"011100001",
  17662=>"111100011",
  17663=>"111001100",
  17664=>"011011000",
  17665=>"110100000",
  17666=>"000101011",
  17667=>"000001000",
  17668=>"001010011",
  17669=>"010111000",
  17670=>"110110100",
  17671=>"000001101",
  17672=>"010101100",
  17673=>"100100100",
  17674=>"100111110",
  17675=>"111100111",
  17676=>"001101001",
  17677=>"000111100",
  17678=>"100110000",
  17679=>"101010010",
  17680=>"101111101",
  17681=>"000110101",
  17682=>"111101001",
  17683=>"100001010",
  17684=>"101111001",
  17685=>"100101111",
  17686=>"110111010",
  17687=>"101000101",
  17688=>"100010000",
  17689=>"111111000",
  17690=>"010001011",
  17691=>"101111110",
  17692=>"110010100",
  17693=>"100001110",
  17694=>"011100001",
  17695=>"010000100",
  17696=>"011000011",
  17697=>"100101100",
  17698=>"111010101",
  17699=>"100000011",
  17700=>"000010011",
  17701=>"001101000",
  17702=>"101101010",
  17703=>"001111110",
  17704=>"000000000",
  17705=>"100000110",
  17706=>"111000011",
  17707=>"010101111",
  17708=>"011110110",
  17709=>"101001011",
  17710=>"010110000",
  17711=>"101001011",
  17712=>"001000010",
  17713=>"110000111",
  17714=>"001111111",
  17715=>"001010111",
  17716=>"100011101",
  17717=>"001100011",
  17718=>"100101000",
  17719=>"010110101",
  17720=>"111100110",
  17721=>"110010111",
  17722=>"000100110",
  17723=>"110110001",
  17724=>"010010001",
  17725=>"111101000",
  17726=>"000111101",
  17727=>"011001110",
  17728=>"010010000",
  17729=>"100011000",
  17730=>"011110100",
  17731=>"000111010",
  17732=>"011011111",
  17733=>"001101001",
  17734=>"110000011",
  17735=>"011010010",
  17736=>"010110010",
  17737=>"000010110",
  17738=>"001001101",
  17739=>"010110100",
  17740=>"111110011",
  17741=>"001100010",
  17742=>"011110000",
  17743=>"100110110",
  17744=>"111000011",
  17745=>"000111001",
  17746=>"010100011",
  17747=>"111100000",
  17748=>"110001110",
  17749=>"011000001",
  17750=>"001010100",
  17751=>"001111101",
  17752=>"010000010",
  17753=>"011001110",
  17754=>"101101101",
  17755=>"010000010",
  17756=>"110101000",
  17757=>"011000001",
  17758=>"110001001",
  17759=>"011100100",
  17760=>"110111100",
  17761=>"001111001",
  17762=>"000110001",
  17763=>"010110000",
  17764=>"000000001",
  17765=>"111110111",
  17766=>"011101000",
  17767=>"111111000",
  17768=>"101011010",
  17769=>"011010001",
  17770=>"110001100",
  17771=>"110010110",
  17772=>"001111010",
  17773=>"111110101",
  17774=>"001000001",
  17775=>"111101110",
  17776=>"000100111",
  17777=>"101001001",
  17778=>"111001001",
  17779=>"011100000",
  17780=>"111110001",
  17781=>"100101110",
  17782=>"010000111",
  17783=>"011001011",
  17784=>"001101011",
  17785=>"111110010",
  17786=>"010110101",
  17787=>"100011011",
  17788=>"111111001",
  17789=>"000010000",
  17790=>"100111010",
  17791=>"000111110",
  17792=>"011000101",
  17793=>"010000000",
  17794=>"000000101",
  17795=>"001101111",
  17796=>"100101110",
  17797=>"000101110",
  17798=>"100110001",
  17799=>"010011000",
  17800=>"000010000",
  17801=>"111100001",
  17802=>"101011110",
  17803=>"001110111",
  17804=>"101001000",
  17805=>"011101100",
  17806=>"000111000",
  17807=>"101000000",
  17808=>"100011111",
  17809=>"100111000",
  17810=>"000111111",
  17811=>"111010100",
  17812=>"011000101",
  17813=>"000000011",
  17814=>"101001101",
  17815=>"111100111",
  17816=>"100011101",
  17817=>"000001001",
  17818=>"110011001",
  17819=>"111001110",
  17820=>"011001111",
  17821=>"000000111",
  17822=>"011011100",
  17823=>"010001101",
  17824=>"000011101",
  17825=>"100010110",
  17826=>"001100110",
  17827=>"101110000",
  17828=>"110111100",
  17829=>"110000111",
  17830=>"011111011",
  17831=>"011001110",
  17832=>"000101110",
  17833=>"001000010",
  17834=>"111100000",
  17835=>"010001110",
  17836=>"110101111",
  17837=>"011011101",
  17838=>"000110000",
  17839=>"100100000",
  17840=>"011001111",
  17841=>"010011001",
  17842=>"111111110",
  17843=>"110000000",
  17844=>"111000100",
  17845=>"111100011",
  17846=>"110110000",
  17847=>"000001011",
  17848=>"001101001",
  17849=>"101101011",
  17850=>"111010101",
  17851=>"100001110",
  17852=>"000000110",
  17853=>"000100100",
  17854=>"100001001",
  17855=>"101111101",
  17856=>"001110110",
  17857=>"100000000",
  17858=>"010110001",
  17859=>"010011100",
  17860=>"000000001",
  17861=>"110011011",
  17862=>"101000110",
  17863=>"000101110",
  17864=>"010111001",
  17865=>"000000010",
  17866=>"101000001",
  17867=>"010000100",
  17868=>"000101011",
  17869=>"000101100",
  17870=>"111101011",
  17871=>"001001001",
  17872=>"011111100",
  17873=>"010111011",
  17874=>"010100001",
  17875=>"010001000",
  17876=>"111110010",
  17877=>"111111011",
  17878=>"000010010",
  17879=>"100001010",
  17880=>"101001011",
  17881=>"100111110",
  17882=>"100100000",
  17883=>"111011010",
  17884=>"101101010",
  17885=>"010101000",
  17886=>"100010110",
  17887=>"110010110",
  17888=>"101000100",
  17889=>"001001111",
  17890=>"000000000",
  17891=>"001011010",
  17892=>"000111100",
  17893=>"011110010",
  17894=>"110101101",
  17895=>"100000111",
  17896=>"001010010",
  17897=>"000010110",
  17898=>"011101101",
  17899=>"010001011",
  17900=>"111011100",
  17901=>"110001111",
  17902=>"000111010",
  17903=>"011000111",
  17904=>"000111111",
  17905=>"011001001",
  17906=>"111100101",
  17907=>"101101100",
  17908=>"001000111",
  17909=>"110111010",
  17910=>"101011110",
  17911=>"001111101",
  17912=>"100101010",
  17913=>"011000101",
  17914=>"001110100",
  17915=>"000111111",
  17916=>"110010100",
  17917=>"111101110",
  17918=>"101111011",
  17919=>"111000100",
  17920=>"100001010",
  17921=>"100010110",
  17922=>"011100010",
  17923=>"011101101",
  17924=>"110111011",
  17925=>"111110111",
  17926=>"110001110",
  17927=>"011001101",
  17928=>"000010101",
  17929=>"010101100",
  17930=>"101010011",
  17931=>"100111100",
  17932=>"101101011",
  17933=>"011011110",
  17934=>"011010000",
  17935=>"110110010",
  17936=>"110111000",
  17937=>"010000101",
  17938=>"001001111",
  17939=>"001010010",
  17940=>"010010111",
  17941=>"110101111",
  17942=>"100100000",
  17943=>"000100010",
  17944=>"011001011",
  17945=>"010000010",
  17946=>"001111110",
  17947=>"110001101",
  17948=>"101000101",
  17949=>"001101111",
  17950=>"000101110",
  17951=>"011000110",
  17952=>"011001111",
  17953=>"101010111",
  17954=>"010111101",
  17955=>"011000000",
  17956=>"100110010",
  17957=>"001000011",
  17958=>"010110100",
  17959=>"100010000",
  17960=>"111001110",
  17961=>"011111010",
  17962=>"000100010",
  17963=>"111111110",
  17964=>"011011011",
  17965=>"110001100",
  17966=>"001111110",
  17967=>"001000000",
  17968=>"111011011",
  17969=>"100001111",
  17970=>"100110111",
  17971=>"001010101",
  17972=>"001001000",
  17973=>"000110111",
  17974=>"111111000",
  17975=>"101000010",
  17976=>"011010100",
  17977=>"111110010",
  17978=>"101011101",
  17979=>"111010101",
  17980=>"011001101",
  17981=>"000010110",
  17982=>"001000001",
  17983=>"000101100",
  17984=>"110010001",
  17985=>"101010110",
  17986=>"011000000",
  17987=>"111100010",
  17988=>"000011110",
  17989=>"010011000",
  17990=>"000001000",
  17991=>"101101000",
  17992=>"101010000",
  17993=>"000011001",
  17994=>"011011000",
  17995=>"111000111",
  17996=>"010111100",
  17997=>"001010111",
  17998=>"001010001",
  17999=>"000100101",
  18000=>"000000000",
  18001=>"001010001",
  18002=>"000010001",
  18003=>"100010001",
  18004=>"000010011",
  18005=>"001110000",
  18006=>"111110111",
  18007=>"110010110",
  18008=>"110110011",
  18009=>"011100011",
  18010=>"001010001",
  18011=>"000101111",
  18012=>"110000011",
  18013=>"100011000",
  18014=>"111000110",
  18015=>"111001010",
  18016=>"100100110",
  18017=>"000111001",
  18018=>"011110101",
  18019=>"011011101",
  18020=>"011001101",
  18021=>"000000101",
  18022=>"001111000",
  18023=>"110110111",
  18024=>"011000110",
  18025=>"001000111",
  18026=>"011110010",
  18027=>"100111111",
  18028=>"100010011",
  18029=>"011011110",
  18030=>"011001100",
  18031=>"010111110",
  18032=>"001110000",
  18033=>"111111001",
  18034=>"110000111",
  18035=>"011001010",
  18036=>"001000111",
  18037=>"011000010",
  18038=>"001011011",
  18039=>"001000000",
  18040=>"110010111",
  18041=>"101110111",
  18042=>"101101001",
  18043=>"011100111",
  18044=>"011001100",
  18045=>"100100010",
  18046=>"110111001",
  18047=>"001000001",
  18048=>"000001101",
  18049=>"001000100",
  18050=>"000010111",
  18051=>"000101101",
  18052=>"010000010",
  18053=>"110101000",
  18054=>"010000101",
  18055=>"101011111",
  18056=>"111011101",
  18057=>"001001011",
  18058=>"111110101",
  18059=>"100100001",
  18060=>"010000110",
  18061=>"100101000",
  18062=>"001111001",
  18063=>"100011111",
  18064=>"110001010",
  18065=>"001101010",
  18066=>"010001010",
  18067=>"000110101",
  18068=>"100010001",
  18069=>"000001000",
  18070=>"011110000",
  18071=>"000101000",
  18072=>"111110111",
  18073=>"100011101",
  18074=>"010010010",
  18075=>"110010101",
  18076=>"001000101",
  18077=>"100111110",
  18078=>"111011101",
  18079=>"111110011",
  18080=>"110010100",
  18081=>"001011100",
  18082=>"011010000",
  18083=>"010001010",
  18084=>"101101001",
  18085=>"001001000",
  18086=>"000101010",
  18087=>"111000000",
  18088=>"110110101",
  18089=>"001110101",
  18090=>"111111110",
  18091=>"010111101",
  18092=>"100001000",
  18093=>"101010001",
  18094=>"101100110",
  18095=>"110011100",
  18096=>"010110010",
  18097=>"101111000",
  18098=>"100111110",
  18099=>"111111101",
  18100=>"011001011",
  18101=>"001110101",
  18102=>"101010110",
  18103=>"011000001",
  18104=>"011111100",
  18105=>"111111110",
  18106=>"110000110",
  18107=>"001110000",
  18108=>"001100010",
  18109=>"100001100",
  18110=>"000100011",
  18111=>"000110100",
  18112=>"010001111",
  18113=>"000010101",
  18114=>"011101100",
  18115=>"011110101",
  18116=>"101111100",
  18117=>"011011110",
  18118=>"110110110",
  18119=>"110101010",
  18120=>"100111011",
  18121=>"010011001",
  18122=>"110110100",
  18123=>"011110111",
  18124=>"101111010",
  18125=>"111100011",
  18126=>"010101010",
  18127=>"110111100",
  18128=>"010111001",
  18129=>"001111001",
  18130=>"111001000",
  18131=>"111011010",
  18132=>"110110111",
  18133=>"001000001",
  18134=>"111011110",
  18135=>"111110001",
  18136=>"100000011",
  18137=>"110110111",
  18138=>"010110000",
  18139=>"011100011",
  18140=>"111010111",
  18141=>"111010111",
  18142=>"110011111",
  18143=>"000110000",
  18144=>"011100111",
  18145=>"100101101",
  18146=>"101101000",
  18147=>"000110001",
  18148=>"100001111",
  18149=>"010000101",
  18150=>"001100001",
  18151=>"110011111",
  18152=>"011000001",
  18153=>"101010101",
  18154=>"011101110",
  18155=>"000111011",
  18156=>"010000000",
  18157=>"001100101",
  18158=>"110111000",
  18159=>"000010100",
  18160=>"000001101",
  18161=>"110000101",
  18162=>"011100010",
  18163=>"010110100",
  18164=>"011100011",
  18165=>"110000000",
  18166=>"000110010",
  18167=>"010110100",
  18168=>"110100000",
  18169=>"001011111",
  18170=>"010000100",
  18171=>"011001001",
  18172=>"110111111",
  18173=>"011110100",
  18174=>"110101111",
  18175=>"011110111",
  18176=>"001100010",
  18177=>"010110010",
  18178=>"001111101",
  18179=>"010010011",
  18180=>"110000101",
  18181=>"101000001",
  18182=>"001000110",
  18183=>"101101101",
  18184=>"100110000",
  18185=>"100010101",
  18186=>"110111101",
  18187=>"000010010",
  18188=>"000011111",
  18189=>"110001001",
  18190=>"101111101",
  18191=>"111011001",
  18192=>"111100101",
  18193=>"000000000",
  18194=>"010010110",
  18195=>"100010010",
  18196=>"011000000",
  18197=>"111111011",
  18198=>"011001011",
  18199=>"010101000",
  18200=>"011010010",
  18201=>"110100010",
  18202=>"100000001",
  18203=>"010101001",
  18204=>"100101010",
  18205=>"001110111",
  18206=>"111011101",
  18207=>"000111011",
  18208=>"101111111",
  18209=>"010000100",
  18210=>"110001000",
  18211=>"100100001",
  18212=>"100000100",
  18213=>"111110010",
  18214=>"111001000",
  18215=>"000000110",
  18216=>"011010101",
  18217=>"100001110",
  18218=>"100100101",
  18219=>"000001001",
  18220=>"010101110",
  18221=>"001000000",
  18222=>"111001010",
  18223=>"100100001",
  18224=>"011010001",
  18225=>"001100101",
  18226=>"000000101",
  18227=>"000100110",
  18228=>"110000011",
  18229=>"101000111",
  18230=>"011011111",
  18231=>"000110100",
  18232=>"001111101",
  18233=>"000100111",
  18234=>"011101011",
  18235=>"011110110",
  18236=>"000100101",
  18237=>"001110000",
  18238=>"011001111",
  18239=>"010011110",
  18240=>"001000101",
  18241=>"101011011",
  18242=>"111011000",
  18243=>"001110011",
  18244=>"110010011",
  18245=>"101110110",
  18246=>"000111100",
  18247=>"110100011",
  18248=>"111111011",
  18249=>"101101110",
  18250=>"100100001",
  18251=>"011001000",
  18252=>"001111001",
  18253=>"001111011",
  18254=>"110111110",
  18255=>"010011110",
  18256=>"001110101",
  18257=>"000010111",
  18258=>"001001001",
  18259=>"001001010",
  18260=>"011000000",
  18261=>"111010000",
  18262=>"011000101",
  18263=>"110111010",
  18264=>"000011000",
  18265=>"110100100",
  18266=>"100011011",
  18267=>"100000000",
  18268=>"111010101",
  18269=>"000001000",
  18270=>"000000100",
  18271=>"110100001",
  18272=>"100001100",
  18273=>"110111011",
  18274=>"001110101",
  18275=>"010011011",
  18276=>"010001001",
  18277=>"100111010",
  18278=>"101001100",
  18279=>"011110111",
  18280=>"101100110",
  18281=>"101010001",
  18282=>"000101101",
  18283=>"100111101",
  18284=>"100011101",
  18285=>"001110111",
  18286=>"101011110",
  18287=>"001001101",
  18288=>"001101110",
  18289=>"110000100",
  18290=>"111101100",
  18291=>"010110111",
  18292=>"010011010",
  18293=>"011000000",
  18294=>"011001001",
  18295=>"110000001",
  18296=>"001010000",
  18297=>"101111111",
  18298=>"001110001",
  18299=>"011110000",
  18300=>"110111001",
  18301=>"111011111",
  18302=>"011110100",
  18303=>"011010011",
  18304=>"101100001",
  18305=>"100001010",
  18306=>"011010110",
  18307=>"000110111",
  18308=>"010000010",
  18309=>"010101101",
  18310=>"000010000",
  18311=>"001001001",
  18312=>"011010100",
  18313=>"111010100",
  18314=>"110110111",
  18315=>"011000110",
  18316=>"001010000",
  18317=>"011100001",
  18318=>"001101101",
  18319=>"001101011",
  18320=>"111011110",
  18321=>"001011111",
  18322=>"110110001",
  18323=>"000101100",
  18324=>"101000100",
  18325=>"001001110",
  18326=>"001100000",
  18327=>"100011100",
  18328=>"010001011",
  18329=>"001100010",
  18330=>"101111011",
  18331=>"010010111",
  18332=>"010000101",
  18333=>"011111011",
  18334=>"001100010",
  18335=>"100001110",
  18336=>"101111001",
  18337=>"010100011",
  18338=>"101000010",
  18339=>"000000111",
  18340=>"100000011",
  18341=>"101101110",
  18342=>"111111000",
  18343=>"011011100",
  18344=>"001100011",
  18345=>"000011000",
  18346=>"111010100",
  18347=>"100000100",
  18348=>"010110010",
  18349=>"110010110",
  18350=>"010011010",
  18351=>"111000101",
  18352=>"001011101",
  18353=>"111001101",
  18354=>"010100010",
  18355=>"110110000",
  18356=>"010011101",
  18357=>"111001111",
  18358=>"101000010",
  18359=>"101011101",
  18360=>"001111111",
  18361=>"001010011",
  18362=>"000101101",
  18363=>"101001001",
  18364=>"110101000",
  18365=>"100010111",
  18366=>"101101100",
  18367=>"000000110",
  18368=>"001010000",
  18369=>"000111001",
  18370=>"011111111",
  18371=>"110111111",
  18372=>"111101100",
  18373=>"011011001",
  18374=>"010010001",
  18375=>"101000111",
  18376=>"010101101",
  18377=>"000010101",
  18378=>"011100110",
  18379=>"110101110",
  18380=>"010101111",
  18381=>"000111101",
  18382=>"000110110",
  18383=>"100001110",
  18384=>"011010010",
  18385=>"011100111",
  18386=>"110011011",
  18387=>"000010001",
  18388=>"111110111",
  18389=>"111111011",
  18390=>"100001110",
  18391=>"111011011",
  18392=>"000111010",
  18393=>"111101110",
  18394=>"000001000",
  18395=>"100100000",
  18396=>"001000011",
  18397=>"000110101",
  18398=>"001011010",
  18399=>"000000101",
  18400=>"000111100",
  18401=>"110101001",
  18402=>"101111011",
  18403=>"110101110",
  18404=>"111000100",
  18405=>"000001111",
  18406=>"101010000",
  18407=>"100010011",
  18408=>"001001110",
  18409=>"111000110",
  18410=>"111011111",
  18411=>"101010101",
  18412=>"110011110",
  18413=>"000000001",
  18414=>"001011111",
  18415=>"011111110",
  18416=>"011011000",
  18417=>"011001100",
  18418=>"110100111",
  18419=>"001001011",
  18420=>"111000101",
  18421=>"001101111",
  18422=>"111100110",
  18423=>"110110011",
  18424=>"101000010",
  18425=>"010100100",
  18426=>"001110000",
  18427=>"101010000",
  18428=>"000000000",
  18429=>"111100100",
  18430=>"010001111",
  18431=>"111000100",
  18432=>"111111011",
  18433=>"101100011",
  18434=>"110011110",
  18435=>"110010001",
  18436=>"110011101",
  18437=>"111000011",
  18438=>"001000110",
  18439=>"111100011",
  18440=>"100101011",
  18441=>"100001110",
  18442=>"001101000",
  18443=>"101100110",
  18444=>"101011000",
  18445=>"111000100",
  18446=>"100101111",
  18447=>"111011111",
  18448=>"101101100",
  18449=>"110110001",
  18450=>"000000101",
  18451=>"100011011",
  18452=>"101111110",
  18453=>"001001110",
  18454=>"100010100",
  18455=>"001010111",
  18456=>"001110011",
  18457=>"000000100",
  18458=>"001011011",
  18459=>"000010100",
  18460=>"110001111",
  18461=>"110011010",
  18462=>"011110101",
  18463=>"010110001",
  18464=>"110110011",
  18465=>"100100010",
  18466=>"010010010",
  18467=>"010010101",
  18468=>"101011111",
  18469=>"001000110",
  18470=>"001011110",
  18471=>"101111011",
  18472=>"110110001",
  18473=>"010011110",
  18474=>"011001110",
  18475=>"101010111",
  18476=>"110101001",
  18477=>"101000111",
  18478=>"110001111",
  18479=>"000001001",
  18480=>"001101101",
  18481=>"100011100",
  18482=>"100011011",
  18483=>"111110010",
  18484=>"101101001",
  18485=>"010000001",
  18486=>"100100101",
  18487=>"110011101",
  18488=>"101000010",
  18489=>"101100011",
  18490=>"010001010",
  18491=>"001011100",
  18492=>"001001011",
  18493=>"011010011",
  18494=>"000111001",
  18495=>"000000011",
  18496=>"101110110",
  18497=>"100001001",
  18498=>"001110110",
  18499=>"010010111",
  18500=>"100101010",
  18501=>"110011010",
  18502=>"010100100",
  18503=>"111001101",
  18504=>"010100110",
  18505=>"011100011",
  18506=>"001000101",
  18507=>"100001100",
  18508=>"010000000",
  18509=>"100011111",
  18510=>"010000011",
  18511=>"010110100",
  18512=>"011100111",
  18513=>"011110111",
  18514=>"001110010",
  18515=>"001010000",
  18516=>"011010010",
  18517=>"011010111",
  18518=>"010011110",
  18519=>"110000000",
  18520=>"110101101",
  18521=>"101101011",
  18522=>"000101000",
  18523=>"000001110",
  18524=>"011010100",
  18525=>"010111011",
  18526=>"110001010",
  18527=>"000011011",
  18528=>"010101101",
  18529=>"101000110",
  18530=>"010100010",
  18531=>"000011100",
  18532=>"000010000",
  18533=>"111011000",
  18534=>"110011000",
  18535=>"010001001",
  18536=>"101001000",
  18537=>"011010111",
  18538=>"010011100",
  18539=>"001001100",
  18540=>"111110110",
  18541=>"100101001",
  18542=>"001010011",
  18543=>"011000000",
  18544=>"111010011",
  18545=>"010010100",
  18546=>"000101110",
  18547=>"000110010",
  18548=>"101001001",
  18549=>"100011010",
  18550=>"111000011",
  18551=>"111110110",
  18552=>"101000001",
  18553=>"000000000",
  18554=>"011011010",
  18555=>"000101001",
  18556=>"010010101",
  18557=>"101111011",
  18558=>"010010000",
  18559=>"011101101",
  18560=>"001110111",
  18561=>"101000000",
  18562=>"111001001",
  18563=>"000000000",
  18564=>"000000100",
  18565=>"111011111",
  18566=>"111001100",
  18567=>"000101100",
  18568=>"001000100",
  18569=>"001011101",
  18570=>"111101000",
  18571=>"001001101",
  18572=>"000111011",
  18573=>"111001100",
  18574=>"100110010",
  18575=>"011011100",
  18576=>"000111101",
  18577=>"110110001",
  18578=>"111000101",
  18579=>"110000000",
  18580=>"000010011",
  18581=>"010001001",
  18582=>"000000000",
  18583=>"111111011",
  18584=>"110100101",
  18585=>"010010010",
  18586=>"101110111",
  18587=>"111000111",
  18588=>"100010000",
  18589=>"110000101",
  18590=>"010100000",
  18591=>"110011011",
  18592=>"111011011",
  18593=>"101100101",
  18594=>"010000110",
  18595=>"100100111",
  18596=>"000111100",
  18597=>"000100111",
  18598=>"011110100",
  18599=>"010010111",
  18600=>"010010110",
  18601=>"110011000",
  18602=>"000110111",
  18603=>"100100110",
  18604=>"011101110",
  18605=>"101001000",
  18606=>"011010010",
  18607=>"010101010",
  18608=>"111100000",
  18609=>"111001100",
  18610=>"110000110",
  18611=>"011011000",
  18612=>"010110010",
  18613=>"111011101",
  18614=>"110100101",
  18615=>"010000111",
  18616=>"001100110",
  18617=>"000101000",
  18618=>"010100010",
  18619=>"010010101",
  18620=>"110101111",
  18621=>"100100001",
  18622=>"000111101",
  18623=>"000111100",
  18624=>"100100100",
  18625=>"100011111",
  18626=>"000000000",
  18627=>"011001000",
  18628=>"010111010",
  18629=>"010000001",
  18630=>"101011110",
  18631=>"100110001",
  18632=>"111010010",
  18633=>"010011001",
  18634=>"110011010",
  18635=>"011010111",
  18636=>"101110000",
  18637=>"000100010",
  18638=>"101001010",
  18639=>"000000100",
  18640=>"000110001",
  18641=>"010110111",
  18642=>"010101100",
  18643=>"000011000",
  18644=>"101110101",
  18645=>"010000110",
  18646=>"111111100",
  18647=>"011111001",
  18648=>"100010110",
  18649=>"111000100",
  18650=>"101111110",
  18651=>"010001110",
  18652=>"100100001",
  18653=>"101010011",
  18654=>"111100010",
  18655=>"100010000",
  18656=>"011010101",
  18657=>"001010100",
  18658=>"100100111",
  18659=>"100010111",
  18660=>"111110101",
  18661=>"010110111",
  18662=>"100110001",
  18663=>"011110111",
  18664=>"110110111",
  18665=>"001101101",
  18666=>"101101101",
  18667=>"000101111",
  18668=>"010110001",
  18669=>"011011010",
  18670=>"101001110",
  18671=>"111000111",
  18672=>"101101111",
  18673=>"111110001",
  18674=>"011010010",
  18675=>"010011000",
  18676=>"111101110",
  18677=>"101011100",
  18678=>"000000111",
  18679=>"010011011",
  18680=>"101010110",
  18681=>"000010001",
  18682=>"001101010",
  18683=>"100110001",
  18684=>"101000011",
  18685=>"101000000",
  18686=>"110100010",
  18687=>"000000111",
  18688=>"110101111",
  18689=>"110001001",
  18690=>"001100111",
  18691=>"100000110",
  18692=>"011100001",
  18693=>"001000101",
  18694=>"000110111",
  18695=>"100001001",
  18696=>"000010000",
  18697=>"000101110",
  18698=>"110011101",
  18699=>"101010110",
  18700=>"110111011",
  18701=>"111011101",
  18702=>"111101110",
  18703=>"100101001",
  18704=>"100101011",
  18705=>"001101011",
  18706=>"100001001",
  18707=>"001100001",
  18708=>"000101101",
  18709=>"001110000",
  18710=>"100101000",
  18711=>"100001100",
  18712=>"010000110",
  18713=>"001111010",
  18714=>"100010001",
  18715=>"011010100",
  18716=>"000101011",
  18717=>"010010011",
  18718=>"101000110",
  18719=>"000100001",
  18720=>"101000010",
  18721=>"101011000",
  18722=>"111101010",
  18723=>"100101010",
  18724=>"110110011",
  18725=>"000111010",
  18726=>"100010000",
  18727=>"001111100",
  18728=>"110100111",
  18729=>"111111110",
  18730=>"101010000",
  18731=>"111010001",
  18732=>"100110000",
  18733=>"100001000",
  18734=>"111101010",
  18735=>"011001101",
  18736=>"101000010",
  18737=>"111010100",
  18738=>"001111110",
  18739=>"000000001",
  18740=>"000010101",
  18741=>"111011000",
  18742=>"100111011",
  18743=>"111010100",
  18744=>"110000001",
  18745=>"011100101",
  18746=>"000000100",
  18747=>"110111000",
  18748=>"011110111",
  18749=>"001010110",
  18750=>"110100100",
  18751=>"001000000",
  18752=>"101010101",
  18753=>"111000001",
  18754=>"110000111",
  18755=>"001010010",
  18756=>"000001100",
  18757=>"110110110",
  18758=>"010110111",
  18759=>"010001101",
  18760=>"110111000",
  18761=>"000101000",
  18762=>"010010000",
  18763=>"000010011",
  18764=>"000110100",
  18765=>"011111111",
  18766=>"101111011",
  18767=>"010000011",
  18768=>"100000100",
  18769=>"010100101",
  18770=>"100010111",
  18771=>"110100100",
  18772=>"100101100",
  18773=>"010101010",
  18774=>"111011111",
  18775=>"000000111",
  18776=>"011001111",
  18777=>"000100110",
  18778=>"001000110",
  18779=>"000110100",
  18780=>"000011001",
  18781=>"110100111",
  18782=>"100001010",
  18783=>"001111010",
  18784=>"101010111",
  18785=>"100101001",
  18786=>"110000101",
  18787=>"000111001",
  18788=>"111111011",
  18789=>"100001101",
  18790=>"101111001",
  18791=>"110011101",
  18792=>"100100101",
  18793=>"001000011",
  18794=>"010110001",
  18795=>"100011101",
  18796=>"101110010",
  18797=>"000000101",
  18798=>"100100110",
  18799=>"001000011",
  18800=>"000011101",
  18801=>"110010101",
  18802=>"000111011",
  18803=>"011001111",
  18804=>"001001010",
  18805=>"000101010",
  18806=>"100110010",
  18807=>"000101111",
  18808=>"000101001",
  18809=>"001010101",
  18810=>"111011010",
  18811=>"010101011",
  18812=>"101101111",
  18813=>"100101011",
  18814=>"001100101",
  18815=>"001001010",
  18816=>"001100111",
  18817=>"000000110",
  18818=>"011001101",
  18819=>"000101100",
  18820=>"000110111",
  18821=>"011000001",
  18822=>"101110011",
  18823=>"001001000",
  18824=>"100100111",
  18825=>"010010001",
  18826=>"010111101",
  18827=>"110010110",
  18828=>"011101000",
  18829=>"011000001",
  18830=>"110101110",
  18831=>"101011101",
  18832=>"110010110",
  18833=>"100110101",
  18834=>"101100101",
  18835=>"000111010",
  18836=>"000100100",
  18837=>"001111111",
  18838=>"101011111",
  18839=>"010111100",
  18840=>"001001100",
  18841=>"010000011",
  18842=>"000011101",
  18843=>"000111010",
  18844=>"110000010",
  18845=>"101010110",
  18846=>"101011100",
  18847=>"110110010",
  18848=>"100100111",
  18849=>"000011100",
  18850=>"001011010",
  18851=>"110101101",
  18852=>"010111011",
  18853=>"010001000",
  18854=>"110001010",
  18855=>"110011111",
  18856=>"100000010",
  18857=>"000100100",
  18858=>"000100110",
  18859=>"111001011",
  18860=>"101101001",
  18861=>"000111001",
  18862=>"011000011",
  18863=>"101111101",
  18864=>"001011111",
  18865=>"011101010",
  18866=>"111111010",
  18867=>"000111000",
  18868=>"010111111",
  18869=>"011110000",
  18870=>"101000100",
  18871=>"011100100",
  18872=>"110101010",
  18873=>"010111010",
  18874=>"111110010",
  18875=>"010100110",
  18876=>"111101000",
  18877=>"001100010",
  18878=>"011100010",
  18879=>"010110001",
  18880=>"011100010",
  18881=>"011001000",
  18882=>"111001110",
  18883=>"101101101",
  18884=>"110000011",
  18885=>"001010010",
  18886=>"100000100",
  18887=>"111010100",
  18888=>"101100001",
  18889=>"001100101",
  18890=>"000110001",
  18891=>"010010001",
  18892=>"010011001",
  18893=>"110001000",
  18894=>"101100101",
  18895=>"110101111",
  18896=>"110010111",
  18897=>"010100010",
  18898=>"101001000",
  18899=>"001101110",
  18900=>"010001011",
  18901=>"001110101",
  18902=>"011001010",
  18903=>"110110100",
  18904=>"110000010",
  18905=>"011000111",
  18906=>"110010110",
  18907=>"110101010",
  18908=>"011101101",
  18909=>"000100000",
  18910=>"001010110",
  18911=>"011101101",
  18912=>"011111010",
  18913=>"110101110",
  18914=>"100010001",
  18915=>"111100000",
  18916=>"000001100",
  18917=>"011111100",
  18918=>"001000011",
  18919=>"101010010",
  18920=>"011110000",
  18921=>"100000110",
  18922=>"100010101",
  18923=>"100001111",
  18924=>"110110111",
  18925=>"010101000",
  18926=>"000101000",
  18927=>"010110011",
  18928=>"010010110",
  18929=>"011101001",
  18930=>"110011011",
  18931=>"010001101",
  18932=>"111001110",
  18933=>"010011010",
  18934=>"000010011",
  18935=>"001001100",
  18936=>"111101011",
  18937=>"011111111",
  18938=>"010101101",
  18939=>"101111111",
  18940=>"000001111",
  18941=>"110011001",
  18942=>"110010010",
  18943=>"110110010",
  18944=>"111111101",
  18945=>"110100100",
  18946=>"010101100",
  18947=>"100000011",
  18948=>"111000001",
  18949=>"000101110",
  18950=>"010101111",
  18951=>"111010111",
  18952=>"011001000",
  18953=>"111001000",
  18954=>"101111010",
  18955=>"011101101",
  18956=>"001011010",
  18957=>"110110111",
  18958=>"000100010",
  18959=>"001110111",
  18960=>"011111111",
  18961=>"000111000",
  18962=>"111001010",
  18963=>"111101011",
  18964=>"100000100",
  18965=>"010010100",
  18966=>"000111100",
  18967=>"111000011",
  18968=>"100110001",
  18969=>"000110010",
  18970=>"000010010",
  18971=>"000011010",
  18972=>"110101110",
  18973=>"100000100",
  18974=>"101010001",
  18975=>"111000110",
  18976=>"100000010",
  18977=>"001000000",
  18978=>"011010100",
  18979=>"011010011",
  18980=>"110001011",
  18981=>"100011100",
  18982=>"100000000",
  18983=>"101011110",
  18984=>"011111101",
  18985=>"011111000",
  18986=>"101111011",
  18987=>"100101101",
  18988=>"101011000",
  18989=>"001011100",
  18990=>"010111100",
  18991=>"100000011",
  18992=>"110001100",
  18993=>"101001100",
  18994=>"001100011",
  18995=>"000000100",
  18996=>"001111000",
  18997=>"010011001",
  18998=>"000001010",
  18999=>"100011101",
  19000=>"101000100",
  19001=>"111100000",
  19002=>"111000111",
  19003=>"010000010",
  19004=>"101010111",
  19005=>"011011010",
  19006=>"001010111",
  19007=>"100010100",
  19008=>"001000010",
  19009=>"111101000",
  19010=>"110010010",
  19011=>"111001101",
  19012=>"000000010",
  19013=>"101011000",
  19014=>"101110011",
  19015=>"110000110",
  19016=>"010001011",
  19017=>"111011111",
  19018=>"011011001",
  19019=>"110010101",
  19020=>"010010111",
  19021=>"100000001",
  19022=>"111101000",
  19023=>"011000011",
  19024=>"100011100",
  19025=>"000101101",
  19026=>"000100001",
  19027=>"110000111",
  19028=>"110111001",
  19029=>"000100011",
  19030=>"001011000",
  19031=>"000011010",
  19032=>"011111110",
  19033=>"000000100",
  19034=>"111101110",
  19035=>"100001111",
  19036=>"110100001",
  19037=>"000110010",
  19038=>"111011011",
  19039=>"111100101",
  19040=>"011010100",
  19041=>"101001100",
  19042=>"101100011",
  19043=>"110001000",
  19044=>"101110111",
  19045=>"011100111",
  19046=>"000010001",
  19047=>"111000101",
  19048=>"111011011",
  19049=>"101010110",
  19050=>"111110111",
  19051=>"001000010",
  19052=>"110100111",
  19053=>"111110011",
  19054=>"100010010",
  19055=>"101111110",
  19056=>"000011110",
  19057=>"111010101",
  19058=>"101111111",
  19059=>"010101101",
  19060=>"000100011",
  19061=>"111100101",
  19062=>"111000101",
  19063=>"001110000",
  19064=>"010010001",
  19065=>"011001111",
  19066=>"110110110",
  19067=>"010000001",
  19068=>"100010101",
  19069=>"101000111",
  19070=>"000001011",
  19071=>"100111001",
  19072=>"010001100",
  19073=>"111110100",
  19074=>"110100001",
  19075=>"101001110",
  19076=>"100100010",
  19077=>"010101001",
  19078=>"000010000",
  19079=>"101010110",
  19080=>"011000001",
  19081=>"101101101",
  19082=>"101010011",
  19083=>"010110111",
  19084=>"110010001",
  19085=>"000010011",
  19086=>"001000010",
  19087=>"100100111",
  19088=>"100100000",
  19089=>"100010101",
  19090=>"101111000",
  19091=>"101101110",
  19092=>"000111110",
  19093=>"010000111",
  19094=>"100110010",
  19095=>"010100010",
  19096=>"010011111",
  19097=>"111101110",
  19098=>"001100011",
  19099=>"100101111",
  19100=>"101011000",
  19101=>"001111000",
  19102=>"001110110",
  19103=>"101010101",
  19104=>"100110000",
  19105=>"100111111",
  19106=>"110001101",
  19107=>"101110001",
  19108=>"110110000",
  19109=>"100011100",
  19110=>"000000100",
  19111=>"000010000",
  19112=>"000100111",
  19113=>"100111010",
  19114=>"100111010",
  19115=>"011110100",
  19116=>"001000111",
  19117=>"111100000",
  19118=>"011111010",
  19119=>"111100100",
  19120=>"001011110",
  19121=>"001000000",
  19122=>"000101001",
  19123=>"000000000",
  19124=>"000110001",
  19125=>"101010100",
  19126=>"000010101",
  19127=>"000011000",
  19128=>"101110101",
  19129=>"111000111",
  19130=>"001000010",
  19131=>"001101011",
  19132=>"000100100",
  19133=>"010101100",
  19134=>"000100000",
  19135=>"000000000",
  19136=>"001101001",
  19137=>"110001010",
  19138=>"000110111",
  19139=>"010100101",
  19140=>"000100101",
  19141=>"000011100",
  19142=>"001111010",
  19143=>"000111000",
  19144=>"110001000",
  19145=>"001000000",
  19146=>"001010101",
  19147=>"110101001",
  19148=>"110011001",
  19149=>"110110001",
  19150=>"000010110",
  19151=>"101000000",
  19152=>"110101111",
  19153=>"101110001",
  19154=>"011101010",
  19155=>"111110001",
  19156=>"010100000",
  19157=>"000010001",
  19158=>"001011110",
  19159=>"110011100",
  19160=>"010001110",
  19161=>"100011011",
  19162=>"100101101",
  19163=>"100100000",
  19164=>"001011100",
  19165=>"001100111",
  19166=>"110111111",
  19167=>"110001101",
  19168=>"100101101",
  19169=>"101110110",
  19170=>"101101111",
  19171=>"010100111",
  19172=>"001001111",
  19173=>"011011110",
  19174=>"011100101",
  19175=>"001111010",
  19176=>"000000100",
  19177=>"000000000",
  19178=>"100010101",
  19179=>"101011010",
  19180=>"010110011",
  19181=>"001100101",
  19182=>"011010111",
  19183=>"011000101",
  19184=>"000111101",
  19185=>"100101001",
  19186=>"110010110",
  19187=>"110111000",
  19188=>"101101111",
  19189=>"100010011",
  19190=>"010010111",
  19191=>"110010100",
  19192=>"000010011",
  19193=>"001101010",
  19194=>"011011010",
  19195=>"101010011",
  19196=>"001010000",
  19197=>"110000111",
  19198=>"110111110",
  19199=>"100110011",
  19200=>"101110001",
  19201=>"110000111",
  19202=>"001101010",
  19203=>"000011110",
  19204=>"001011010",
  19205=>"110011010",
  19206=>"011110110",
  19207=>"110000101",
  19208=>"001001001",
  19209=>"010010101",
  19210=>"000010001",
  19211=>"111100010",
  19212=>"011111100",
  19213=>"101101111",
  19214=>"001111110",
  19215=>"100000110",
  19216=>"000100011",
  19217=>"010011000",
  19218=>"100010000",
  19219=>"010001011",
  19220=>"001100000",
  19221=>"111001001",
  19222=>"111011000",
  19223=>"100110011",
  19224=>"110011100",
  19225=>"111010000",
  19226=>"000011011",
  19227=>"000010001",
  19228=>"010011001",
  19229=>"110011111",
  19230=>"010100100",
  19231=>"110110100",
  19232=>"110001110",
  19233=>"101001101",
  19234=>"110011101",
  19235=>"011011100",
  19236=>"011001010",
  19237=>"000001001",
  19238=>"001101100",
  19239=>"010000110",
  19240=>"100101001",
  19241=>"011111000",
  19242=>"111100010",
  19243=>"011100100",
  19244=>"001101111",
  19245=>"100100011",
  19246=>"100000001",
  19247=>"011100001",
  19248=>"110111111",
  19249=>"001011110",
  19250=>"000100111",
  19251=>"011101011",
  19252=>"110110110",
  19253=>"100100000",
  19254=>"100000011",
  19255=>"000100010",
  19256=>"101111111",
  19257=>"010110100",
  19258=>"110000101",
  19259=>"000011100",
  19260=>"100000011",
  19261=>"100001001",
  19262=>"001000001",
  19263=>"000110101",
  19264=>"100111111",
  19265=>"110110111",
  19266=>"110110110",
  19267=>"001101000",
  19268=>"000010011",
  19269=>"000100110",
  19270=>"011000000",
  19271=>"101001011",
  19272=>"100001011",
  19273=>"011001001",
  19274=>"010110001",
  19275=>"110000101",
  19276=>"011000010",
  19277=>"011001010",
  19278=>"111010101",
  19279=>"110000101",
  19280=>"111011011",
  19281=>"100010001",
  19282=>"101011111",
  19283=>"010110011",
  19284=>"001101011",
  19285=>"011001111",
  19286=>"001000001",
  19287=>"011010000",
  19288=>"111010011",
  19289=>"011100001",
  19290=>"111110101",
  19291=>"101101001",
  19292=>"111110011",
  19293=>"001110000",
  19294=>"100101001",
  19295=>"000101001",
  19296=>"101111011",
  19297=>"100000111",
  19298=>"101000011",
  19299=>"001000111",
  19300=>"000100010",
  19301=>"000100000",
  19302=>"110101011",
  19303=>"001011010",
  19304=>"111010010",
  19305=>"101100111",
  19306=>"000001100",
  19307=>"010000001",
  19308=>"011001011",
  19309=>"111101100",
  19310=>"101010001",
  19311=>"100001111",
  19312=>"101101010",
  19313=>"011010111",
  19314=>"001110011",
  19315=>"110100100",
  19316=>"100000011",
  19317=>"010111110",
  19318=>"111011110",
  19319=>"110011110",
  19320=>"010110010",
  19321=>"110010101",
  19322=>"111110101",
  19323=>"101000110",
  19324=>"100101000",
  19325=>"001010100",
  19326=>"000110100",
  19327=>"110101100",
  19328=>"110111010",
  19329=>"101101001",
  19330=>"011101000",
  19331=>"101010000",
  19332=>"111010111",
  19333=>"111000011",
  19334=>"011011110",
  19335=>"001001011",
  19336=>"100001111",
  19337=>"011000100",
  19338=>"100011100",
  19339=>"101111110",
  19340=>"111101001",
  19341=>"011110011",
  19342=>"111000101",
  19343=>"111110000",
  19344=>"110010001",
  19345=>"110011011",
  19346=>"000011010",
  19347=>"111011000",
  19348=>"111000101",
  19349=>"100011111",
  19350=>"000100101",
  19351=>"000011001",
  19352=>"010011110",
  19353=>"010111011",
  19354=>"001000010",
  19355=>"110100101",
  19356=>"111110010",
  19357=>"111000000",
  19358=>"010101001",
  19359=>"011000000",
  19360=>"000011000",
  19361=>"000100100",
  19362=>"001010000",
  19363=>"101111001",
  19364=>"100010001",
  19365=>"101010101",
  19366=>"001110011",
  19367=>"110010010",
  19368=>"111100110",
  19369=>"000110100",
  19370=>"100101101",
  19371=>"011010001",
  19372=>"100001100",
  19373=>"011011000",
  19374=>"010001110",
  19375=>"001010000",
  19376=>"001100011",
  19377=>"000001010",
  19378=>"011111010",
  19379=>"001111000",
  19380=>"111111100",
  19381=>"111110000",
  19382=>"100010110",
  19383=>"010011001",
  19384=>"111001110",
  19385=>"000010011",
  19386=>"111111100",
  19387=>"110100011",
  19388=>"101001111",
  19389=>"110110000",
  19390=>"110011100",
  19391=>"101000100",
  19392=>"000100011",
  19393=>"001001101",
  19394=>"111100111",
  19395=>"100001101",
  19396=>"111101110",
  19397=>"011100101",
  19398=>"100010101",
  19399=>"000001110",
  19400=>"111111010",
  19401=>"101101111",
  19402=>"010010010",
  19403=>"010001000",
  19404=>"111000100",
  19405=>"010001001",
  19406=>"111000101",
  19407=>"011110011",
  19408=>"111000001",
  19409=>"010111011",
  19410=>"100010001",
  19411=>"011110110",
  19412=>"001101100",
  19413=>"110111000",
  19414=>"101010010",
  19415=>"101000111",
  19416=>"011101100",
  19417=>"011101010",
  19418=>"101111111",
  19419=>"111001010",
  19420=>"110000100",
  19421=>"101001011",
  19422=>"011011111",
  19423=>"101111001",
  19424=>"001010000",
  19425=>"000010111",
  19426=>"010000110",
  19427=>"110001000",
  19428=>"110000000",
  19429=>"110010000",
  19430=>"110001111",
  19431=>"110010010",
  19432=>"000100000",
  19433=>"000011010",
  19434=>"001001110",
  19435=>"111011011",
  19436=>"110110100",
  19437=>"111100101",
  19438=>"000100100",
  19439=>"111000010",
  19440=>"100110100",
  19441=>"100111101",
  19442=>"001000000",
  19443=>"111110001",
  19444=>"010010101",
  19445=>"000100010",
  19446=>"111011000",
  19447=>"010000011",
  19448=>"000011011",
  19449=>"101001110",
  19450=>"010100000",
  19451=>"001010001",
  19452=>"100011010",
  19453=>"111100010",
  19454=>"001100000",
  19455=>"000001001",
  19456=>"000110011",
  19457=>"010101011",
  19458=>"110100001",
  19459=>"111000110",
  19460=>"010101000",
  19461=>"011101011",
  19462=>"110011000",
  19463=>"001001001",
  19464=>"111011111",
  19465=>"010101011",
  19466=>"111001100",
  19467=>"110001000",
  19468=>"101101101",
  19469=>"110001010",
  19470=>"101100001",
  19471=>"110001010",
  19472=>"111110101",
  19473=>"100001101",
  19474=>"010000111",
  19475=>"101101110",
  19476=>"101000000",
  19477=>"001111110",
  19478=>"011000000",
  19479=>"101000010",
  19480=>"000011000",
  19481=>"000011100",
  19482=>"100100111",
  19483=>"101010111",
  19484=>"010101110",
  19485=>"101110000",
  19486=>"000010100",
  19487=>"111101011",
  19488=>"110000010",
  19489=>"000011101",
  19490=>"011010001",
  19491=>"010010101",
  19492=>"011010100",
  19493=>"011100000",
  19494=>"101011100",
  19495=>"111010011",
  19496=>"110101111",
  19497=>"100101101",
  19498=>"010110100",
  19499=>"000011011",
  19500=>"001000000",
  19501=>"110101000",
  19502=>"000000110",
  19503=>"000000000",
  19504=>"011111001",
  19505=>"101110111",
  19506=>"011100111",
  19507=>"011110010",
  19508=>"100010001",
  19509=>"000110010",
  19510=>"011110110",
  19511=>"010111111",
  19512=>"111000110",
  19513=>"000001101",
  19514=>"000000111",
  19515=>"000100001",
  19516=>"101001010",
  19517=>"011011111",
  19518=>"000001010",
  19519=>"001100100",
  19520=>"110100000",
  19521=>"000010101",
  19522=>"100101001",
  19523=>"000110101",
  19524=>"010101100",
  19525=>"011101110",
  19526=>"000100001",
  19527=>"000000000",
  19528=>"101000101",
  19529=>"111111110",
  19530=>"011001000",
  19531=>"011111011",
  19532=>"100011100",
  19533=>"111010100",
  19534=>"101110001",
  19535=>"011101011",
  19536=>"111100010",
  19537=>"100101000",
  19538=>"111111011",
  19539=>"111000100",
  19540=>"000111011",
  19541=>"111011000",
  19542=>"010101010",
  19543=>"000011000",
  19544=>"000101110",
  19545=>"001101000",
  19546=>"111110001",
  19547=>"101000000",
  19548=>"010101000",
  19549=>"001010110",
  19550=>"100111010",
  19551=>"100011001",
  19552=>"011011111",
  19553=>"011011100",
  19554=>"000001000",
  19555=>"110010011",
  19556=>"001011100",
  19557=>"000111010",
  19558=>"010110000",
  19559=>"001010110",
  19560=>"101111011",
  19561=>"011010110",
  19562=>"110001000",
  19563=>"001110000",
  19564=>"011101000",
  19565=>"111110010",
  19566=>"111001011",
  19567=>"000010000",
  19568=>"100100001",
  19569=>"001101100",
  19570=>"001010100",
  19571=>"100011100",
  19572=>"110100101",
  19573=>"110111110",
  19574=>"000000111",
  19575=>"100100100",
  19576=>"001111000",
  19577=>"110101010",
  19578=>"101100110",
  19579=>"111010111",
  19580=>"110111110",
  19581=>"111101110",
  19582=>"011111110",
  19583=>"100100001",
  19584=>"000010110",
  19585=>"110111100",
  19586=>"010101101",
  19587=>"111011000",
  19588=>"000101000",
  19589=>"010100111",
  19590=>"001000110",
  19591=>"100110100",
  19592=>"111110111",
  19593=>"101001000",
  19594=>"000000010",
  19595=>"111011100",
  19596=>"101111100",
  19597=>"101111100",
  19598=>"111000011",
  19599=>"100010111",
  19600=>"111101001",
  19601=>"001101000",
  19602=>"111011111",
  19603=>"111101100",
  19604=>"100000001",
  19605=>"110010101",
  19606=>"111101100",
  19607=>"001011100",
  19608=>"111010111",
  19609=>"111111100",
  19610=>"000010100",
  19611=>"001110110",
  19612=>"000100101",
  19613=>"011100011",
  19614=>"001110001",
  19615=>"111010001",
  19616=>"001011011",
  19617=>"010100110",
  19618=>"101100001",
  19619=>"000001101",
  19620=>"100000000",
  19621=>"111111111",
  19622=>"101100000",
  19623=>"101010111",
  19624=>"101010010",
  19625=>"000101011",
  19626=>"010110111",
  19627=>"111100111",
  19628=>"110011011",
  19629=>"000000001",
  19630=>"101100111",
  19631=>"110011111",
  19632=>"001011110",
  19633=>"100111000",
  19634=>"110100110",
  19635=>"110100001",
  19636=>"111001111",
  19637=>"000101110",
  19638=>"100001110",
  19639=>"010011110",
  19640=>"100110101",
  19641=>"101001010",
  19642=>"001001111",
  19643=>"111100111",
  19644=>"010101001",
  19645=>"011000011",
  19646=>"000111111",
  19647=>"001010001",
  19648=>"100100111",
  19649=>"100001100",
  19650=>"001010111",
  19651=>"001001111",
  19652=>"101001000",
  19653=>"011111101",
  19654=>"110101110",
  19655=>"000001101",
  19656=>"110001111",
  19657=>"101011010",
  19658=>"100010000",
  19659=>"101001001",
  19660=>"110101111",
  19661=>"010111101",
  19662=>"101010110",
  19663=>"001110001",
  19664=>"110100110",
  19665=>"001101100",
  19666=>"000001100",
  19667=>"011101011",
  19668=>"001011110",
  19669=>"001100111",
  19670=>"001101001",
  19671=>"001110001",
  19672=>"000111100",
  19673=>"101000001",
  19674=>"110111110",
  19675=>"100000100",
  19676=>"111111000",
  19677=>"100101001",
  19678=>"110110101",
  19679=>"110000101",
  19680=>"010110101",
  19681=>"110000000",
  19682=>"011001000",
  19683=>"101110101",
  19684=>"011000010",
  19685=>"101010011",
  19686=>"100000010",
  19687=>"111110000",
  19688=>"100001100",
  19689=>"000101011",
  19690=>"001110010",
  19691=>"000111111",
  19692=>"110011011",
  19693=>"000011101",
  19694=>"010000001",
  19695=>"001010010",
  19696=>"100110010",
  19697=>"100110110",
  19698=>"001001111",
  19699=>"010100000",
  19700=>"101100011",
  19701=>"101101000",
  19702=>"011110111",
  19703=>"001010010",
  19704=>"111100011",
  19705=>"000101101",
  19706=>"010001010",
  19707=>"011001011",
  19708=>"000101100",
  19709=>"110010000",
  19710=>"001101110",
  19711=>"010100011",
  19712=>"001001000",
  19713=>"110100111",
  19714=>"101010000",
  19715=>"000001100",
  19716=>"011001100",
  19717=>"001000100",
  19718=>"011110100",
  19719=>"010000011",
  19720=>"010011100",
  19721=>"001000100",
  19722=>"000011010",
  19723=>"101100100",
  19724=>"101101011",
  19725=>"000110101",
  19726=>"111101110",
  19727=>"110000100",
  19728=>"000010010",
  19729=>"101100111",
  19730=>"011000000",
  19731=>"100001011",
  19732=>"100011111",
  19733=>"111101010",
  19734=>"001011110",
  19735=>"100011110",
  19736=>"010110000",
  19737=>"001001001",
  19738=>"010111111",
  19739=>"001100111",
  19740=>"101000011",
  19741=>"011101000",
  19742=>"110000111",
  19743=>"110010001",
  19744=>"001000111",
  19745=>"001111101",
  19746=>"101111000",
  19747=>"110000101",
  19748=>"011111101",
  19749=>"110110000",
  19750=>"101000111",
  19751=>"011111101",
  19752=>"000010001",
  19753=>"100101111",
  19754=>"101100001",
  19755=>"010000000",
  19756=>"111100101",
  19757=>"110111001",
  19758=>"000011001",
  19759=>"100111100",
  19760=>"100000111",
  19761=>"000000010",
  19762=>"011111101",
  19763=>"010000110",
  19764=>"100111100",
  19765=>"000110001",
  19766=>"001111100",
  19767=>"001011010",
  19768=>"001010111",
  19769=>"010100100",
  19770=>"100111111",
  19771=>"000000010",
  19772=>"010011011",
  19773=>"100111110",
  19774=>"001100101",
  19775=>"111011001",
  19776=>"100110000",
  19777=>"101100100",
  19778=>"000111111",
  19779=>"011100101",
  19780=>"000101100",
  19781=>"000101100",
  19782=>"111001010",
  19783=>"000001011",
  19784=>"100010111",
  19785=>"000000011",
  19786=>"011001000",
  19787=>"010101000",
  19788=>"010100111",
  19789=>"010110010",
  19790=>"001100001",
  19791=>"000110011",
  19792=>"000111010",
  19793=>"100011101",
  19794=>"011010000",
  19795=>"001110111",
  19796=>"010100000",
  19797=>"000000010",
  19798=>"001100010",
  19799=>"110010111",
  19800=>"011001110",
  19801=>"010000011",
  19802=>"101110000",
  19803=>"111001000",
  19804=>"101011000",
  19805=>"110000110",
  19806=>"001011011",
  19807=>"110110100",
  19808=>"010101111",
  19809=>"111011100",
  19810=>"001111100",
  19811=>"001010101",
  19812=>"001100110",
  19813=>"100000100",
  19814=>"101000011",
  19815=>"100101000",
  19816=>"010011010",
  19817=>"100010011",
  19818=>"001011010",
  19819=>"011011100",
  19820=>"010011110",
  19821=>"010100110",
  19822=>"001101101",
  19823=>"001101011",
  19824=>"110010001",
  19825=>"001111110",
  19826=>"100010001",
  19827=>"011110001",
  19828=>"110011100",
  19829=>"111111101",
  19830=>"000011111",
  19831=>"110100110",
  19832=>"100001111",
  19833=>"110011101",
  19834=>"110011110",
  19835=>"101000000",
  19836=>"001100010",
  19837=>"000110100",
  19838=>"110010010",
  19839=>"001100100",
  19840=>"101011101",
  19841=>"001010100",
  19842=>"101010100",
  19843=>"100101100",
  19844=>"101001000",
  19845=>"110101111",
  19846=>"110111111",
  19847=>"101011001",
  19848=>"000110011",
  19849=>"011110001",
  19850=>"111010100",
  19851=>"110101011",
  19852=>"000000011",
  19853=>"000010011",
  19854=>"110010110",
  19855=>"011101010",
  19856=>"010010001",
  19857=>"011001111",
  19858=>"101100101",
  19859=>"110111001",
  19860=>"011000011",
  19861=>"101000101",
  19862=>"011010110",
  19863=>"111111001",
  19864=>"101110110",
  19865=>"110000111",
  19866=>"000011111",
  19867=>"011011101",
  19868=>"111011010",
  19869=>"001110000",
  19870=>"111000101",
  19871=>"100000001",
  19872=>"010011011",
  19873=>"011000111",
  19874=>"010000001",
  19875=>"001000110",
  19876=>"111011100",
  19877=>"000001110",
  19878=>"010101110",
  19879=>"011000101",
  19880=>"000010001",
  19881=>"000100001",
  19882=>"101100001",
  19883=>"010001111",
  19884=>"100010110",
  19885=>"011101101",
  19886=>"011101110",
  19887=>"101000010",
  19888=>"010111010",
  19889=>"000110100",
  19890=>"101100101",
  19891=>"010000110",
  19892=>"111110011",
  19893=>"010001011",
  19894=>"111011101",
  19895=>"101110101",
  19896=>"101100110",
  19897=>"000011011",
  19898=>"100101000",
  19899=>"111101000",
  19900=>"000110111",
  19901=>"101100000",
  19902=>"010010100",
  19903=>"111001010",
  19904=>"011011011",
  19905=>"011011100",
  19906=>"101010010",
  19907=>"100011110",
  19908=>"010001111",
  19909=>"010100011",
  19910=>"001111110",
  19911=>"100010010",
  19912=>"010101110",
  19913=>"000110101",
  19914=>"111011111",
  19915=>"011100111",
  19916=>"111111110",
  19917=>"010000110",
  19918=>"011001011",
  19919=>"011101000",
  19920=>"000100001",
  19921=>"001111011",
  19922=>"001000001",
  19923=>"110000111",
  19924=>"011100110",
  19925=>"001110011",
  19926=>"110011001",
  19927=>"000000011",
  19928=>"000001000",
  19929=>"101011101",
  19930=>"001001100",
  19931=>"001010101",
  19932=>"001000010",
  19933=>"000011011",
  19934=>"001000100",
  19935=>"011101110",
  19936=>"001011111",
  19937=>"010011010",
  19938=>"000000100",
  19939=>"110010101",
  19940=>"100001101",
  19941=>"100011111",
  19942=>"001101101",
  19943=>"000100011",
  19944=>"010101011",
  19945=>"100111101",
  19946=>"100101100",
  19947=>"001100111",
  19948=>"101001011",
  19949=>"101001100",
  19950=>"000000000",
  19951=>"100110011",
  19952=>"011010011",
  19953=>"111101000",
  19954=>"010110000",
  19955=>"001101110",
  19956=>"010110110",
  19957=>"111100111",
  19958=>"100111000",
  19959=>"000100010",
  19960=>"000000100",
  19961=>"110100011",
  19962=>"100010100",
  19963=>"100001000",
  19964=>"000111010",
  19965=>"111111111",
  19966=>"100000111",
  19967=>"110100010",
  19968=>"011001010",
  19969=>"101011110",
  19970=>"101010001",
  19971=>"111100111",
  19972=>"010011010",
  19973=>"000110000",
  19974=>"110110010",
  19975=>"100100101",
  19976=>"000100110",
  19977=>"001101111",
  19978=>"100110101",
  19979=>"100000100",
  19980=>"010101011",
  19981=>"011111110",
  19982=>"001111111",
  19983=>"001010010",
  19984=>"010101011",
  19985=>"100000100",
  19986=>"101010111",
  19987=>"011110011",
  19988=>"000100100",
  19989=>"101001101",
  19990=>"111111010",
  19991=>"111010010",
  19992=>"001000101",
  19993=>"111011110",
  19994=>"001011001",
  19995=>"111111110",
  19996=>"100010010",
  19997=>"011111101",
  19998=>"101101010",
  19999=>"100100010",
  20000=>"010101001",
  20001=>"000001011",
  20002=>"000001000",
  20003=>"011001110",
  20004=>"101010100",
  20005=>"001101000",
  20006=>"001110101",
  20007=>"010111011",
  20008=>"001010010",
  20009=>"001011001",
  20010=>"011001110",
  20011=>"100011000",
  20012=>"110010111",
  20013=>"111001001",
  20014=>"101010111",
  20015=>"001110111",
  20016=>"111011001",
  20017=>"100100111",
  20018=>"111001011",
  20019=>"010111101",
  20020=>"001100000",
  20021=>"001011101",
  20022=>"101000101",
  20023=>"110010011",
  20024=>"001001111",
  20025=>"011110001",
  20026=>"110110110",
  20027=>"001110111",
  20028=>"111111010",
  20029=>"000000001",
  20030=>"001101100",
  20031=>"100011101",
  20032=>"011101100",
  20033=>"010100111",
  20034=>"100110101",
  20035=>"110101011",
  20036=>"101100001",
  20037=>"101111110",
  20038=>"010001011",
  20039=>"111010011",
  20040=>"010000100",
  20041=>"110000000",
  20042=>"001011100",
  20043=>"101111100",
  20044=>"000110110",
  20045=>"010101000",
  20046=>"001101011",
  20047=>"111101010",
  20048=>"010110011",
  20049=>"111001110",
  20050=>"110001111",
  20051=>"101000100",
  20052=>"000100101",
  20053=>"000001001",
  20054=>"001001100",
  20055=>"000111011",
  20056=>"100011001",
  20057=>"111100110",
  20058=>"001111101",
  20059=>"101010101",
  20060=>"000101101",
  20061=>"000011000",
  20062=>"001001101",
  20063=>"101101101",
  20064=>"011010000",
  20065=>"110011111",
  20066=>"110100110",
  20067=>"001100010",
  20068=>"111110000",
  20069=>"100001000",
  20070=>"010110110",
  20071=>"101011111",
  20072=>"000100100",
  20073=>"101010000",
  20074=>"000000100",
  20075=>"101010001",
  20076=>"101000101",
  20077=>"010110100",
  20078=>"111000111",
  20079=>"100010010",
  20080=>"111000110",
  20081=>"000100001",
  20082=>"100000110",
  20083=>"100011100",
  20084=>"101100011",
  20085=>"000001111",
  20086=>"000001001",
  20087=>"101101000",
  20088=>"101110000",
  20089=>"111100000",
  20090=>"100110101",
  20091=>"010111100",
  20092=>"101110000",
  20093=>"110010111",
  20094=>"000110000",
  20095=>"111101101",
  20096=>"101110111",
  20097=>"101110111",
  20098=>"110001000",
  20099=>"111101011",
  20100=>"000110000",
  20101=>"001000011",
  20102=>"011010000",
  20103=>"111100010",
  20104=>"001100101",
  20105=>"011001111",
  20106=>"000001011",
  20107=>"111100010",
  20108=>"110100001",
  20109=>"011101111",
  20110=>"011000101",
  20111=>"000100000",
  20112=>"100110000",
  20113=>"010101100",
  20114=>"001110000",
  20115=>"001100011",
  20116=>"011101001",
  20117=>"110011100",
  20118=>"000001111",
  20119=>"110000011",
  20120=>"000100001",
  20121=>"110101001",
  20122=>"100110010",
  20123=>"010110110",
  20124=>"111011011",
  20125=>"110111101",
  20126=>"000101101",
  20127=>"011101011",
  20128=>"100111000",
  20129=>"100010011",
  20130=>"000000011",
  20131=>"101100110",
  20132=>"001110001",
  20133=>"010010010",
  20134=>"100001111",
  20135=>"000001001",
  20136=>"001100011",
  20137=>"001110100",
  20138=>"000001110",
  20139=>"110010110",
  20140=>"011000111",
  20141=>"010000100",
  20142=>"001111010",
  20143=>"111101001",
  20144=>"001001101",
  20145=>"010100101",
  20146=>"001011001",
  20147=>"011001111",
  20148=>"100100111",
  20149=>"001101111",
  20150=>"010100001",
  20151=>"000011000",
  20152=>"011000111",
  20153=>"110010110",
  20154=>"000110000",
  20155=>"100110100",
  20156=>"000110000",
  20157=>"011000110",
  20158=>"010011111",
  20159=>"101011001",
  20160=>"001011001",
  20161=>"101101010",
  20162=>"111111010",
  20163=>"001010001",
  20164=>"110110110",
  20165=>"011011000",
  20166=>"000101001",
  20167=>"100100101",
  20168=>"010101111",
  20169=>"000100010",
  20170=>"000011011",
  20171=>"101001011",
  20172=>"000110111",
  20173=>"111101001",
  20174=>"110001001",
  20175=>"101011111",
  20176=>"110101000",
  20177=>"110001101",
  20178=>"011100101",
  20179=>"111010001",
  20180=>"000001101",
  20181=>"110000000",
  20182=>"110000100",
  20183=>"010110100",
  20184=>"011000110",
  20185=>"101010111",
  20186=>"110001101",
  20187=>"101011111",
  20188=>"011111010",
  20189=>"110000010",
  20190=>"000110110",
  20191=>"010111000",
  20192=>"110011110",
  20193=>"100000000",
  20194=>"001011000",
  20195=>"001111001",
  20196=>"010001000",
  20197=>"100100110",
  20198=>"010100110",
  20199=>"110111000",
  20200=>"011011111",
  20201=>"000110100",
  20202=>"011101101",
  20203=>"100100011",
  20204=>"000110100",
  20205=>"100010010",
  20206=>"010101001",
  20207=>"101111111",
  20208=>"110111110",
  20209=>"011111111",
  20210=>"010000110",
  20211=>"110101110",
  20212=>"011001010",
  20213=>"100110101",
  20214=>"000100101",
  20215=>"101101101",
  20216=>"010010000",
  20217=>"000100001",
  20218=>"000011111",
  20219=>"000010011",
  20220=>"101010100",
  20221=>"110110110",
  20222=>"011000100",
  20223=>"100001000",
  20224=>"001110100",
  20225=>"001111001",
  20226=>"010001010",
  20227=>"001011111",
  20228=>"011001011",
  20229=>"010000000",
  20230=>"110111101",
  20231=>"111001110",
  20232=>"110001101",
  20233=>"000110010",
  20234=>"000010101",
  20235=>"000111000",
  20236=>"101101101",
  20237=>"110111110",
  20238=>"110011010",
  20239=>"110111101",
  20240=>"110001010",
  20241=>"101000000",
  20242=>"100010100",
  20243=>"010100100",
  20244=>"010111110",
  20245=>"001101000",
  20246=>"011001111",
  20247=>"010100111",
  20248=>"111111101",
  20249=>"100011101",
  20250=>"011011000",
  20251=>"100010110",
  20252=>"000011010",
  20253=>"010110100",
  20254=>"100111110",
  20255=>"010010110",
  20256=>"100101101",
  20257=>"111110001",
  20258=>"101000000",
  20259=>"000110110",
  20260=>"000000010",
  20261=>"011001111",
  20262=>"010111110",
  20263=>"000110000",
  20264=>"100100011",
  20265=>"100000001",
  20266=>"100001011",
  20267=>"111111000",
  20268=>"011100001",
  20269=>"010010010",
  20270=>"000110001",
  20271=>"010011011",
  20272=>"000010001",
  20273=>"111110110",
  20274=>"110000011",
  20275=>"011000010",
  20276=>"100100101",
  20277=>"110111010",
  20278=>"001000001",
  20279=>"000111001",
  20280=>"010010000",
  20281=>"010001000",
  20282=>"101101011",
  20283=>"000100001",
  20284=>"010101010",
  20285=>"100010000",
  20286=>"000110111",
  20287=>"110011100",
  20288=>"111111110",
  20289=>"101100111",
  20290=>"011110111",
  20291=>"000101100",
  20292=>"010000101",
  20293=>"101100011",
  20294=>"000010011",
  20295=>"001110111",
  20296=>"111011101",
  20297=>"100101011",
  20298=>"001100111",
  20299=>"001101010",
  20300=>"010010101",
  20301=>"101111011",
  20302=>"001000011",
  20303=>"001011010",
  20304=>"010001110",
  20305=>"000000111",
  20306=>"001001111",
  20307=>"000001101",
  20308=>"011100110",
  20309=>"011110011",
  20310=>"000100011",
  20311=>"100110010",
  20312=>"110011010",
  20313=>"000001110",
  20314=>"010001001",
  20315=>"010011010",
  20316=>"110000011",
  20317=>"011000101",
  20318=>"110010111",
  20319=>"101001101",
  20320=>"111110011",
  20321=>"001111100",
  20322=>"111110110",
  20323=>"000011101",
  20324=>"010111111",
  20325=>"111111111",
  20326=>"110000000",
  20327=>"001101010",
  20328=>"110011010",
  20329=>"101011010",
  20330=>"101101100",
  20331=>"001100100",
  20332=>"100000101",
  20333=>"111110101",
  20334=>"000001001",
  20335=>"100011011",
  20336=>"110101000",
  20337=>"011101000",
  20338=>"111000110",
  20339=>"001010001",
  20340=>"000110010",
  20341=>"011000101",
  20342=>"000011000",
  20343=>"000000100",
  20344=>"010111000",
  20345=>"111000101",
  20346=>"111110111",
  20347=>"100011101",
  20348=>"001000000",
  20349=>"001110100",
  20350=>"111100001",
  20351=>"111000010",
  20352=>"111001100",
  20353=>"011011100",
  20354=>"100010011",
  20355=>"010000100",
  20356=>"100000011",
  20357=>"100101000",
  20358=>"010111010",
  20359=>"001101010",
  20360=>"001000110",
  20361=>"110100011",
  20362=>"011000001",
  20363=>"100011011",
  20364=>"011001100",
  20365=>"100100010",
  20366=>"111111110",
  20367=>"110110000",
  20368=>"011110100",
  20369=>"110111001",
  20370=>"000010110",
  20371=>"010110011",
  20372=>"001110111",
  20373=>"011001010",
  20374=>"101110000",
  20375=>"001111111",
  20376=>"100000100",
  20377=>"001000001",
  20378=>"100011000",
  20379=>"101000100",
  20380=>"100111111",
  20381=>"101100101",
  20382=>"011100110",
  20383=>"111001000",
  20384=>"000001011",
  20385=>"010100111",
  20386=>"001110011",
  20387=>"110001000",
  20388=>"001000001",
  20389=>"101000110",
  20390=>"101011001",
  20391=>"011000001",
  20392=>"110100000",
  20393=>"000110010",
  20394=>"001001011",
  20395=>"011101111",
  20396=>"000100100",
  20397=>"001011110",
  20398=>"111100100",
  20399=>"000000111",
  20400=>"111010100",
  20401=>"111110111",
  20402=>"101011101",
  20403=>"111011010",
  20404=>"111101000",
  20405=>"110011101",
  20406=>"011000111",
  20407=>"000001100",
  20408=>"111001101",
  20409=>"001111011",
  20410=>"110011100",
  20411=>"100001111",
  20412=>"100101001",
  20413=>"001110000",
  20414=>"001010110",
  20415=>"001011001",
  20416=>"000101010",
  20417=>"101101110",
  20418=>"100111111",
  20419=>"000010010",
  20420=>"110010111",
  20421=>"110000001",
  20422=>"011010111",
  20423=>"110010111",
  20424=>"000000010",
  20425=>"101101010",
  20426=>"101001101",
  20427=>"110101010",
  20428=>"000000010",
  20429=>"100110101",
  20430=>"001011010",
  20431=>"111001000",
  20432=>"011101101",
  20433=>"011011001",
  20434=>"100100000",
  20435=>"010001001",
  20436=>"110001001",
  20437=>"100110111",
  20438=>"000110100",
  20439=>"000000000",
  20440=>"111000010",
  20441=>"111100001",
  20442=>"011000110",
  20443=>"011111101",
  20444=>"111001001",
  20445=>"111011100",
  20446=>"000101101",
  20447=>"111110011",
  20448=>"010001100",
  20449=>"100001010",
  20450=>"100011011",
  20451=>"101001101",
  20452=>"000000001",
  20453=>"101100001",
  20454=>"111111001",
  20455=>"110000010",
  20456=>"110111111",
  20457=>"110111000",
  20458=>"101101001",
  20459=>"011111011",
  20460=>"000100001",
  20461=>"100001001",
  20462=>"100110010",
  20463=>"000101000",
  20464=>"100001101",
  20465=>"100100010",
  20466=>"101110000",
  20467=>"111101101",
  20468=>"110011111",
  20469=>"100011110",
  20470=>"011001101",
  20471=>"101111100",
  20472=>"010100001",
  20473=>"101100110",
  20474=>"001101111",
  20475=>"011010001",
  20476=>"111100101",
  20477=>"010111011",
  20478=>"000001110",
  20479=>"000111101",
  20480=>"101001110",
  20481=>"000110011",
  20482=>"010110100",
  20483=>"010010111",
  20484=>"101001001",
  20485=>"110011100",
  20486=>"000010011",
  20487=>"111101000",
  20488=>"011001010",
  20489=>"011110011",
  20490=>"101000111",
  20491=>"100011110",
  20492=>"001100011",
  20493=>"011000100",
  20494=>"000111110",
  20495=>"010100010",
  20496=>"100110010",
  20497=>"001100001",
  20498=>"101011000",
  20499=>"011110001",
  20500=>"010100100",
  20501=>"101101111",
  20502=>"111111110",
  20503=>"100000000",
  20504=>"010101000",
  20505=>"001001110",
  20506=>"000101110",
  20507=>"000001100",
  20508=>"111101101",
  20509=>"011000101",
  20510=>"110001101",
  20511=>"000111011",
  20512=>"001001111",
  20513=>"011101011",
  20514=>"110101110",
  20515=>"001011110",
  20516=>"010011010",
  20517=>"010011101",
  20518=>"000110001",
  20519=>"110101111",
  20520=>"110111000",
  20521=>"011000110",
  20522=>"010010110",
  20523=>"001001001",
  20524=>"101011001",
  20525=>"101111010",
  20526=>"011100100",
  20527=>"001101110",
  20528=>"001011110",
  20529=>"010100100",
  20530=>"111010010",
  20531=>"110010101",
  20532=>"111001111",
  20533=>"101101000",
  20534=>"110111011",
  20535=>"001001101",
  20536=>"011000001",
  20537=>"010100101",
  20538=>"100111111",
  20539=>"010001011",
  20540=>"000001000",
  20541=>"101100011",
  20542=>"101100111",
  20543=>"000001101",
  20544=>"010011100",
  20545=>"101000000",
  20546=>"100010100",
  20547=>"001011010",
  20548=>"111100101",
  20549=>"111101101",
  20550=>"100010110",
  20551=>"101010100",
  20552=>"001011101",
  20553=>"010011000",
  20554=>"100110010",
  20555=>"110000100",
  20556=>"100000010",
  20557=>"100011010",
  20558=>"111111111",
  20559=>"101100001",
  20560=>"011110011",
  20561=>"110100110",
  20562=>"010111111",
  20563=>"100110001",
  20564=>"000000100",
  20565=>"111010000",
  20566=>"000000110",
  20567=>"110111010",
  20568=>"010101111",
  20569=>"110101001",
  20570=>"011111000",
  20571=>"101000011",
  20572=>"000010010",
  20573=>"010000100",
  20574=>"000001000",
  20575=>"000001111",
  20576=>"100000001",
  20577=>"011001001",
  20578=>"011110101",
  20579=>"010010111",
  20580=>"011111011",
  20581=>"100111101",
  20582=>"111011000",
  20583=>"100001000",
  20584=>"000101110",
  20585=>"100010010",
  20586=>"001101100",
  20587=>"110111111",
  20588=>"111100101",
  20589=>"111101101",
  20590=>"000110000",
  20591=>"111100001",
  20592=>"110111010",
  20593=>"000110010",
  20594=>"010110011",
  20595=>"111101111",
  20596=>"100001001",
  20597=>"111100010",
  20598=>"001001001",
  20599=>"101110000",
  20600=>"000111011",
  20601=>"111000011",
  20602=>"111111001",
  20603=>"101100101",
  20604=>"110000000",
  20605=>"010000111",
  20606=>"110000011",
  20607=>"010001110",
  20608=>"011100001",
  20609=>"001111101",
  20610=>"000011000",
  20611=>"000100100",
  20612=>"001001101",
  20613=>"001100010",
  20614=>"001011111",
  20615=>"101001100",
  20616=>"101011011",
  20617=>"111011100",
  20618=>"101111000",
  20619=>"010011001",
  20620=>"110101001",
  20621=>"001111100",
  20622=>"110100010",
  20623=>"010101111",
  20624=>"110100111",
  20625=>"000110011",
  20626=>"110110101",
  20627=>"101011001",
  20628=>"000010100",
  20629=>"001110000",
  20630=>"001011000",
  20631=>"111110111",
  20632=>"011010010",
  20633=>"111101101",
  20634=>"010111000",
  20635=>"010010100",
  20636=>"001010010",
  20637=>"101100111",
  20638=>"100011001",
  20639=>"010000010",
  20640=>"111111001",
  20641=>"101110110",
  20642=>"100110100",
  20643=>"001011110",
  20644=>"101001010",
  20645=>"010000110",
  20646=>"110110110",
  20647=>"111100000",
  20648=>"010010100",
  20649=>"110101001",
  20650=>"100100110",
  20651=>"001100110",
  20652=>"100000111",
  20653=>"110001100",
  20654=>"110001110",
  20655=>"010011110",
  20656=>"001100100",
  20657=>"000101001",
  20658=>"000000011",
  20659=>"000001100",
  20660=>"001111000",
  20661=>"111010100",
  20662=>"110011100",
  20663=>"101101010",
  20664=>"011000010",
  20665=>"000100100",
  20666=>"110101001",
  20667=>"001111001",
  20668=>"011110100",
  20669=>"001010111",
  20670=>"001000100",
  20671=>"011010111",
  20672=>"101111011",
  20673=>"000010100",
  20674=>"011101000",
  20675=>"000001100",
  20676=>"111110110",
  20677=>"110000000",
  20678=>"101010110",
  20679=>"010010101",
  20680=>"011011110",
  20681=>"000111101",
  20682=>"111001101",
  20683=>"101101011",
  20684=>"101111000",
  20685=>"101111110",
  20686=>"000000011",
  20687=>"000110001",
  20688=>"100000010",
  20689=>"011010001",
  20690=>"110011000",
  20691=>"000110001",
  20692=>"101001001",
  20693=>"111001000",
  20694=>"101000000",
  20695=>"100010101",
  20696=>"011000000",
  20697=>"111011010",
  20698=>"000001001",
  20699=>"000011100",
  20700=>"001101011",
  20701=>"111110010",
  20702=>"000000000",
  20703=>"010111100",
  20704=>"101000010",
  20705=>"000100000",
  20706=>"111111111",
  20707=>"000111101",
  20708=>"011111110",
  20709=>"010100001",
  20710=>"010000100",
  20711=>"110101011",
  20712=>"010000010",
  20713=>"011011100",
  20714=>"010000100",
  20715=>"110010100",
  20716=>"101000001",
  20717=>"011001100",
  20718=>"100001010",
  20719=>"110001011",
  20720=>"010000110",
  20721=>"000101100",
  20722=>"010101000",
  20723=>"111001111",
  20724=>"110011111",
  20725=>"001110101",
  20726=>"100100010",
  20727=>"010101000",
  20728=>"100001000",
  20729=>"111110100",
  20730=>"011110011",
  20731=>"010101010",
  20732=>"110100011",
  20733=>"111111010",
  20734=>"000001111",
  20735=>"010010111",
  20736=>"101111001",
  20737=>"110010010",
  20738=>"000110000",
  20739=>"111001011",
  20740=>"101111110",
  20741=>"010110000",
  20742=>"110101010",
  20743=>"010110000",
  20744=>"001101000",
  20745=>"010100000",
  20746=>"010011111",
  20747=>"111100111",
  20748=>"110010001",
  20749=>"111001011",
  20750=>"010111101",
  20751=>"001011100",
  20752=>"011000001",
  20753=>"101110101",
  20754=>"010011110",
  20755=>"101110101",
  20756=>"100101110",
  20757=>"011001110",
  20758=>"001010010",
  20759=>"100001101",
  20760=>"011010101",
  20761=>"111010001",
  20762=>"001100001",
  20763=>"111101011",
  20764=>"000110010",
  20765=>"111110010",
  20766=>"111011001",
  20767=>"100010100",
  20768=>"010000110",
  20769=>"001011100",
  20770=>"000010000",
  20771=>"110110111",
  20772=>"011010000",
  20773=>"110001001",
  20774=>"111101010",
  20775=>"100110000",
  20776=>"100100001",
  20777=>"111111101",
  20778=>"010111101",
  20779=>"111010001",
  20780=>"100001010",
  20781=>"100001110",
  20782=>"111110011",
  20783=>"101010010",
  20784=>"000110100",
  20785=>"100111111",
  20786=>"000000110",
  20787=>"110000010",
  20788=>"111001100",
  20789=>"111001110",
  20790=>"111100110",
  20791=>"010001111",
  20792=>"000101100",
  20793=>"110111011",
  20794=>"011110100",
  20795=>"011000100",
  20796=>"001011100",
  20797=>"011011110",
  20798=>"100010100",
  20799=>"011001000",
  20800=>"111100100",
  20801=>"011000100",
  20802=>"011010101",
  20803=>"100110010",
  20804=>"000110000",
  20805=>"100101010",
  20806=>"110011000",
  20807=>"010000110",
  20808=>"100011100",
  20809=>"101000000",
  20810=>"011110101",
  20811=>"001010110",
  20812=>"000011011",
  20813=>"010111001",
  20814=>"111010100",
  20815=>"010101001",
  20816=>"111110011",
  20817=>"101001011",
  20818=>"011010100",
  20819=>"000001000",
  20820=>"001101111",
  20821=>"110001100",
  20822=>"011101111",
  20823=>"000001001",
  20824=>"100010010",
  20825=>"111000011",
  20826=>"111101110",
  20827=>"111101101",
  20828=>"011110100",
  20829=>"000000111",
  20830=>"110001110",
  20831=>"111010101",
  20832=>"101000100",
  20833=>"101010101",
  20834=>"111100000",
  20835=>"001001001",
  20836=>"010010000",
  20837=>"110110001",
  20838=>"111111100",
  20839=>"010010001",
  20840=>"110111111",
  20841=>"001010110",
  20842=>"110111100",
  20843=>"011101000",
  20844=>"001100000",
  20845=>"011100110",
  20846=>"000010011",
  20847=>"111011100",
  20848=>"110100111",
  20849=>"101000000",
  20850=>"111101001",
  20851=>"000111010",
  20852=>"001000001",
  20853=>"111110111",
  20854=>"101110101",
  20855=>"001000000",
  20856=>"000100101",
  20857=>"101010001",
  20858=>"110000011",
  20859=>"011101101",
  20860=>"110110001",
  20861=>"011101111",
  20862=>"010111101",
  20863=>"000010001",
  20864=>"010010000",
  20865=>"110001001",
  20866=>"110100010",
  20867=>"010100001",
  20868=>"011100110",
  20869=>"000000010",
  20870=>"110110011",
  20871=>"101000110",
  20872=>"100000010",
  20873=>"000110100",
  20874=>"000100110",
  20875=>"000100111",
  20876=>"001101001",
  20877=>"001100100",
  20878=>"000001110",
  20879=>"010101100",
  20880=>"100010011",
  20881=>"000000000",
  20882=>"010110111",
  20883=>"011001001",
  20884=>"111110111",
  20885=>"001100000",
  20886=>"110010100",
  20887=>"111000000",
  20888=>"010000110",
  20889=>"000100001",
  20890=>"001100000",
  20891=>"111011011",
  20892=>"111111100",
  20893=>"010100110",
  20894=>"001100100",
  20895=>"001000110",
  20896=>"111011011",
  20897=>"010101101",
  20898=>"100111011",
  20899=>"011001001",
  20900=>"111110010",
  20901=>"100101011",
  20902=>"101111111",
  20903=>"011111001",
  20904=>"111101000",
  20905=>"001110110",
  20906=>"000000100",
  20907=>"010000001",
  20908=>"000000000",
  20909=>"111101100",
  20910=>"110000100",
  20911=>"000000001",
  20912=>"101110111",
  20913=>"111101000",
  20914=>"000000110",
  20915=>"001110111",
  20916=>"111101110",
  20917=>"101111001",
  20918=>"000000101",
  20919=>"101101001",
  20920=>"001010111",
  20921=>"110000001",
  20922=>"101000010",
  20923=>"101101101",
  20924=>"100111100",
  20925=>"011101101",
  20926=>"101001000",
  20927=>"111011101",
  20928=>"000001000",
  20929=>"100101110",
  20930=>"110111101",
  20931=>"011000111",
  20932=>"010111010",
  20933=>"101111011",
  20934=>"101010011",
  20935=>"100010101",
  20936=>"000001000",
  20937=>"000100000",
  20938=>"010100000",
  20939=>"000001011",
  20940=>"001000100",
  20941=>"011001010",
  20942=>"011011010",
  20943=>"100101110",
  20944=>"111001011",
  20945=>"100000000",
  20946=>"000000101",
  20947=>"011110110",
  20948=>"010110000",
  20949=>"000101100",
  20950=>"000110101",
  20951=>"011100100",
  20952=>"110100010",
  20953=>"110010001",
  20954=>"010010100",
  20955=>"100010100",
  20956=>"000101000",
  20957=>"111101001",
  20958=>"010110111",
  20959=>"000111000",
  20960=>"111010100",
  20961=>"000110101",
  20962=>"011100001",
  20963=>"100111011",
  20964=>"111010010",
  20965=>"111010001",
  20966=>"011011111",
  20967=>"010100110",
  20968=>"000011101",
  20969=>"000011110",
  20970=>"101010110",
  20971=>"001001010",
  20972=>"110001100",
  20973=>"100110100",
  20974=>"011011100",
  20975=>"100101011",
  20976=>"110100011",
  20977=>"011111111",
  20978=>"101010011",
  20979=>"000011011",
  20980=>"111000010",
  20981=>"011100110",
  20982=>"100000101",
  20983=>"011100111",
  20984=>"001001100",
  20985=>"000110000",
  20986=>"101111001",
  20987=>"111111000",
  20988=>"010100110",
  20989=>"101011011",
  20990=>"111011001",
  20991=>"011011101",
  20992=>"010111100",
  20993=>"001101111",
  20994=>"110100101",
  20995=>"010010001",
  20996=>"010000011",
  20997=>"010110000",
  20998=>"011000000",
  20999=>"011011001",
  21000=>"101001100",
  21001=>"010000000",
  21002=>"111010101",
  21003=>"100000101",
  21004=>"000000110",
  21005=>"001110010",
  21006=>"111001000",
  21007=>"100100111",
  21008=>"111011101",
  21009=>"000011110",
  21010=>"000011111",
  21011=>"011010111",
  21012=>"100010101",
  21013=>"111101011",
  21014=>"100001000",
  21015=>"000011000",
  21016=>"000010111",
  21017=>"110001111",
  21018=>"000100000",
  21019=>"101011111",
  21020=>"010101000",
  21021=>"100010011",
  21022=>"011100010",
  21023=>"000110110",
  21024=>"111010011",
  21025=>"101110000",
  21026=>"011010110",
  21027=>"111001001",
  21028=>"110110000",
  21029=>"111110100",
  21030=>"000011000",
  21031=>"111100111",
  21032=>"010001101",
  21033=>"011111101",
  21034=>"010111001",
  21035=>"101000101",
  21036=>"000100110",
  21037=>"100010001",
  21038=>"010001101",
  21039=>"000000000",
  21040=>"101100011",
  21041=>"010011111",
  21042=>"101101100",
  21043=>"111101110",
  21044=>"010101100",
  21045=>"111001000",
  21046=>"110000100",
  21047=>"100000100",
  21048=>"110101010",
  21049=>"111010110",
  21050=>"001001010",
  21051=>"010000100",
  21052=>"010101001",
  21053=>"000111010",
  21054=>"101101000",
  21055=>"011111011",
  21056=>"110000001",
  21057=>"011010001",
  21058=>"011011010",
  21059=>"110111100",
  21060=>"110100101",
  21061=>"010111101",
  21062=>"100000000",
  21063=>"011010110",
  21064=>"011110110",
  21065=>"110001100",
  21066=>"110010101",
  21067=>"101001000",
  21068=>"000011101",
  21069=>"010000101",
  21070=>"100101101",
  21071=>"000001100",
  21072=>"110000111",
  21073=>"100101111",
  21074=>"010111110",
  21075=>"000110000",
  21076=>"101100110",
  21077=>"010001010",
  21078=>"100010010",
  21079=>"101110000",
  21080=>"101011011",
  21081=>"100011010",
  21082=>"100010111",
  21083=>"101000101",
  21084=>"011001111",
  21085=>"001100100",
  21086=>"101100101",
  21087=>"101111011",
  21088=>"011000010",
  21089=>"011010000",
  21090=>"101110111",
  21091=>"111100100",
  21092=>"000010000",
  21093=>"011111111",
  21094=>"110010010",
  21095=>"001100011",
  21096=>"000000010",
  21097=>"000010000",
  21098=>"101110011",
  21099=>"011001001",
  21100=>"000110001",
  21101=>"100110111",
  21102=>"110100011",
  21103=>"111110000",
  21104=>"000001001",
  21105=>"110110011",
  21106=>"010010111",
  21107=>"011000111",
  21108=>"100000111",
  21109=>"101011000",
  21110=>"100010011",
  21111=>"110100110",
  21112=>"101100011",
  21113=>"100011001",
  21114=>"001111000",
  21115=>"100011110",
  21116=>"111000110",
  21117=>"000010110",
  21118=>"111001000",
  21119=>"011010001",
  21120=>"011011010",
  21121=>"111110000",
  21122=>"110111000",
  21123=>"001001001",
  21124=>"110000111",
  21125=>"000110101",
  21126=>"010110001",
  21127=>"101111110",
  21128=>"111111101",
  21129=>"110010001",
  21130=>"011010100",
  21131=>"011011010",
  21132=>"000100000",
  21133=>"010110101",
  21134=>"010000010",
  21135=>"111000100",
  21136=>"000110110",
  21137=>"101101101",
  21138=>"100100001",
  21139=>"101100011",
  21140=>"010100001",
  21141=>"111110010",
  21142=>"101011010",
  21143=>"011101110",
  21144=>"010111100",
  21145=>"100010110",
  21146=>"111100111",
  21147=>"011010111",
  21148=>"110101010",
  21149=>"010111100",
  21150=>"011101000",
  21151=>"110101101",
  21152=>"001110111",
  21153=>"111100101",
  21154=>"011101110",
  21155=>"010100010",
  21156=>"100000111",
  21157=>"011111001",
  21158=>"011000100",
  21159=>"000000000",
  21160=>"000001010",
  21161=>"000010100",
  21162=>"010101111",
  21163=>"100000100",
  21164=>"000111000",
  21165=>"101001111",
  21166=>"111101111",
  21167=>"010101000",
  21168=>"100000101",
  21169=>"100111000",
  21170=>"010011000",
  21171=>"100001101",
  21172=>"000110000",
  21173=>"011100110",
  21174=>"110111101",
  21175=>"010001010",
  21176=>"100111100",
  21177=>"011000110",
  21178=>"111000101",
  21179=>"000101100",
  21180=>"110000100",
  21181=>"000010010",
  21182=>"110011110",
  21183=>"010110010",
  21184=>"001001010",
  21185=>"111101010",
  21186=>"000011010",
  21187=>"111110001",
  21188=>"010101100",
  21189=>"001110101",
  21190=>"111110101",
  21191=>"101001000",
  21192=>"000101010",
  21193=>"111000111",
  21194=>"110101011",
  21195=>"011001010",
  21196=>"000011101",
  21197=>"101111010",
  21198=>"001101111",
  21199=>"010001000",
  21200=>"001011001",
  21201=>"110110111",
  21202=>"000110011",
  21203=>"001111011",
  21204=>"010101001",
  21205=>"010010111",
  21206=>"101100010",
  21207=>"000001011",
  21208=>"001111101",
  21209=>"001011011",
  21210=>"001111101",
  21211=>"111001011",
  21212=>"111100000",
  21213=>"101101110",
  21214=>"000000101",
  21215=>"110011000",
  21216=>"000000001",
  21217=>"111110011",
  21218=>"110011100",
  21219=>"111000111",
  21220=>"011000000",
  21221=>"110100111",
  21222=>"001011111",
  21223=>"000000011",
  21224=>"100001110",
  21225=>"111100100",
  21226=>"001000110",
  21227=>"000001001",
  21228=>"000010010",
  21229=>"100101011",
  21230=>"101011111",
  21231=>"010101000",
  21232=>"010100011",
  21233=>"100101000",
  21234=>"111111001",
  21235=>"110001010",
  21236=>"010010100",
  21237=>"001100000",
  21238=>"100100010",
  21239=>"011001011",
  21240=>"101010100",
  21241=>"010010100",
  21242=>"100000011",
  21243=>"110111011",
  21244=>"001100111",
  21245=>"000110111",
  21246=>"101100100",
  21247=>"111000001",
  21248=>"110000100",
  21249=>"000100010",
  21250=>"111100111",
  21251=>"111000011",
  21252=>"100100101",
  21253=>"100100100",
  21254=>"010101100",
  21255=>"011001010",
  21256=>"110000101",
  21257=>"101001111",
  21258=>"111110001",
  21259=>"011000011",
  21260=>"010100110",
  21261=>"001010110",
  21262=>"000101010",
  21263=>"101000101",
  21264=>"101010100",
  21265=>"111000011",
  21266=>"000010101",
  21267=>"011010101",
  21268=>"001101001",
  21269=>"001100101",
  21270=>"010010101",
  21271=>"100100110",
  21272=>"010011000",
  21273=>"001010010",
  21274=>"000011100",
  21275=>"011100100",
  21276=>"011111000",
  21277=>"100111001",
  21278=>"111100100",
  21279=>"100010011",
  21280=>"001100000",
  21281=>"000100100",
  21282=>"000001111",
  21283=>"010010010",
  21284=>"010111000",
  21285=>"111001000",
  21286=>"011100111",
  21287=>"011100100",
  21288=>"011000101",
  21289=>"111001010",
  21290=>"111111100",
  21291=>"011100111",
  21292=>"100000010",
  21293=>"101001000",
  21294=>"101000110",
  21295=>"110000001",
  21296=>"101100101",
  21297=>"001101000",
  21298=>"111110101",
  21299=>"010000101",
  21300=>"110101111",
  21301=>"001000011",
  21302=>"010011000",
  21303=>"110011001",
  21304=>"001000110",
  21305=>"010001011",
  21306=>"010011101",
  21307=>"010010001",
  21308=>"010100100",
  21309=>"111111110",
  21310=>"111110110",
  21311=>"010100110",
  21312=>"111010010",
  21313=>"110000111",
  21314=>"111111101",
  21315=>"011110000",
  21316=>"001010001",
  21317=>"100101110",
  21318=>"011011001",
  21319=>"101111101",
  21320=>"010100000",
  21321=>"010111001",
  21322=>"100001110",
  21323=>"011110000",
  21324=>"010111101",
  21325=>"110111111",
  21326=>"010100011",
  21327=>"000111101",
  21328=>"101110001",
  21329=>"111010100",
  21330=>"110110100",
  21331=>"110000100",
  21332=>"100000000",
  21333=>"100000011",
  21334=>"110101010",
  21335=>"110111101",
  21336=>"100000000",
  21337=>"110111110",
  21338=>"110100010",
  21339=>"111110111",
  21340=>"101011111",
  21341=>"100111010",
  21342=>"010110001",
  21343=>"000010100",
  21344=>"011101101",
  21345=>"111111010",
  21346=>"000110100",
  21347=>"110100101",
  21348=>"100111011",
  21349=>"110110010",
  21350=>"110110001",
  21351=>"011011111",
  21352=>"000010001",
  21353=>"111000110",
  21354=>"010100010",
  21355=>"001111110",
  21356=>"100111101",
  21357=>"011001111",
  21358=>"001100011",
  21359=>"011111001",
  21360=>"101101011",
  21361=>"100111000",
  21362=>"010011111",
  21363=>"011110100",
  21364=>"011000100",
  21365=>"001010111",
  21366=>"001111110",
  21367=>"101011000",
  21368=>"110100000",
  21369=>"001000000",
  21370=>"001100000",
  21371=>"010001001",
  21372=>"110100000",
  21373=>"000000111",
  21374=>"001101111",
  21375=>"000100100",
  21376=>"110011111",
  21377=>"011100111",
  21378=>"000000001",
  21379=>"001000000",
  21380=>"100110111",
  21381=>"111000110",
  21382=>"001010110",
  21383=>"101010110",
  21384=>"001111111",
  21385=>"110110111",
  21386=>"011101100",
  21387=>"000000011",
  21388=>"111000100",
  21389=>"111101101",
  21390=>"000101001",
  21391=>"100101000",
  21392=>"010011000",
  21393=>"100101001",
  21394=>"110010000",
  21395=>"001101100",
  21396=>"100100101",
  21397=>"011000011",
  21398=>"101000101",
  21399=>"101010011",
  21400=>"000011000",
  21401=>"001011000",
  21402=>"010111110",
  21403=>"110100100",
  21404=>"111111001",
  21405=>"101101000",
  21406=>"100000010",
  21407=>"101010000",
  21408=>"110100011",
  21409=>"001111101",
  21410=>"111000110",
  21411=>"010000000",
  21412=>"110000001",
  21413=>"010011100",
  21414=>"101101110",
  21415=>"011101110",
  21416=>"010000001",
  21417=>"110110010",
  21418=>"001111110",
  21419=>"100100000",
  21420=>"010000000",
  21421=>"010100110",
  21422=>"111110101",
  21423=>"011011100",
  21424=>"010010010",
  21425=>"100111010",
  21426=>"001110110",
  21427=>"000001011",
  21428=>"100111010",
  21429=>"010001000",
  21430=>"011000111",
  21431=>"101011011",
  21432=>"010110000",
  21433=>"001000001",
  21434=>"110101100",
  21435=>"011011111",
  21436=>"001100011",
  21437=>"101011011",
  21438=>"100111110",
  21439=>"110010001",
  21440=>"001001001",
  21441=>"010010010",
  21442=>"011101110",
  21443=>"010111011",
  21444=>"000100010",
  21445=>"111110111",
  21446=>"101001001",
  21447=>"001010000",
  21448=>"101100110",
  21449=>"100100001",
  21450=>"111110011",
  21451=>"100111110",
  21452=>"000100111",
  21453=>"001100000",
  21454=>"100000010",
  21455=>"111011110",
  21456=>"010110111",
  21457=>"001000000",
  21458=>"110111100",
  21459=>"110101101",
  21460=>"010101010",
  21461=>"111101100",
  21462=>"001111011",
  21463=>"100001110",
  21464=>"000111100",
  21465=>"001001101",
  21466=>"000100111",
  21467=>"000101100",
  21468=>"111101000",
  21469=>"011111101",
  21470=>"101011100",
  21471=>"011101011",
  21472=>"000100000",
  21473=>"010010101",
  21474=>"010101011",
  21475=>"111001110",
  21476=>"000000011",
  21477=>"001011101",
  21478=>"111100010",
  21479=>"000110010",
  21480=>"011000010",
  21481=>"101100111",
  21482=>"000111000",
  21483=>"110101000",
  21484=>"111111001",
  21485=>"101101101",
  21486=>"001110100",
  21487=>"111010001",
  21488=>"010010101",
  21489=>"101011100",
  21490=>"000100001",
  21491=>"101111101",
  21492=>"001111110",
  21493=>"010101001",
  21494=>"110011000",
  21495=>"001000000",
  21496=>"100100000",
  21497=>"010000111",
  21498=>"111000001",
  21499=>"110000001",
  21500=>"011100100",
  21501=>"111011101",
  21502=>"100010110",
  21503=>"100010100",
  21504=>"001000010",
  21505=>"100111000",
  21506=>"010000011",
  21507=>"100100110",
  21508=>"100100001",
  21509=>"100111000",
  21510=>"100111111",
  21511=>"100011011",
  21512=>"001010011",
  21513=>"011001111",
  21514=>"100000000",
  21515=>"111100111",
  21516=>"101100011",
  21517=>"011110100",
  21518=>"001001011",
  21519=>"010010101",
  21520=>"001101010",
  21521=>"011110110",
  21522=>"000000001",
  21523=>"101100111",
  21524=>"000010000",
  21525=>"000100110",
  21526=>"001100110",
  21527=>"100111010",
  21528=>"111101010",
  21529=>"000000001",
  21530=>"111101110",
  21531=>"010000110",
  21532=>"111101000",
  21533=>"011100010",
  21534=>"011110110",
  21535=>"110100101",
  21536=>"110010010",
  21537=>"010001111",
  21538=>"111111011",
  21539=>"100011100",
  21540=>"101001000",
  21541=>"010111010",
  21542=>"110101111",
  21543=>"001001001",
  21544=>"111010011",
  21545=>"100110011",
  21546=>"101001110",
  21547=>"110010011",
  21548=>"011011101",
  21549=>"000000111",
  21550=>"110101011",
  21551=>"011000101",
  21552=>"000011001",
  21553=>"011100100",
  21554=>"111011010",
  21555=>"101011001",
  21556=>"001001100",
  21557=>"101100100",
  21558=>"111110100",
  21559=>"110010000",
  21560=>"100001001",
  21561=>"100101001",
  21562=>"110101111",
  21563=>"011011100",
  21564=>"011000100",
  21565=>"011000111",
  21566=>"111000000",
  21567=>"011000101",
  21568=>"011000010",
  21569=>"000000000",
  21570=>"100000000",
  21571=>"101001100",
  21572=>"100011111",
  21573=>"011011100",
  21574=>"111101100",
  21575=>"010000010",
  21576=>"001001011",
  21577=>"010001011",
  21578=>"101101110",
  21579=>"011011000",
  21580=>"101100101",
  21581=>"111001000",
  21582=>"101100001",
  21583=>"010010111",
  21584=>"101111000",
  21585=>"111001011",
  21586=>"010010000",
  21587=>"010111111",
  21588=>"111100100",
  21589=>"110001001",
  21590=>"111101000",
  21591=>"111111001",
  21592=>"110111011",
  21593=>"100010011",
  21594=>"111000101",
  21595=>"000000010",
  21596=>"000000110",
  21597=>"111011010",
  21598=>"000001001",
  21599=>"101000010",
  21600=>"001000001",
  21601=>"011100001",
  21602=>"111111111",
  21603=>"000010001",
  21604=>"010111001",
  21605=>"101000110",
  21606=>"010010000",
  21607=>"111010001",
  21608=>"011001001",
  21609=>"101101011",
  21610=>"110101010",
  21611=>"101110011",
  21612=>"011011001",
  21613=>"100111110",
  21614=>"000010000",
  21615=>"011011110",
  21616=>"010001101",
  21617=>"110110111",
  21618=>"110111110",
  21619=>"111011100",
  21620=>"010101000",
  21621=>"100000011",
  21622=>"100011011",
  21623=>"110111010",
  21624=>"110000111",
  21625=>"101010101",
  21626=>"101011011",
  21627=>"010110010",
  21628=>"100100010",
  21629=>"100100011",
  21630=>"100000100",
  21631=>"001110101",
  21632=>"110111101",
  21633=>"000000111",
  21634=>"111110110",
  21635=>"001101010",
  21636=>"110111011",
  21637=>"000100100",
  21638=>"001111111",
  21639=>"011101011",
  21640=>"110111010",
  21641=>"010011100",
  21642=>"011110011",
  21643=>"111010000",
  21644=>"001011110",
  21645=>"001010100",
  21646=>"010101010",
  21647=>"101101110",
  21648=>"001001011",
  21649=>"101011000",
  21650=>"011100000",
  21651=>"111000110",
  21652=>"010010011",
  21653=>"101001110",
  21654=>"111010000",
  21655=>"011011010",
  21656=>"000100100",
  21657=>"000110100",
  21658=>"010010001",
  21659=>"101011000",
  21660=>"000110010",
  21661=>"000001001",
  21662=>"101110001",
  21663=>"100101000",
  21664=>"001100010",
  21665=>"110110100",
  21666=>"000101010",
  21667=>"000110101",
  21668=>"101001111",
  21669=>"110100011",
  21670=>"110111011",
  21671=>"001011111",
  21672=>"001010111",
  21673=>"111011011",
  21674=>"011101111",
  21675=>"100100001",
  21676=>"111110111",
  21677=>"111100001",
  21678=>"100111101",
  21679=>"111111111",
  21680=>"111110001",
  21681=>"001001011",
  21682=>"111010100",
  21683=>"011101100",
  21684=>"100010101",
  21685=>"101010001",
  21686=>"011010010",
  21687=>"111000000",
  21688=>"111111011",
  21689=>"001100110",
  21690=>"101010101",
  21691=>"010111101",
  21692=>"010001100",
  21693=>"011011011",
  21694=>"010010001",
  21695=>"000111110",
  21696=>"110010111",
  21697=>"100111111",
  21698=>"001010001",
  21699=>"001010011",
  21700=>"111010101",
  21701=>"110001011",
  21702=>"011111000",
  21703=>"110100110",
  21704=>"101011101",
  21705=>"100101101",
  21706=>"011101001",
  21707=>"010101101",
  21708=>"001011111",
  21709=>"010101110",
  21710=>"110111011",
  21711=>"101011000",
  21712=>"011001001",
  21713=>"111100100",
  21714=>"001000101",
  21715=>"011001001",
  21716=>"001001110",
  21717=>"010001010",
  21718=>"010010000",
  21719=>"100110101",
  21720=>"100100010",
  21721=>"100001000",
  21722=>"011001001",
  21723=>"110100101",
  21724=>"001111100",
  21725=>"001111000",
  21726=>"010010001",
  21727=>"100001111",
  21728=>"110011001",
  21729=>"110101111",
  21730=>"011101000",
  21731=>"001100001",
  21732=>"001110111",
  21733=>"111011011",
  21734=>"110000111",
  21735=>"011000111",
  21736=>"011110111",
  21737=>"010111111",
  21738=>"111101101",
  21739=>"010110010",
  21740=>"000010111",
  21741=>"011011011",
  21742=>"101000000",
  21743=>"110000000",
  21744=>"011010100",
  21745=>"101111011",
  21746=>"011011001",
  21747=>"111010110",
  21748=>"110111111",
  21749=>"010101111",
  21750=>"101101000",
  21751=>"110110001",
  21752=>"101000101",
  21753=>"010101111",
  21754=>"000110011",
  21755=>"010010101",
  21756=>"111010011",
  21757=>"101101010",
  21758=>"010101000",
  21759=>"010010000",
  21760=>"001001101",
  21761=>"111111111",
  21762=>"000010111",
  21763=>"010010111",
  21764=>"110101010",
  21765=>"000101001",
  21766=>"001100110",
  21767=>"011101010",
  21768=>"101000000",
  21769=>"000011111",
  21770=>"000001001",
  21771=>"100100011",
  21772=>"111000001",
  21773=>"100101001",
  21774=>"100001010",
  21775=>"100000111",
  21776=>"110110001",
  21777=>"111110110",
  21778=>"000000001",
  21779=>"000000011",
  21780=>"110111110",
  21781=>"001110110",
  21782=>"111101011",
  21783=>"011101111",
  21784=>"110011100",
  21785=>"101000100",
  21786=>"001011101",
  21787=>"001000001",
  21788=>"011011011",
  21789=>"000010011",
  21790=>"110011111",
  21791=>"000000010",
  21792=>"011100111",
  21793=>"000011000",
  21794=>"010111111",
  21795=>"011000001",
  21796=>"010001101",
  21797=>"110010110",
  21798=>"001111000",
  21799=>"000010111",
  21800=>"000100100",
  21801=>"010011010",
  21802=>"100011110",
  21803=>"101101000",
  21804=>"100000010",
  21805=>"110000111",
  21806=>"000010101",
  21807=>"100100000",
  21808=>"000100100",
  21809=>"001100011",
  21810=>"111101111",
  21811=>"101010001",
  21812=>"000010010",
  21813=>"010000001",
  21814=>"001101001",
  21815=>"101000000",
  21816=>"100010011",
  21817=>"110111111",
  21818=>"111010000",
  21819=>"010011010",
  21820=>"010001111",
  21821=>"000100101",
  21822=>"000010101",
  21823=>"001110100",
  21824=>"110011010",
  21825=>"010001001",
  21826=>"111011111",
  21827=>"001011110",
  21828=>"100110110",
  21829=>"010100000",
  21830=>"111011011",
  21831=>"101011000",
  21832=>"011101010",
  21833=>"000111100",
  21834=>"001110011",
  21835=>"000001000",
  21836=>"100111101",
  21837=>"010001000",
  21838=>"110110111",
  21839=>"001111110",
  21840=>"000100111",
  21841=>"111100110",
  21842=>"101110001",
  21843=>"011011100",
  21844=>"000010011",
  21845=>"111110110",
  21846=>"000000010",
  21847=>"001000110",
  21848=>"001010101",
  21849=>"111101010",
  21850=>"101100101",
  21851=>"101101000",
  21852=>"100010111",
  21853=>"111111101",
  21854=>"110100100",
  21855=>"001110000",
  21856=>"010100001",
  21857=>"100000111",
  21858=>"111101011",
  21859=>"010100000",
  21860=>"000001010",
  21861=>"111010100",
  21862=>"101111100",
  21863=>"010011101",
  21864=>"111101010",
  21865=>"000001000",
  21866=>"101101011",
  21867=>"100100001",
  21868=>"011110111",
  21869=>"111101010",
  21870=>"011000011",
  21871=>"111010100",
  21872=>"001010111",
  21873=>"110111110",
  21874=>"000111100",
  21875=>"011001100",
  21876=>"001111010",
  21877=>"111010010",
  21878=>"110011110",
  21879=>"010110000",
  21880=>"010111111",
  21881=>"011010111",
  21882=>"111110011",
  21883=>"100110001",
  21884=>"111011100",
  21885=>"111100011",
  21886=>"011001100",
  21887=>"110100011",
  21888=>"100101101",
  21889=>"101111100",
  21890=>"001000111",
  21891=>"100101101",
  21892=>"011010010",
  21893=>"101100111",
  21894=>"100111100",
  21895=>"101011010",
  21896=>"111111010",
  21897=>"101011111",
  21898=>"101110001",
  21899=>"100000011",
  21900=>"100010010",
  21901=>"011101101",
  21902=>"101001000",
  21903=>"100100100",
  21904=>"000001010",
  21905=>"000000001",
  21906=>"010110101",
  21907=>"010010000",
  21908=>"000001010",
  21909=>"100100111",
  21910=>"011000010",
  21911=>"101010110",
  21912=>"001001110",
  21913=>"110000000",
  21914=>"010101110",
  21915=>"100001101",
  21916=>"111011001",
  21917=>"100011000",
  21918=>"101001100",
  21919=>"100101001",
  21920=>"011000001",
  21921=>"000010110",
  21922=>"001101110",
  21923=>"111010000",
  21924=>"001000101",
  21925=>"100011101",
  21926=>"001000010",
  21927=>"100100111",
  21928=>"110110011",
  21929=>"111111110",
  21930=>"000100000",
  21931=>"111101110",
  21932=>"110001101",
  21933=>"110101000",
  21934=>"001010100",
  21935=>"111111000",
  21936=>"101110100",
  21937=>"111111101",
  21938=>"110101100",
  21939=>"111111000",
  21940=>"101010100",
  21941=>"110110111",
  21942=>"100011110",
  21943=>"110010111",
  21944=>"000001110",
  21945=>"001111110",
  21946=>"110001110",
  21947=>"100111101",
  21948=>"101000011",
  21949=>"111101111",
  21950=>"100001111",
  21951=>"011001010",
  21952=>"011010100",
  21953=>"110000010",
  21954=>"000110111",
  21955=>"010010011",
  21956=>"011000010",
  21957=>"101001000",
  21958=>"110010100",
  21959=>"010101100",
  21960=>"000100001",
  21961=>"000101011",
  21962=>"010011010",
  21963=>"011100110",
  21964=>"100011110",
  21965=>"001001110",
  21966=>"100101001",
  21967=>"011111011",
  21968=>"100111100",
  21969=>"101011000",
  21970=>"010110101",
  21971=>"000101100",
  21972=>"111111010",
  21973=>"011011110",
  21974=>"101111010",
  21975=>"000000111",
  21976=>"010000000",
  21977=>"001100011",
  21978=>"011000000",
  21979=>"001101010",
  21980=>"001111100",
  21981=>"111111010",
  21982=>"111001000",
  21983=>"000010100",
  21984=>"010111110",
  21985=>"001011111",
  21986=>"111110101",
  21987=>"010000101",
  21988=>"000000010",
  21989=>"110101111",
  21990=>"110111000",
  21991=>"010001010",
  21992=>"110111010",
  21993=>"000101001",
  21994=>"000000100",
  21995=>"111011111",
  21996=>"010110110",
  21997=>"010111100",
  21998=>"100000100",
  21999=>"101111000",
  22000=>"000100010",
  22001=>"010011111",
  22002=>"010000101",
  22003=>"000000101",
  22004=>"010000000",
  22005=>"110111101",
  22006=>"100100011",
  22007=>"111010010",
  22008=>"000100010",
  22009=>"100101101",
  22010=>"001111000",
  22011=>"111001111",
  22012=>"001010010",
  22013=>"011011100",
  22014=>"111000110",
  22015=>"100110111",
  22016=>"100000111",
  22017=>"111001100",
  22018=>"111110100",
  22019=>"111110001",
  22020=>"010011101",
  22021=>"000111110",
  22022=>"001001000",
  22023=>"010000001",
  22024=>"000011011",
  22025=>"011111000",
  22026=>"101011111",
  22027=>"101100000",
  22028=>"110101101",
  22029=>"101001100",
  22030=>"000100100",
  22031=>"011011001",
  22032=>"000111001",
  22033=>"011101110",
  22034=>"111011101",
  22035=>"111110110",
  22036=>"010000010",
  22037=>"100101001",
  22038=>"101000100",
  22039=>"011101001",
  22040=>"111010111",
  22041=>"111001010",
  22042=>"111010001",
  22043=>"010010100",
  22044=>"010101000",
  22045=>"010101111",
  22046=>"000101100",
  22047=>"010110110",
  22048=>"011101111",
  22049=>"001101101",
  22050=>"001011000",
  22051=>"000110010",
  22052=>"100111110",
  22053=>"000111111",
  22054=>"010001000",
  22055=>"001101000",
  22056=>"011000000",
  22057=>"110101100",
  22058=>"000001000",
  22059=>"101001011",
  22060=>"111011000",
  22061=>"011000101",
  22062=>"101101110",
  22063=>"001101100",
  22064=>"001111001",
  22065=>"000011111",
  22066=>"101001011",
  22067=>"110011100",
  22068=>"000111000",
  22069=>"011010101",
  22070=>"111101101",
  22071=>"010001001",
  22072=>"101110101",
  22073=>"010011101",
  22074=>"010000011",
  22075=>"101001111",
  22076=>"011111000",
  22077=>"111111101",
  22078=>"001111001",
  22079=>"000100000",
  22080=>"000001101",
  22081=>"001101001",
  22082=>"110010000",
  22083=>"111110000",
  22084=>"111100000",
  22085=>"010000010",
  22086=>"000110010",
  22087=>"010100001",
  22088=>"100010011",
  22089=>"000110111",
  22090=>"101110101",
  22091=>"011110000",
  22092=>"000100001",
  22093=>"011001100",
  22094=>"010110110",
  22095=>"000011011",
  22096=>"011000110",
  22097=>"010010011",
  22098=>"010011010",
  22099=>"001111101",
  22100=>"000110101",
  22101=>"100110111",
  22102=>"001111110",
  22103=>"000011100",
  22104=>"100110011",
  22105=>"000011100",
  22106=>"011000001",
  22107=>"110100011",
  22108=>"011011110",
  22109=>"011010010",
  22110=>"100110110",
  22111=>"101100010",
  22112=>"000111000",
  22113=>"111111111",
  22114=>"100001010",
  22115=>"001100111",
  22116=>"010011010",
  22117=>"110011111",
  22118=>"000110011",
  22119=>"100110100",
  22120=>"100001001",
  22121=>"101000000",
  22122=>"111000111",
  22123=>"010001011",
  22124=>"100001001",
  22125=>"111010111",
  22126=>"111110010",
  22127=>"111111101",
  22128=>"000111110",
  22129=>"110101000",
  22130=>"001101100",
  22131=>"111011111",
  22132=>"100000011",
  22133=>"011001101",
  22134=>"000100110",
  22135=>"110000110",
  22136=>"110011000",
  22137=>"100101110",
  22138=>"010000100",
  22139=>"101010000",
  22140=>"000101000",
  22141=>"110000010",
  22142=>"100100000",
  22143=>"111101010",
  22144=>"010010110",
  22145=>"111010011",
  22146=>"000001101",
  22147=>"100000011",
  22148=>"000110010",
  22149=>"101001011",
  22150=>"010011111",
  22151=>"100110000",
  22152=>"100100001",
  22153=>"010011000",
  22154=>"110011110",
  22155=>"110001011",
  22156=>"100001001",
  22157=>"101011000",
  22158=>"110011010",
  22159=>"000011101",
  22160=>"001001001",
  22161=>"100011010",
  22162=>"111111111",
  22163=>"011000001",
  22164=>"011110111",
  22165=>"101011001",
  22166=>"011100010",
  22167=>"110010100",
  22168=>"010110101",
  22169=>"001011100",
  22170=>"111100101",
  22171=>"010111111",
  22172=>"001100001",
  22173=>"001001101",
  22174=>"001001011",
  22175=>"011100111",
  22176=>"110110101",
  22177=>"011100100",
  22178=>"000010100",
  22179=>"000100110",
  22180=>"010110111",
  22181=>"100011010",
  22182=>"011010010",
  22183=>"010111110",
  22184=>"000011110",
  22185=>"001111101",
  22186=>"010001001",
  22187=>"001000111",
  22188=>"100111111",
  22189=>"111011001",
  22190=>"111111010",
  22191=>"111110101",
  22192=>"001001011",
  22193=>"111110001",
  22194=>"001001100",
  22195=>"111110111",
  22196=>"111111010",
  22197=>"100101000",
  22198=>"101000111",
  22199=>"010010011",
  22200=>"101001011",
  22201=>"001011101",
  22202=>"111111111",
  22203=>"100111011",
  22204=>"000110100",
  22205=>"111110100",
  22206=>"001110101",
  22207=>"100001110",
  22208=>"111000110",
  22209=>"000000100",
  22210=>"110011111",
  22211=>"000100000",
  22212=>"100100000",
  22213=>"100100111",
  22214=>"000111110",
  22215=>"001011110",
  22216=>"101100110",
  22217=>"101010110",
  22218=>"110100000",
  22219=>"000000000",
  22220=>"000000011",
  22221=>"111100101",
  22222=>"101011000",
  22223=>"101111110",
  22224=>"001111111",
  22225=>"100001011",
  22226=>"101010101",
  22227=>"101111110",
  22228=>"010111100",
  22229=>"010010000",
  22230=>"111110011",
  22231=>"110010010",
  22232=>"000110101",
  22233=>"101011111",
  22234=>"011111110",
  22235=>"111100000",
  22236=>"010000011",
  22237=>"101010001",
  22238=>"111011011",
  22239=>"000010111",
  22240=>"101010101",
  22241=>"001101111",
  22242=>"001001000",
  22243=>"100000000",
  22244=>"100001000",
  22245=>"111100101",
  22246=>"001001010",
  22247=>"110110001",
  22248=>"001001111",
  22249=>"111000100",
  22250=>"001111010",
  22251=>"101111001",
  22252=>"010111011",
  22253=>"111110110",
  22254=>"011100001",
  22255=>"000011111",
  22256=>"000010011",
  22257=>"011000011",
  22258=>"010011010",
  22259=>"000011101",
  22260=>"100111111",
  22261=>"001001010",
  22262=>"010111001",
  22263=>"001100111",
  22264=>"101101000",
  22265=>"111001010",
  22266=>"001111111",
  22267=>"100001010",
  22268=>"110011010",
  22269=>"101000111",
  22270=>"000001100",
  22271=>"001101011",
  22272=>"011011001",
  22273=>"000001111",
  22274=>"000011010",
  22275=>"001101001",
  22276=>"101100010",
  22277=>"010010100",
  22278=>"001111001",
  22279=>"010000100",
  22280=>"000100010",
  22281=>"001110111",
  22282=>"000001010",
  22283=>"100100100",
  22284=>"110000010",
  22285=>"001000101",
  22286=>"000100101",
  22287=>"000000010",
  22288=>"011101111",
  22289=>"100000011",
  22290=>"011011101",
  22291=>"110010000",
  22292=>"011001000",
  22293=>"110011000",
  22294=>"101010100",
  22295=>"000110111",
  22296=>"001011100",
  22297=>"000101011",
  22298=>"000010111",
  22299=>"001111101",
  22300=>"000111001",
  22301=>"100000001",
  22302=>"010001011",
  22303=>"100110101",
  22304=>"001101100",
  22305=>"010000000",
  22306=>"110001000",
  22307=>"110011101",
  22308=>"100011010",
  22309=>"111010001",
  22310=>"101010100",
  22311=>"101010011",
  22312=>"000011110",
  22313=>"100011001",
  22314=>"001011011",
  22315=>"001110011",
  22316=>"111010000",
  22317=>"100101100",
  22318=>"111011010",
  22319=>"010001001",
  22320=>"001101111",
  22321=>"000101010",
  22322=>"000000000",
  22323=>"000010000",
  22324=>"010011110",
  22325=>"001001011",
  22326=>"100111101",
  22327=>"010011011",
  22328=>"000011000",
  22329=>"111100010",
  22330=>"110111100",
  22331=>"100111001",
  22332=>"011000001",
  22333=>"000100100",
  22334=>"000001111",
  22335=>"000011101",
  22336=>"001100001",
  22337=>"001001110",
  22338=>"111000101",
  22339=>"111100100",
  22340=>"010011110",
  22341=>"100101111",
  22342=>"101111011",
  22343=>"001011110",
  22344=>"110011011",
  22345=>"100101110",
  22346=>"000100100",
  22347=>"010110111",
  22348=>"001000110",
  22349=>"000011001",
  22350=>"000010001",
  22351=>"001010100",
  22352=>"000110010",
  22353=>"111011111",
  22354=>"110100000",
  22355=>"001001000",
  22356=>"001001010",
  22357=>"110101110",
  22358=>"100011101",
  22359=>"100100110",
  22360=>"010110000",
  22361=>"100100000",
  22362=>"100111110",
  22363=>"010100101",
  22364=>"000011011",
  22365=>"101100111",
  22366=>"111100100",
  22367=>"110100010",
  22368=>"110010010",
  22369=>"000000110",
  22370=>"011011011",
  22371=>"000110000",
  22372=>"010100110",
  22373=>"111011011",
  22374=>"000110011",
  22375=>"101111011",
  22376=>"000011001",
  22377=>"110111111",
  22378=>"010100010",
  22379=>"011011011",
  22380=>"001110000",
  22381=>"100010001",
  22382=>"010011111",
  22383=>"101011111",
  22384=>"011000010",
  22385=>"001101000",
  22386=>"001110011",
  22387=>"110010000",
  22388=>"000010111",
  22389=>"010010011",
  22390=>"111010000",
  22391=>"011100000",
  22392=>"011001001",
  22393=>"000010100",
  22394=>"000011110",
  22395=>"010000000",
  22396=>"101010111",
  22397=>"110111000",
  22398=>"010000100",
  22399=>"101110101",
  22400=>"101110110",
  22401=>"000000100",
  22402=>"110000101",
  22403=>"101110011",
  22404=>"101101000",
  22405=>"010010111",
  22406=>"010110101",
  22407=>"110111010",
  22408=>"010001111",
  22409=>"100110111",
  22410=>"000000110",
  22411=>"100110100",
  22412=>"110110000",
  22413=>"011000110",
  22414=>"010010001",
  22415=>"100001011",
  22416=>"101001110",
  22417=>"000110101",
  22418=>"010100111",
  22419=>"111111110",
  22420=>"000001000",
  22421=>"111001100",
  22422=>"001110101",
  22423=>"110010000",
  22424=>"111111010",
  22425=>"111001100",
  22426=>"010010010",
  22427=>"110010010",
  22428=>"000010101",
  22429=>"011101000",
  22430=>"011001110",
  22431=>"100000010",
  22432=>"000000000",
  22433=>"100110101",
  22434=>"010110111",
  22435=>"000010100",
  22436=>"001110111",
  22437=>"010110001",
  22438=>"000001110",
  22439=>"000110100",
  22440=>"101000000",
  22441=>"001011000",
  22442=>"110011111",
  22443=>"001000000",
  22444=>"000011011",
  22445=>"000101111",
  22446=>"001100010",
  22447=>"010101010",
  22448=>"000001001",
  22449=>"010111100",
  22450=>"110101000",
  22451=>"000010001",
  22452=>"000000111",
  22453=>"110110000",
  22454=>"110001111",
  22455=>"001100001",
  22456=>"001010011",
  22457=>"010111000",
  22458=>"011111110",
  22459=>"010100100",
  22460=>"100001101",
  22461=>"101001100",
  22462=>"101101101",
  22463=>"110011000",
  22464=>"010011010",
  22465=>"111011010",
  22466=>"111111100",
  22467=>"110000101",
  22468=>"111111100",
  22469=>"001101001",
  22470=>"101011001",
  22471=>"110001000",
  22472=>"110100010",
  22473=>"101000000",
  22474=>"111001010",
  22475=>"010010101",
  22476=>"111011101",
  22477=>"001111111",
  22478=>"000000111",
  22479=>"100101011",
  22480=>"101110011",
  22481=>"100100111",
  22482=>"100001111",
  22483=>"010001100",
  22484=>"001100111",
  22485=>"000001111",
  22486=>"011100001",
  22487=>"110010111",
  22488=>"111000101",
  22489=>"010111010",
  22490=>"110110110",
  22491=>"010010110",
  22492=>"000000001",
  22493=>"010000001",
  22494=>"011000000",
  22495=>"100101000",
  22496=>"111111011",
  22497=>"111001011",
  22498=>"101110111",
  22499=>"011010101",
  22500=>"001100011",
  22501=>"001011001",
  22502=>"111001011",
  22503=>"011111110",
  22504=>"010010110",
  22505=>"111001011",
  22506=>"010110001",
  22507=>"001100010",
  22508=>"110000100",
  22509=>"000000100",
  22510=>"101111001",
  22511=>"100101101",
  22512=>"001000111",
  22513=>"001000110",
  22514=>"000011010",
  22515=>"000100101",
  22516=>"010101101",
  22517=>"100101000",
  22518=>"011010110",
  22519=>"111100000",
  22520=>"011010110",
  22521=>"001001011",
  22522=>"000101010",
  22523=>"111000110",
  22524=>"010010001",
  22525=>"000011001",
  22526=>"010101010",
  22527=>"111101100",
  22528=>"101010101",
  22529=>"010110001",
  22530=>"010011011",
  22531=>"110100100",
  22532=>"010010011",
  22533=>"000111111",
  22534=>"010111110",
  22535=>"000010110",
  22536=>"101110101",
  22537=>"110000000",
  22538=>"100000111",
  22539=>"110101111",
  22540=>"011001001",
  22541=>"110011001",
  22542=>"011011110",
  22543=>"010001100",
  22544=>"110100100",
  22545=>"100100001",
  22546=>"011001001",
  22547=>"001000000",
  22548=>"001010101",
  22549=>"101101111",
  22550=>"000110000",
  22551=>"100000111",
  22552=>"000100111",
  22553=>"001011100",
  22554=>"010010110",
  22555=>"011010010",
  22556=>"110101010",
  22557=>"000110011",
  22558=>"001011010",
  22559=>"000111111",
  22560=>"000001100",
  22561=>"000110100",
  22562=>"110100100",
  22563=>"101010101",
  22564=>"011111110",
  22565=>"011000011",
  22566=>"111101110",
  22567=>"000110100",
  22568=>"001001011",
  22569=>"101110111",
  22570=>"010110110",
  22571=>"011011000",
  22572=>"101010110",
  22573=>"110101111",
  22574=>"010110100",
  22575=>"101101101",
  22576=>"101001010",
  22577=>"000111001",
  22578=>"100110100",
  22579=>"011111111",
  22580=>"100001001",
  22581=>"011101000",
  22582=>"000100010",
  22583=>"010010110",
  22584=>"100001100",
  22585=>"000111011",
  22586=>"101011010",
  22587=>"100110010",
  22588=>"011111111",
  22589=>"110110011",
  22590=>"000001101",
  22591=>"000110000",
  22592=>"001111110",
  22593=>"000110000",
  22594=>"111001011",
  22595=>"001000000",
  22596=>"011011100",
  22597=>"001001001",
  22598=>"101111101",
  22599=>"110101011",
  22600=>"010011010",
  22601=>"110110111",
  22602=>"001010000",
  22603=>"010010001",
  22604=>"101101011",
  22605=>"000010101",
  22606=>"000111010",
  22607=>"111111110",
  22608=>"111010110",
  22609=>"111111100",
  22610=>"001011110",
  22611=>"001010000",
  22612=>"010000100",
  22613=>"101100111",
  22614=>"000011101",
  22615=>"001001001",
  22616=>"010001111",
  22617=>"001101011",
  22618=>"101100111",
  22619=>"011100010",
  22620=>"100110000",
  22621=>"000100010",
  22622=>"000011111",
  22623=>"010001101",
  22624=>"111110000",
  22625=>"111101001",
  22626=>"000001010",
  22627=>"110101110",
  22628=>"010010100",
  22629=>"111001001",
  22630=>"110110011",
  22631=>"111011101",
  22632=>"111101000",
  22633=>"111101110",
  22634=>"010011011",
  22635=>"001110000",
  22636=>"001000010",
  22637=>"110000101",
  22638=>"110111101",
  22639=>"001010111",
  22640=>"000111110",
  22641=>"101110011",
  22642=>"101001000",
  22643=>"000010101",
  22644=>"010011101",
  22645=>"101010000",
  22646=>"100111110",
  22647=>"100000111",
  22648=>"110110000",
  22649=>"111101000",
  22650=>"111001111",
  22651=>"111111110",
  22652=>"000111001",
  22653=>"101101100",
  22654=>"010100101",
  22655=>"000001101",
  22656=>"001110100",
  22657=>"001000000",
  22658=>"000001000",
  22659=>"100010000",
  22660=>"001001111",
  22661=>"000111001",
  22662=>"100111001",
  22663=>"000110011",
  22664=>"011001011",
  22665=>"011001101",
  22666=>"001010110",
  22667=>"011000111",
  22668=>"000011110",
  22669=>"100011001",
  22670=>"110000000",
  22671=>"111010011",
  22672=>"101010100",
  22673=>"111000010",
  22674=>"000010111",
  22675=>"000101100",
  22676=>"101110111",
  22677=>"001111111",
  22678=>"111101000",
  22679=>"110011110",
  22680=>"000100101",
  22681=>"111101001",
  22682=>"001011100",
  22683=>"011101100",
  22684=>"001110000",
  22685=>"101101101",
  22686=>"001011000",
  22687=>"100001100",
  22688=>"000101010",
  22689=>"001010011",
  22690=>"111111111",
  22691=>"110010101",
  22692=>"010110111",
  22693=>"011010100",
  22694=>"010011010",
  22695=>"111101110",
  22696=>"100111000",
  22697=>"111100101",
  22698=>"111000010",
  22699=>"100101110",
  22700=>"101011111",
  22701=>"101100010",
  22702=>"011100000",
  22703=>"110011111",
  22704=>"000100111",
  22705=>"111110010",
  22706=>"010110111",
  22707=>"000001011",
  22708=>"111101011",
  22709=>"100110001",
  22710=>"101101011",
  22711=>"110110000",
  22712=>"010100001",
  22713=>"000001110",
  22714=>"111011110",
  22715=>"011101101",
  22716=>"001011011",
  22717=>"100100010",
  22718=>"011011001",
  22719=>"101000001",
  22720=>"111010100",
  22721=>"011010100",
  22722=>"000000011",
  22723=>"100111010",
  22724=>"000110010",
  22725=>"111011011",
  22726=>"100010000",
  22727=>"011010111",
  22728=>"011101010",
  22729=>"111110111",
  22730=>"100001011",
  22731=>"010011000",
  22732=>"101100111",
  22733=>"101110101",
  22734=>"000011111",
  22735=>"011111011",
  22736=>"110001101",
  22737=>"111001101",
  22738=>"000000111",
  22739=>"011001100",
  22740=>"001100101",
  22741=>"011111001",
  22742=>"001110111",
  22743=>"111110010",
  22744=>"100000001",
  22745=>"101110010",
  22746=>"000110110",
  22747=>"101000101",
  22748=>"011110111",
  22749=>"110001001",
  22750=>"011010011",
  22751=>"110001100",
  22752=>"111100001",
  22753=>"110111111",
  22754=>"001100010",
  22755=>"001001010",
  22756=>"110110111",
  22757=>"101011001",
  22758=>"111101110",
  22759=>"010010101",
  22760=>"111101010",
  22761=>"111100001",
  22762=>"010110110",
  22763=>"001101001",
  22764=>"111001111",
  22765=>"101001111",
  22766=>"000001001",
  22767=>"000010000",
  22768=>"010001001",
  22769=>"000100000",
  22770=>"010010100",
  22771=>"100001000",
  22772=>"000001100",
  22773=>"000000000",
  22774=>"100001011",
  22775=>"110001010",
  22776=>"001010000",
  22777=>"000001100",
  22778=>"111000111",
  22779=>"001000010",
  22780=>"000001010",
  22781=>"010110110",
  22782=>"001001110",
  22783=>"010000110",
  22784=>"111111110",
  22785=>"001011111",
  22786=>"101110111",
  22787=>"110010111",
  22788=>"111111011",
  22789=>"000001110",
  22790=>"000111001",
  22791=>"010111100",
  22792=>"001110011",
  22793=>"100010001",
  22794=>"001101000",
  22795=>"101100111",
  22796=>"100001001",
  22797=>"000001101",
  22798=>"101110110",
  22799=>"000010000",
  22800=>"110110010",
  22801=>"010010000",
  22802=>"101110111",
  22803=>"110011100",
  22804=>"100010101",
  22805=>"010000001",
  22806=>"111110101",
  22807=>"010011101",
  22808=>"110111100",
  22809=>"010100010",
  22810=>"100110001",
  22811=>"111001000",
  22812=>"000011110",
  22813=>"001000110",
  22814=>"110111100",
  22815=>"011001111",
  22816=>"001001001",
  22817=>"110110101",
  22818=>"011101111",
  22819=>"110000001",
  22820=>"011101011",
  22821=>"111010011",
  22822=>"101001001",
  22823=>"110100110",
  22824=>"001110010",
  22825=>"000110111",
  22826=>"001011111",
  22827=>"001110101",
  22828=>"011111101",
  22829=>"010100110",
  22830=>"001000011",
  22831=>"011001110",
  22832=>"101011101",
  22833=>"111010110",
  22834=>"010101101",
  22835=>"010110011",
  22836=>"100100000",
  22837=>"001101101",
  22838=>"101111000",
  22839=>"010010000",
  22840=>"001000000",
  22841=>"001001011",
  22842=>"111001010",
  22843=>"011010010",
  22844=>"001000010",
  22845=>"100000010",
  22846=>"111100110",
  22847=>"111011100",
  22848=>"000101110",
  22849=>"111010010",
  22850=>"101001011",
  22851=>"011110000",
  22852=>"000000011",
  22853=>"101010100",
  22854=>"000101110",
  22855=>"111000000",
  22856=>"110110011",
  22857=>"000010010",
  22858=>"001101111",
  22859=>"100011000",
  22860=>"011000000",
  22861=>"001011011",
  22862=>"000000000",
  22863=>"101110111",
  22864=>"001000000",
  22865=>"100111111",
  22866=>"001010100",
  22867=>"000111100",
  22868=>"100001010",
  22869=>"000111110",
  22870=>"011110101",
  22871=>"001100101",
  22872=>"010111111",
  22873=>"000100100",
  22874=>"100111101",
  22875=>"000101000",
  22876=>"000110001",
  22877=>"111111001",
  22878=>"001101100",
  22879=>"100000010",
  22880=>"100100101",
  22881=>"010011010",
  22882=>"010010110",
  22883=>"001111110",
  22884=>"100110000",
  22885=>"110111000",
  22886=>"000011010",
  22887=>"110101010",
  22888=>"100011111",
  22889=>"011100001",
  22890=>"000011101",
  22891=>"001111101",
  22892=>"101011010",
  22893=>"010101011",
  22894=>"001111101",
  22895=>"001000101",
  22896=>"000110010",
  22897=>"111011111",
  22898=>"101010000",
  22899=>"010000010",
  22900=>"001011110",
  22901=>"110010000",
  22902=>"000000101",
  22903=>"111101000",
  22904=>"011100100",
  22905=>"110010000",
  22906=>"111011110",
  22907=>"001100000",
  22908=>"110110110",
  22909=>"100001010",
  22910=>"110100111",
  22911=>"101100001",
  22912=>"000100100",
  22913=>"110011111",
  22914=>"100011100",
  22915=>"010010101",
  22916=>"100110101",
  22917=>"111111011",
  22918=>"011111110",
  22919=>"101011111",
  22920=>"001011110",
  22921=>"111100110",
  22922=>"011100110",
  22923=>"111010011",
  22924=>"111011110",
  22925=>"111010011",
  22926=>"000111001",
  22927=>"101100000",
  22928=>"111110111",
  22929=>"001011100",
  22930=>"110000110",
  22931=>"001001100",
  22932=>"010011000",
  22933=>"000111000",
  22934=>"101000010",
  22935=>"100111101",
  22936=>"010000101",
  22937=>"011100111",
  22938=>"101101110",
  22939=>"101110111",
  22940=>"100111111",
  22941=>"001111011",
  22942=>"100001011",
  22943=>"111111101",
  22944=>"001001111",
  22945=>"001000010",
  22946=>"010000011",
  22947=>"101000010",
  22948=>"111110111",
  22949=>"101001011",
  22950=>"010010000",
  22951=>"001100011",
  22952=>"000010111",
  22953=>"000010011",
  22954=>"000001001",
  22955=>"100000010",
  22956=>"000010011",
  22957=>"001100111",
  22958=>"011100011",
  22959=>"101110111",
  22960=>"001110100",
  22961=>"111000000",
  22962=>"001110000",
  22963=>"011001011",
  22964=>"011000011",
  22965=>"011100001",
  22966=>"100111101",
  22967=>"000010010",
  22968=>"100000001",
  22969=>"000101011",
  22970=>"001100100",
  22971=>"101000100",
  22972=>"011110111",
  22973=>"011100101",
  22974=>"001001011",
  22975=>"000101000",
  22976=>"000010010",
  22977=>"100111111",
  22978=>"010111100",
  22979=>"000101111",
  22980=>"111000001",
  22981=>"010110100",
  22982=>"001010100",
  22983=>"100000101",
  22984=>"111111111",
  22985=>"000000001",
  22986=>"000111101",
  22987=>"000101010",
  22988=>"000110110",
  22989=>"101101101",
  22990=>"000100110",
  22991=>"100001010",
  22992=>"011010000",
  22993=>"011101101",
  22994=>"000011010",
  22995=>"010001010",
  22996=>"000100001",
  22997=>"100100100",
  22998=>"010010110",
  22999=>"110001110",
  23000=>"000010001",
  23001=>"010101111",
  23002=>"111101001",
  23003=>"100000111",
  23004=>"111101111",
  23005=>"110001010",
  23006=>"101001100",
  23007=>"110110000",
  23008=>"111110100",
  23009=>"100001111",
  23010=>"110101010",
  23011=>"001001011",
  23012=>"000100001",
  23013=>"001111000",
  23014=>"100000010",
  23015=>"011001101",
  23016=>"010110111",
  23017=>"110110111",
  23018=>"000100100",
  23019=>"010110000",
  23020=>"000001111",
  23021=>"111000111",
  23022=>"101111111",
  23023=>"110001011",
  23024=>"001101111",
  23025=>"000111010",
  23026=>"100101000",
  23027=>"101011010",
  23028=>"110011100",
  23029=>"101000110",
  23030=>"011010000",
  23031=>"000001101",
  23032=>"000111001",
  23033=>"111000110",
  23034=>"101101011",
  23035=>"010101010",
  23036=>"101010001",
  23037=>"110001000",
  23038=>"010011010",
  23039=>"101110000",
  23040=>"010101000",
  23041=>"011000000",
  23042=>"111011010",
  23043=>"011000001",
  23044=>"000100010",
  23045=>"000101101",
  23046=>"110010100",
  23047=>"110111110",
  23048=>"110100000",
  23049=>"011010111",
  23050=>"110011001",
  23051=>"010101000",
  23052=>"100111110",
  23053=>"000101000",
  23054=>"010100110",
  23055=>"100010011",
  23056=>"010011000",
  23057=>"100010000",
  23058=>"100100100",
  23059=>"110011111",
  23060=>"110101000",
  23061=>"111000000",
  23062=>"111100100",
  23063=>"100010011",
  23064=>"100011100",
  23065=>"001010001",
  23066=>"001110110",
  23067=>"001111101",
  23068=>"101100011",
  23069=>"100000100",
  23070=>"011111001",
  23071=>"000010011",
  23072=>"010110001",
  23073=>"000000010",
  23074=>"001000010",
  23075=>"100000100",
  23076=>"100111111",
  23077=>"000001010",
  23078=>"000000011",
  23079=>"000101100",
  23080=>"000010100",
  23081=>"001100010",
  23082=>"011110010",
  23083=>"001010101",
  23084=>"011000100",
  23085=>"000011011",
  23086=>"001000010",
  23087=>"000000111",
  23088=>"111000010",
  23089=>"011111000",
  23090=>"101000001",
  23091=>"101100011",
  23092=>"100110000",
  23093=>"000001000",
  23094=>"100111010",
  23095=>"011100011",
  23096=>"011001110",
  23097=>"011101011",
  23098=>"110110111",
  23099=>"110010100",
  23100=>"000010011",
  23101=>"110100010",
  23102=>"000001001",
  23103=>"101101010",
  23104=>"110111010",
  23105=>"111011001",
  23106=>"111101000",
  23107=>"010110011",
  23108=>"110100100",
  23109=>"010100101",
  23110=>"001111110",
  23111=>"100110010",
  23112=>"010001100",
  23113=>"110001011",
  23114=>"011011001",
  23115=>"101010000",
  23116=>"010110100",
  23117=>"100001010",
  23118=>"001010100",
  23119=>"001110000",
  23120=>"101111011",
  23121=>"111000000",
  23122=>"101110001",
  23123=>"010100001",
  23124=>"100100100",
  23125=>"000011100",
  23126=>"101100101",
  23127=>"110110111",
  23128=>"001000111",
  23129=>"000110001",
  23130=>"101111000",
  23131=>"001010101",
  23132=>"100100001",
  23133=>"000100000",
  23134=>"000101100",
  23135=>"100100110",
  23136=>"011101000",
  23137=>"011101010",
  23138=>"110011111",
  23139=>"010000001",
  23140=>"101110001",
  23141=>"100101000",
  23142=>"110000000",
  23143=>"100000000",
  23144=>"010110010",
  23145=>"010001011",
  23146=>"000011101",
  23147=>"100110011",
  23148=>"000110101",
  23149=>"110010100",
  23150=>"000101010",
  23151=>"101011100",
  23152=>"000101001",
  23153=>"000000111",
  23154=>"000011001",
  23155=>"111000111",
  23156=>"111101110",
  23157=>"001001101",
  23158=>"101111101",
  23159=>"111100111",
  23160=>"100011110",
  23161=>"110110010",
  23162=>"100111000",
  23163=>"111010110",
  23164=>"010111101",
  23165=>"000100101",
  23166=>"100000100",
  23167=>"101001010",
  23168=>"111010101",
  23169=>"101100100",
  23170=>"000000001",
  23171=>"101000100",
  23172=>"000101110",
  23173=>"111111011",
  23174=>"011010010",
  23175=>"110101010",
  23176=>"000001011",
  23177=>"011000101",
  23178=>"011001111",
  23179=>"110100100",
  23180=>"111011110",
  23181=>"111111101",
  23182=>"011110010",
  23183=>"011101110",
  23184=>"010110001",
  23185=>"110010111",
  23186=>"001010101",
  23187=>"011100010",
  23188=>"001011000",
  23189=>"000000101",
  23190=>"001111010",
  23191=>"111001001",
  23192=>"110001001",
  23193=>"000101101",
  23194=>"110100111",
  23195=>"011001000",
  23196=>"111110110",
  23197=>"111011110",
  23198=>"111011000",
  23199=>"101000000",
  23200=>"001110111",
  23201=>"001110101",
  23202=>"001000010",
  23203=>"110100111",
  23204=>"110011100",
  23205=>"111100110",
  23206=>"000011100",
  23207=>"101101000",
  23208=>"101111011",
  23209=>"001110101",
  23210=>"001100110",
  23211=>"011001011",
  23212=>"100110111",
  23213=>"100001001",
  23214=>"110101000",
  23215=>"010100011",
  23216=>"000010000",
  23217=>"100010100",
  23218=>"001010000",
  23219=>"110110010",
  23220=>"000100001",
  23221=>"110101110",
  23222=>"111010010",
  23223=>"010110111",
  23224=>"011000010",
  23225=>"110000111",
  23226=>"011001110",
  23227=>"111010000",
  23228=>"000001000",
  23229=>"011111101",
  23230=>"001100010",
  23231=>"100110010",
  23232=>"011011110",
  23233=>"011110001",
  23234=>"011011010",
  23235=>"110011101",
  23236=>"100110111",
  23237=>"110100111",
  23238=>"110011011",
  23239=>"001100011",
  23240=>"001001101",
  23241=>"110110111",
  23242=>"011010000",
  23243=>"010101100",
  23244=>"010001110",
  23245=>"101010000",
  23246=>"101111001",
  23247=>"110111000",
  23248=>"110000000",
  23249=>"101100101",
  23250=>"000001000",
  23251=>"001000001",
  23252=>"000111010",
  23253=>"000000101",
  23254=>"010110010",
  23255=>"111011101",
  23256=>"000110001",
  23257=>"111100111",
  23258=>"111010101",
  23259=>"111110100",
  23260=>"001110001",
  23261=>"010111001",
  23262=>"111110010",
  23263=>"100010110",
  23264=>"110010011",
  23265=>"101011001",
  23266=>"111100000",
  23267=>"010110001",
  23268=>"000011001",
  23269=>"001010111",
  23270=>"010100110",
  23271=>"111101000",
  23272=>"100100111",
  23273=>"000000010",
  23274=>"000101010",
  23275=>"100001110",
  23276=>"001000001",
  23277=>"010110101",
  23278=>"100101101",
  23279=>"000100101",
  23280=>"110010101",
  23281=>"011100010",
  23282=>"111000000",
  23283=>"100101000",
  23284=>"001100101",
  23285=>"001101001",
  23286=>"011010101",
  23287=>"110010011",
  23288=>"111110100",
  23289=>"111110110",
  23290=>"011000001",
  23291=>"111000001",
  23292=>"100100001",
  23293=>"100101010",
  23294=>"001010101",
  23295=>"000010000",
  23296=>"111001100",
  23297=>"101111111",
  23298=>"100111001",
  23299=>"000111000",
  23300=>"000010011",
  23301=>"000110100",
  23302=>"000110110",
  23303=>"100111010",
  23304=>"011011111",
  23305=>"000011011",
  23306=>"100000101",
  23307=>"001111110",
  23308=>"110110111",
  23309=>"110010000",
  23310=>"111001010",
  23311=>"010000010",
  23312=>"011100100",
  23313=>"010101010",
  23314=>"001111100",
  23315=>"010001010",
  23316=>"010000000",
  23317=>"010010010",
  23318=>"111001011",
  23319=>"100110011",
  23320=>"101101011",
  23321=>"100101000",
  23322=>"100110001",
  23323=>"011000001",
  23324=>"111001110",
  23325=>"000001110",
  23326=>"111001011",
  23327=>"111000110",
  23328=>"100100001",
  23329=>"110010100",
  23330=>"110001110",
  23331=>"110000111",
  23332=>"111011111",
  23333=>"111001110",
  23334=>"001100100",
  23335=>"010100111",
  23336=>"111011010",
  23337=>"001110001",
  23338=>"011110010",
  23339=>"000001100",
  23340=>"111110101",
  23341=>"000000010",
  23342=>"110101100",
  23343=>"101111111",
  23344=>"000001111",
  23345=>"000110110",
  23346=>"011101101",
  23347=>"000100101",
  23348=>"000000000",
  23349=>"111001011",
  23350=>"101001101",
  23351=>"001111000",
  23352=>"000100100",
  23353=>"100001010",
  23354=>"101100010",
  23355=>"100001000",
  23356=>"100111101",
  23357=>"000101100",
  23358=>"010000011",
  23359=>"000111111",
  23360=>"011000111",
  23361=>"111111110",
  23362=>"100110110",
  23363=>"101010111",
  23364=>"110101110",
  23365=>"010001011",
  23366=>"110101100",
  23367=>"000000110",
  23368=>"110111010",
  23369=>"110010011",
  23370=>"010011111",
  23371=>"001010010",
  23372=>"011101011",
  23373=>"000001010",
  23374=>"000011010",
  23375=>"101011100",
  23376=>"111011001",
  23377=>"001111111",
  23378=>"011110101",
  23379=>"100011011",
  23380=>"101100011",
  23381=>"110100011",
  23382=>"000110000",
  23383=>"000010111",
  23384=>"010110000",
  23385=>"100011010",
  23386=>"011001011",
  23387=>"010010111",
  23388=>"010011011",
  23389=>"100010011",
  23390=>"111110011",
  23391=>"101100110",
  23392=>"000000011",
  23393=>"001001100",
  23394=>"111110100",
  23395=>"110100000",
  23396=>"111110011",
  23397=>"100000101",
  23398=>"111101100",
  23399=>"001111111",
  23400=>"110111010",
  23401=>"000001110",
  23402=>"111011111",
  23403=>"110001001",
  23404=>"100101010",
  23405=>"111011101",
  23406=>"001000000",
  23407=>"000101000",
  23408=>"100101100",
  23409=>"010100101",
  23410=>"111010111",
  23411=>"011001101",
  23412=>"000101001",
  23413=>"110011001",
  23414=>"110111110",
  23415=>"001010010",
  23416=>"011001001",
  23417=>"100010100",
  23418=>"011001101",
  23419=>"010100000",
  23420=>"001000011",
  23421=>"100011101",
  23422=>"110100110",
  23423=>"010011110",
  23424=>"110101100",
  23425=>"000100111",
  23426=>"011110101",
  23427=>"100001010",
  23428=>"100001100",
  23429=>"000101011",
  23430=>"010011011",
  23431=>"101001001",
  23432=>"101101011",
  23433=>"100100111",
  23434=>"000100001",
  23435=>"000010010",
  23436=>"010111001",
  23437=>"000111000",
  23438=>"100010110",
  23439=>"001110011",
  23440=>"100100000",
  23441=>"011011101",
  23442=>"001100001",
  23443=>"100101010",
  23444=>"111011100",
  23445=>"000011101",
  23446=>"111011111",
  23447=>"111101101",
  23448=>"001011010",
  23449=>"111100110",
  23450=>"011000000",
  23451=>"111011001",
  23452=>"111010100",
  23453=>"000001001",
  23454=>"001101100",
  23455=>"101000111",
  23456=>"010001111",
  23457=>"111111001",
  23458=>"011000011",
  23459=>"000001001",
  23460=>"011001111",
  23461=>"001100111",
  23462=>"001110000",
  23463=>"010010110",
  23464=>"101100000",
  23465=>"000010100",
  23466=>"000000000",
  23467=>"011110100",
  23468=>"001111010",
  23469=>"111011111",
  23470=>"100010000",
  23471=>"010101100",
  23472=>"101011000",
  23473=>"110110011",
  23474=>"001101100",
  23475=>"000000000",
  23476=>"000100000",
  23477=>"110010011",
  23478=>"101100000",
  23479=>"110001000",
  23480=>"100011010",
  23481=>"001000011",
  23482=>"000011110",
  23483=>"000001100",
  23484=>"000001001",
  23485=>"100010010",
  23486=>"110010101",
  23487=>"011010101",
  23488=>"001110011",
  23489=>"101111100",
  23490=>"000100010",
  23491=>"110111000",
  23492=>"100111010",
  23493=>"010111000",
  23494=>"010111010",
  23495=>"111010100",
  23496=>"100000011",
  23497=>"000010000",
  23498=>"011011000",
  23499=>"111111011",
  23500=>"001010001",
  23501=>"100000011",
  23502=>"111000100",
  23503=>"110111001",
  23504=>"001000110",
  23505=>"001101000",
  23506=>"110110100",
  23507=>"110000010",
  23508=>"111111011",
  23509=>"111111110",
  23510=>"001010100",
  23511=>"000100001",
  23512=>"110000101",
  23513=>"110101110",
  23514=>"101001101",
  23515=>"111100100",
  23516=>"011100110",
  23517=>"101010100",
  23518=>"001010110",
  23519=>"110010101",
  23520=>"110011101",
  23521=>"101000001",
  23522=>"001110000",
  23523=>"110011011",
  23524=>"010001011",
  23525=>"000010100",
  23526=>"000000110",
  23527=>"110101111",
  23528=>"010001100",
  23529=>"011110100",
  23530=>"011110111",
  23531=>"000110001",
  23532=>"100111000",
  23533=>"000110001",
  23534=>"110000100",
  23535=>"000100100",
  23536=>"000101011",
  23537=>"001011100",
  23538=>"000110010",
  23539=>"111100010",
  23540=>"001100011",
  23541=>"100001010",
  23542=>"010111011",
  23543=>"101111100",
  23544=>"100101000",
  23545=>"000110100",
  23546=>"000100000",
  23547=>"111110011",
  23548=>"001000011",
  23549=>"100011100",
  23550=>"000100000",
  23551=>"111101010",
  23552=>"110101110",
  23553=>"001110001",
  23554=>"010010001",
  23555=>"010111110",
  23556=>"001010010",
  23557=>"011001110",
  23558=>"111000110",
  23559=>"100100100",
  23560=>"000010100",
  23561=>"010111010",
  23562=>"111100001",
  23563=>"001100110",
  23564=>"010100101",
  23565=>"111100011",
  23566=>"110010011",
  23567=>"111111001",
  23568=>"001110000",
  23569=>"110100110",
  23570=>"011010001",
  23571=>"100100010",
  23572=>"100010000",
  23573=>"110111000",
  23574=>"000011101",
  23575=>"111101010",
  23576=>"000110100",
  23577=>"100001110",
  23578=>"011110010",
  23579=>"011001101",
  23580=>"001011111",
  23581=>"000000000",
  23582=>"111101001",
  23583=>"010110101",
  23584=>"010011100",
  23585=>"110001110",
  23586=>"000000000",
  23587=>"010000000",
  23588=>"011011010",
  23589=>"011100001",
  23590=>"010100010",
  23591=>"011010100",
  23592=>"110101101",
  23593=>"100110111",
  23594=>"010100010",
  23595=>"101101111",
  23596=>"111111101",
  23597=>"100010010",
  23598=>"011101100",
  23599=>"000011001",
  23600=>"111010000",
  23601=>"001101011",
  23602=>"000010010",
  23603=>"100111000",
  23604=>"001011010",
  23605=>"101100111",
  23606=>"001011000",
  23607=>"010111101",
  23608=>"000100110",
  23609=>"111110011",
  23610=>"100010000",
  23611=>"000001001",
  23612=>"101100110",
  23613=>"100111100",
  23614=>"111001101",
  23615=>"101100010",
  23616=>"011100101",
  23617=>"000000010",
  23618=>"000111101",
  23619=>"101111100",
  23620=>"100111100",
  23621=>"111010101",
  23622=>"101001011",
  23623=>"110010010",
  23624=>"110000011",
  23625=>"000110100",
  23626=>"100000000",
  23627=>"111011110",
  23628=>"111001001",
  23629=>"111010111",
  23630=>"100001001",
  23631=>"110100010",
  23632=>"100000101",
  23633=>"011100010",
  23634=>"111011111",
  23635=>"101111001",
  23636=>"011101100",
  23637=>"100000100",
  23638=>"001010111",
  23639=>"001011010",
  23640=>"110011111",
  23641=>"001010011",
  23642=>"000010011",
  23643=>"011010111",
  23644=>"110011010",
  23645=>"000100000",
  23646=>"000001011",
  23647=>"000010001",
  23648=>"001101101",
  23649=>"111010001",
  23650=>"001111011",
  23651=>"000000101",
  23652=>"000001011",
  23653=>"110010101",
  23654=>"001100101",
  23655=>"001010010",
  23656=>"000011010",
  23657=>"000011010",
  23658=>"001110100",
  23659=>"110000011",
  23660=>"111000101",
  23661=>"010011011",
  23662=>"100111010",
  23663=>"111010110",
  23664=>"100101001",
  23665=>"000010001",
  23666=>"010010110",
  23667=>"011110101",
  23668=>"011100001",
  23669=>"000000111",
  23670=>"000010000",
  23671=>"101000000",
  23672=>"000011101",
  23673=>"001011101",
  23674=>"001011101",
  23675=>"101010110",
  23676=>"010001110",
  23677=>"100000000",
  23678=>"001100000",
  23679=>"100100000",
  23680=>"100111101",
  23681=>"111110000",
  23682=>"011101000",
  23683=>"000001011",
  23684=>"101110001",
  23685=>"010001110",
  23686=>"100111111",
  23687=>"000000110",
  23688=>"011100110",
  23689=>"100101100",
  23690=>"011000100",
  23691=>"001001000",
  23692=>"001110011",
  23693=>"110000110",
  23694=>"101110100",
  23695=>"101011111",
  23696=>"010010011",
  23697=>"010101000",
  23698=>"000110010",
  23699=>"111001100",
  23700=>"100011000",
  23701=>"011001101",
  23702=>"011001000",
  23703=>"100111001",
  23704=>"010000011",
  23705=>"110011001",
  23706=>"010000100",
  23707=>"000101101",
  23708=>"010010000",
  23709=>"010110000",
  23710=>"111100011",
  23711=>"101011110",
  23712=>"001000000",
  23713=>"100011000",
  23714=>"011010100",
  23715=>"100100001",
  23716=>"011011111",
  23717=>"111110111",
  23718=>"101010110",
  23719=>"111010101",
  23720=>"110100011",
  23721=>"000101100",
  23722=>"101010100",
  23723=>"001100011",
  23724=>"111111010",
  23725=>"111101011",
  23726=>"111011111",
  23727=>"001000100",
  23728=>"101110100",
  23729=>"111011111",
  23730=>"101110010",
  23731=>"100000100",
  23732=>"011001100",
  23733=>"000101111",
  23734=>"100101001",
  23735=>"101111101",
  23736=>"010010111",
  23737=>"001001100",
  23738=>"000001000",
  23739=>"111000110",
  23740=>"110011111",
  23741=>"101010111",
  23742=>"011111011",
  23743=>"101000011",
  23744=>"111110111",
  23745=>"011100011",
  23746=>"101000001",
  23747=>"000110000",
  23748=>"000001111",
  23749=>"000001111",
  23750=>"010101010",
  23751=>"111111111",
  23752=>"001110010",
  23753=>"001011101",
  23754=>"000011000",
  23755=>"110001000",
  23756=>"011010001",
  23757=>"010110010",
  23758=>"101101111",
  23759=>"010000100",
  23760=>"011100110",
  23761=>"001100000",
  23762=>"000011001",
  23763=>"100000110",
  23764=>"110000011",
  23765=>"001101111",
  23766=>"111011110",
  23767=>"000001101",
  23768=>"101111100",
  23769=>"100010111",
  23770=>"101110101",
  23771=>"100001001",
  23772=>"000010111",
  23773=>"110111000",
  23774=>"000100100",
  23775=>"110011000",
  23776=>"100010001",
  23777=>"111100011",
  23778=>"110101010",
  23779=>"000110101",
  23780=>"100000000",
  23781=>"000001010",
  23782=>"100000110",
  23783=>"000001011",
  23784=>"000011111",
  23785=>"011111001",
  23786=>"111001001",
  23787=>"110011001",
  23788=>"111101000",
  23789=>"001000111",
  23790=>"101110000",
  23791=>"011001001",
  23792=>"011101000",
  23793=>"111111001",
  23794=>"100000001",
  23795=>"101000000",
  23796=>"010000001",
  23797=>"101110110",
  23798=>"010010011",
  23799=>"101101101",
  23800=>"011111001",
  23801=>"100000011",
  23802=>"011101110",
  23803=>"001010101",
  23804=>"010000000",
  23805=>"111010010",
  23806=>"011000100",
  23807=>"110000101",
  23808=>"110001010",
  23809=>"100101101",
  23810=>"001001111",
  23811=>"100000111",
  23812=>"010010000",
  23813=>"001101101",
  23814=>"011010101",
  23815=>"110110001",
  23816=>"110010011",
  23817=>"000001111",
  23818=>"001110010",
  23819=>"110000110",
  23820=>"000100101",
  23821=>"101001000",
  23822=>"010000111",
  23823=>"001001001",
  23824=>"000000001",
  23825=>"010101101",
  23826=>"100101010",
  23827=>"010001011",
  23828=>"100001011",
  23829=>"010000101",
  23830=>"110111111",
  23831=>"010100111",
  23832=>"100101110",
  23833=>"010101110",
  23834=>"101000101",
  23835=>"101011100",
  23836=>"101000001",
  23837=>"001001100",
  23838=>"010111000",
  23839=>"010000100",
  23840=>"011110100",
  23841=>"101100001",
  23842=>"110010001",
  23843=>"001100100",
  23844=>"001011110",
  23845=>"001011001",
  23846=>"001001000",
  23847=>"101001001",
  23848=>"001111010",
  23849=>"111001000",
  23850=>"011100010",
  23851=>"011111001",
  23852=>"100000101",
  23853=>"000111101",
  23854=>"110010111",
  23855=>"011000100",
  23856=>"001111110",
  23857=>"011001100",
  23858=>"001100100",
  23859=>"011110111",
  23860=>"001010000",
  23861=>"100000101",
  23862=>"010101011",
  23863=>"000001110",
  23864=>"000011101",
  23865=>"010010010",
  23866=>"111001110",
  23867=>"011110100",
  23868=>"000011011",
  23869=>"001110001",
  23870=>"011001001",
  23871=>"001011001",
  23872=>"000011111",
  23873=>"001001111",
  23874=>"011101101",
  23875=>"111101000",
  23876=>"000101111",
  23877=>"001011111",
  23878=>"000011010",
  23879=>"000001011",
  23880=>"000111111",
  23881=>"111100100",
  23882=>"111111000",
  23883=>"100100000",
  23884=>"011010101",
  23885=>"101011111",
  23886=>"111010010",
  23887=>"101100001",
  23888=>"101101101",
  23889=>"000100101",
  23890=>"101011110",
  23891=>"100101011",
  23892=>"100011001",
  23893=>"011010010",
  23894=>"101100010",
  23895=>"110100001",
  23896=>"111000110",
  23897=>"011010000",
  23898=>"001001101",
  23899=>"100010010",
  23900=>"011011001",
  23901=>"000000110",
  23902=>"101001010",
  23903=>"000110100",
  23904=>"000010010",
  23905=>"111000111",
  23906=>"000010101",
  23907=>"100110110",
  23908=>"001001000",
  23909=>"111111011",
  23910=>"100010010",
  23911=>"110001010",
  23912=>"001000010",
  23913=>"011101101",
  23914=>"000011101",
  23915=>"011101000",
  23916=>"111011101",
  23917=>"100001111",
  23918=>"101010010",
  23919=>"001011000",
  23920=>"011011100",
  23921=>"111000110",
  23922=>"000110110",
  23923=>"010100000",
  23924=>"100100111",
  23925=>"000101100",
  23926=>"011001011",
  23927=>"111110110",
  23928=>"001000100",
  23929=>"101100000",
  23930=>"010010011",
  23931=>"010010100",
  23932=>"100010001",
  23933=>"010101011",
  23934=>"010101001",
  23935=>"101001010",
  23936=>"111101100",
  23937=>"000000001",
  23938=>"100001101",
  23939=>"111010101",
  23940=>"111101010",
  23941=>"100111110",
  23942=>"111011010",
  23943=>"010000110",
  23944=>"001111001",
  23945=>"011001010",
  23946=>"100111010",
  23947=>"010110110",
  23948=>"011000100",
  23949=>"111100110",
  23950=>"111101011",
  23951=>"000000000",
  23952=>"001100000",
  23953=>"100101110",
  23954=>"011100001",
  23955=>"010000110",
  23956=>"100111000",
  23957=>"010000001",
  23958=>"000110110",
  23959=>"010100111",
  23960=>"000101110",
  23961=>"010110011",
  23962=>"011000011",
  23963=>"100000111",
  23964=>"101000000",
  23965=>"111111111",
  23966=>"110110100",
  23967=>"001000100",
  23968=>"011001000",
  23969=>"111100100",
  23970=>"001001000",
  23971=>"100011110",
  23972=>"011010101",
  23973=>"100100010",
  23974=>"001110011",
  23975=>"010010101",
  23976=>"100110100",
  23977=>"010101100",
  23978=>"001000110",
  23979=>"100100101",
  23980=>"001100110",
  23981=>"001000110",
  23982=>"000001111",
  23983=>"010010000",
  23984=>"000101001",
  23985=>"000111011",
  23986=>"101111111",
  23987=>"101001101",
  23988=>"010000001",
  23989=>"001001001",
  23990=>"111111110",
  23991=>"000000010",
  23992=>"110101000",
  23993=>"000100011",
  23994=>"011000100",
  23995=>"101001011",
  23996=>"111100011",
  23997=>"000111011",
  23998=>"111100001",
  23999=>"110000000",
  24000=>"100000001",
  24001=>"001110111",
  24002=>"001101110",
  24003=>"111001001",
  24004=>"100101001",
  24005=>"101001001",
  24006=>"001100101",
  24007=>"111011100",
  24008=>"101110001",
  24009=>"101111001",
  24010=>"100001110",
  24011=>"101101111",
  24012=>"111001010",
  24013=>"000010011",
  24014=>"011100000",
  24015=>"001111011",
  24016=>"101000110",
  24017=>"001111100",
  24018=>"010000001",
  24019=>"100000001",
  24020=>"100101100",
  24021=>"100101010",
  24022=>"010001011",
  24023=>"011101000",
  24024=>"111111101",
  24025=>"100111011",
  24026=>"101100010",
  24027=>"011010101",
  24028=>"000111111",
  24029=>"011001001",
  24030=>"111011110",
  24031=>"000000000",
  24032=>"111001110",
  24033=>"000001100",
  24034=>"010111000",
  24035=>"100001000",
  24036=>"101100000",
  24037=>"001111001",
  24038=>"101100100",
  24039=>"101100000",
  24040=>"101011000",
  24041=>"100101010",
  24042=>"010101101",
  24043=>"110001110",
  24044=>"010110000",
  24045=>"010001011",
  24046=>"001001001",
  24047=>"100100000",
  24048=>"001100101",
  24049=>"010011010",
  24050=>"010000001",
  24051=>"101100110",
  24052=>"110010100",
  24053=>"101110010",
  24054=>"101100100",
  24055=>"110101011",
  24056=>"010011110",
  24057=>"100010100",
  24058=>"011100101",
  24059=>"000110010",
  24060=>"001010001",
  24061=>"100000111",
  24062=>"111110101",
  24063=>"010000010",
  24064=>"001000000",
  24065=>"010011100",
  24066=>"111000101",
  24067=>"111001001",
  24068=>"010100001",
  24069=>"111011111",
  24070=>"110101001",
  24071=>"111111101",
  24072=>"101101000",
  24073=>"011100000",
  24074=>"100111110",
  24075=>"011100101",
  24076=>"110010111",
  24077=>"011110001",
  24078=>"111000101",
  24079=>"101010000",
  24080=>"100100100",
  24081=>"000010010",
  24082=>"001001111",
  24083=>"010110001",
  24084=>"001010000",
  24085=>"001111110",
  24086=>"011001010",
  24087=>"000100100",
  24088=>"100101100",
  24089=>"000011010",
  24090=>"110100010",
  24091=>"011101000",
  24092=>"000011100",
  24093=>"001100111",
  24094=>"110000111",
  24095=>"101000111",
  24096=>"000011001",
  24097=>"000000100",
  24098=>"100010011",
  24099=>"100010000",
  24100=>"011101001",
  24101=>"010101111",
  24102=>"100001011",
  24103=>"110111010",
  24104=>"010000111",
  24105=>"001001010",
  24106=>"010111101",
  24107=>"100111010",
  24108=>"101010011",
  24109=>"000110101",
  24110=>"001010001",
  24111=>"011001011",
  24112=>"010100001",
  24113=>"000110110",
  24114=>"010001000",
  24115=>"001111111",
  24116=>"000110000",
  24117=>"101011011",
  24118=>"001010101",
  24119=>"100001000",
  24120=>"101110101",
  24121=>"000101110",
  24122=>"101111101",
  24123=>"100100110",
  24124=>"101101110",
  24125=>"001001001",
  24126=>"101100000",
  24127=>"100100010",
  24128=>"000000110",
  24129=>"011011010",
  24130=>"111101101",
  24131=>"001101010",
  24132=>"111001111",
  24133=>"101111111",
  24134=>"011111010",
  24135=>"001010010",
  24136=>"000101010",
  24137=>"100001001",
  24138=>"010111000",
  24139=>"101010101",
  24140=>"010111111",
  24141=>"100111011",
  24142=>"101111111",
  24143=>"100001010",
  24144=>"010010011",
  24145=>"011111101",
  24146=>"011010011",
  24147=>"000001001",
  24148=>"010000001",
  24149=>"100001001",
  24150=>"110111100",
  24151=>"001110111",
  24152=>"000100111",
  24153=>"110001101",
  24154=>"111110111",
  24155=>"001010000",
  24156=>"001011000",
  24157=>"010101001",
  24158=>"000010111",
  24159=>"000010000",
  24160=>"000010100",
  24161=>"011000110",
  24162=>"101101111",
  24163=>"001000110",
  24164=>"110000111",
  24165=>"000001000",
  24166=>"010101100",
  24167=>"010011111",
  24168=>"011000111",
  24169=>"010110010",
  24170=>"110100000",
  24171=>"110110010",
  24172=>"101010100",
  24173=>"110100000",
  24174=>"111000011",
  24175=>"011100011",
  24176=>"100000001",
  24177=>"000101111",
  24178=>"111101111",
  24179=>"101111011",
  24180=>"001010111",
  24181=>"011010001",
  24182=>"101011010",
  24183=>"010100111",
  24184=>"000010010",
  24185=>"111011101",
  24186=>"000000001",
  24187=>"101100011",
  24188=>"111100010",
  24189=>"010111001",
  24190=>"110110001",
  24191=>"000010101",
  24192=>"011110110",
  24193=>"111101100",
  24194=>"001011001",
  24195=>"000001101",
  24196=>"001111000",
  24197=>"100101101",
  24198=>"011001000",
  24199=>"000010110",
  24200=>"000000101",
  24201=>"010101001",
  24202=>"000110111",
  24203=>"001100010",
  24204=>"001000000",
  24205=>"100011000",
  24206=>"101110001",
  24207=>"101010111",
  24208=>"011010100",
  24209=>"010011000",
  24210=>"001011001",
  24211=>"010101110",
  24212=>"101010000",
  24213=>"011000110",
  24214=>"110000110",
  24215=>"011101001",
  24216=>"111011001",
  24217=>"010010110",
  24218=>"110001100",
  24219=>"101101011",
  24220=>"011001110",
  24221=>"000000101",
  24222=>"101111110",
  24223=>"011101001",
  24224=>"110011111",
  24225=>"100000100",
  24226=>"010000010",
  24227=>"010110000",
  24228=>"111110111",
  24229=>"000011100",
  24230=>"000010000",
  24231=>"011010010",
  24232=>"111110101",
  24233=>"110100111",
  24234=>"011110000",
  24235=>"010011100",
  24236=>"111000101",
  24237=>"110101001",
  24238=>"110110111",
  24239=>"111001100",
  24240=>"010011100",
  24241=>"001000110",
  24242=>"111001000",
  24243=>"100011011",
  24244=>"011100000",
  24245=>"100111100",
  24246=>"100101100",
  24247=>"110010010",
  24248=>"101101010",
  24249=>"010001101",
  24250=>"111011111",
  24251=>"000100001",
  24252=>"100000011",
  24253=>"011101100",
  24254=>"001101101",
  24255=>"001100001",
  24256=>"110111011",
  24257=>"101000011",
  24258=>"111100000",
  24259=>"010100011",
  24260=>"101101011",
  24261=>"011011100",
  24262=>"100011111",
  24263=>"110010110",
  24264=>"010001001",
  24265=>"001010101",
  24266=>"111000011",
  24267=>"100011001",
  24268=>"010110100",
  24269=>"010101110",
  24270=>"011110010",
  24271=>"111110010",
  24272=>"011111110",
  24273=>"111101101",
  24274=>"100001101",
  24275=>"001111001",
  24276=>"010001000",
  24277=>"010111110",
  24278=>"110111010",
  24279=>"010100111",
  24280=>"101111000",
  24281=>"001001010",
  24282=>"111001001",
  24283=>"000000111",
  24284=>"000000001",
  24285=>"111111111",
  24286=>"000111011",
  24287=>"011110101",
  24288=>"000000101",
  24289=>"001100001",
  24290=>"101110000",
  24291=>"101010010",
  24292=>"000001100",
  24293=>"001110110",
  24294=>"110001100",
  24295=>"001111010",
  24296=>"110011110",
  24297=>"010010110",
  24298=>"111111010",
  24299=>"010010100",
  24300=>"101001011",
  24301=>"000101111",
  24302=>"000000110",
  24303=>"110011010",
  24304=>"011101111",
  24305=>"001100010",
  24306=>"110010110",
  24307=>"111011001",
  24308=>"101110001",
  24309=>"111110011",
  24310=>"111110100",
  24311=>"010001010",
  24312=>"101000011",
  24313=>"111111011",
  24314=>"000111011",
  24315=>"000111000",
  24316=>"111101011",
  24317=>"011101010",
  24318=>"110101000",
  24319=>"100101000",
  24320=>"111111011",
  24321=>"111011110",
  24322=>"010110110",
  24323=>"011100110",
  24324=>"010010011",
  24325=>"101001110",
  24326=>"110010000",
  24327=>"100000000",
  24328=>"111000011",
  24329=>"111011010",
  24330=>"011111011",
  24331=>"000110100",
  24332=>"100101100",
  24333=>"011001110",
  24334=>"110100000",
  24335=>"000000100",
  24336=>"011101000",
  24337=>"001100111",
  24338=>"011010101",
  24339=>"110000010",
  24340=>"101000110",
  24341=>"111110000",
  24342=>"010010010",
  24343=>"110110111",
  24344=>"101000111",
  24345=>"011001111",
  24346=>"000000101",
  24347=>"001101110",
  24348=>"101100011",
  24349=>"111001110",
  24350=>"111100100",
  24351=>"111111000",
  24352=>"110100000",
  24353=>"111011011",
  24354=>"001000001",
  24355=>"101101010",
  24356=>"010000010",
  24357=>"111110001",
  24358=>"100001011",
  24359=>"110100101",
  24360=>"110011001",
  24361=>"001000110",
  24362=>"110010010",
  24363=>"101000001",
  24364=>"011100111",
  24365=>"000000011",
  24366=>"101111110",
  24367=>"101110101",
  24368=>"100001111",
  24369=>"110110000",
  24370=>"010111100",
  24371=>"110010101",
  24372=>"100010111",
  24373=>"000010101",
  24374=>"110111011",
  24375=>"101101101",
  24376=>"110111100",
  24377=>"001010011",
  24378=>"011110001",
  24379=>"001101010",
  24380=>"110010110",
  24381=>"001101011",
  24382=>"100000011",
  24383=>"100110010",
  24384=>"100001101",
  24385=>"111011100",
  24386=>"011110001",
  24387=>"101101001",
  24388=>"100010001",
  24389=>"100101110",
  24390=>"110101101",
  24391=>"111101111",
  24392=>"010011111",
  24393=>"000010011",
  24394=>"100101001",
  24395=>"011000001",
  24396=>"100010100",
  24397=>"000001011",
  24398=>"111111011",
  24399=>"100110000",
  24400=>"101101110",
  24401=>"110111010",
  24402=>"000100000",
  24403=>"000100000",
  24404=>"001011010",
  24405=>"000000001",
  24406=>"100111100",
  24407=>"110111000",
  24408=>"110010001",
  24409=>"110000111",
  24410=>"010001111",
  24411=>"001101011",
  24412=>"101010000",
  24413=>"011010100",
  24414=>"101011000",
  24415=>"000101111",
  24416=>"011000010",
  24417=>"011111100",
  24418=>"001000100",
  24419=>"101010110",
  24420=>"100001110",
  24421=>"001110101",
  24422=>"100011111",
  24423=>"110010011",
  24424=>"001000011",
  24425=>"010100000",
  24426=>"000101000",
  24427=>"111110010",
  24428=>"010000011",
  24429=>"000100100",
  24430=>"001000110",
  24431=>"111001101",
  24432=>"111000010",
  24433=>"110111101",
  24434=>"110110101",
  24435=>"000011100",
  24436=>"010001100",
  24437=>"001011111",
  24438=>"101011101",
  24439=>"000000011",
  24440=>"010110100",
  24441=>"011010101",
  24442=>"111111000",
  24443=>"011111010",
  24444=>"100100111",
  24445=>"000101001",
  24446=>"000111011",
  24447=>"110100001",
  24448=>"110000101",
  24449=>"011110101",
  24450=>"100110110",
  24451=>"000111001",
  24452=>"100110110",
  24453=>"111000100",
  24454=>"111000100",
  24455=>"001010000",
  24456=>"111010111",
  24457=>"111101101",
  24458=>"110100000",
  24459=>"000100001",
  24460=>"001000000",
  24461=>"100110100",
  24462=>"111001100",
  24463=>"111101001",
  24464=>"111101011",
  24465=>"010110011",
  24466=>"101100100",
  24467=>"101000000",
  24468=>"000011110",
  24469=>"000100110",
  24470=>"010010000",
  24471=>"011110101",
  24472=>"000101000",
  24473=>"011111000",
  24474=>"111010100",
  24475=>"000010111",
  24476=>"001011011",
  24477=>"001010000",
  24478=>"000000000",
  24479=>"111100010",
  24480=>"001101011",
  24481=>"100100011",
  24482=>"111111011",
  24483=>"010101111",
  24484=>"000010111",
  24485=>"110000010",
  24486=>"101011101",
  24487=>"000010100",
  24488=>"011010011",
  24489=>"010000010",
  24490=>"111001100",
  24491=>"100000111",
  24492=>"001110000",
  24493=>"101111010",
  24494=>"111011100",
  24495=>"100100001",
  24496=>"000000110",
  24497=>"101110000",
  24498=>"111001010",
  24499=>"100111100",
  24500=>"100010110",
  24501=>"000111111",
  24502=>"001001111",
  24503=>"100100110",
  24504=>"001000001",
  24505=>"101100111",
  24506=>"001010011",
  24507=>"110111000",
  24508=>"101111010",
  24509=>"101101111",
  24510=>"001111011",
  24511=>"000011001",
  24512=>"000110000",
  24513=>"001000001",
  24514=>"110111000",
  24515=>"010100101",
  24516=>"111011000",
  24517=>"001000010",
  24518=>"010010111",
  24519=>"101110000",
  24520=>"011110000",
  24521=>"100100010",
  24522=>"111010000",
  24523=>"111110101",
  24524=>"110100110",
  24525=>"101100111",
  24526=>"110001101",
  24527=>"101111111",
  24528=>"011011000",
  24529=>"101100001",
  24530=>"100010010",
  24531=>"111111100",
  24532=>"111001111",
  24533=>"110100110",
  24534=>"011010110",
  24535=>"001001101",
  24536=>"010111100",
  24537=>"001111000",
  24538=>"000110111",
  24539=>"010100111",
  24540=>"010101010",
  24541=>"100000011",
  24542=>"101000111",
  24543=>"100110000",
  24544=>"110100000",
  24545=>"100100110",
  24546=>"001001001",
  24547=>"101110111",
  24548=>"011111111",
  24549=>"000111000",
  24550=>"000000101",
  24551=>"001101010",
  24552=>"001010111",
  24553=>"010000000",
  24554=>"101101000",
  24555=>"101110001",
  24556=>"111010010",
  24557=>"001111001",
  24558=>"101110100",
  24559=>"110110011",
  24560=>"001011010",
  24561=>"011011001",
  24562=>"000100111",
  24563=>"011000111",
  24564=>"111000111",
  24565=>"100111001",
  24566=>"111010011",
  24567=>"010000111",
  24568=>"000001010",
  24569=>"011100000",
  24570=>"010100010",
  24571=>"001110011",
  24572=>"100001101",
  24573=>"111100010",
  24574=>"000101110",
  24575=>"011000011",
  24576=>"100000000",
  24577=>"000010001",
  24578=>"111101100",
  24579=>"101100101",
  24580=>"101010011",
  24581=>"011100101",
  24582=>"110101111",
  24583=>"010010110",
  24584=>"010100000",
  24585=>"001110101",
  24586=>"101010111",
  24587=>"110010010",
  24588=>"000101010",
  24589=>"000001110",
  24590=>"100001100",
  24591=>"001001101",
  24592=>"001010011",
  24593=>"101000010",
  24594=>"110010101",
  24595=>"111010101",
  24596=>"001000011",
  24597=>"000110100",
  24598=>"111011111",
  24599=>"011110100",
  24600=>"110100010",
  24601=>"010100101",
  24602=>"001101000",
  24603=>"001011001",
  24604=>"101101011",
  24605=>"110011001",
  24606=>"010100110",
  24607=>"111111000",
  24608=>"010101010",
  24609=>"100010100",
  24610=>"001100001",
  24611=>"010001000",
  24612=>"100001000",
  24613=>"110111100",
  24614=>"000100010",
  24615=>"000010110",
  24616=>"001001000",
  24617=>"100111010",
  24618=>"001000011",
  24619=>"101010010",
  24620=>"101000010",
  24621=>"000010010",
  24622=>"011010110",
  24623=>"000111011",
  24624=>"001110110",
  24625=>"111111111",
  24626=>"110010100",
  24627=>"110001011",
  24628=>"111101100",
  24629=>"110001111",
  24630=>"110001111",
  24631=>"100110110",
  24632=>"111100110",
  24633=>"100011001",
  24634=>"001011111",
  24635=>"111010101",
  24636=>"010010111",
  24637=>"110100000",
  24638=>"000101100",
  24639=>"111010100",
  24640=>"001001111",
  24641=>"010010011",
  24642=>"101101100",
  24643=>"100101011",
  24644=>"110010100",
  24645=>"000110010",
  24646=>"100100101",
  24647=>"100100100",
  24648=>"001101010",
  24649=>"101000010",
  24650=>"111001111",
  24651=>"110000111",
  24652=>"111011111",
  24653=>"011001100",
  24654=>"110011010",
  24655=>"111111010",
  24656=>"111111001",
  24657=>"011011010",
  24658=>"000000011",
  24659=>"010111100",
  24660=>"011111000",
  24661=>"011010100",
  24662=>"000101011",
  24663=>"100101001",
  24664=>"110111101",
  24665=>"101001010",
  24666=>"010111100",
  24667=>"011111011",
  24668=>"101111010",
  24669=>"100101101",
  24670=>"110101001",
  24671=>"100100111",
  24672=>"101111111",
  24673=>"111000101",
  24674=>"001101110",
  24675=>"101101100",
  24676=>"110001110",
  24677=>"010011011",
  24678=>"000001110",
  24679=>"100100101",
  24680=>"100101110",
  24681=>"110011101",
  24682=>"011110111",
  24683=>"101010011",
  24684=>"100101111",
  24685=>"011111101",
  24686=>"110000010",
  24687=>"010011001",
  24688=>"010000000",
  24689=>"010110101",
  24690=>"001101110",
  24691=>"110010110",
  24692=>"111101010",
  24693=>"101110000",
  24694=>"111100000",
  24695=>"111011001",
  24696=>"110111001",
  24697=>"010000100",
  24698=>"001000101",
  24699=>"000010111",
  24700=>"101000111",
  24701=>"000100010",
  24702=>"000011000",
  24703=>"110100111",
  24704=>"110001010",
  24705=>"000011111",
  24706=>"000101101",
  24707=>"011100011",
  24708=>"000000101",
  24709=>"011010000",
  24710=>"011001100",
  24711=>"010010000",
  24712=>"110100110",
  24713=>"011011010",
  24714=>"101010000",
  24715=>"010010111",
  24716=>"100101010",
  24717=>"010111011",
  24718=>"111110101",
  24719=>"010110011",
  24720=>"000100000",
  24721=>"111111011",
  24722=>"111011110",
  24723=>"010000101",
  24724=>"001000010",
  24725=>"000111100",
  24726=>"000000100",
  24727=>"011101110",
  24728=>"010010010",
  24729=>"000011000",
  24730=>"111011111",
  24731=>"100111101",
  24732=>"001011100",
  24733=>"110001111",
  24734=>"110001100",
  24735=>"000001110",
  24736=>"001000000",
  24737=>"000111111",
  24738=>"000000111",
  24739=>"110111001",
  24740=>"010011111",
  24741=>"001011000",
  24742=>"000111011",
  24743=>"111110001",
  24744=>"011111000",
  24745=>"011011110",
  24746=>"111110010",
  24747=>"010011011",
  24748=>"001000111",
  24749=>"010100010",
  24750=>"111101100",
  24751=>"110010000",
  24752=>"111111111",
  24753=>"010100010",
  24754=>"001111100",
  24755=>"111000100",
  24756=>"101001011",
  24757=>"000011001",
  24758=>"110011101",
  24759=>"011011111",
  24760=>"001110001",
  24761=>"000101001",
  24762=>"001001100",
  24763=>"000011000",
  24764=>"110010000",
  24765=>"011011001",
  24766=>"100011100",
  24767=>"010001000",
  24768=>"111001100",
  24769=>"100100111",
  24770=>"100001111",
  24771=>"101111101",
  24772=>"010100111",
  24773=>"000110111",
  24774=>"110000100",
  24775=>"100011010",
  24776=>"110011110",
  24777=>"000001000",
  24778=>"000110101",
  24779=>"101100010",
  24780=>"100011111",
  24781=>"011100011",
  24782=>"111000011",
  24783=>"100010001",
  24784=>"111100000",
  24785=>"110001011",
  24786=>"111011011",
  24787=>"111010011",
  24788=>"000011000",
  24789=>"001001001",
  24790=>"011101111",
  24791=>"010100000",
  24792=>"010001001",
  24793=>"111011001",
  24794=>"100010010",
  24795=>"111100011",
  24796=>"110001010",
  24797=>"110101011",
  24798=>"000110000",
  24799=>"110001011",
  24800=>"101000111",
  24801=>"101011111",
  24802=>"110001010",
  24803=>"000000100",
  24804=>"010100100",
  24805=>"011000011",
  24806=>"000001001",
  24807=>"111001010",
  24808=>"100010111",
  24809=>"101001111",
  24810=>"000100100",
  24811=>"111110110",
  24812=>"001110000",
  24813=>"011101101",
  24814=>"110101100",
  24815=>"010000001",
  24816=>"011111011",
  24817=>"001100001",
  24818=>"101001000",
  24819=>"110001101",
  24820=>"110111011",
  24821=>"010110011",
  24822=>"001011011",
  24823=>"111101000",
  24824=>"111001110",
  24825=>"000110011",
  24826=>"100010000",
  24827=>"011001010",
  24828=>"110111101",
  24829=>"011000011",
  24830=>"100001110",
  24831=>"011110111",
  24832=>"101110111",
  24833=>"111100111",
  24834=>"100001110",
  24835=>"011100100",
  24836=>"010010101",
  24837=>"000110001",
  24838=>"011100111",
  24839=>"101101110",
  24840=>"010010010",
  24841=>"011010111",
  24842=>"011100101",
  24843=>"111101011",
  24844=>"100001001",
  24845=>"100111110",
  24846=>"011001101",
  24847=>"000101100",
  24848=>"111100101",
  24849=>"111000111",
  24850=>"001010100",
  24851=>"000101010",
  24852=>"010000110",
  24853=>"000101000",
  24854=>"000111000",
  24855=>"001011000",
  24856=>"001001010",
  24857=>"101100001",
  24858=>"101100000",
  24859=>"011011000",
  24860=>"011100000",
  24861=>"111001111",
  24862=>"001010000",
  24863=>"001000011",
  24864=>"000101000",
  24865=>"000101110",
  24866=>"000101111",
  24867=>"011110110",
  24868=>"111011010",
  24869=>"101011001",
  24870=>"010010111",
  24871=>"011000110",
  24872=>"111100011",
  24873=>"101000100",
  24874=>"101100111",
  24875=>"010001110",
  24876=>"011011000",
  24877=>"101111110",
  24878=>"001100111",
  24879=>"010011000",
  24880=>"000000000",
  24881=>"010110111",
  24882=>"101001011",
  24883=>"011101011",
  24884=>"110000000",
  24885=>"001000000",
  24886=>"110011110",
  24887=>"101110111",
  24888=>"001011111",
  24889=>"000011001",
  24890=>"011000000",
  24891=>"001100101",
  24892=>"101100100",
  24893=>"110110101",
  24894=>"110111111",
  24895=>"000001110",
  24896=>"010011011",
  24897=>"000100100",
  24898=>"011000000",
  24899=>"000001100",
  24900=>"000001001",
  24901=>"101111110",
  24902=>"000000111",
  24903=>"000111111",
  24904=>"101110010",
  24905=>"001010101",
  24906=>"111001111",
  24907=>"111001001",
  24908=>"111010000",
  24909=>"010110111",
  24910=>"011010101",
  24911=>"101110000",
  24912=>"110101101",
  24913=>"101010110",
  24914=>"111111111",
  24915=>"111101010",
  24916=>"000101000",
  24917=>"001000100",
  24918=>"011111011",
  24919=>"110010000",
  24920=>"010101011",
  24921=>"000101010",
  24922=>"000101001",
  24923=>"010110000",
  24924=>"111101101",
  24925=>"011111100",
  24926=>"110100011",
  24927=>"000011000",
  24928=>"101110001",
  24929=>"000000110",
  24930=>"100100111",
  24931=>"110011001",
  24932=>"010001110",
  24933=>"010010000",
  24934=>"000001101",
  24935=>"010110010",
  24936=>"010011000",
  24937=>"011101100",
  24938=>"100000101",
  24939=>"100110110",
  24940=>"101100100",
  24941=>"101110000",
  24942=>"101000100",
  24943=>"001111010",
  24944=>"001111111",
  24945=>"111001000",
  24946=>"111111100",
  24947=>"110000111",
  24948=>"000000010",
  24949=>"010110000",
  24950=>"001110111",
  24951=>"110111001",
  24952=>"011111000",
  24953=>"001001111",
  24954=>"010011110",
  24955=>"111000100",
  24956=>"101101100",
  24957=>"101011110",
  24958=>"000111100",
  24959=>"010010011",
  24960=>"100111101",
  24961=>"011101100",
  24962=>"010010101",
  24963=>"000101110",
  24964=>"011010001",
  24965=>"111100010",
  24966=>"000001101",
  24967=>"011101011",
  24968=>"110001110",
  24969=>"011100101",
  24970=>"010010110",
  24971=>"010001000",
  24972=>"000001101",
  24973=>"110001111",
  24974=>"100001000",
  24975=>"000100111",
  24976=>"110011110",
  24977=>"001000001",
  24978=>"011000011",
  24979=>"110110101",
  24980=>"010001010",
  24981=>"111111111",
  24982=>"101101010",
  24983=>"111010101",
  24984=>"100110101",
  24985=>"001100110",
  24986=>"011001100",
  24987=>"100010000",
  24988=>"101101000",
  24989=>"010111100",
  24990=>"111111010",
  24991=>"111111100",
  24992=>"101101101",
  24993=>"111101111",
  24994=>"011110100",
  24995=>"000000001",
  24996=>"011111110",
  24997=>"000010001",
  24998=>"010110011",
  24999=>"001101101",
  25000=>"100111111",
  25001=>"110000010",
  25002=>"111011010",
  25003=>"010100011",
  25004=>"111110111",
  25005=>"001011111",
  25006=>"101111101",
  25007=>"000010101",
  25008=>"011001001",
  25009=>"101011001",
  25010=>"100011010",
  25011=>"000111001",
  25012=>"101011100",
  25013=>"011001011",
  25014=>"101100001",
  25015=>"110011101",
  25016=>"111111100",
  25017=>"000000001",
  25018=>"011001010",
  25019=>"010000011",
  25020=>"101010011",
  25021=>"001111000",
  25022=>"011010100",
  25023=>"000001100",
  25024=>"000000000",
  25025=>"000011111",
  25026=>"001110110",
  25027=>"111011101",
  25028=>"110010011",
  25029=>"010010100",
  25030=>"001010111",
  25031=>"101001101",
  25032=>"010101000",
  25033=>"101001100",
  25034=>"011001011",
  25035=>"101100000",
  25036=>"101001101",
  25037=>"000101001",
  25038=>"100000101",
  25039=>"001110010",
  25040=>"011110011",
  25041=>"100010100",
  25042=>"011101000",
  25043=>"110011011",
  25044=>"000111100",
  25045=>"000100001",
  25046=>"111001000",
  25047=>"010111010",
  25048=>"110001101",
  25049=>"111100001",
  25050=>"100001111",
  25051=>"111001011",
  25052=>"101110001",
  25053=>"111011101",
  25054=>"010000111",
  25055=>"010000000",
  25056=>"111100011",
  25057=>"101001100",
  25058=>"001111010",
  25059=>"110100011",
  25060=>"110110100",
  25061=>"100100000",
  25062=>"110101101",
  25063=>"010100110",
  25064=>"000110111",
  25065=>"010111101",
  25066=>"000001000",
  25067=>"100111001",
  25068=>"000001011",
  25069=>"010000001",
  25070=>"110101101",
  25071=>"000100110",
  25072=>"100011001",
  25073=>"111110101",
  25074=>"011010000",
  25075=>"101100010",
  25076=>"001000010",
  25077=>"010000010",
  25078=>"101110111",
  25079=>"010101001",
  25080=>"101111000",
  25081=>"111001001",
  25082=>"100000110",
  25083=>"000111111",
  25084=>"001101011",
  25085=>"011111010",
  25086=>"010100010",
  25087=>"100010001",
  25088=>"111111010",
  25089=>"011011001",
  25090=>"101001011",
  25091=>"111100010",
  25092=>"101100101",
  25093=>"010000010",
  25094=>"100011010",
  25095=>"010010100",
  25096=>"001101101",
  25097=>"011101111",
  25098=>"110000111",
  25099=>"100010000",
  25100=>"001010001",
  25101=>"101100010",
  25102=>"001101100",
  25103=>"000011100",
  25104=>"001001100",
  25105=>"100001101",
  25106=>"000001110",
  25107=>"101110011",
  25108=>"001011011",
  25109=>"110100110",
  25110=>"111000101",
  25111=>"110010100",
  25112=>"110000000",
  25113=>"010111010",
  25114=>"100001101",
  25115=>"100001011",
  25116=>"111001010",
  25117=>"000110000",
  25118=>"011101000",
  25119=>"101111111",
  25120=>"101011011",
  25121=>"111110011",
  25122=>"011000000",
  25123=>"100111010",
  25124=>"001000000",
  25125=>"000000111",
  25126=>"000100110",
  25127=>"111100101",
  25128=>"100010000",
  25129=>"010001011",
  25130=>"100110000",
  25131=>"011100011",
  25132=>"011101001",
  25133=>"110001000",
  25134=>"100010100",
  25135=>"100110000",
  25136=>"000111100",
  25137=>"110101000",
  25138=>"000100110",
  25139=>"100000000",
  25140=>"000111000",
  25141=>"111111011",
  25142=>"101101000",
  25143=>"110000111",
  25144=>"110110001",
  25145=>"111100011",
  25146=>"100001000",
  25147=>"100111011",
  25148=>"010010100",
  25149=>"110110111",
  25150=>"001010000",
  25151=>"001001101",
  25152=>"000001000",
  25153=>"101101111",
  25154=>"000011100",
  25155=>"111010000",
  25156=>"001011010",
  25157=>"010111011",
  25158=>"111101011",
  25159=>"001000001",
  25160=>"101001000",
  25161=>"000101110",
  25162=>"110010111",
  25163=>"100101101",
  25164=>"000110100",
  25165=>"100101001",
  25166=>"000001101",
  25167=>"011000011",
  25168=>"100011110",
  25169=>"111000100",
  25170=>"001000000",
  25171=>"101010110",
  25172=>"001001010",
  25173=>"000111000",
  25174=>"100010000",
  25175=>"001001010",
  25176=>"011001110",
  25177=>"101011001",
  25178=>"001001110",
  25179=>"100101000",
  25180=>"000111111",
  25181=>"011111101",
  25182=>"011111111",
  25183=>"100000011",
  25184=>"101000101",
  25185=>"010000101",
  25186=>"101000001",
  25187=>"011001010",
  25188=>"000000110",
  25189=>"110001011",
  25190=>"101001111",
  25191=>"110111110",
  25192=>"000100011",
  25193=>"110000011",
  25194=>"111101011",
  25195=>"101010001",
  25196=>"111001010",
  25197=>"111111001",
  25198=>"101100011",
  25199=>"111100000",
  25200=>"011011001",
  25201=>"101101001",
  25202=>"011010100",
  25203=>"111011000",
  25204=>"100001111",
  25205=>"000000110",
  25206=>"111100100",
  25207=>"000001111",
  25208=>"110101100",
  25209=>"000011111",
  25210=>"110101000",
  25211=>"110000010",
  25212=>"110001000",
  25213=>"110111011",
  25214=>"010001010",
  25215=>"110111111",
  25216=>"010001001",
  25217=>"000100011",
  25218=>"000000111",
  25219=>"001011000",
  25220=>"110001111",
  25221=>"001101001",
  25222=>"110001010",
  25223=>"101110010",
  25224=>"100110010",
  25225=>"010000010",
  25226=>"101111011",
  25227=>"110101010",
  25228=>"001001001",
  25229=>"011101000",
  25230=>"001110000",
  25231=>"110001000",
  25232=>"001011001",
  25233=>"111110010",
  25234=>"101000001",
  25235=>"000011100",
  25236=>"000111001",
  25237=>"111100000",
  25238=>"110011100",
  25239=>"010100011",
  25240=>"000111110",
  25241=>"111110011",
  25242=>"101101000",
  25243=>"001000001",
  25244=>"011010111",
  25245=>"110110110",
  25246=>"010101101",
  25247=>"111111011",
  25248=>"110000100",
  25249=>"111111100",
  25250=>"101000001",
  25251=>"001110001",
  25252=>"111101010",
  25253=>"101011110",
  25254=>"100101111",
  25255=>"011101100",
  25256=>"011111110",
  25257=>"101000100",
  25258=>"010010010",
  25259=>"001001110",
  25260=>"110000011",
  25261=>"001111101",
  25262=>"111000010",
  25263=>"110011010",
  25264=>"000100110",
  25265=>"110101000",
  25266=>"011011100",
  25267=>"110010000",
  25268=>"100101010",
  25269=>"111000010",
  25270=>"110001000",
  25271=>"001110010",
  25272=>"100100100",
  25273=>"100001100",
  25274=>"010011011",
  25275=>"010110101",
  25276=>"111010000",
  25277=>"111111100",
  25278=>"000000101",
  25279=>"001101000",
  25280=>"111110101",
  25281=>"011100111",
  25282=>"100110000",
  25283=>"111100100",
  25284=>"000011000",
  25285=>"000001101",
  25286=>"110011110",
  25287=>"001100100",
  25288=>"100111000",
  25289=>"000001100",
  25290=>"100110101",
  25291=>"010100100",
  25292=>"001111101",
  25293=>"001110101",
  25294=>"000101000",
  25295=>"010001011",
  25296=>"101011000",
  25297=>"011101110",
  25298=>"101100001",
  25299=>"001001010",
  25300=>"000100000",
  25301=>"010110011",
  25302=>"101101010",
  25303=>"000111101",
  25304=>"111001010",
  25305=>"100000001",
  25306=>"011111001",
  25307=>"101110000",
  25308=>"001001110",
  25309=>"001101001",
  25310=>"101001001",
  25311=>"000111000",
  25312=>"011010100",
  25313=>"100001010",
  25314=>"000111110",
  25315=>"101100010",
  25316=>"000100011",
  25317=>"011011111",
  25318=>"010100010",
  25319=>"000001110",
  25320=>"101001001",
  25321=>"101010001",
  25322=>"111110100",
  25323=>"100110101",
  25324=>"000000011",
  25325=>"110000110",
  25326=>"110000000",
  25327=>"011110100",
  25328=>"001011001",
  25329=>"101000001",
  25330=>"101001111",
  25331=>"101011111",
  25332=>"000100000",
  25333=>"111100111",
  25334=>"010101000",
  25335=>"010110010",
  25336=>"000100101",
  25337=>"110000110",
  25338=>"100100100",
  25339=>"101110001",
  25340=>"001110001",
  25341=>"000000110",
  25342=>"101111110",
  25343=>"100000100",
  25344=>"001001010",
  25345=>"001010111",
  25346=>"001001100",
  25347=>"000100011",
  25348=>"100010010",
  25349=>"000011111",
  25350=>"100010011",
  25351=>"101111110",
  25352=>"101101000",
  25353=>"010100100",
  25354=>"011000111",
  25355=>"101001100",
  25356=>"110010010",
  25357=>"111010011",
  25358=>"000111000",
  25359=>"001001111",
  25360=>"110011110",
  25361=>"001101011",
  25362=>"001000010",
  25363=>"101111110",
  25364=>"010010010",
  25365=>"010110101",
  25366=>"100100000",
  25367=>"100000011",
  25368=>"110001001",
  25369=>"001000100",
  25370=>"001101000",
  25371=>"111010000",
  25372=>"011100100",
  25373=>"010111101",
  25374=>"110110001",
  25375=>"100101000",
  25376=>"000100001",
  25377=>"110111001",
  25378=>"011000101",
  25379=>"100100011",
  25380=>"110011000",
  25381=>"011010111",
  25382=>"001101101",
  25383=>"101111111",
  25384=>"100101000",
  25385=>"110001000",
  25386=>"111111101",
  25387=>"101111111",
  25388=>"011100111",
  25389=>"111011110",
  25390=>"010100110",
  25391=>"110111111",
  25392=>"011010010",
  25393=>"101000001",
  25394=>"111011111",
  25395=>"000011110",
  25396=>"011011100",
  25397=>"111000001",
  25398=>"111001011",
  25399=>"100100101",
  25400=>"001010101",
  25401=>"110110000",
  25402=>"011010110",
  25403=>"000001010",
  25404=>"101001010",
  25405=>"001001010",
  25406=>"111001100",
  25407=>"000110110",
  25408=>"100101011",
  25409=>"100000111",
  25410=>"101010011",
  25411=>"011101001",
  25412=>"101100000",
  25413=>"100101000",
  25414=>"001011110",
  25415=>"110001010",
  25416=>"100001001",
  25417=>"110001010",
  25418=>"001011110",
  25419=>"110101011",
  25420=>"111111111",
  25421=>"000001011",
  25422=>"011001011",
  25423=>"110010100",
  25424=>"101101010",
  25425=>"101000000",
  25426=>"111101011",
  25427=>"010100101",
  25428=>"110101011",
  25429=>"011010010",
  25430=>"001100101",
  25431=>"011100100",
  25432=>"000000010",
  25433=>"101100000",
  25434=>"111010001",
  25435=>"111001010",
  25436=>"011111100",
  25437=>"000101001",
  25438=>"100111011",
  25439=>"000010001",
  25440=>"001100100",
  25441=>"101101111",
  25442=>"101111000",
  25443=>"111011001",
  25444=>"011111001",
  25445=>"001100111",
  25446=>"011100001",
  25447=>"001111111",
  25448=>"011110111",
  25449=>"100101001",
  25450=>"010101110",
  25451=>"111010010",
  25452=>"011010001",
  25453=>"101110010",
  25454=>"111000100",
  25455=>"001101100",
  25456=>"000001110",
  25457=>"001010100",
  25458=>"101010111",
  25459=>"111101100",
  25460=>"110010001",
  25461=>"001000100",
  25462=>"000111101",
  25463=>"000101101",
  25464=>"100110111",
  25465=>"110001010",
  25466=>"011010010",
  25467=>"000001111",
  25468=>"010010110",
  25469=>"000101011",
  25470=>"100000110",
  25471=>"000101010",
  25472=>"000011000",
  25473=>"101001010",
  25474=>"111000000",
  25475=>"000001010",
  25476=>"110111110",
  25477=>"101111011",
  25478=>"001000011",
  25479=>"010000001",
  25480=>"111111000",
  25481=>"110100111",
  25482=>"110110100",
  25483=>"111101111",
  25484=>"100001000",
  25485=>"011010000",
  25486=>"000110111",
  25487=>"101111110",
  25488=>"100011110",
  25489=>"001010111",
  25490=>"001100010",
  25491=>"011100111",
  25492=>"101001011",
  25493=>"000100101",
  25494=>"011010001",
  25495=>"000100011",
  25496=>"000111011",
  25497=>"000001110",
  25498=>"000100101",
  25499=>"010100011",
  25500=>"100011111",
  25501=>"000101101",
  25502=>"101101101",
  25503=>"101101011",
  25504=>"011110001",
  25505=>"111011000",
  25506=>"111010000",
  25507=>"101000100",
  25508=>"101000010",
  25509=>"100011100",
  25510=>"100011110",
  25511=>"010110101",
  25512=>"000001011",
  25513=>"111101111",
  25514=>"001001010",
  25515=>"001001110",
  25516=>"101010111",
  25517=>"101110010",
  25518=>"000111000",
  25519=>"010001000",
  25520=>"001100101",
  25521=>"111010101",
  25522=>"111111100",
  25523=>"010000000",
  25524=>"111111101",
  25525=>"110000001",
  25526=>"010001010",
  25527=>"100000010",
  25528=>"000110001",
  25529=>"001001010",
  25530=>"100100100",
  25531=>"110011010",
  25532=>"110001010",
  25533=>"101010000",
  25534=>"001010010",
  25535=>"001011101",
  25536=>"001101101",
  25537=>"101010001",
  25538=>"101000110",
  25539=>"111001011",
  25540=>"001100001",
  25541=>"111100111",
  25542=>"111100010",
  25543=>"110011001",
  25544=>"011010001",
  25545=>"110111110",
  25546=>"111010100",
  25547=>"011000101",
  25548=>"111111001",
  25549=>"101100101",
  25550=>"010011111",
  25551=>"100100100",
  25552=>"100110110",
  25553=>"111110011",
  25554=>"011000110",
  25555=>"110010100",
  25556=>"111110010",
  25557=>"011010010",
  25558=>"010011110",
  25559=>"000000000",
  25560=>"100110101",
  25561=>"101101111",
  25562=>"101001111",
  25563=>"000110111",
  25564=>"101111110",
  25565=>"010001010",
  25566=>"111011001",
  25567=>"100100111",
  25568=>"111110011",
  25569=>"111101101",
  25570=>"110000110",
  25571=>"100111010",
  25572=>"000011011",
  25573=>"000001011",
  25574=>"000111110",
  25575=>"011100001",
  25576=>"001101110",
  25577=>"011010110",
  25578=>"001010011",
  25579=>"000000100",
  25580=>"011101001",
  25581=>"010011010",
  25582=>"011001101",
  25583=>"011101111",
  25584=>"000100100",
  25585=>"001011110",
  25586=>"000001010",
  25587=>"010010011",
  25588=>"111100000",
  25589=>"101110100",
  25590=>"100101111",
  25591=>"010001110",
  25592=>"000101010",
  25593=>"100111110",
  25594=>"111011110",
  25595=>"000111101",
  25596=>"010100010",
  25597=>"111001111",
  25598=>"111101111",
  25599=>"011011011",
  25600=>"011111010",
  25601=>"111000011",
  25602=>"010101001",
  25603=>"000100101",
  25604=>"001111111",
  25605=>"011011001",
  25606=>"011010111",
  25607=>"101111100",
  25608=>"000111001",
  25609=>"000111111",
  25610=>"001000100",
  25611=>"110011011",
  25612=>"011000000",
  25613=>"000100010",
  25614=>"110100010",
  25615=>"001010011",
  25616=>"010111110",
  25617=>"001011111",
  25618=>"101111110",
  25619=>"011001011",
  25620=>"011001110",
  25621=>"000100001",
  25622=>"111111111",
  25623=>"001100000",
  25624=>"010111111",
  25625=>"001011010",
  25626=>"000001000",
  25627=>"011010010",
  25628=>"010011000",
  25629=>"100010100",
  25630=>"111100100",
  25631=>"011100000",
  25632=>"110111011",
  25633=>"110101101",
  25634=>"010100000",
  25635=>"101011110",
  25636=>"100111010",
  25637=>"100100011",
  25638=>"001100011",
  25639=>"011011101",
  25640=>"110110001",
  25641=>"001000001",
  25642=>"000000111",
  25643=>"100111110",
  25644=>"010111010",
  25645=>"110101000",
  25646=>"000000011",
  25647=>"100101001",
  25648=>"111011111",
  25649=>"001111111",
  25650=>"010011000",
  25651=>"110000100",
  25652=>"100000011",
  25653=>"000110011",
  25654=>"000011010",
  25655=>"011101111",
  25656=>"001000101",
  25657=>"001000000",
  25658=>"010010111",
  25659=>"101100000",
  25660=>"110011010",
  25661=>"111111101",
  25662=>"000000000",
  25663=>"001100010",
  25664=>"111000000",
  25665=>"000100101",
  25666=>"010101011",
  25667=>"010101110",
  25668=>"010000001",
  25669=>"000111101",
  25670=>"001100111",
  25671=>"001100111",
  25672=>"010010001",
  25673=>"101110000",
  25674=>"101110011",
  25675=>"001011010",
  25676=>"110010011",
  25677=>"010001000",
  25678=>"100110111",
  25679=>"101010110",
  25680=>"111101000",
  25681=>"000111000",
  25682=>"010000111",
  25683=>"001001011",
  25684=>"001101110",
  25685=>"110111111",
  25686=>"001011110",
  25687=>"111110110",
  25688=>"010111010",
  25689=>"010000101",
  25690=>"101111101",
  25691=>"000100010",
  25692=>"110110010",
  25693=>"000110001",
  25694=>"100000011",
  25695=>"011100111",
  25696=>"000001010",
  25697=>"111111100",
  25698=>"101001111",
  25699=>"010001111",
  25700=>"010010100",
  25701=>"110111101",
  25702=>"001000110",
  25703=>"010011110",
  25704=>"101110000",
  25705=>"111101010",
  25706=>"011000100",
  25707=>"011001010",
  25708=>"011001011",
  25709=>"101110101",
  25710=>"111010101",
  25711=>"010110100",
  25712=>"110000101",
  25713=>"011111111",
  25714=>"001010110",
  25715=>"010010101",
  25716=>"000001010",
  25717=>"101010001",
  25718=>"101100111",
  25719=>"000010110",
  25720=>"110001100",
  25721=>"010001110",
  25722=>"111110101",
  25723=>"010010010",
  25724=>"001000111",
  25725=>"101100011",
  25726=>"110000001",
  25727=>"000111010",
  25728=>"110110001",
  25729=>"011010101",
  25730=>"100010101",
  25731=>"101011100",
  25732=>"101111010",
  25733=>"101010101",
  25734=>"111110011",
  25735=>"001000011",
  25736=>"011110000",
  25737=>"110010001",
  25738=>"011101110",
  25739=>"111111001",
  25740=>"111100010",
  25741=>"011001001",
  25742=>"010010010",
  25743=>"101011010",
  25744=>"110011110",
  25745=>"010100000",
  25746=>"001100110",
  25747=>"011001010",
  25748=>"000010100",
  25749=>"000000010",
  25750=>"110011010",
  25751=>"000000010",
  25752=>"010010100",
  25753=>"000111100",
  25754=>"100000011",
  25755=>"101110100",
  25756=>"110001111",
  25757=>"111101101",
  25758=>"011011110",
  25759=>"000110110",
  25760=>"000011100",
  25761=>"011101100",
  25762=>"000110101",
  25763=>"111000110",
  25764=>"000000101",
  25765=>"000110111",
  25766=>"100101000",
  25767=>"101000111",
  25768=>"000111100",
  25769=>"111110100",
  25770=>"011100011",
  25771=>"100101111",
  25772=>"110101111",
  25773=>"000001011",
  25774=>"000000010",
  25775=>"010000000",
  25776=>"011011001",
  25777=>"111001101",
  25778=>"010110010",
  25779=>"001101111",
  25780=>"111110010",
  25781=>"011110000",
  25782=>"111001101",
  25783=>"000011110",
  25784=>"010110110",
  25785=>"001111111",
  25786=>"101001111",
  25787=>"110110011",
  25788=>"110111010",
  25789=>"000111000",
  25790=>"000011111",
  25791=>"111010101",
  25792=>"001111111",
  25793=>"100110111",
  25794=>"100110000",
  25795=>"110001110",
  25796=>"110010010",
  25797=>"011010110",
  25798=>"111100010",
  25799=>"110001101",
  25800=>"111110110",
  25801=>"001100011",
  25802=>"011010111",
  25803=>"000101101",
  25804=>"101101110",
  25805=>"001110000",
  25806=>"110000011",
  25807=>"101000101",
  25808=>"111100101",
  25809=>"010011011",
  25810=>"100111001",
  25811=>"001100000",
  25812=>"111111001",
  25813=>"001001111",
  25814=>"101010000",
  25815=>"111101010",
  25816=>"101110000",
  25817=>"110100001",
  25818=>"100000010",
  25819=>"100000010",
  25820=>"010010000",
  25821=>"111001110",
  25822=>"111010100",
  25823=>"000000111",
  25824=>"110100010",
  25825=>"000000010",
  25826=>"010100101",
  25827=>"001100000",
  25828=>"001110000",
  25829=>"100111111",
  25830=>"010111111",
  25831=>"100101001",
  25832=>"001110000",
  25833=>"001101100",
  25834=>"010100001",
  25835=>"000110100",
  25836=>"110101110",
  25837=>"011000011",
  25838=>"101100110",
  25839=>"001011111",
  25840=>"111011111",
  25841=>"000100110",
  25842=>"011011010",
  25843=>"110111011",
  25844=>"100001100",
  25845=>"001000111",
  25846=>"001101110",
  25847=>"100011010",
  25848=>"010111001",
  25849=>"001010000",
  25850=>"101011011",
  25851=>"101110000",
  25852=>"110101110",
  25853=>"111101100",
  25854=>"110011100",
  25855=>"101001011",
  25856=>"010000110",
  25857=>"100001100",
  25858=>"001110100",
  25859=>"110001110",
  25860=>"111000010",
  25861=>"001011111",
  25862=>"100110101",
  25863=>"100111100",
  25864=>"101000011",
  25865=>"100001111",
  25866=>"100000111",
  25867=>"101101111",
  25868=>"010101010",
  25869=>"001100100",
  25870=>"111100101",
  25871=>"000100001",
  25872=>"000001100",
  25873=>"010010010",
  25874=>"000001100",
  25875=>"010111010",
  25876=>"010110000",
  25877=>"011110001",
  25878=>"000001101",
  25879=>"001000000",
  25880=>"100110100",
  25881=>"110000110",
  25882=>"000001100",
  25883=>"010111000",
  25884=>"001001100",
  25885=>"011101000",
  25886=>"001001100",
  25887=>"010111101",
  25888=>"000101000",
  25889=>"011011000",
  25890=>"110101001",
  25891=>"111100111",
  25892=>"101000111",
  25893=>"111001100",
  25894=>"000100111",
  25895=>"110010100",
  25896=>"101101001",
  25897=>"011000000",
  25898=>"101010001",
  25899=>"100010000",
  25900=>"110010010",
  25901=>"011001000",
  25902=>"001001001",
  25903=>"000011101",
  25904=>"010111001",
  25905=>"100011011",
  25906=>"100011111",
  25907=>"001011110",
  25908=>"000011010",
  25909=>"111111101",
  25910=>"100010011",
  25911=>"101111011",
  25912=>"011011000",
  25913=>"111101111",
  25914=>"100101100",
  25915=>"111011100",
  25916=>"000100111",
  25917=>"001001001",
  25918=>"011010001",
  25919=>"101000000",
  25920=>"010111111",
  25921=>"100000111",
  25922=>"011110000",
  25923=>"111011110",
  25924=>"001110000",
  25925=>"001001010",
  25926=>"011100000",
  25927=>"011001001",
  25928=>"010110100",
  25929=>"000001010",
  25930=>"011110100",
  25931=>"001010000",
  25932=>"111111100",
  25933=>"000011100",
  25934=>"100110000",
  25935=>"101010111",
  25936=>"111110111",
  25937=>"010110111",
  25938=>"001000100",
  25939=>"101010010",
  25940=>"100111010",
  25941=>"010010011",
  25942=>"000000011",
  25943=>"101110101",
  25944=>"111010000",
  25945=>"100101100",
  25946=>"101100011",
  25947=>"110001100",
  25948=>"011011000",
  25949=>"101010110",
  25950=>"001110011",
  25951=>"111010000",
  25952=>"000100000",
  25953=>"010010000",
  25954=>"011101101",
  25955=>"111010001",
  25956=>"110000011",
  25957=>"100111100",
  25958=>"011010111",
  25959=>"000000101",
  25960=>"111011110",
  25961=>"111011110",
  25962=>"110001100",
  25963=>"011000110",
  25964=>"100100100",
  25965=>"110110000",
  25966=>"010000101",
  25967=>"001110110",
  25968=>"000110011",
  25969=>"011101001",
  25970=>"000110100",
  25971=>"011110000",
  25972=>"001011100",
  25973=>"001001110",
  25974=>"010001001",
  25975=>"000111010",
  25976=>"100101110",
  25977=>"001001110",
  25978=>"111100101",
  25979=>"000101010",
  25980=>"001101000",
  25981=>"111111000",
  25982=>"000011110",
  25983=>"111100010",
  25984=>"001111110",
  25985=>"001011101",
  25986=>"001011011",
  25987=>"101010111",
  25988=>"111111101",
  25989=>"111000011",
  25990=>"101111110",
  25991=>"110101000",
  25992=>"011100110",
  25993=>"101101000",
  25994=>"110111100",
  25995=>"000000100",
  25996=>"101000101",
  25997=>"100011100",
  25998=>"111111000",
  25999=>"001100100",
  26000=>"010111101",
  26001=>"101000010",
  26002=>"010000010",
  26003=>"000100100",
  26004=>"100011001",
  26005=>"111011001",
  26006=>"110101000",
  26007=>"111111001",
  26008=>"101000010",
  26009=>"100110011",
  26010=>"101011101",
  26011=>"001110001",
  26012=>"100101110",
  26013=>"010010110",
  26014=>"110011010",
  26015=>"100100011",
  26016=>"101010010",
  26017=>"110101010",
  26018=>"100100010",
  26019=>"110011111",
  26020=>"110101000",
  26021=>"111000000",
  26022=>"111001000",
  26023=>"010111010",
  26024=>"110101111",
  26025=>"110001011",
  26026=>"100001111",
  26027=>"010010111",
  26028=>"000000111",
  26029=>"011100110",
  26030=>"100000111",
  26031=>"101000010",
  26032=>"010101000",
  26033=>"111011010",
  26034=>"101101011",
  26035=>"000000100",
  26036=>"000101100",
  26037=>"000000111",
  26038=>"110011111",
  26039=>"101111101",
  26040=>"110001101",
  26041=>"000110000",
  26042=>"111111111",
  26043=>"001000000",
  26044=>"011001111",
  26045=>"001001110",
  26046=>"001111011",
  26047=>"010010000",
  26048=>"000100100",
  26049=>"010100111",
  26050=>"001011000",
  26051=>"101100001",
  26052=>"010000100",
  26053=>"110000010",
  26054=>"100011100",
  26055=>"110000000",
  26056=>"111001111",
  26057=>"100001010",
  26058=>"001010000",
  26059=>"101101110",
  26060=>"001110000",
  26061=>"101101101",
  26062=>"010100100",
  26063=>"011111011",
  26064=>"011010100",
  26065=>"010001110",
  26066=>"100010111",
  26067=>"001001010",
  26068=>"010101111",
  26069=>"110101010",
  26070=>"010000011",
  26071=>"111000100",
  26072=>"001110011",
  26073=>"001110110",
  26074=>"010111010",
  26075=>"000111010",
  26076=>"010100001",
  26077=>"101100100",
  26078=>"101010001",
  26079=>"011111110",
  26080=>"101000000",
  26081=>"000001000",
  26082=>"111000100",
  26083=>"001100110",
  26084=>"111100010",
  26085=>"101001101",
  26086=>"110100101",
  26087=>"011001100",
  26088=>"111001000",
  26089=>"111111011",
  26090=>"001011011",
  26091=>"100101101",
  26092=>"110011111",
  26093=>"011000011",
  26094=>"110011000",
  26095=>"101001011",
  26096=>"110111101",
  26097=>"001111000",
  26098=>"010010000",
  26099=>"110001100",
  26100=>"001001100",
  26101=>"011010101",
  26102=>"001101100",
  26103=>"100000101",
  26104=>"110000011",
  26105=>"011010000",
  26106=>"100110011",
  26107=>"110101011",
  26108=>"011100111",
  26109=>"000101100",
  26110=>"110000111",
  26111=>"010001111",
  26112=>"110111001",
  26113=>"010011011",
  26114=>"111011101",
  26115=>"111011111",
  26116=>"010010001",
  26117=>"100101111",
  26118=>"001010100",
  26119=>"011010010",
  26120=>"000101011",
  26121=>"001110111",
  26122=>"010011101",
  26123=>"000001101",
  26124=>"001010011",
  26125=>"000101001",
  26126=>"111000100",
  26127=>"110101010",
  26128=>"011011111",
  26129=>"010010010",
  26130=>"110010000",
  26131=>"100011111",
  26132=>"010010001",
  26133=>"101110100",
  26134=>"010110110",
  26135=>"000111011",
  26136=>"011101001",
  26137=>"101100111",
  26138=>"100111000",
  26139=>"101000001",
  26140=>"111000000",
  26141=>"101110001",
  26142=>"100101010",
  26143=>"011110101",
  26144=>"101100110",
  26145=>"011010011",
  26146=>"000000010",
  26147=>"110001001",
  26148=>"001100101",
  26149=>"110010101",
  26150=>"111110001",
  26151=>"100111001",
  26152=>"110110010",
  26153=>"110001001",
  26154=>"010011011",
  26155=>"110111010",
  26156=>"001100111",
  26157=>"100101111",
  26158=>"011011011",
  26159=>"011101011",
  26160=>"110010000",
  26161=>"011101001",
  26162=>"101010101",
  26163=>"111101001",
  26164=>"011101101",
  26165=>"111100100",
  26166=>"001000010",
  26167=>"011100001",
  26168=>"011101010",
  26169=>"011100110",
  26170=>"001101011",
  26171=>"000101100",
  26172=>"010100101",
  26173=>"010110000",
  26174=>"010011010",
  26175=>"010110110",
  26176=>"111000110",
  26177=>"001110010",
  26178=>"000001110",
  26179=>"010001000",
  26180=>"100101010",
  26181=>"100000011",
  26182=>"111010010",
  26183=>"100000100",
  26184=>"110100111",
  26185=>"010000111",
  26186=>"101000010",
  26187=>"010001010",
  26188=>"110001100",
  26189=>"101101010",
  26190=>"011001101",
  26191=>"111010010",
  26192=>"011111000",
  26193=>"010010011",
  26194=>"101010101",
  26195=>"001111011",
  26196=>"000001111",
  26197=>"100000011",
  26198=>"111110110",
  26199=>"011000011",
  26200=>"001000000",
  26201=>"011001011",
  26202=>"110110010",
  26203=>"001001010",
  26204=>"001100010",
  26205=>"010101100",
  26206=>"101011100",
  26207=>"111110000",
  26208=>"111011111",
  26209=>"010110111",
  26210=>"111010001",
  26211=>"011001011",
  26212=>"001110101",
  26213=>"001100100",
  26214=>"111100000",
  26215=>"111011111",
  26216=>"100110011",
  26217=>"101101110",
  26218=>"100101111",
  26219=>"000011001",
  26220=>"000011011",
  26221=>"111011010",
  26222=>"001111011",
  26223=>"000100110",
  26224=>"000011100",
  26225=>"000001000",
  26226=>"100010101",
  26227=>"011101011",
  26228=>"101010101",
  26229=>"011100011",
  26230=>"111111001",
  26231=>"000010111",
  26232=>"000111010",
  26233=>"110111011",
  26234=>"100111110",
  26235=>"111110101",
  26236=>"111111000",
  26237=>"011000001",
  26238=>"011010001",
  26239=>"000010111",
  26240=>"110111111",
  26241=>"101001111",
  26242=>"010101011",
  26243=>"110010000",
  26244=>"010110001",
  26245=>"100000000",
  26246=>"000110111",
  26247=>"001101101",
  26248=>"011010110",
  26249=>"111010111",
  26250=>"001100010",
  26251=>"011100001",
  26252=>"001111000",
  26253=>"100100111",
  26254=>"100100010",
  26255=>"100110111",
  26256=>"000010011",
  26257=>"101111100",
  26258=>"010110100",
  26259=>"100100110",
  26260=>"101011100",
  26261=>"111110101",
  26262=>"000111111",
  26263=>"101111001",
  26264=>"000111011",
  26265=>"010000110",
  26266=>"000000000",
  26267=>"011110000",
  26268=>"001100110",
  26269=>"010011111",
  26270=>"001111110",
  26271=>"011001011",
  26272=>"110101101",
  26273=>"100011000",
  26274=>"101100000",
  26275=>"110110100",
  26276=>"111111111",
  26277=>"000010001",
  26278=>"111000111",
  26279=>"111001010",
  26280=>"111110101",
  26281=>"100101001",
  26282=>"111000011",
  26283=>"011110100",
  26284=>"111110110",
  26285=>"000011001",
  26286=>"111000010",
  26287=>"101101111",
  26288=>"110100110",
  26289=>"101011001",
  26290=>"000010110",
  26291=>"001011101",
  26292=>"001101010",
  26293=>"111100001",
  26294=>"001010010",
  26295=>"110101011",
  26296=>"000111000",
  26297=>"000010101",
  26298=>"011001111",
  26299=>"001001001",
  26300=>"010011101",
  26301=>"001000001",
  26302=>"100110010",
  26303=>"010001111",
  26304=>"111011011",
  26305=>"110010101",
  26306=>"011110010",
  26307=>"001000000",
  26308=>"100110001",
  26309=>"110100011",
  26310=>"001110000",
  26311=>"100110010",
  26312=>"011000110",
  26313=>"010100110",
  26314=>"100000100",
  26315=>"000000101",
  26316=>"100000001",
  26317=>"111110000",
  26318=>"111110100",
  26319=>"111010111",
  26320=>"001111000",
  26321=>"101100010",
  26322=>"110010001",
  26323=>"000111100",
  26324=>"100011101",
  26325=>"100110000",
  26326=>"000000101",
  26327=>"000110110",
  26328=>"001001111",
  26329=>"001010111",
  26330=>"111100011",
  26331=>"110110010",
  26332=>"111101111",
  26333=>"010011011",
  26334=>"011100001",
  26335=>"001001111",
  26336=>"000000101",
  26337=>"001010111",
  26338=>"010101111",
  26339=>"011111111",
  26340=>"100111111",
  26341=>"000100101",
  26342=>"110101111",
  26343=>"010010111",
  26344=>"000101000",
  26345=>"110000100",
  26346=>"110100101",
  26347=>"011011111",
  26348=>"010111110",
  26349=>"000110000",
  26350=>"000000101",
  26351=>"111101110",
  26352=>"001100001",
  26353=>"000110001",
  26354=>"001001110",
  26355=>"001010001",
  26356=>"010101110",
  26357=>"010110110",
  26358=>"110101110",
  26359=>"111111101",
  26360=>"111100010",
  26361=>"110001011",
  26362=>"100000001",
  26363=>"100000100",
  26364=>"000001000",
  26365=>"010111010",
  26366=>"100100101",
  26367=>"001011111",
  26368=>"000110111",
  26369=>"010011111",
  26370=>"100111111",
  26371=>"001111000",
  26372=>"011001000",
  26373=>"101010101",
  26374=>"101001100",
  26375=>"001110110",
  26376=>"000110100",
  26377=>"011001101",
  26378=>"111000000",
  26379=>"101000100",
  26380=>"100101000",
  26381=>"001100101",
  26382=>"010010101",
  26383=>"001001010",
  26384=>"111111000",
  26385=>"000001001",
  26386=>"101001011",
  26387=>"101010101",
  26388=>"101101010",
  26389=>"100010011",
  26390=>"000110010",
  26391=>"111001110",
  26392=>"111011001",
  26393=>"111011010",
  26394=>"000100001",
  26395=>"000110011",
  26396=>"010100101",
  26397=>"001110000",
  26398=>"101001000",
  26399=>"111101101",
  26400=>"111110111",
  26401=>"100010100",
  26402=>"110100101",
  26403=>"010000100",
  26404=>"001100000",
  26405=>"000101100",
  26406=>"000110101",
  26407=>"010010010",
  26408=>"111111010",
  26409=>"111011100",
  26410=>"000001000",
  26411=>"110001001",
  26412=>"100000011",
  26413=>"100010000",
  26414=>"011111100",
  26415=>"111101010",
  26416=>"011011111",
  26417=>"000100100",
  26418=>"100001001",
  26419=>"010101110",
  26420=>"110001000",
  26421=>"111110010",
  26422=>"100010110",
  26423=>"001111101",
  26424=>"010110000",
  26425=>"110111101",
  26426=>"100000000",
  26427=>"100110100",
  26428=>"111111111",
  26429=>"101101110",
  26430=>"000001100",
  26431=>"000010101",
  26432=>"100110101",
  26433=>"000111010",
  26434=>"110110010",
  26435=>"111001110",
  26436=>"101110101",
  26437=>"001000011",
  26438=>"101110000",
  26439=>"010010000",
  26440=>"101100110",
  26441=>"100111110",
  26442=>"100000010",
  26443=>"100000001",
  26444=>"010111000",
  26445=>"111000110",
  26446=>"110000111",
  26447=>"010100001",
  26448=>"100001010",
  26449=>"001110101",
  26450=>"010010110",
  26451=>"110000111",
  26452=>"010100010",
  26453=>"110101100",
  26454=>"111111000",
  26455=>"000110110",
  26456=>"111110100",
  26457=>"101011010",
  26458=>"101011100",
  26459=>"111101101",
  26460=>"101011001",
  26461=>"101001110",
  26462=>"111000011",
  26463=>"001100111",
  26464=>"010000000",
  26465=>"100000110",
  26466=>"010011111",
  26467=>"100111100",
  26468=>"001100111",
  26469=>"000110110",
  26470=>"000000100",
  26471=>"100000110",
  26472=>"011011001",
  26473=>"100011000",
  26474=>"101111110",
  26475=>"110001101",
  26476=>"111000110",
  26477=>"111100110",
  26478=>"000011110",
  26479=>"010101110",
  26480=>"101011111",
  26481=>"000111101",
  26482=>"101100000",
  26483=>"110010110",
  26484=>"011000110",
  26485=>"000010111",
  26486=>"010111111",
  26487=>"001010000",
  26488=>"000110001",
  26489=>"110000101",
  26490=>"101001011",
  26491=>"000110010",
  26492=>"010000010",
  26493=>"101110001",
  26494=>"001010111",
  26495=>"100000001",
  26496=>"010111000",
  26497=>"001110010",
  26498=>"101101000",
  26499=>"001101000",
  26500=>"111110111",
  26501=>"101111100",
  26502=>"000011111",
  26503=>"011101000",
  26504=>"111011000",
  26505=>"000001010",
  26506=>"011001110",
  26507=>"000010001",
  26508=>"100101000",
  26509=>"110011011",
  26510=>"010101011",
  26511=>"011101000",
  26512=>"001100100",
  26513=>"010001100",
  26514=>"000001111",
  26515=>"111111111",
  26516=>"101110011",
  26517=>"001001000",
  26518=>"010110111",
  26519=>"100111010",
  26520=>"010111001",
  26521=>"011011000",
  26522=>"111100011",
  26523=>"101001000",
  26524=>"111110011",
  26525=>"110011011",
  26526=>"000000101",
  26527=>"110011101",
  26528=>"111100010",
  26529=>"111100100",
  26530=>"001011110",
  26531=>"000000100",
  26532=>"011000111",
  26533=>"111110111",
  26534=>"001010101",
  26535=>"110001100",
  26536=>"010000011",
  26537=>"000001010",
  26538=>"100101111",
  26539=>"101001110",
  26540=>"101011101",
  26541=>"001100000",
  26542=>"100001101",
  26543=>"011001011",
  26544=>"001110110",
  26545=>"111000000",
  26546=>"100001100",
  26547=>"101010000",
  26548=>"011010000",
  26549=>"111100000",
  26550=>"001011001",
  26551=>"100101011",
  26552=>"101011011",
  26553=>"010110000",
  26554=>"000000011",
  26555=>"001000001",
  26556=>"111000000",
  26557=>"100101001",
  26558=>"001010111",
  26559=>"111001000",
  26560=>"110101011",
  26561=>"110101000",
  26562=>"111101111",
  26563=>"100111110",
  26564=>"101111111",
  26565=>"001110101",
  26566=>"101001000",
  26567=>"000000110",
  26568=>"000010100",
  26569=>"110100001",
  26570=>"110111001",
  26571=>"011100101",
  26572=>"010010101",
  26573=>"001001000",
  26574=>"100000010",
  26575=>"010000011",
  26576=>"010111110",
  26577=>"000000101",
  26578=>"101011011",
  26579=>"001000000",
  26580=>"000010010",
  26581=>"011110110",
  26582=>"001001010",
  26583=>"001100111",
  26584=>"001111011",
  26585=>"100110111",
  26586=>"110000100",
  26587=>"000000011",
  26588=>"110000001",
  26589=>"101010111",
  26590=>"011110000",
  26591=>"110011111",
  26592=>"111000111",
  26593=>"111100110",
  26594=>"100010001",
  26595=>"011111111",
  26596=>"110100000",
  26597=>"010110010",
  26598=>"000010100",
  26599=>"100001010",
  26600=>"101110010",
  26601=>"110110011",
  26602=>"010000011",
  26603=>"001001101",
  26604=>"000000010",
  26605=>"010001000",
  26606=>"110010100",
  26607=>"110111011",
  26608=>"001000101",
  26609=>"010000110",
  26610=>"010110000",
  26611=>"110110111",
  26612=>"001101001",
  26613=>"010000111",
  26614=>"001100111",
  26615=>"101000001",
  26616=>"100001000",
  26617=>"001110000",
  26618=>"001100110",
  26619=>"111000001",
  26620=>"000000000",
  26621=>"010001011",
  26622=>"011100011",
  26623=>"101110111",
  26624=>"011001101",
  26625=>"011000010",
  26626=>"100010011",
  26627=>"010010000",
  26628=>"111000110",
  26629=>"110000110",
  26630=>"101000100",
  26631=>"100100001",
  26632=>"111110011",
  26633=>"011100011",
  26634=>"111000101",
  26635=>"111101000",
  26636=>"100111000",
  26637=>"011011101",
  26638=>"011111101",
  26639=>"000100010",
  26640=>"101011111",
  26641=>"011010011",
  26642=>"001110110",
  26643=>"010110110",
  26644=>"011101100",
  26645=>"101100111",
  26646=>"101111000",
  26647=>"010110011",
  26648=>"101100110",
  26649=>"101110011",
  26650=>"111000010",
  26651=>"101000001",
  26652=>"010111101",
  26653=>"100000101",
  26654=>"011000000",
  26655=>"100010111",
  26656=>"001100001",
  26657=>"100101011",
  26658=>"011111011",
  26659=>"000111110",
  26660=>"011010000",
  26661=>"110100011",
  26662=>"110101011",
  26663=>"010100001",
  26664=>"000101111",
  26665=>"111111010",
  26666=>"010100100",
  26667=>"011010000",
  26668=>"001111011",
  26669=>"110000110",
  26670=>"111011010",
  26671=>"000000000",
  26672=>"110110110",
  26673=>"000101001",
  26674=>"011011110",
  26675=>"000111000",
  26676=>"110011001",
  26677=>"011100001",
  26678=>"001001011",
  26679=>"010111011",
  26680=>"101101011",
  26681=>"000000000",
  26682=>"110100001",
  26683=>"001101001",
  26684=>"011001010",
  26685=>"111010111",
  26686=>"110111011",
  26687=>"000111111",
  26688=>"111100000",
  26689=>"011010000",
  26690=>"111110111",
  26691=>"001010100",
  26692=>"101011101",
  26693=>"010011001",
  26694=>"001000011",
  26695=>"100100100",
  26696=>"000001010",
  26697=>"001011100",
  26698=>"100111111",
  26699=>"010000001",
  26700=>"010110110",
  26701=>"110011000",
  26702=>"100101001",
  26703=>"110001101",
  26704=>"011000101",
  26705=>"000000101",
  26706=>"001011010",
  26707=>"100011110",
  26708=>"111110100",
  26709=>"001101100",
  26710=>"010111110",
  26711=>"100001101",
  26712=>"000100010",
  26713=>"101001011",
  26714=>"111100111",
  26715=>"100000001",
  26716=>"001110110",
  26717=>"000101001",
  26718=>"100001110",
  26719=>"010100100",
  26720=>"000010010",
  26721=>"001000110",
  26722=>"001101001",
  26723=>"000101011",
  26724=>"100101001",
  26725=>"010101000",
  26726=>"001011000",
  26727=>"111000110",
  26728=>"000110011",
  26729=>"101100011",
  26730=>"011000011",
  26731=>"111111011",
  26732=>"110001000",
  26733=>"001100101",
  26734=>"011000110",
  26735=>"100110001",
  26736=>"100110111",
  26737=>"111100000",
  26738=>"000110110",
  26739=>"010101001",
  26740=>"000000110",
  26741=>"001110101",
  26742=>"010010001",
  26743=>"000010110",
  26744=>"111011001",
  26745=>"000000110",
  26746=>"101011011",
  26747=>"101100100",
  26748=>"111011110",
  26749=>"001000111",
  26750=>"000111111",
  26751=>"101001100",
  26752=>"000101101",
  26753=>"110101010",
  26754=>"101001101",
  26755=>"110100111",
  26756=>"001001011",
  26757=>"111001101",
  26758=>"101110001",
  26759=>"010000100",
  26760=>"110111011",
  26761=>"100100110",
  26762=>"011101001",
  26763=>"011101110",
  26764=>"101100011",
  26765=>"000110001",
  26766=>"110111010",
  26767=>"010010000",
  26768=>"100011110",
  26769=>"001000110",
  26770=>"001001110",
  26771=>"111000010",
  26772=>"001110010",
  26773=>"000011001",
  26774=>"011010011",
  26775=>"111101011",
  26776=>"101101110",
  26777=>"001001010",
  26778=>"001011101",
  26779=>"111001110",
  26780=>"111000010",
  26781=>"100010000",
  26782=>"110101011",
  26783=>"011110111",
  26784=>"010101111",
  26785=>"011011101",
  26786=>"011000011",
  26787=>"101110000",
  26788=>"101110001",
  26789=>"110101110",
  26790=>"101111010",
  26791=>"111111001",
  26792=>"101100010",
  26793=>"001000100",
  26794=>"100010111",
  26795=>"100111011",
  26796=>"011110110",
  26797=>"110011011",
  26798=>"010010000",
  26799=>"000110101",
  26800=>"111111010",
  26801=>"000110011",
  26802=>"001001000",
  26803=>"011000000",
  26804=>"101010101",
  26805=>"100011001",
  26806=>"000111011",
  26807=>"110011010",
  26808=>"000111001",
  26809=>"101101100",
  26810=>"010010011",
  26811=>"100001011",
  26812=>"010111110",
  26813=>"001010000",
  26814=>"101001110",
  26815=>"110010011",
  26816=>"100010111",
  26817=>"101110101",
  26818=>"110100011",
  26819=>"011111111",
  26820=>"001001001",
  26821=>"000000001",
  26822=>"000000101",
  26823=>"101100010",
  26824=>"001011101",
  26825=>"010010000",
  26826=>"001011111",
  26827=>"110001101",
  26828=>"110101100",
  26829=>"110010110",
  26830=>"000101001",
  26831=>"010101101",
  26832=>"010000000",
  26833=>"101001001",
  26834=>"001101000",
  26835=>"101111100",
  26836=>"011001000",
  26837=>"110010011",
  26838=>"011110101",
  26839=>"000001011",
  26840=>"000011000",
  26841=>"111001000",
  26842=>"010001010",
  26843=>"111111101",
  26844=>"000110000",
  26845=>"110010111",
  26846=>"101010000",
  26847=>"000010000",
  26848=>"011110011",
  26849=>"101101011",
  26850=>"000101110",
  26851=>"000100001",
  26852=>"111000010",
  26853=>"010000111",
  26854=>"010010111",
  26855=>"011000111",
  26856=>"001101101",
  26857=>"011100101",
  26858=>"000100100",
  26859=>"000110011",
  26860=>"110111001",
  26861=>"100001001",
  26862=>"000101101",
  26863=>"010100110",
  26864=>"101111100",
  26865=>"001011100",
  26866=>"000101000",
  26867=>"011111001",
  26868=>"000110010",
  26869=>"000111111",
  26870=>"100110101",
  26871=>"110110101",
  26872=>"111110000",
  26873=>"101110101",
  26874=>"100111111",
  26875=>"100100100",
  26876=>"000000110",
  26877=>"011111000",
  26878=>"000101110",
  26879=>"000111111",
  26880=>"011111010",
  26881=>"011111111",
  26882=>"111110110",
  26883=>"111111010",
  26884=>"101011111",
  26885=>"110101101",
  26886=>"000011001",
  26887=>"100000001",
  26888=>"000100101",
  26889=>"111111101",
  26890=>"001101000",
  26891=>"111000101",
  26892=>"101110010",
  26893=>"000100001",
  26894=>"010111010",
  26895=>"000001111",
  26896=>"000000101",
  26897=>"111011011",
  26898=>"011000111",
  26899=>"100100110",
  26900=>"000011101",
  26901=>"100011010",
  26902=>"110010101",
  26903=>"000111111",
  26904=>"110001110",
  26905=>"101111011",
  26906=>"111001110",
  26907=>"100101110",
  26908=>"000010001",
  26909=>"011100101",
  26910=>"000111001",
  26911=>"001001001",
  26912=>"000011000",
  26913=>"100111101",
  26914=>"110010101",
  26915=>"110011100",
  26916=>"111111001",
  26917=>"100001011",
  26918=>"110101110",
  26919=>"001111110",
  26920=>"111000011",
  26921=>"100000010",
  26922=>"110000010",
  26923=>"111101000",
  26924=>"010011101",
  26925=>"011100100",
  26926=>"000011011",
  26927=>"010101110",
  26928=>"000001000",
  26929=>"101001111",
  26930=>"001000011",
  26931=>"010001110",
  26932=>"101111011",
  26933=>"001001010",
  26934=>"110010101",
  26935=>"000111011",
  26936=>"100101110",
  26937=>"011101011",
  26938=>"000100010",
  26939=>"001101010",
  26940=>"010000101",
  26941=>"100011111",
  26942=>"101101000",
  26943=>"000111101",
  26944=>"011100001",
  26945=>"110100001",
  26946=>"011000011",
  26947=>"011110110",
  26948=>"110010101",
  26949=>"000110011",
  26950=>"111010100",
  26951=>"010011111",
  26952=>"010110001",
  26953=>"111000111",
  26954=>"011111100",
  26955=>"000001111",
  26956=>"001111100",
  26957=>"110101011",
  26958=>"001100010",
  26959=>"100100110",
  26960=>"010101110",
  26961=>"111100010",
  26962=>"111111110",
  26963=>"010001001",
  26964=>"000010001",
  26965=>"111000010",
  26966=>"011011000",
  26967=>"100110100",
  26968=>"011100010",
  26969=>"000111111",
  26970=>"010011000",
  26971=>"100100000",
  26972=>"110001001",
  26973=>"010000011",
  26974=>"101110111",
  26975=>"010100101",
  26976=>"111001000",
  26977=>"011001000",
  26978=>"001011111",
  26979=>"100000000",
  26980=>"000011111",
  26981=>"111010010",
  26982=>"011110101",
  26983=>"011010111",
  26984=>"011010011",
  26985=>"000000011",
  26986=>"011000101",
  26987=>"101101010",
  26988=>"010100110",
  26989=>"100111110",
  26990=>"101001000",
  26991=>"011111100",
  26992=>"110000111",
  26993=>"000011011",
  26994=>"111111100",
  26995=>"100000011",
  26996=>"101001011",
  26997=>"000010011",
  26998=>"110010001",
  26999=>"000001110",
  27000=>"100110111",
  27001=>"011011010",
  27002=>"100011111",
  27003=>"010011000",
  27004=>"101111010",
  27005=>"110010101",
  27006=>"001101011",
  27007=>"110101100",
  27008=>"101001011",
  27009=>"000010000",
  27010=>"001001001",
  27011=>"010111110",
  27012=>"011000011",
  27013=>"100011111",
  27014=>"101101110",
  27015=>"111111100",
  27016=>"110100000",
  27017=>"101001011",
  27018=>"111010110",
  27019=>"100100111",
  27020=>"000010001",
  27021=>"111110111",
  27022=>"100110010",
  27023=>"110011001",
  27024=>"001011110",
  27025=>"001000110",
  27026=>"001110010",
  27027=>"110001011",
  27028=>"100111001",
  27029=>"000101010",
  27030=>"100110000",
  27031=>"100011000",
  27032=>"010100001",
  27033=>"001001111",
  27034=>"001111101",
  27035=>"010010011",
  27036=>"111011000",
  27037=>"101011001",
  27038=>"111000000",
  27039=>"111010110",
  27040=>"111110100",
  27041=>"100001010",
  27042=>"111101000",
  27043=>"110000011",
  27044=>"110101110",
  27045=>"000011001",
  27046=>"010101111",
  27047=>"010101010",
  27048=>"110010001",
  27049=>"100011000",
  27050=>"001101000",
  27051=>"011011010",
  27052=>"111001101",
  27053=>"110111110",
  27054=>"111111100",
  27055=>"010101010",
  27056=>"000110010",
  27057=>"011000010",
  27058=>"000011000",
  27059=>"011110010",
  27060=>"001100011",
  27061=>"111100011",
  27062=>"000111001",
  27063=>"111101111",
  27064=>"010000101",
  27065=>"111100011",
  27066=>"011000100",
  27067=>"001001000",
  27068=>"101001001",
  27069=>"000000001",
  27070=>"100010110",
  27071=>"111001101",
  27072=>"100000001",
  27073=>"110000000",
  27074=>"101110110",
  27075=>"010011100",
  27076=>"111010111",
  27077=>"001010010",
  27078=>"000100011",
  27079=>"111001000",
  27080=>"011100100",
  27081=>"001001000",
  27082=>"000000100",
  27083=>"011111111",
  27084=>"100110010",
  27085=>"000000100",
  27086=>"001100000",
  27087=>"111100110",
  27088=>"101111110",
  27089=>"110011000",
  27090=>"000011001",
  27091=>"101100111",
  27092=>"001100011",
  27093=>"010100011",
  27094=>"110100101",
  27095=>"011100011",
  27096=>"010000000",
  27097=>"110111011",
  27098=>"001000010",
  27099=>"000111000",
  27100=>"110011000",
  27101=>"001011101",
  27102=>"001110111",
  27103=>"010001110",
  27104=>"111011101",
  27105=>"001000011",
  27106=>"010010000",
  27107=>"000011000",
  27108=>"011101111",
  27109=>"111000110",
  27110=>"100001011",
  27111=>"011111011",
  27112=>"001100111",
  27113=>"000001100",
  27114=>"011001001",
  27115=>"110111111",
  27116=>"001100000",
  27117=>"011000001",
  27118=>"111010110",
  27119=>"101101000",
  27120=>"011010000",
  27121=>"101000000",
  27122=>"111101010",
  27123=>"000010101",
  27124=>"000010100",
  27125=>"000110001",
  27126=>"111111111",
  27127=>"011010001",
  27128=>"101110001",
  27129=>"110011000",
  27130=>"000100001",
  27131=>"110000001",
  27132=>"001000100",
  27133=>"111010101",
  27134=>"110100101",
  27135=>"000110101",
  27136=>"010111110",
  27137=>"001000110",
  27138=>"011110101",
  27139=>"000110101",
  27140=>"101101000",
  27141=>"101000110",
  27142=>"111100011",
  27143=>"010100001",
  27144=>"011001110",
  27145=>"001001001",
  27146=>"001100011",
  27147=>"001000101",
  27148=>"100101110",
  27149=>"010001111",
  27150=>"111101001",
  27151=>"101101000",
  27152=>"110000110",
  27153=>"000000111",
  27154=>"111010000",
  27155=>"001101110",
  27156=>"101001000",
  27157=>"001111100",
  27158=>"010111000",
  27159=>"110111111",
  27160=>"111101001",
  27161=>"010001111",
  27162=>"111101000",
  27163=>"100110001",
  27164=>"011111111",
  27165=>"110010011",
  27166=>"110110110",
  27167=>"000101110",
  27168=>"010001111",
  27169=>"010110111",
  27170=>"011011111",
  27171=>"000010001",
  27172=>"000001000",
  27173=>"000000110",
  27174=>"000001111",
  27175=>"000100101",
  27176=>"010000001",
  27177=>"000111111",
  27178=>"111011000",
  27179=>"101011011",
  27180=>"100010000",
  27181=>"100111111",
  27182=>"010100000",
  27183=>"010101100",
  27184=>"010011110",
  27185=>"110010010",
  27186=>"001101000",
  27187=>"101011100",
  27188=>"010001001",
  27189=>"000111100",
  27190=>"000101000",
  27191=>"000110110",
  27192=>"111001100",
  27193=>"010001111",
  27194=>"100010000",
  27195=>"101111010",
  27196=>"100001010",
  27197=>"011010001",
  27198=>"100100100",
  27199=>"011001010",
  27200=>"100100101",
  27201=>"001101000",
  27202=>"010100011",
  27203=>"000111111",
  27204=>"101001001",
  27205=>"100010100",
  27206=>"111010000",
  27207=>"101011001",
  27208=>"100100011",
  27209=>"000101001",
  27210=>"110111100",
  27211=>"000001000",
  27212=>"001010010",
  27213=>"000010010",
  27214=>"100011110",
  27215=>"011100011",
  27216=>"110101001",
  27217=>"111001000",
  27218=>"000101010",
  27219=>"000110010",
  27220=>"001010011",
  27221=>"100010101",
  27222=>"001011111",
  27223=>"001111010",
  27224=>"010111000",
  27225=>"111001111",
  27226=>"110010100",
  27227=>"001001001",
  27228=>"010000000",
  27229=>"101100100",
  27230=>"001010101",
  27231=>"010010000",
  27232=>"001001010",
  27233=>"010000001",
  27234=>"111101100",
  27235=>"011000011",
  27236=>"101010111",
  27237=>"100011010",
  27238=>"101010011",
  27239=>"000111100",
  27240=>"110000110",
  27241=>"001110000",
  27242=>"101011011",
  27243=>"101000011",
  27244=>"001101001",
  27245=>"010101100",
  27246=>"001101100",
  27247=>"001011010",
  27248=>"011100101",
  27249=>"010001000",
  27250=>"011000000",
  27251=>"001101100",
  27252=>"100010100",
  27253=>"100110010",
  27254=>"011011010",
  27255=>"100101001",
  27256=>"101010111",
  27257=>"110000101",
  27258=>"110000101",
  27259=>"111000001",
  27260=>"001010100",
  27261=>"011100010",
  27262=>"001100110",
  27263=>"111101011",
  27264=>"111111010",
  27265=>"110101001",
  27266=>"011111110",
  27267=>"101010010",
  27268=>"001111100",
  27269=>"000000000",
  27270=>"101110101",
  27271=>"111111111",
  27272=>"111101011",
  27273=>"010000000",
  27274=>"011010110",
  27275=>"010001001",
  27276=>"001111100",
  27277=>"011100000",
  27278=>"111000001",
  27279=>"111110101",
  27280=>"000011111",
  27281=>"010010110",
  27282=>"101110111",
  27283=>"100111110",
  27284=>"101111111",
  27285=>"100101111",
  27286=>"101111010",
  27287=>"100100100",
  27288=>"101001100",
  27289=>"010110000",
  27290=>"101010010",
  27291=>"011001000",
  27292=>"010011010",
  27293=>"110001101",
  27294=>"000011101",
  27295=>"100011011",
  27296=>"100011100",
  27297=>"010001001",
  27298=>"001000001",
  27299=>"101001101",
  27300=>"001111111",
  27301=>"110000000",
  27302=>"100000011",
  27303=>"100111110",
  27304=>"001001001",
  27305=>"100001001",
  27306=>"001100000",
  27307=>"011100010",
  27308=>"000110010",
  27309=>"101100001",
  27310=>"101011111",
  27311=>"110010110",
  27312=>"100110111",
  27313=>"101011001",
  27314=>"010110010",
  27315=>"100100100",
  27316=>"010100100",
  27317=>"000010101",
  27318=>"010011111",
  27319=>"011011100",
  27320=>"010001110",
  27321=>"111010110",
  27322=>"111110011",
  27323=>"100100011",
  27324=>"101111101",
  27325=>"100110010",
  27326=>"001001100",
  27327=>"101010110",
  27328=>"101001110",
  27329=>"000010110",
  27330=>"110001010",
  27331=>"010111010",
  27332=>"110011010",
  27333=>"110111000",
  27334=>"101010000",
  27335=>"000100000",
  27336=>"111001110",
  27337=>"000011000",
  27338=>"000101100",
  27339=>"000001001",
  27340=>"111001111",
  27341=>"110100000",
  27342=>"000001001",
  27343=>"000001110",
  27344=>"110101001",
  27345=>"010110001",
  27346=>"110111110",
  27347=>"111001000",
  27348=>"010010000",
  27349=>"000101001",
  27350=>"100110101",
  27351=>"001110111",
  27352=>"010011011",
  27353=>"110010100",
  27354=>"000111000",
  27355=>"101101101",
  27356=>"101101101",
  27357=>"101101010",
  27358=>"100101111",
  27359=>"010101011",
  27360=>"101111001",
  27361=>"111000100",
  27362=>"010010110",
  27363=>"101000111",
  27364=>"010010010",
  27365=>"111100010",
  27366=>"001100100",
  27367=>"100010001",
  27368=>"001001101",
  27369=>"111111111",
  27370=>"000110100",
  27371=>"100100110",
  27372=>"000000100",
  27373=>"101101101",
  27374=>"011010010",
  27375=>"110100011",
  27376=>"110101100",
  27377=>"100000110",
  27378=>"101010010",
  27379=>"100111010",
  27380=>"100111000",
  27381=>"001000010",
  27382=>"111011001",
  27383=>"000011111",
  27384=>"010000010",
  27385=>"000010011",
  27386=>"001100110",
  27387=>"001011000",
  27388=>"110110000",
  27389=>"000000101",
  27390=>"010001001",
  27391=>"010101101",
  27392=>"101010010",
  27393=>"001110011",
  27394=>"001101010",
  27395=>"101101100",
  27396=>"101000100",
  27397=>"000100110",
  27398=>"110100000",
  27399=>"110101110",
  27400=>"000010011",
  27401=>"110101100",
  27402=>"001000101",
  27403=>"110111000",
  27404=>"000001110",
  27405=>"110101111",
  27406=>"111000100",
  27407=>"011011000",
  27408=>"011001100",
  27409=>"011000011",
  27410=>"110101101",
  27411=>"001010011",
  27412=>"111100101",
  27413=>"000010010",
  27414=>"100011000",
  27415=>"110001110",
  27416=>"000101001",
  27417=>"011010000",
  27418=>"000100100",
  27419=>"100100011",
  27420=>"010001101",
  27421=>"111100010",
  27422=>"110100101",
  27423=>"010110110",
  27424=>"111010111",
  27425=>"010001001",
  27426=>"111010010",
  27427=>"111100011",
  27428=>"110010010",
  27429=>"000100000",
  27430=>"111110011",
  27431=>"111010100",
  27432=>"010010100",
  27433=>"011001000",
  27434=>"111101110",
  27435=>"111010001",
  27436=>"100100001",
  27437=>"000001110",
  27438=>"001101000",
  27439=>"100110011",
  27440=>"000101001",
  27441=>"001001000",
  27442=>"110001101",
  27443=>"000100100",
  27444=>"001011111",
  27445=>"100111001",
  27446=>"011100010",
  27447=>"111001000",
  27448=>"001111101",
  27449=>"110011110",
  27450=>"110011100",
  27451=>"100100010",
  27452=>"011000000",
  27453=>"001011001",
  27454=>"101111000",
  27455=>"100111111",
  27456=>"110110010",
  27457=>"000011110",
  27458=>"100111011",
  27459=>"100101001",
  27460=>"001101001",
  27461=>"101011111",
  27462=>"011110011",
  27463=>"011101000",
  27464=>"011011111",
  27465=>"100110100",
  27466=>"101001100",
  27467=>"111101000",
  27468=>"000010011",
  27469=>"101110111",
  27470=>"011111011",
  27471=>"001000000",
  27472=>"111011001",
  27473=>"010001111",
  27474=>"001001011",
  27475=>"000010001",
  27476=>"100011110",
  27477=>"110100000",
  27478=>"111111001",
  27479=>"001011001",
  27480=>"000000010",
  27481=>"001001011",
  27482=>"011101001",
  27483=>"001110001",
  27484=>"000011101",
  27485=>"100000001",
  27486=>"100011001",
  27487=>"001010001",
  27488=>"000100001",
  27489=>"011010001",
  27490=>"001100100",
  27491=>"110100110",
  27492=>"011001100",
  27493=>"000111101",
  27494=>"000000010",
  27495=>"011010101",
  27496=>"001001101",
  27497=>"011000100",
  27498=>"100001101",
  27499=>"101100110",
  27500=>"010000110",
  27501=>"001001001",
  27502=>"111111011",
  27503=>"111101001",
  27504=>"001101110",
  27505=>"001010100",
  27506=>"010010010",
  27507=>"111101101",
  27508=>"000010100",
  27509=>"010001001",
  27510=>"110000100",
  27511=>"110010000",
  27512=>"000000000",
  27513=>"111000111",
  27514=>"011101111",
  27515=>"001000010",
  27516=>"010110100",
  27517=>"010111100",
  27518=>"101001010",
  27519=>"001110110",
  27520=>"010110110",
  27521=>"101111010",
  27522=>"000100000",
  27523=>"111100011",
  27524=>"000010110",
  27525=>"110000011",
  27526=>"101101101",
  27527=>"101101011",
  27528=>"110110110",
  27529=>"000110100",
  27530=>"011111010",
  27531=>"110101000",
  27532=>"010110111",
  27533=>"000100011",
  27534=>"000010100",
  27535=>"100010010",
  27536=>"001010000",
  27537=>"110111000",
  27538=>"101110000",
  27539=>"011000011",
  27540=>"101010000",
  27541=>"100000000",
  27542=>"001110110",
  27543=>"101011011",
  27544=>"111011101",
  27545=>"000110100",
  27546=>"001111100",
  27547=>"110001011",
  27548=>"101101111",
  27549=>"101110101",
  27550=>"000111110",
  27551=>"100000011",
  27552=>"110000011",
  27553=>"010000011",
  27554=>"011100110",
  27555=>"011111101",
  27556=>"000110010",
  27557=>"000011010",
  27558=>"001001000",
  27559=>"110101111",
  27560=>"100111111",
  27561=>"110000101",
  27562=>"100100000",
  27563=>"010110001",
  27564=>"000100001",
  27565=>"100110111",
  27566=>"110001010",
  27567=>"001001000",
  27568=>"110110011",
  27569=>"111111101",
  27570=>"000110111",
  27571=>"101110100",
  27572=>"011010100",
  27573=>"001010100",
  27574=>"101110010",
  27575=>"111010110",
  27576=>"011101000",
  27577=>"111111101",
  27578=>"110001000",
  27579=>"100111000",
  27580=>"110100001",
  27581=>"011111110",
  27582=>"001010111",
  27583=>"101111011",
  27584=>"001101111",
  27585=>"000110000",
  27586=>"000010001",
  27587=>"111111010",
  27588=>"001110100",
  27589=>"011101101",
  27590=>"010001101",
  27591=>"110111100",
  27592=>"001110011",
  27593=>"001000110",
  27594=>"111001000",
  27595=>"001100000",
  27596=>"101100111",
  27597=>"111000000",
  27598=>"110011011",
  27599=>"011110001",
  27600=>"110000110",
  27601=>"110010100",
  27602=>"001010001",
  27603=>"010001110",
  27604=>"101001111",
  27605=>"101101011",
  27606=>"111101100",
  27607=>"010010011",
  27608=>"010100000",
  27609=>"110000100",
  27610=>"111111001",
  27611=>"110011000",
  27612=>"011001010",
  27613=>"110100011",
  27614=>"111000001",
  27615=>"110100100",
  27616=>"010001100",
  27617=>"101100001",
  27618=>"000011011",
  27619=>"000111000",
  27620=>"010010001",
  27621=>"010000011",
  27622=>"010101001",
  27623=>"101101101",
  27624=>"000001000",
  27625=>"011010001",
  27626=>"011100100",
  27627=>"100010111",
  27628=>"000111001",
  27629=>"100001000",
  27630=>"000011010",
  27631=>"000011000",
  27632=>"001010001",
  27633=>"000000101",
  27634=>"001111000",
  27635=>"100001111",
  27636=>"111110110",
  27637=>"000111011",
  27638=>"100110011",
  27639=>"001000000",
  27640=>"111100000",
  27641=>"010000001",
  27642=>"100100100",
  27643=>"000000001",
  27644=>"011100100",
  27645=>"011110001",
  27646=>"001100110",
  27647=>"110001111",
  27648=>"010111011",
  27649=>"001110000",
  27650=>"110111111",
  27651=>"111100111",
  27652=>"110011010",
  27653=>"000100101",
  27654=>"011111001",
  27655=>"110000101",
  27656=>"111011010",
  27657=>"000110111",
  27658=>"001110001",
  27659=>"000011101",
  27660=>"001110110",
  27661=>"101110001",
  27662=>"010000100",
  27663=>"000011011",
  27664=>"001000011",
  27665=>"010010010",
  27666=>"101111000",
  27667=>"001000011",
  27668=>"110110011",
  27669=>"010011110",
  27670=>"010100110",
  27671=>"011100001",
  27672=>"101100011",
  27673=>"110110010",
  27674=>"101111101",
  27675=>"101100111",
  27676=>"110111011",
  27677=>"010101010",
  27678=>"000100110",
  27679=>"010110000",
  27680=>"111110100",
  27681=>"101111100",
  27682=>"000001111",
  27683=>"010011100",
  27684=>"000110100",
  27685=>"100001011",
  27686=>"000110110",
  27687=>"011110111",
  27688=>"010100001",
  27689=>"100001100",
  27690=>"110011111",
  27691=>"111001100",
  27692=>"001111000",
  27693=>"110011011",
  27694=>"001000111",
  27695=>"101110001",
  27696=>"011001110",
  27697=>"100110001",
  27698=>"000111110",
  27699=>"101100110",
  27700=>"110110100",
  27701=>"000111000",
  27702=>"100011011",
  27703=>"101111100",
  27704=>"010111000",
  27705=>"101001001",
  27706=>"111101010",
  27707=>"101000011",
  27708=>"001010010",
  27709=>"111100000",
  27710=>"100000101",
  27711=>"101101011",
  27712=>"010010101",
  27713=>"001000011",
  27714=>"110100111",
  27715=>"110010101",
  27716=>"101000011",
  27717=>"101001011",
  27718=>"110000110",
  27719=>"110001010",
  27720=>"111100000",
  27721=>"111100001",
  27722=>"101110011",
  27723=>"010000010",
  27724=>"001100101",
  27725=>"100100001",
  27726=>"101011010",
  27727=>"100000101",
  27728=>"011111110",
  27729=>"010111111",
  27730=>"000000001",
  27731=>"101001101",
  27732=>"110100011",
  27733=>"001110010",
  27734=>"000110101",
  27735=>"011011011",
  27736=>"010011101",
  27737=>"101101001",
  27738=>"001011110",
  27739=>"010101100",
  27740=>"100011010",
  27741=>"111101000",
  27742=>"100101110",
  27743=>"010101010",
  27744=>"001110001",
  27745=>"010110101",
  27746=>"110101100",
  27747=>"010100010",
  27748=>"111100011",
  27749=>"101001010",
  27750=>"001111101",
  27751=>"010010100",
  27752=>"100110110",
  27753=>"000001000",
  27754=>"000000111",
  27755=>"101001001",
  27756=>"111001010",
  27757=>"000001101",
  27758=>"000111101",
  27759=>"111001001",
  27760=>"110111010",
  27761=>"011011001",
  27762=>"110101001",
  27763=>"001110110",
  27764=>"100011111",
  27765=>"101101110",
  27766=>"001100100",
  27767=>"111010110",
  27768=>"111010000",
  27769=>"010000001",
  27770=>"110110111",
  27771=>"111101100",
  27772=>"110010001",
  27773=>"111101100",
  27774=>"111100101",
  27775=>"000011011",
  27776=>"100001000",
  27777=>"111011010",
  27778=>"000000000",
  27779=>"010011101",
  27780=>"001001001",
  27781=>"111011000",
  27782=>"001111010",
  27783=>"100111100",
  27784=>"111101001",
  27785=>"011100011",
  27786=>"111000101",
  27787=>"000111000",
  27788=>"011100111",
  27789=>"100100101",
  27790=>"100110000",
  27791=>"111111001",
  27792=>"101001100",
  27793=>"001111010",
  27794=>"000001001",
  27795=>"110111100",
  27796=>"101100010",
  27797=>"111101010",
  27798=>"001100000",
  27799=>"110110001",
  27800=>"111011001",
  27801=>"111101101",
  27802=>"100000100",
  27803=>"000100001",
  27804=>"101100000",
  27805=>"111001111",
  27806=>"010010101",
  27807=>"010111101",
  27808=>"100011100",
  27809=>"110111101",
  27810=>"001101001",
  27811=>"111010100",
  27812=>"010111101",
  27813=>"100010001",
  27814=>"001100010",
  27815=>"100110001",
  27816=>"010100000",
  27817=>"011110000",
  27818=>"010010010",
  27819=>"011010011",
  27820=>"110001001",
  27821=>"111111010",
  27822=>"100111111",
  27823=>"100000110",
  27824=>"010111111",
  27825=>"110001101",
  27826=>"110111100",
  27827=>"100100000",
  27828=>"001101011",
  27829=>"111111111",
  27830=>"010010100",
  27831=>"011110110",
  27832=>"001100101",
  27833=>"101000001",
  27834=>"100011001",
  27835=>"011111010",
  27836=>"111010001",
  27837=>"001000001",
  27838=>"001011001",
  27839=>"001100110",
  27840=>"010101101",
  27841=>"000011000",
  27842=>"110011101",
  27843=>"010010010",
  27844=>"001101001",
  27845=>"101000111",
  27846=>"110011001",
  27847=>"011110010",
  27848=>"010011100",
  27849=>"011000000",
  27850=>"111010110",
  27851=>"001011100",
  27852=>"001100110",
  27853=>"001000010",
  27854=>"111111111",
  27855=>"101010111",
  27856=>"001101010",
  27857=>"011000010",
  27858=>"110011011",
  27859=>"110100011",
  27860=>"010000100",
  27861=>"110010111",
  27862=>"001001011",
  27863=>"100000100",
  27864=>"001100000",
  27865=>"000000010",
  27866=>"100000011",
  27867=>"010101011",
  27868=>"110000011",
  27869=>"110111000",
  27870=>"101111001",
  27871=>"011111111",
  27872=>"010110100",
  27873=>"011000111",
  27874=>"010010111",
  27875=>"001000100",
  27876=>"011001110",
  27877=>"101110110",
  27878=>"111100001",
  27879=>"100001011",
  27880=>"100001110",
  27881=>"010010110",
  27882=>"011010011",
  27883=>"001010110",
  27884=>"110110011",
  27885=>"010011000",
  27886=>"000100110",
  27887=>"110000010",
  27888=>"111001001",
  27889=>"111111111",
  27890=>"010010010",
  27891=>"100100100",
  27892=>"111000111",
  27893=>"110011111",
  27894=>"111110110",
  27895=>"000000100",
  27896=>"000100000",
  27897=>"011111010",
  27898=>"000101011",
  27899=>"011111110",
  27900=>"010110000",
  27901=>"001111100",
  27902=>"010111001",
  27903=>"101110000",
  27904=>"100100000",
  27905=>"011000100",
  27906=>"111000110",
  27907=>"101101100",
  27908=>"000100111",
  27909=>"101010101",
  27910=>"001011001",
  27911=>"101000111",
  27912=>"100001001",
  27913=>"100100111",
  27914=>"011101111",
  27915=>"111001110",
  27916=>"100110100",
  27917=>"010101100",
  27918=>"111110000",
  27919=>"001011110",
  27920=>"110011010",
  27921=>"100011101",
  27922=>"011011001",
  27923=>"110101100",
  27924=>"110110010",
  27925=>"010110000",
  27926=>"100101110",
  27927=>"101001000",
  27928=>"100101111",
  27929=>"101100010",
  27930=>"011000000",
  27931=>"010001001",
  27932=>"011001101",
  27933=>"110100100",
  27934=>"001001101",
  27935=>"000011000",
  27936=>"111110010",
  27937=>"001011000",
  27938=>"100110100",
  27939=>"100100011",
  27940=>"001110000",
  27941=>"000100001",
  27942=>"000011111",
  27943=>"111100011",
  27944=>"101010000",
  27945=>"101111111",
  27946=>"010001100",
  27947=>"111010111",
  27948=>"100011000",
  27949=>"110001101",
  27950=>"110111110",
  27951=>"110110101",
  27952=>"001001011",
  27953=>"101101010",
  27954=>"100000000",
  27955=>"100011010",
  27956=>"001100100",
  27957=>"001110100",
  27958=>"011010101",
  27959=>"111110100",
  27960=>"100001010",
  27961=>"010101100",
  27962=>"101110110",
  27963=>"100001110",
  27964=>"001011001",
  27965=>"100110110",
  27966=>"000001101",
  27967=>"000010000",
  27968=>"111101111",
  27969=>"001101100",
  27970=>"110011101",
  27971=>"000100001",
  27972=>"110000110",
  27973=>"100000010",
  27974=>"000011001",
  27975=>"000010010",
  27976=>"011010110",
  27977=>"100111011",
  27978=>"101110110",
  27979=>"100010001",
  27980=>"010011110",
  27981=>"000010111",
  27982=>"110010110",
  27983=>"110100000",
  27984=>"101000100",
  27985=>"011101110",
  27986=>"100101101",
  27987=>"001001010",
  27988=>"000000000",
  27989=>"110111101",
  27990=>"101100001",
  27991=>"010001101",
  27992=>"100000101",
  27993=>"001001010",
  27994=>"001100011",
  27995=>"111100101",
  27996=>"111010010",
  27997=>"001110001",
  27998=>"101110111",
  27999=>"001100100",
  28000=>"110110101",
  28001=>"100001111",
  28002=>"001100000",
  28003=>"010010101",
  28004=>"001100110",
  28005=>"010111000",
  28006=>"101100011",
  28007=>"000101000",
  28008=>"101000001",
  28009=>"001011101",
  28010=>"111110001",
  28011=>"010000011",
  28012=>"001000100",
  28013=>"001000111",
  28014=>"000101010",
  28015=>"010000011",
  28016=>"010000001",
  28017=>"001101100",
  28018=>"100010101",
  28019=>"000101011",
  28020=>"100000111",
  28021=>"011110100",
  28022=>"110000001",
  28023=>"001111101",
  28024=>"011101100",
  28025=>"000000000",
  28026=>"010101010",
  28027=>"010110111",
  28028=>"000011011",
  28029=>"111110010",
  28030=>"111111011",
  28031=>"000101010",
  28032=>"010100100",
  28033=>"100100101",
  28034=>"000111110",
  28035=>"101101011",
  28036=>"010111001",
  28037=>"100000101",
  28038=>"001001000",
  28039=>"100110101",
  28040=>"000100100",
  28041=>"001010100",
  28042=>"000010101",
  28043=>"111111111",
  28044=>"011000111",
  28045=>"111000011",
  28046=>"110011100",
  28047=>"111001010",
  28048=>"100001000",
  28049=>"110011101",
  28050=>"011011111",
  28051=>"000010111",
  28052=>"000110001",
  28053=>"010000010",
  28054=>"010000011",
  28055=>"001111010",
  28056=>"011001011",
  28057=>"111011011",
  28058=>"000011010",
  28059=>"010000000",
  28060=>"111111110",
  28061=>"000100010",
  28062=>"011010101",
  28063=>"110110111",
  28064=>"001001000",
  28065=>"101101111",
  28066=>"001001110",
  28067=>"101111101",
  28068=>"101100101",
  28069=>"000001011",
  28070=>"111000101",
  28071=>"001010011",
  28072=>"110010110",
  28073=>"100111000",
  28074=>"011000010",
  28075=>"000011100",
  28076=>"110110100",
  28077=>"010000101",
  28078=>"110100100",
  28079=>"100000101",
  28080=>"000111010",
  28081=>"111010011",
  28082=>"001001110",
  28083=>"100111111",
  28084=>"111000101",
  28085=>"000111110",
  28086=>"000001111",
  28087=>"010111011",
  28088=>"011010110",
  28089=>"111000000",
  28090=>"000100110",
  28091=>"101111110",
  28092=>"101001100",
  28093=>"010111111",
  28094=>"011001010",
  28095=>"100000001",
  28096=>"000100111",
  28097=>"011000100",
  28098=>"111001011",
  28099=>"000000011",
  28100=>"100110010",
  28101=>"001010101",
  28102=>"011001100",
  28103=>"111000010",
  28104=>"110001100",
  28105=>"011100100",
  28106=>"011000111",
  28107=>"101111111",
  28108=>"110010110",
  28109=>"011001100",
  28110=>"000100010",
  28111=>"100101000",
  28112=>"010100010",
  28113=>"011011011",
  28114=>"101000010",
  28115=>"011000111",
  28116=>"100110101",
  28117=>"010010010",
  28118=>"000001010",
  28119=>"011001000",
  28120=>"111101011",
  28121=>"011111111",
  28122=>"111100001",
  28123=>"010110010",
  28124=>"110000110",
  28125=>"101010001",
  28126=>"111011001",
  28127=>"111010000",
  28128=>"010000001",
  28129=>"010100100",
  28130=>"111100000",
  28131=>"100010000",
  28132=>"001000000",
  28133=>"100100011",
  28134=>"101111110",
  28135=>"101001010",
  28136=>"011010010",
  28137=>"000110010",
  28138=>"001111010",
  28139=>"011011011",
  28140=>"010100000",
  28141=>"011110000",
  28142=>"110110101",
  28143=>"110000010",
  28144=>"101110000",
  28145=>"011100010",
  28146=>"010101001",
  28147=>"001011111",
  28148=>"111010100",
  28149=>"100101000",
  28150=>"110100110",
  28151=>"101000101",
  28152=>"110100001",
  28153=>"000100101",
  28154=>"010011111",
  28155=>"100011110",
  28156=>"100101011",
  28157=>"010010011",
  28158=>"100100110",
  28159=>"110111011",
  28160=>"000010010",
  28161=>"000101011",
  28162=>"110000000",
  28163=>"111010111",
  28164=>"101101100",
  28165=>"111101001",
  28166=>"101100011",
  28167=>"000000011",
  28168=>"010001011",
  28169=>"101010100",
  28170=>"011100000",
  28171=>"100101100",
  28172=>"010100101",
  28173=>"110111011",
  28174=>"100110111",
  28175=>"110111111",
  28176=>"110100101",
  28177=>"111101101",
  28178=>"000011001",
  28179=>"001000011",
  28180=>"111101011",
  28181=>"110110010",
  28182=>"001110110",
  28183=>"000110100",
  28184=>"100101111",
  28185=>"000000011",
  28186=>"011110110",
  28187=>"011001100",
  28188=>"110010100",
  28189=>"110111011",
  28190=>"011111000",
  28191=>"011111111",
  28192=>"010101101",
  28193=>"110001010",
  28194=>"000000111",
  28195=>"101111011",
  28196=>"001110101",
  28197=>"111011101",
  28198=>"101111110",
  28199=>"101100011",
  28200=>"100001101",
  28201=>"001010111",
  28202=>"001001111",
  28203=>"101110001",
  28204=>"010100100",
  28205=>"011000000",
  28206=>"101100001",
  28207=>"100001100",
  28208=>"100100110",
  28209=>"111111100",
  28210=>"110110101",
  28211=>"101000111",
  28212=>"001011010",
  28213=>"000011000",
  28214=>"001100101",
  28215=>"001100111",
  28216=>"110111000",
  28217=>"111111010",
  28218=>"001101101",
  28219=>"110101001",
  28220=>"011110000",
  28221=>"001010111",
  28222=>"001000001",
  28223=>"000101111",
  28224=>"111100101",
  28225=>"000100001",
  28226=>"111100010",
  28227=>"010100000",
  28228=>"101001010",
  28229=>"100100000",
  28230=>"000101111",
  28231=>"100010100",
  28232=>"100111101",
  28233=>"011010001",
  28234=>"000101101",
  28235=>"001101101",
  28236=>"010001011",
  28237=>"000100100",
  28238=>"111010110",
  28239=>"011110010",
  28240=>"000000011",
  28241=>"011110000",
  28242=>"110001101",
  28243=>"001111001",
  28244=>"001010110",
  28245=>"100001100",
  28246=>"000000000",
  28247=>"111111111",
  28248=>"111111111",
  28249=>"100110100",
  28250=>"001010100",
  28251=>"110000100",
  28252=>"010110010",
  28253=>"100100100",
  28254=>"001111101",
  28255=>"010100001",
  28256=>"100010010",
  28257=>"101001101",
  28258=>"000000110",
  28259=>"010000100",
  28260=>"101010001",
  28261=>"111101111",
  28262=>"001011110",
  28263=>"011001011",
  28264=>"011111110",
  28265=>"011010111",
  28266=>"000101110",
  28267=>"110010011",
  28268=>"100100110",
  28269=>"110001100",
  28270=>"111111000",
  28271=>"011001111",
  28272=>"100011000",
  28273=>"000000000",
  28274=>"000101001",
  28275=>"100011111",
  28276=>"001110000",
  28277=>"111110110",
  28278=>"110100011",
  28279=>"001100001",
  28280=>"100000011",
  28281=>"011110101",
  28282=>"010101110",
  28283=>"100101011",
  28284=>"010010111",
  28285=>"110011111",
  28286=>"001110110",
  28287=>"111001100",
  28288=>"010111000",
  28289=>"110100010",
  28290=>"110101111",
  28291=>"010110011",
  28292=>"011111110",
  28293=>"100011011",
  28294=>"010100011",
  28295=>"001101110",
  28296=>"101000010",
  28297=>"111111011",
  28298=>"011001110",
  28299=>"110011110",
  28300=>"011010011",
  28301=>"110000000",
  28302=>"011010010",
  28303=>"111111101",
  28304=>"000110000",
  28305=>"110111001",
  28306=>"001100000",
  28307=>"010101000",
  28308=>"111111101",
  28309=>"101010101",
  28310=>"011011010",
  28311=>"000101110",
  28312=>"000110000",
  28313=>"110000000",
  28314=>"000000011",
  28315=>"000011110",
  28316=>"001001000",
  28317=>"111110110",
  28318=>"100101111",
  28319=>"000000110",
  28320=>"001111100",
  28321=>"110010110",
  28322=>"011100100",
  28323=>"001010001",
  28324=>"001101100",
  28325=>"010100010",
  28326=>"111101100",
  28327=>"001010010",
  28328=>"010010100",
  28329=>"101010010",
  28330=>"000110011",
  28331=>"001010101",
  28332=>"010010101",
  28333=>"100100111",
  28334=>"001000110",
  28335=>"010010000",
  28336=>"110011001",
  28337=>"100000001",
  28338=>"101001101",
  28339=>"000101100",
  28340=>"010111000",
  28341=>"111101110",
  28342=>"000001011",
  28343=>"000011110",
  28344=>"100111010",
  28345=>"001001010",
  28346=>"011111101",
  28347=>"101011111",
  28348=>"000101011",
  28349=>"011001000",
  28350=>"100111111",
  28351=>"000010011",
  28352=>"010010100",
  28353=>"011111000",
  28354=>"000011011",
  28355=>"100011101",
  28356=>"100011001",
  28357=>"011100101",
  28358=>"111101101",
  28359=>"111100111",
  28360=>"001001010",
  28361=>"011010001",
  28362=>"011111110",
  28363=>"101001011",
  28364=>"011001110",
  28365=>"000110101",
  28366=>"011000011",
  28367=>"110110101",
  28368=>"100101001",
  28369=>"101001000",
  28370=>"110110000",
  28371=>"000010011",
  28372=>"001111100",
  28373=>"110011000",
  28374=>"000001110",
  28375=>"000100101",
  28376=>"010001110",
  28377=>"111101011",
  28378=>"100011011",
  28379=>"010011000",
  28380=>"011111001",
  28381=>"110011110",
  28382=>"001011011",
  28383=>"010110111",
  28384=>"000111000",
  28385=>"010100110",
  28386=>"010101010",
  28387=>"000000000",
  28388=>"010000111",
  28389=>"000000000",
  28390=>"100011010",
  28391=>"110111000",
  28392=>"111011100",
  28393=>"001100011",
  28394=>"110000000",
  28395=>"001001011",
  28396=>"000000000",
  28397=>"000001100",
  28398=>"011010001",
  28399=>"100001011",
  28400=>"111000000",
  28401=>"010110000",
  28402=>"100001010",
  28403=>"111101101",
  28404=>"111101110",
  28405=>"100111011",
  28406=>"101000111",
  28407=>"110010010",
  28408=>"111100001",
  28409=>"101000100",
  28410=>"010001010",
  28411=>"010100101",
  28412=>"100100110",
  28413=>"100110111",
  28414=>"000110011",
  28415=>"111100101",
  28416=>"000011110",
  28417=>"010000010",
  28418=>"100001001",
  28419=>"101001011",
  28420=>"100011101",
  28421=>"001100101",
  28422=>"110000111",
  28423=>"100010000",
  28424=>"110101010",
  28425=>"111000001",
  28426=>"101111110",
  28427=>"010111001",
  28428=>"010010111",
  28429=>"001101010",
  28430=>"100011101",
  28431=>"001001110",
  28432=>"000101001",
  28433=>"000101111",
  28434=>"101010000",
  28435=>"001000011",
  28436=>"001100000",
  28437=>"000101000",
  28438=>"011110101",
  28439=>"100011000",
  28440=>"001011110",
  28441=>"101100110",
  28442=>"011111010",
  28443=>"010100101",
  28444=>"010001101",
  28445=>"001000101",
  28446=>"101110001",
  28447=>"001011100",
  28448=>"011101100",
  28449=>"100001001",
  28450=>"110110101",
  28451=>"001101001",
  28452=>"001010011",
  28453=>"010111011",
  28454=>"101010001",
  28455=>"010010100",
  28456=>"111111110",
  28457=>"111001011",
  28458=>"110011111",
  28459=>"111101001",
  28460=>"001010001",
  28461=>"000110101",
  28462=>"010001000",
  28463=>"011101010",
  28464=>"111010010",
  28465=>"100010001",
  28466=>"010111010",
  28467=>"111000110",
  28468=>"111100011",
  28469=>"010101100",
  28470=>"110100000",
  28471=>"111011101",
  28472=>"110110101",
  28473=>"001100010",
  28474=>"011101000",
  28475=>"110010011",
  28476=>"110000111",
  28477=>"111011111",
  28478=>"010011001",
  28479=>"011110110",
  28480=>"001101000",
  28481=>"100100101",
  28482=>"100100001",
  28483=>"111100100",
  28484=>"101000001",
  28485=>"011010000",
  28486=>"110100011",
  28487=>"111101100",
  28488=>"110011001",
  28489=>"001100001",
  28490=>"111010100",
  28491=>"001110100",
  28492=>"010101100",
  28493=>"000011111",
  28494=>"100000010",
  28495=>"100111110",
  28496=>"100011110",
  28497=>"110011011",
  28498=>"010001110",
  28499=>"111111100",
  28500=>"000111110",
  28501=>"011101001",
  28502=>"101010101",
  28503=>"010011100",
  28504=>"010010011",
  28505=>"100110010",
  28506=>"110101000",
  28507=>"101000110",
  28508=>"001111000",
  28509=>"101001011",
  28510=>"000100001",
  28511=>"100101101",
  28512=>"000100000",
  28513=>"110000011",
  28514=>"000011101",
  28515=>"110000001",
  28516=>"011011011",
  28517=>"101111100",
  28518=>"001011011",
  28519=>"111000001",
  28520=>"111110101",
  28521=>"101011101",
  28522=>"000000000",
  28523=>"111001000",
  28524=>"011000001",
  28525=>"001110010",
  28526=>"110001110",
  28527=>"100110110",
  28528=>"111011011",
  28529=>"010010011",
  28530=>"111000101",
  28531=>"110000010",
  28532=>"010100010",
  28533=>"011011011",
  28534=>"000101010",
  28535=>"101100000",
  28536=>"110100111",
  28537=>"001001001",
  28538=>"101000111",
  28539=>"010111011",
  28540=>"001001000",
  28541=>"110001111",
  28542=>"111111100",
  28543=>"010000011",
  28544=>"110100101",
  28545=>"111110101",
  28546=>"010111110",
  28547=>"000100001",
  28548=>"000010111",
  28549=>"001111100",
  28550=>"101100001",
  28551=>"111001101",
  28552=>"100101100",
  28553=>"010101101",
  28554=>"010001011",
  28555=>"000100011",
  28556=>"011001100",
  28557=>"111101101",
  28558=>"000000101",
  28559=>"100101010",
  28560=>"000011000",
  28561=>"110101111",
  28562=>"011110100",
  28563=>"110101111",
  28564=>"111011000",
  28565=>"101101111",
  28566=>"111101101",
  28567=>"100000000",
  28568=>"010111111",
  28569=>"011111100",
  28570=>"111011100",
  28571=>"101100011",
  28572=>"100101111",
  28573=>"001000001",
  28574=>"011110001",
  28575=>"000001001",
  28576=>"001110001",
  28577=>"110000011",
  28578=>"000001110",
  28579=>"001000011",
  28580=>"100010001",
  28581=>"111101100",
  28582=>"100010011",
  28583=>"010010010",
  28584=>"101010100",
  28585=>"010001000",
  28586=>"011100100",
  28587=>"000100000",
  28588=>"010110000",
  28589=>"010100110",
  28590=>"010000101",
  28591=>"001011101",
  28592=>"101000001",
  28593=>"010010100",
  28594=>"000101100",
  28595=>"011100111",
  28596=>"011000110",
  28597=>"101001100",
  28598=>"101101100",
  28599=>"111001110",
  28600=>"001100001",
  28601=>"000000001",
  28602=>"110111011",
  28603=>"000111001",
  28604=>"110100011",
  28605=>"110001001",
  28606=>"010001110",
  28607=>"011010001",
  28608=>"111000001",
  28609=>"110100000",
  28610=>"111001110",
  28611=>"001010101",
  28612=>"111011011",
  28613=>"010110010",
  28614=>"110000001",
  28615=>"011110110",
  28616=>"000011001",
  28617=>"010110110",
  28618=>"111100100",
  28619=>"011001010",
  28620=>"000000001",
  28621=>"101101000",
  28622=>"110000101",
  28623=>"010100001",
  28624=>"011001000",
  28625=>"010010100",
  28626=>"111001111",
  28627=>"010000111",
  28628=>"010111101",
  28629=>"001101100",
  28630=>"011001100",
  28631=>"111011011",
  28632=>"001011011",
  28633=>"101111100",
  28634=>"010001001",
  28635=>"010000000",
  28636=>"101100010",
  28637=>"010111000",
  28638=>"010100010",
  28639=>"010000010",
  28640=>"001010100",
  28641=>"101000001",
  28642=>"010010101",
  28643=>"000111001",
  28644=>"010111010",
  28645=>"000010000",
  28646=>"110111011",
  28647=>"001111101",
  28648=>"000001100",
  28649=>"011111101",
  28650=>"101001100",
  28651=>"010110100",
  28652=>"100100011",
  28653=>"001100011",
  28654=>"110000100",
  28655=>"001001111",
  28656=>"000101101",
  28657=>"110010111",
  28658=>"101010100",
  28659=>"001101101",
  28660=>"010011000",
  28661=>"111011111",
  28662=>"101000100",
  28663=>"000010010",
  28664=>"000011001",
  28665=>"000111000",
  28666=>"010101000",
  28667=>"110111001",
  28668=>"001101011",
  28669=>"001010110",
  28670=>"001100100",
  28671=>"000001101",
  28672=>"001100000",
  28673=>"001010000",
  28674=>"100110011",
  28675=>"111110111",
  28676=>"110111100",
  28677=>"100101001",
  28678=>"110000000",
  28679=>"010101001",
  28680=>"110101010",
  28681=>"001110011",
  28682=>"101110111",
  28683=>"111000000",
  28684=>"001001000",
  28685=>"001011110",
  28686=>"001011111",
  28687=>"101010110",
  28688=>"011001001",
  28689=>"011110110",
  28690=>"011100111",
  28691=>"111000111",
  28692=>"000000010",
  28693=>"000001001",
  28694=>"010011101",
  28695=>"000110010",
  28696=>"110000000",
  28697=>"111001110",
  28698=>"111011110",
  28699=>"000010010",
  28700=>"111011010",
  28701=>"010101111",
  28702=>"000101100",
  28703=>"110010101",
  28704=>"101010010",
  28705=>"101100001",
  28706=>"110010010",
  28707=>"111101001",
  28708=>"110111010",
  28709=>"100110011",
  28710=>"101010101",
  28711=>"110001010",
  28712=>"100110010",
  28713=>"000000110",
  28714=>"011011111",
  28715=>"001011111",
  28716=>"011000000",
  28717=>"100000000",
  28718=>"111100111",
  28719=>"101101011",
  28720=>"011110100",
  28721=>"011001011",
  28722=>"111011001",
  28723=>"110010000",
  28724=>"001000101",
  28725=>"111001101",
  28726=>"110010101",
  28727=>"010100000",
  28728=>"101110110",
  28729=>"101001110",
  28730=>"000010110",
  28731=>"110100000",
  28732=>"101111111",
  28733=>"000111001",
  28734=>"100100001",
  28735=>"110000010",
  28736=>"101010010",
  28737=>"000110111",
  28738=>"100001101",
  28739=>"001011001",
  28740=>"111111101",
  28741=>"011010010",
  28742=>"111111011",
  28743=>"001100001",
  28744=>"011001100",
  28745=>"111001010",
  28746=>"000101100",
  28747=>"100111111",
  28748=>"110010001",
  28749=>"001101010",
  28750=>"110111000",
  28751=>"100110111",
  28752=>"000010100",
  28753=>"110110111",
  28754=>"110100100",
  28755=>"000000000",
  28756=>"000110111",
  28757=>"110101110",
  28758=>"010010111",
  28759=>"110100010",
  28760=>"010011001",
  28761=>"010000100",
  28762=>"111011110",
  28763=>"011001010",
  28764=>"110110000",
  28765=>"001001010",
  28766=>"001001010",
  28767=>"101101111",
  28768=>"011100100",
  28769=>"011010001",
  28770=>"000111111",
  28771=>"100000100",
  28772=>"110010001",
  28773=>"001001001",
  28774=>"110101101",
  28775=>"111110011",
  28776=>"011000100",
  28777=>"111111001",
  28778=>"111111111",
  28779=>"010000001",
  28780=>"100001111",
  28781=>"011111101",
  28782=>"110010000",
  28783=>"110000001",
  28784=>"010100111",
  28785=>"010101000",
  28786=>"011010100",
  28787=>"010100000",
  28788=>"010001101",
  28789=>"000101010",
  28790=>"011110000",
  28791=>"011000100",
  28792=>"011001110",
  28793=>"000111000",
  28794=>"101110010",
  28795=>"001111000",
  28796=>"000010111",
  28797=>"010111011",
  28798=>"001100010",
  28799=>"100101111",
  28800=>"100101100",
  28801=>"000010011",
  28802=>"000111101",
  28803=>"110010000",
  28804=>"110100100",
  28805=>"011100010",
  28806=>"111110111",
  28807=>"000110110",
  28808=>"101000000",
  28809=>"000101010",
  28810=>"110000100",
  28811=>"110010001",
  28812=>"100000011",
  28813=>"011000000",
  28814=>"001101010",
  28815=>"111110110",
  28816=>"111011100",
  28817=>"011010001",
  28818=>"100000011",
  28819=>"011100100",
  28820=>"101101110",
  28821=>"011001011",
  28822=>"011000001",
  28823=>"010010101",
  28824=>"010011010",
  28825=>"101111010",
  28826=>"100100111",
  28827=>"111011001",
  28828=>"100010100",
  28829=>"011110101",
  28830=>"010110101",
  28831=>"001101101",
  28832=>"100000001",
  28833=>"110000110",
  28834=>"110110001",
  28835=>"010100011",
  28836=>"011011110",
  28837=>"111111110",
  28838=>"000000001",
  28839=>"000010001",
  28840=>"011001001",
  28841=>"100010110",
  28842=>"001110000",
  28843=>"000010000",
  28844=>"001000001",
  28845=>"111010011",
  28846=>"010101011",
  28847=>"001110010",
  28848=>"101011010",
  28849=>"001001000",
  28850=>"001100011",
  28851=>"100111000",
  28852=>"100000011",
  28853=>"101101110",
  28854=>"101110011",
  28855=>"100100001",
  28856=>"000000011",
  28857=>"001000000",
  28858=>"101010010",
  28859=>"100010111",
  28860=>"111010001",
  28861=>"001111001",
  28862=>"001000100",
  28863=>"010100001",
  28864=>"110000011",
  28865=>"101111001",
  28866=>"010101111",
  28867=>"001111011",
  28868=>"010011011",
  28869=>"101011001",
  28870=>"101001001",
  28871=>"100010000",
  28872=>"101000111",
  28873=>"110000111",
  28874=>"110011100",
  28875=>"100111100",
  28876=>"000010011",
  28877=>"010110011",
  28878=>"101011111",
  28879=>"010011100",
  28880=>"010111100",
  28881=>"011100001",
  28882=>"100010100",
  28883=>"100101101",
  28884=>"100001010",
  28885=>"000001101",
  28886=>"100101111",
  28887=>"011011111",
  28888=>"001101101",
  28889=>"100101111",
  28890=>"000000100",
  28891=>"100110001",
  28892=>"001011001",
  28893=>"001010110",
  28894=>"111111100",
  28895=>"111101001",
  28896=>"010011100",
  28897=>"010111011",
  28898=>"011111111",
  28899=>"010100000",
  28900=>"101011101",
  28901=>"001111101",
  28902=>"000010001",
  28903=>"010111010",
  28904=>"100110110",
  28905=>"000001100",
  28906=>"111110100",
  28907=>"010101100",
  28908=>"000101101",
  28909=>"010110001",
  28910=>"000000101",
  28911=>"010000110",
  28912=>"000100000",
  28913=>"000011000",
  28914=>"111000011",
  28915=>"011111000",
  28916=>"110111000",
  28917=>"010000001",
  28918=>"111000111",
  28919=>"010100000",
  28920=>"110010100",
  28921=>"111101101",
  28922=>"010010101",
  28923=>"000000100",
  28924=>"010000000",
  28925=>"001101001",
  28926=>"100100110",
  28927=>"111111110",
  28928=>"101001101",
  28929=>"010000010",
  28930=>"011110111",
  28931=>"001010101",
  28932=>"111010110",
  28933=>"110000101",
  28934=>"011011000",
  28935=>"010100111",
  28936=>"101001100",
  28937=>"100001001",
  28938=>"111001111",
  28939=>"111100110",
  28940=>"000101100",
  28941=>"111110000",
  28942=>"010011100",
  28943=>"100010001",
  28944=>"101001011",
  28945=>"000001101",
  28946=>"010110111",
  28947=>"101101101",
  28948=>"111011001",
  28949=>"011001000",
  28950=>"000010000",
  28951=>"100101001",
  28952=>"001111110",
  28953=>"001111110",
  28954=>"111110010",
  28955=>"001101101",
  28956=>"111101100",
  28957=>"010000010",
  28958=>"011011010",
  28959=>"000000001",
  28960=>"101000010",
  28961=>"101100010",
  28962=>"010111000",
  28963=>"110001010",
  28964=>"100110001",
  28965=>"110001001",
  28966=>"011000011",
  28967=>"110010001",
  28968=>"110000011",
  28969=>"011110101",
  28970=>"100100111",
  28971=>"011001110",
  28972=>"100100110",
  28973=>"100111100",
  28974=>"001001110",
  28975=>"011011100",
  28976=>"011011101",
  28977=>"100001100",
  28978=>"010100101",
  28979=>"001001011",
  28980=>"110000111",
  28981=>"000111001",
  28982=>"010100101",
  28983=>"011110111",
  28984=>"000010010",
  28985=>"010011111",
  28986=>"000111000",
  28987=>"000011001",
  28988=>"111100100",
  28989=>"100111001",
  28990=>"000111111",
  28991=>"101111011",
  28992=>"111001110",
  28993=>"111111001",
  28994=>"001001111",
  28995=>"100101011",
  28996=>"101101001",
  28997=>"100110010",
  28998=>"010100011",
  28999=>"110111001",
  29000=>"011110001",
  29001=>"000100000",
  29002=>"101000100",
  29003=>"011000011",
  29004=>"000101100",
  29005=>"101011100",
  29006=>"100111101",
  29007=>"101111110",
  29008=>"110111100",
  29009=>"101110011",
  29010=>"010100111",
  29011=>"110100000",
  29012=>"100000100",
  29013=>"101100001",
  29014=>"111010100",
  29015=>"110000010",
  29016=>"111101000",
  29017=>"100010001",
  29018=>"010110011",
  29019=>"000000111",
  29020=>"100101011",
  29021=>"011011100",
  29022=>"001001010",
  29023=>"110100101",
  29024=>"100010011",
  29025=>"010000001",
  29026=>"001000100",
  29027=>"110001000",
  29028=>"110011110",
  29029=>"000101111",
  29030=>"010011100",
  29031=>"010100101",
  29032=>"101101000",
  29033=>"010001111",
  29034=>"101110000",
  29035=>"001110111",
  29036=>"101001011",
  29037=>"110101010",
  29038=>"111100000",
  29039=>"010110111",
  29040=>"110011101",
  29041=>"111100111",
  29042=>"000100101",
  29043=>"100000111",
  29044=>"110001100",
  29045=>"011110101",
  29046=>"011011000",
  29047=>"100111110",
  29048=>"100001011",
  29049=>"011111111",
  29050=>"110100011",
  29051=>"111101000",
  29052=>"001111010",
  29053=>"001011011",
  29054=>"001000101",
  29055=>"110101101",
  29056=>"000110000",
  29057=>"000000110",
  29058=>"001110011",
  29059=>"101111011",
  29060=>"110001110",
  29061=>"011110000",
  29062=>"111110101",
  29063=>"000100101",
  29064=>"100101111",
  29065=>"000011000",
  29066=>"101000100",
  29067=>"111101101",
  29068=>"110100110",
  29069=>"101001011",
  29070=>"000001001",
  29071=>"111001010",
  29072=>"111010110",
  29073=>"111001100",
  29074=>"101100100",
  29075=>"110110111",
  29076=>"110000010",
  29077=>"010010111",
  29078=>"101011100",
  29079=>"100101000",
  29080=>"100010011",
  29081=>"100000001",
  29082=>"000100110",
  29083=>"001100101",
  29084=>"110111101",
  29085=>"110110000",
  29086=>"010100010",
  29087=>"011010001",
  29088=>"001101011",
  29089=>"111001011",
  29090=>"101010010",
  29091=>"010010010",
  29092=>"100010010",
  29093=>"100000000",
  29094=>"011011001",
  29095=>"011111000",
  29096=>"000111101",
  29097=>"010100001",
  29098=>"000000111",
  29099=>"000110111",
  29100=>"001111110",
  29101=>"000000010",
  29102=>"111110101",
  29103=>"110110010",
  29104=>"000011110",
  29105=>"001010101",
  29106=>"111111111",
  29107=>"010010111",
  29108=>"111011011",
  29109=>"010000011",
  29110=>"110011101",
  29111=>"101110001",
  29112=>"001000001",
  29113=>"011000010",
  29114=>"000100000",
  29115=>"100010011",
  29116=>"101000111",
  29117=>"010101100",
  29118=>"010101111",
  29119=>"101011111",
  29120=>"110000000",
  29121=>"110011000",
  29122=>"000100011",
  29123=>"100100000",
  29124=>"000000110",
  29125=>"110101111",
  29126=>"101101101",
  29127=>"100001001",
  29128=>"001010010",
  29129=>"110111001",
  29130=>"001000000",
  29131=>"111110001",
  29132=>"001100110",
  29133=>"100010110",
  29134=>"011010000",
  29135=>"000011001",
  29136=>"001110111",
  29137=>"010011111",
  29138=>"001100111",
  29139=>"110100111",
  29140=>"100101110",
  29141=>"110000011",
  29142=>"011100001",
  29143=>"111111001",
  29144=>"101010000",
  29145=>"110011010",
  29146=>"110001001",
  29147=>"101101001",
  29148=>"110001111",
  29149=>"110101001",
  29150=>"010110001",
  29151=>"111011110",
  29152=>"011101100",
  29153=>"001000101",
  29154=>"100001010",
  29155=>"101101111",
  29156=>"111101110",
  29157=>"000101111",
  29158=>"110110010",
  29159=>"111100000",
  29160=>"110110111",
  29161=>"010000011",
  29162=>"001100010",
  29163=>"010110111",
  29164=>"010001000",
  29165=>"111000001",
  29166=>"000110010",
  29167=>"010101001",
  29168=>"000010000",
  29169=>"000101001",
  29170=>"100000000",
  29171=>"100101010",
  29172=>"111101000",
  29173=>"000100011",
  29174=>"011110111",
  29175=>"100011101",
  29176=>"011100001",
  29177=>"100010000",
  29178=>"001100100",
  29179=>"111100011",
  29180=>"111100010",
  29181=>"111100110",
  29182=>"110011001",
  29183=>"111010001",
  29184=>"001111001",
  29185=>"101101010",
  29186=>"001111110",
  29187=>"110001010",
  29188=>"101101000",
  29189=>"110010011",
  29190=>"110110110",
  29191=>"010111001",
  29192=>"100000110",
  29193=>"100110000",
  29194=>"001101101",
  29195=>"101100111",
  29196=>"001001001",
  29197=>"001011000",
  29198=>"011100111",
  29199=>"010001111",
  29200=>"110001011",
  29201=>"010111010",
  29202=>"110111010",
  29203=>"111111110",
  29204=>"100100000",
  29205=>"111100000",
  29206=>"000001011",
  29207=>"111101100",
  29208=>"101000100",
  29209=>"000000000",
  29210=>"010101100",
  29211=>"010110010",
  29212=>"010000010",
  29213=>"101000110",
  29214=>"100110101",
  29215=>"101010011",
  29216=>"110011000",
  29217=>"011101010",
  29218=>"001000101",
  29219=>"110000000",
  29220=>"010000101",
  29221=>"100101011",
  29222=>"100101110",
  29223=>"101011110",
  29224=>"110010101",
  29225=>"000011010",
  29226=>"011001010",
  29227=>"000110101",
  29228=>"000000111",
  29229=>"001000101",
  29230=>"110011001",
  29231=>"100000100",
  29232=>"110100010",
  29233=>"111011010",
  29234=>"101101111",
  29235=>"100000111",
  29236=>"110000011",
  29237=>"111110000",
  29238=>"001000110",
  29239=>"111000111",
  29240=>"011101000",
  29241=>"010000001",
  29242=>"010001010",
  29243=>"010111010",
  29244=>"001101101",
  29245=>"000111011",
  29246=>"101010000",
  29247=>"011110000",
  29248=>"001001010",
  29249=>"110010101",
  29250=>"110011111",
  29251=>"100000001",
  29252=>"000100010",
  29253=>"011000001",
  29254=>"001001000",
  29255=>"111000011",
  29256=>"110001100",
  29257=>"111100000",
  29258=>"111010110",
  29259=>"110110111",
  29260=>"101001000",
  29261=>"000100000",
  29262=>"101010101",
  29263=>"100011000",
  29264=>"100101101",
  29265=>"110000000",
  29266=>"010001111",
  29267=>"111101000",
  29268=>"010000110",
  29269=>"011110001",
  29270=>"100010011",
  29271=>"011001010",
  29272=>"011111110",
  29273=>"011011101",
  29274=>"100100110",
  29275=>"010011001",
  29276=>"000110111",
  29277=>"110000101",
  29278=>"010100010",
  29279=>"001101001",
  29280=>"111101100",
  29281=>"010100001",
  29282=>"000110001",
  29283=>"000110000",
  29284=>"010100011",
  29285=>"100001100",
  29286=>"011110011",
  29287=>"000111101",
  29288=>"001001010",
  29289=>"101000000",
  29290=>"000001010",
  29291=>"010011111",
  29292=>"100000111",
  29293=>"110001001",
  29294=>"100100101",
  29295=>"101010010",
  29296=>"111000100",
  29297=>"000001110",
  29298=>"110101110",
  29299=>"100011100",
  29300=>"011100011",
  29301=>"000000101",
  29302=>"010111111",
  29303=>"111111001",
  29304=>"011100010",
  29305=>"111110110",
  29306=>"111000011",
  29307=>"110100000",
  29308=>"110101001",
  29309=>"100001100",
  29310=>"101011101",
  29311=>"110001100",
  29312=>"110010110",
  29313=>"100100110",
  29314=>"011101100",
  29315=>"110000110",
  29316=>"101000011",
  29317=>"101100101",
  29318=>"001010101",
  29319=>"011111011",
  29320=>"111100000",
  29321=>"011001101",
  29322=>"111111111",
  29323=>"110110000",
  29324=>"111011111",
  29325=>"110111101",
  29326=>"001001010",
  29327=>"100001111",
  29328=>"000001011",
  29329=>"010101101",
  29330=>"110101001",
  29331=>"000110010",
  29332=>"100100100",
  29333=>"000111110",
  29334=>"101001110",
  29335=>"010010101",
  29336=>"010011111",
  29337=>"100101010",
  29338=>"100001011",
  29339=>"111110000",
  29340=>"101110011",
  29341=>"110111100",
  29342=>"110101001",
  29343=>"100100111",
  29344=>"011111011",
  29345=>"011010011",
  29346=>"101010000",
  29347=>"100000111",
  29348=>"101101110",
  29349=>"101101111",
  29350=>"110000000",
  29351=>"000000000",
  29352=>"011111100",
  29353=>"101000101",
  29354=>"110000110",
  29355=>"011110000",
  29356=>"101001111",
  29357=>"000100111",
  29358=>"011001010",
  29359=>"101000100",
  29360=>"011000100",
  29361=>"001001111",
  29362=>"001011010",
  29363=>"000010000",
  29364=>"000101101",
  29365=>"000000000",
  29366=>"101010000",
  29367=>"111101100",
  29368=>"110000111",
  29369=>"111110010",
  29370=>"100010110",
  29371=>"100110011",
  29372=>"100010011",
  29373=>"000000000",
  29374=>"101010111",
  29375=>"010000010",
  29376=>"011000000",
  29377=>"100001000",
  29378=>"001011101",
  29379=>"110101100",
  29380=>"100001010",
  29381=>"010101100",
  29382=>"011000001",
  29383=>"001101010",
  29384=>"101101011",
  29385=>"011010111",
  29386=>"000011101",
  29387=>"100111011",
  29388=>"000101111",
  29389=>"100111010",
  29390=>"010000101",
  29391=>"000111000",
  29392=>"001000010",
  29393=>"011011100",
  29394=>"000101001",
  29395=>"110000100",
  29396=>"011011000",
  29397=>"100010111",
  29398=>"010111110",
  29399=>"010010010",
  29400=>"110011101",
  29401=>"010110011",
  29402=>"011000101",
  29403=>"001000100",
  29404=>"101101101",
  29405=>"001011111",
  29406=>"110110111",
  29407=>"111010100",
  29408=>"000001000",
  29409=>"010011011",
  29410=>"111010000",
  29411=>"010000111",
  29412=>"101001011",
  29413=>"010110110",
  29414=>"110100011",
  29415=>"110011110",
  29416=>"110100101",
  29417=>"011010001",
  29418=>"010001000",
  29419=>"000100110",
  29420=>"100000110",
  29421=>"000111010",
  29422=>"000111111",
  29423=>"111000111",
  29424=>"110001011",
  29425=>"000001100",
  29426=>"010011001",
  29427=>"011000110",
  29428=>"010010001",
  29429=>"111101111",
  29430=>"101101011",
  29431=>"111110010",
  29432=>"111110001",
  29433=>"001001111",
  29434=>"110100010",
  29435=>"111100001",
  29436=>"110001001",
  29437=>"101110000",
  29438=>"111111011",
  29439=>"100111110",
  29440=>"110111000",
  29441=>"111101010",
  29442=>"110100110",
  29443=>"111101000",
  29444=>"011110101",
  29445=>"011000111",
  29446=>"111100101",
  29447=>"011111001",
  29448=>"010110101",
  29449=>"010000101",
  29450=>"110011111",
  29451=>"111011111",
  29452=>"110101100",
  29453=>"010000000",
  29454=>"000111001",
  29455=>"011011001",
  29456=>"111000000",
  29457=>"111111000",
  29458=>"001000110",
  29459=>"110010111",
  29460=>"001011011",
  29461=>"110110001",
  29462=>"110101101",
  29463=>"000000010",
  29464=>"110111001",
  29465=>"101001110",
  29466=>"111011100",
  29467=>"011011110",
  29468=>"101010000",
  29469=>"010011011",
  29470=>"001001001",
  29471=>"111001000",
  29472=>"011111100",
  29473=>"101000001",
  29474=>"001100111",
  29475=>"010111110",
  29476=>"011000001",
  29477=>"011010111",
  29478=>"100001001",
  29479=>"001001100",
  29480=>"000100001",
  29481=>"010101000",
  29482=>"111111111",
  29483=>"000001100",
  29484=>"111110011",
  29485=>"101001000",
  29486=>"100110000",
  29487=>"000010000",
  29488=>"000000111",
  29489=>"110011001",
  29490=>"000100111",
  29491=>"100011111",
  29492=>"010101100",
  29493=>"111011011",
  29494=>"110011111",
  29495=>"100000011",
  29496=>"001100110",
  29497=>"000111000",
  29498=>"101110011",
  29499=>"000101000",
  29500=>"111100100",
  29501=>"000111111",
  29502=>"100000001",
  29503=>"111001100",
  29504=>"101110000",
  29505=>"110001000",
  29506=>"101100101",
  29507=>"011110010",
  29508=>"100101100",
  29509=>"111111101",
  29510=>"100111101",
  29511=>"101000110",
  29512=>"010100101",
  29513=>"010001000",
  29514=>"011010000",
  29515=>"011000101",
  29516=>"011100001",
  29517=>"010100001",
  29518=>"001111011",
  29519=>"110011011",
  29520=>"000101110",
  29521=>"100101100",
  29522=>"000000011",
  29523=>"000110011",
  29524=>"011011110",
  29525=>"000111000",
  29526=>"001000101",
  29527=>"110010110",
  29528=>"101110011",
  29529=>"110101100",
  29530=>"011110101",
  29531=>"101111100",
  29532=>"100101100",
  29533=>"101111111",
  29534=>"000011110",
  29535=>"110011000",
  29536=>"011001101",
  29537=>"110110000",
  29538=>"110101110",
  29539=>"101110111",
  29540=>"001000000",
  29541=>"100110111",
  29542=>"110010101",
  29543=>"001100001",
  29544=>"111010100",
  29545=>"001111010",
  29546=>"111100001",
  29547=>"000000111",
  29548=>"011010001",
  29549=>"001111001",
  29550=>"000010011",
  29551=>"011110101",
  29552=>"111110110",
  29553=>"110011010",
  29554=>"000110000",
  29555=>"101001000",
  29556=>"110101111",
  29557=>"100001100",
  29558=>"011000111",
  29559=>"111011101",
  29560=>"111000100",
  29561=>"101000010",
  29562=>"110010110",
  29563=>"111000000",
  29564=>"000010001",
  29565=>"101110111",
  29566=>"011000001",
  29567=>"011010001",
  29568=>"011100001",
  29569=>"100101111",
  29570=>"011111101",
  29571=>"101101100",
  29572=>"110000100",
  29573=>"110101011",
  29574=>"101100111",
  29575=>"000001011",
  29576=>"001001010",
  29577=>"011110000",
  29578=>"101010100",
  29579=>"111001101",
  29580=>"000001100",
  29581=>"001001011",
  29582=>"101110100",
  29583=>"011110110",
  29584=>"100010000",
  29585=>"100100000",
  29586=>"000001111",
  29587=>"110001010",
  29588=>"011010010",
  29589=>"111010111",
  29590=>"111111001",
  29591=>"101001010",
  29592=>"001101000",
  29593=>"010000101",
  29594=>"000000111",
  29595=>"000001101",
  29596=>"101001000",
  29597=>"001010100",
  29598=>"000110011",
  29599=>"110101100",
  29600=>"101110001",
  29601=>"111001011",
  29602=>"010011011",
  29603=>"101111011",
  29604=>"011000000",
  29605=>"011110110",
  29606=>"101000111",
  29607=>"110100001",
  29608=>"010110011",
  29609=>"000111001",
  29610=>"100010101",
  29611=>"000000010",
  29612=>"001010001",
  29613=>"000010101",
  29614=>"000100000",
  29615=>"010101000",
  29616=>"111110101",
  29617=>"111111010",
  29618=>"110000111",
  29619=>"011100110",
  29620=>"101000010",
  29621=>"001000110",
  29622=>"000011000",
  29623=>"000010101",
  29624=>"111011100",
  29625=>"001100111",
  29626=>"110010010",
  29627=>"100001001",
  29628=>"001001000",
  29629=>"100101111",
  29630=>"010001100",
  29631=>"100001011",
  29632=>"001110101",
  29633=>"001000001",
  29634=>"000010101",
  29635=>"000110111",
  29636=>"000110010",
  29637=>"101100100",
  29638=>"100111100",
  29639=>"101101111",
  29640=>"000101111",
  29641=>"110110101",
  29642=>"010101001",
  29643=>"001110000",
  29644=>"110101000",
  29645=>"110100111",
  29646=>"000000001",
  29647=>"010011000",
  29648=>"011100011",
  29649=>"001111001",
  29650=>"001001000",
  29651=>"011010000",
  29652=>"110011110",
  29653=>"111101111",
  29654=>"001000000",
  29655=>"101010101",
  29656=>"110101000",
  29657=>"101100111",
  29658=>"010010010",
  29659=>"000101000",
  29660=>"011011011",
  29661=>"010000001",
  29662=>"111110011",
  29663=>"010010101",
  29664=>"000010110",
  29665=>"001111110",
  29666=>"111111100",
  29667=>"110101100",
  29668=>"010110010",
  29669=>"111001100",
  29670=>"001111111",
  29671=>"011110100",
  29672=>"001000100",
  29673=>"001110001",
  29674=>"101000101",
  29675=>"101101111",
  29676=>"000011000",
  29677=>"000001110",
  29678=>"110000011",
  29679=>"100111110",
  29680=>"101000111",
  29681=>"000011001",
  29682=>"111000110",
  29683=>"110100000",
  29684=>"100010010",
  29685=>"000001101",
  29686=>"101010010",
  29687=>"101011010",
  29688=>"000101111",
  29689=>"110010001",
  29690=>"111101110",
  29691=>"100010001",
  29692=>"000010000",
  29693=>"110110110",
  29694=>"101010010",
  29695=>"101110011",
  29696=>"101111000",
  29697=>"001111110",
  29698=>"100000001",
  29699=>"011101111",
  29700=>"001111000",
  29701=>"100011000",
  29702=>"000011111",
  29703=>"111000111",
  29704=>"110011000",
  29705=>"011011011",
  29706=>"000001011",
  29707=>"000010111",
  29708=>"000100000",
  29709=>"011101111",
  29710=>"010101011",
  29711=>"010101010",
  29712=>"101101010",
  29713=>"001111010",
  29714=>"011110010",
  29715=>"010000010",
  29716=>"111011111",
  29717=>"101100000",
  29718=>"111101100",
  29719=>"111111111",
  29720=>"110101010",
  29721=>"010110100",
  29722=>"001001010",
  29723=>"011111101",
  29724=>"000100000",
  29725=>"111111100",
  29726=>"111111010",
  29727=>"000111111",
  29728=>"111101000",
  29729=>"101111101",
  29730=>"010011110",
  29731=>"111011111",
  29732=>"000110101",
  29733=>"010101000",
  29734=>"101111100",
  29735=>"000010010",
  29736=>"011011011",
  29737=>"110011110",
  29738=>"100101101",
  29739=>"000110010",
  29740=>"000011110",
  29741=>"010010101",
  29742=>"010101010",
  29743=>"100111110",
  29744=>"100001011",
  29745=>"111010010",
  29746=>"100010101",
  29747=>"001111111",
  29748=>"001101111",
  29749=>"010010000",
  29750=>"101000011",
  29751=>"101101010",
  29752=>"000100010",
  29753=>"110100000",
  29754=>"001110010",
  29755=>"010011110",
  29756=>"011010001",
  29757=>"100010101",
  29758=>"010000010",
  29759=>"001001011",
  29760=>"001111101",
  29761=>"000110010",
  29762=>"000000000",
  29763=>"001101011",
  29764=>"000000001",
  29765=>"100010001",
  29766=>"110101110",
  29767=>"011000001",
  29768=>"111100001",
  29769=>"000011101",
  29770=>"011000000",
  29771=>"110001000",
  29772=>"100110110",
  29773=>"101111110",
  29774=>"111110000",
  29775=>"010011000",
  29776=>"000000010",
  29777=>"000100000",
  29778=>"111101010",
  29779=>"101101111",
  29780=>"011110000",
  29781=>"010110010",
  29782=>"111011100",
  29783=>"011100011",
  29784=>"100001101",
  29785=>"001000010",
  29786=>"100010100",
  29787=>"100110101",
  29788=>"101000111",
  29789=>"000001100",
  29790=>"011110010",
  29791=>"001000001",
  29792=>"111101011",
  29793=>"100010101",
  29794=>"000011101",
  29795=>"101101011",
  29796=>"010111010",
  29797=>"001111111",
  29798=>"010111110",
  29799=>"001001000",
  29800=>"100011110",
  29801=>"011110101",
  29802=>"111101101",
  29803=>"111010011",
  29804=>"101100111",
  29805=>"010100000",
  29806=>"101110111",
  29807=>"100010010",
  29808=>"000000100",
  29809=>"101001001",
  29810=>"000111000",
  29811=>"010101010",
  29812=>"101000111",
  29813=>"111101001",
  29814=>"000111111",
  29815=>"111001110",
  29816=>"111101001",
  29817=>"001100111",
  29818=>"010000100",
  29819=>"101100111",
  29820=>"010011010",
  29821=>"000000001",
  29822=>"000011011",
  29823=>"100011101",
  29824=>"000101101",
  29825=>"110100100",
  29826=>"011000010",
  29827=>"100000110",
  29828=>"000000001",
  29829=>"100011110",
  29830=>"011000111",
  29831=>"010011111",
  29832=>"101100101",
  29833=>"001000011",
  29834=>"111011010",
  29835=>"010100101",
  29836=>"111001100",
  29837=>"010001001",
  29838=>"111010000",
  29839=>"110110010",
  29840=>"011000111",
  29841=>"110011111",
  29842=>"011011000",
  29843=>"110010101",
  29844=>"000010000",
  29845=>"000100111",
  29846=>"110011000",
  29847=>"100000110",
  29848=>"010111011",
  29849=>"001011000",
  29850=>"101000000",
  29851=>"101111010",
  29852=>"101101001",
  29853=>"111100010",
  29854=>"100011111",
  29855=>"111111000",
  29856=>"010101111",
  29857=>"110111010",
  29858=>"010110111",
  29859=>"000000100",
  29860=>"011011110",
  29861=>"000100001",
  29862=>"000111001",
  29863=>"000010111",
  29864=>"110101000",
  29865=>"000000101",
  29866=>"000100011",
  29867=>"011100001",
  29868=>"001111111",
  29869=>"100100101",
  29870=>"000100010",
  29871=>"010110011",
  29872=>"100101110",
  29873=>"010111110",
  29874=>"111100100",
  29875=>"011000100",
  29876=>"110110001",
  29877=>"110100001",
  29878=>"110001011",
  29879=>"010000101",
  29880=>"100011111",
  29881=>"001101110",
  29882=>"111010001",
  29883=>"101010100",
  29884=>"001001011",
  29885=>"110110111",
  29886=>"000010000",
  29887=>"010001000",
  29888=>"110011110",
  29889=>"101101111",
  29890=>"010010111",
  29891=>"011100010",
  29892=>"111111110",
  29893=>"001010010",
  29894=>"110100110",
  29895=>"000010110",
  29896=>"101100111",
  29897=>"011000010",
  29898=>"000101101",
  29899=>"011111010",
  29900=>"100001111",
  29901=>"000011111",
  29902=>"001011000",
  29903=>"001000101",
  29904=>"001010101",
  29905=>"010111101",
  29906=>"101100110",
  29907=>"001100111",
  29908=>"110010110",
  29909=>"100011111",
  29910=>"111011110",
  29911=>"100111000",
  29912=>"100111010",
  29913=>"110101011",
  29914=>"010111101",
  29915=>"000110110",
  29916=>"000101010",
  29917=>"100101100",
  29918=>"000010000",
  29919=>"100111101",
  29920=>"000100000",
  29921=>"000101001",
  29922=>"110000011",
  29923=>"100101100",
  29924=>"001011011",
  29925=>"110000100",
  29926=>"111110001",
  29927=>"111110101",
  29928=>"001000011",
  29929=>"000000000",
  29930=>"000011011",
  29931=>"101111111",
  29932=>"000001000",
  29933=>"100100110",
  29934=>"100011100",
  29935=>"100000100",
  29936=>"101110011",
  29937=>"010101101",
  29938=>"011001010",
  29939=>"111001000",
  29940=>"110001110",
  29941=>"000011000",
  29942=>"010001100",
  29943=>"011100000",
  29944=>"100011011",
  29945=>"100111100",
  29946=>"101110110",
  29947=>"110001110",
  29948=>"101110101",
  29949=>"001110011",
  29950=>"001010101",
  29951=>"110100001",
  29952=>"110000011",
  29953=>"010001110",
  29954=>"010101010",
  29955=>"100011001",
  29956=>"000010101",
  29957=>"010000100",
  29958=>"000010010",
  29959=>"101011101",
  29960=>"111110101",
  29961=>"111011001",
  29962=>"101011001",
  29963=>"011110110",
  29964=>"011110111",
  29965=>"110010010",
  29966=>"001110010",
  29967=>"000000101",
  29968=>"011110100",
  29969=>"001100001",
  29970=>"000100011",
  29971=>"011011100",
  29972=>"000011100",
  29973=>"010100000",
  29974=>"001000011",
  29975=>"100001011",
  29976=>"110110110",
  29977=>"110101011",
  29978=>"101101111",
  29979=>"110010010",
  29980=>"001001110",
  29981=>"011110111",
  29982=>"000010001",
  29983=>"000111101",
  29984=>"010010010",
  29985=>"000110110",
  29986=>"101111111",
  29987=>"101101111",
  29988=>"011001110",
  29989=>"010010001",
  29990=>"000100110",
  29991=>"110110100",
  29992=>"010111101",
  29993=>"100110010",
  29994=>"101010110",
  29995=>"100000100",
  29996=>"111010010",
  29997=>"101100110",
  29998=>"001000011",
  29999=>"101011101",
  30000=>"110101000",
  30001=>"101100110",
  30002=>"101000000",
  30003=>"101111000",
  30004=>"001011111",
  30005=>"100001000",
  30006=>"011011111",
  30007=>"100010110",
  30008=>"010101110",
  30009=>"010100011",
  30010=>"111011111",
  30011=>"100000001",
  30012=>"100100111",
  30013=>"100111000",
  30014=>"111100011",
  30015=>"111011011",
  30016=>"111110101",
  30017=>"101001100",
  30018=>"010100001",
  30019=>"011111010",
  30020=>"000001000",
  30021=>"100001110",
  30022=>"000101100",
  30023=>"110101001",
  30024=>"110010010",
  30025=>"000001100",
  30026=>"101010000",
  30027=>"011011110",
  30028=>"100010101",
  30029=>"010010110",
  30030=>"011110101",
  30031=>"111101111",
  30032=>"001111010",
  30033=>"010111001",
  30034=>"000011100",
  30035=>"001000001",
  30036=>"101111101",
  30037=>"100110111",
  30038=>"110100111",
  30039=>"000000011",
  30040=>"010100101",
  30041=>"101001100",
  30042=>"110001111",
  30043=>"000000011",
  30044=>"100000111",
  30045=>"010001010",
  30046=>"110111101",
  30047=>"001010010",
  30048=>"110001110",
  30049=>"010101010",
  30050=>"111100000",
  30051=>"011111111",
  30052=>"000010000",
  30053=>"010100010",
  30054=>"000010100",
  30055=>"000000110",
  30056=>"001101010",
  30057=>"000000101",
  30058=>"011001111",
  30059=>"000000101",
  30060=>"000011000",
  30061=>"110110110",
  30062=>"001000011",
  30063=>"101010101",
  30064=>"011001010",
  30065=>"100000001",
  30066=>"011110010",
  30067=>"110001000",
  30068=>"111110110",
  30069=>"101100000",
  30070=>"111111111",
  30071=>"110110101",
  30072=>"011110100",
  30073=>"010000100",
  30074=>"100100101",
  30075=>"001001011",
  30076=>"010110101",
  30077=>"100010011",
  30078=>"011011010",
  30079=>"011100110",
  30080=>"010100110",
  30081=>"010110101",
  30082=>"111110111",
  30083=>"111110001",
  30084=>"001101001",
  30085=>"000111001",
  30086=>"111111111",
  30087=>"110101011",
  30088=>"110110001",
  30089=>"110111111",
  30090=>"000110001",
  30091=>"000000100",
  30092=>"001011000",
  30093=>"000110010",
  30094=>"001101110",
  30095=>"001101010",
  30096=>"111001010",
  30097=>"000001001",
  30098=>"101111001",
  30099=>"000000010",
  30100=>"111000110",
  30101=>"111011000",
  30102=>"110111111",
  30103=>"111111100",
  30104=>"101011111",
  30105=>"000110111",
  30106=>"101000010",
  30107=>"111111010",
  30108=>"011001111",
  30109=>"000000101",
  30110=>"001111110",
  30111=>"100001000",
  30112=>"100111100",
  30113=>"100000000",
  30114=>"110010000",
  30115=>"011000101",
  30116=>"011000110",
  30117=>"001111011",
  30118=>"000100111",
  30119=>"111111110",
  30120=>"111011011",
  30121=>"111101110",
  30122=>"001100000",
  30123=>"111010110",
  30124=>"101111011",
  30125=>"000011101",
  30126=>"000001011",
  30127=>"011011101",
  30128=>"011110111",
  30129=>"010011001",
  30130=>"000011100",
  30131=>"011010111",
  30132=>"000110001",
  30133=>"000111111",
  30134=>"100011001",
  30135=>"001100001",
  30136=>"001000101",
  30137=>"001011101",
  30138=>"000100000",
  30139=>"111001000",
  30140=>"110000100",
  30141=>"110110010",
  30142=>"001000000",
  30143=>"111101011",
  30144=>"000000010",
  30145=>"011000100",
  30146=>"000111000",
  30147=>"111111000",
  30148=>"001011010",
  30149=>"011100011",
  30150=>"000011100",
  30151=>"111100101",
  30152=>"111011110",
  30153=>"111101111",
  30154=>"111100101",
  30155=>"101110110",
  30156=>"111110101",
  30157=>"000010111",
  30158=>"101010011",
  30159=>"111100000",
  30160=>"010100011",
  30161=>"100010110",
  30162=>"110111101",
  30163=>"101111010",
  30164=>"101101100",
  30165=>"000001100",
  30166=>"000101001",
  30167=>"010010001",
  30168=>"100001010",
  30169=>"000011110",
  30170=>"101000101",
  30171=>"000010101",
  30172=>"010110100",
  30173=>"101011111",
  30174=>"001011001",
  30175=>"011110100",
  30176=>"100010111",
  30177=>"111011101",
  30178=>"001010000",
  30179=>"101101101",
  30180=>"110110010",
  30181=>"010101010",
  30182=>"111001110",
  30183=>"100001111",
  30184=>"100101011",
  30185=>"111000011",
  30186=>"011000011",
  30187=>"000101101",
  30188=>"001000101",
  30189=>"011010100",
  30190=>"110111111",
  30191=>"001010000",
  30192=>"011001101",
  30193=>"101010000",
  30194=>"101110111",
  30195=>"111001001",
  30196=>"000110110",
  30197=>"100101110",
  30198=>"110000010",
  30199=>"111101100",
  30200=>"010011111",
  30201=>"001101111",
  30202=>"101001101",
  30203=>"011101000",
  30204=>"110101101",
  30205=>"010010000",
  30206=>"010110100",
  30207=>"110000000",
  30208=>"011111110",
  30209=>"010010111",
  30210=>"000101000",
  30211=>"010010111",
  30212=>"111100010",
  30213=>"111100000",
  30214=>"101010010",
  30215=>"111101101",
  30216=>"111010000",
  30217=>"110111111",
  30218=>"000101010",
  30219=>"100101000",
  30220=>"111010011",
  30221=>"010001101",
  30222=>"000101000",
  30223=>"110001111",
  30224=>"110000100",
  30225=>"001011111",
  30226=>"010111010",
  30227=>"001101011",
  30228=>"000100000",
  30229=>"101101111",
  30230=>"100101011",
  30231=>"001110101",
  30232=>"011010000",
  30233=>"100001101",
  30234=>"000011100",
  30235=>"001101100",
  30236=>"001000000",
  30237=>"111100001",
  30238=>"000010101",
  30239=>"100101011",
  30240=>"001011011",
  30241=>"000010011",
  30242=>"110100111",
  30243=>"110000010",
  30244=>"110001000",
  30245=>"001001111",
  30246=>"100010100",
  30247=>"001111101",
  30248=>"000101101",
  30249=>"000101001",
  30250=>"001001111",
  30251=>"111100110",
  30252=>"001001101",
  30253=>"000000101",
  30254=>"101111011",
  30255=>"000010101",
  30256=>"010000100",
  30257=>"100101011",
  30258=>"110111101",
  30259=>"010100111",
  30260=>"100101011",
  30261=>"100010101",
  30262=>"100011100",
  30263=>"010011111",
  30264=>"111111101",
  30265=>"110111110",
  30266=>"110000000",
  30267=>"111011000",
  30268=>"100100101",
  30269=>"001011000",
  30270=>"101001010",
  30271=>"101101001",
  30272=>"111100101",
  30273=>"110100100",
  30274=>"010001100",
  30275=>"000010000",
  30276=>"111010010",
  30277=>"101000010",
  30278=>"101010000",
  30279=>"111111001",
  30280=>"000000001",
  30281=>"111010110",
  30282=>"110111001",
  30283=>"011100111",
  30284=>"011000100",
  30285=>"101000000",
  30286=>"001110100",
  30287=>"101011010",
  30288=>"101101110",
  30289=>"010011010",
  30290=>"001111110",
  30291=>"001110110",
  30292=>"101111001",
  30293=>"001011100",
  30294=>"010000101",
  30295=>"011010011",
  30296=>"001101000",
  30297=>"000100101",
  30298=>"100101010",
  30299=>"000001010",
  30300=>"011011111",
  30301=>"110110111",
  30302=>"100010000",
  30303=>"000011111",
  30304=>"100001010",
  30305=>"111001000",
  30306=>"001100101",
  30307=>"000100101",
  30308=>"111111110",
  30309=>"101111001",
  30310=>"000011001",
  30311=>"100110101",
  30312=>"000001001",
  30313=>"100111110",
  30314=>"101000011",
  30315=>"010101000",
  30316=>"001101011",
  30317=>"100000010",
  30318=>"010001001",
  30319=>"100111001",
  30320=>"111011011",
  30321=>"110110011",
  30322=>"001011010",
  30323=>"001010011",
  30324=>"000110111",
  30325=>"011111001",
  30326=>"011101010",
  30327=>"110100011",
  30328=>"011010100",
  30329=>"110011101",
  30330=>"111101010",
  30331=>"110101100",
  30332=>"011010000",
  30333=>"001011001",
  30334=>"111101111",
  30335=>"011111011",
  30336=>"001001111",
  30337=>"011101001",
  30338=>"011101100",
  30339=>"101010100",
  30340=>"111011010",
  30341=>"100000100",
  30342=>"101011110",
  30343=>"110000011",
  30344=>"000001100",
  30345=>"100001000",
  30346=>"101100000",
  30347=>"111100100",
  30348=>"011000000",
  30349=>"011001001",
  30350=>"011011011",
  30351=>"111111101",
  30352=>"110111010",
  30353=>"011011110",
  30354=>"000110110",
  30355=>"001111011",
  30356=>"010000101",
  30357=>"010011110",
  30358=>"000100100",
  30359=>"101101010",
  30360=>"111000100",
  30361=>"001010000",
  30362=>"100101010",
  30363=>"001110000",
  30364=>"111010001",
  30365=>"010000101",
  30366=>"110111100",
  30367=>"010111101",
  30368=>"101110001",
  30369=>"111010101",
  30370=>"010110101",
  30371=>"111110011",
  30372=>"111001000",
  30373=>"100111110",
  30374=>"111111100",
  30375=>"111001010",
  30376=>"100111110",
  30377=>"000001010",
  30378=>"001101100",
  30379=>"001100000",
  30380=>"111001010",
  30381=>"110000011",
  30382=>"000011011",
  30383=>"000001000",
  30384=>"001101100",
  30385=>"001100110",
  30386=>"011010000",
  30387=>"011111001",
  30388=>"010000001",
  30389=>"001110100",
  30390=>"000010011",
  30391=>"111101100",
  30392=>"000000111",
  30393=>"110101011",
  30394=>"010000000",
  30395=>"011010010",
  30396=>"000101101",
  30397=>"001000111",
  30398=>"000100010",
  30399=>"101110101",
  30400=>"101111111",
  30401=>"101011101",
  30402=>"111010011",
  30403=>"000010100",
  30404=>"111001110",
  30405=>"010010001",
  30406=>"001111001",
  30407=>"000111010",
  30408=>"010101001",
  30409=>"001011110",
  30410=>"101010101",
  30411=>"110101111",
  30412=>"111111000",
  30413=>"011000000",
  30414=>"001110010",
  30415=>"110110101",
  30416=>"111111000",
  30417=>"111101101",
  30418=>"101001010",
  30419=>"000000111",
  30420=>"000111010",
  30421=>"100001001",
  30422=>"000001110",
  30423=>"101110110",
  30424=>"101000010",
  30425=>"000000010",
  30426=>"111111111",
  30427=>"001001001",
  30428=>"111001101",
  30429=>"111100101",
  30430=>"011010000",
  30431=>"111011011",
  30432=>"000111001",
  30433=>"100001011",
  30434=>"000110111",
  30435=>"101101101",
  30436=>"011000100",
  30437=>"100011111",
  30438=>"000011111",
  30439=>"110111101",
  30440=>"101010100",
  30441=>"000100100",
  30442=>"001000000",
  30443=>"000001110",
  30444=>"001011011",
  30445=>"110100101",
  30446=>"010100001",
  30447=>"100001101",
  30448=>"010000100",
  30449=>"111010001",
  30450=>"101001111",
  30451=>"100010010",
  30452=>"000100000",
  30453=>"111011010",
  30454=>"111111011",
  30455=>"001110100",
  30456=>"011100101",
  30457=>"101101110",
  30458=>"100001110",
  30459=>"000011101",
  30460=>"110110110",
  30461=>"010100100",
  30462=>"000001101",
  30463=>"101100100",
  30464=>"010110000",
  30465=>"001110110",
  30466=>"111010010",
  30467=>"100010000",
  30468=>"100011010",
  30469=>"000101111",
  30470=>"010101010",
  30471=>"000001100",
  30472=>"011000101",
  30473=>"111100101",
  30474=>"101001011",
  30475=>"100111111",
  30476=>"011100001",
  30477=>"010000111",
  30478=>"110001000",
  30479=>"111110010",
  30480=>"000111100",
  30481=>"001010000",
  30482=>"100000110",
  30483=>"000000000",
  30484=>"000001100",
  30485=>"110011101",
  30486=>"111101000",
  30487=>"111111010",
  30488=>"111110010",
  30489=>"011010111",
  30490=>"110100001",
  30491=>"000001101",
  30492=>"001111010",
  30493=>"101000101",
  30494=>"000100010",
  30495=>"100011011",
  30496=>"111101001",
  30497=>"001100001",
  30498=>"000111111",
  30499=>"111111101",
  30500=>"010001110",
  30501=>"001101000",
  30502=>"101011100",
  30503=>"111001100",
  30504=>"110010111",
  30505=>"111110010",
  30506=>"111101000",
  30507=>"101000100",
  30508=>"111101100",
  30509=>"110001001",
  30510=>"110010100",
  30511=>"010010001",
  30512=>"011111101",
  30513=>"000000101",
  30514=>"000100111",
  30515=>"110110001",
  30516=>"000110001",
  30517=>"010000011",
  30518=>"110010000",
  30519=>"111011011",
  30520=>"110100110",
  30521=>"001110000",
  30522=>"010001011",
  30523=>"000000011",
  30524=>"000000100",
  30525=>"000010100",
  30526=>"011010010",
  30527=>"111111011",
  30528=>"101010000",
  30529=>"110100101",
  30530=>"100010010",
  30531=>"011110111",
  30532=>"001011101",
  30533=>"100101001",
  30534=>"000010110",
  30535=>"001111010",
  30536=>"101100110",
  30537=>"000010010",
  30538=>"111110111",
  30539=>"001110111",
  30540=>"100111110",
  30541=>"000100101",
  30542=>"110000010",
  30543=>"010100011",
  30544=>"110000011",
  30545=>"001011101",
  30546=>"001110101",
  30547=>"000100001",
  30548=>"011100001",
  30549=>"011101001",
  30550=>"011011111",
  30551=>"100100000",
  30552=>"011110001",
  30553=>"011101101",
  30554=>"111011100",
  30555=>"100110011",
  30556=>"110111100",
  30557=>"000001110",
  30558=>"101100001",
  30559=>"000010101",
  30560=>"011001011",
  30561=>"000111000",
  30562=>"110000100",
  30563=>"100100111",
  30564=>"010001010",
  30565=>"011101001",
  30566=>"000010111",
  30567=>"100111011",
  30568=>"001000100",
  30569=>"110110101",
  30570=>"000100110",
  30571=>"010001001",
  30572=>"000101011",
  30573=>"010110000",
  30574=>"100011110",
  30575=>"111000000",
  30576=>"000001001",
  30577=>"110100111",
  30578=>"101011111",
  30579=>"100000111",
  30580=>"111010011",
  30581=>"100000101",
  30582=>"011011001",
  30583=>"110001011",
  30584=>"011000000",
  30585=>"000011001",
  30586=>"001001000",
  30587=>"101011000",
  30588=>"010110001",
  30589=>"000100110",
  30590=>"001010010",
  30591=>"111101111",
  30592=>"100000011",
  30593=>"100100100",
  30594=>"111000100",
  30595=>"010001010",
  30596=>"101000010",
  30597=>"110001110",
  30598=>"000100010",
  30599=>"001100111",
  30600=>"000101100",
  30601=>"001101000",
  30602=>"010000101",
  30603=>"000101001",
  30604=>"000010011",
  30605=>"000001010",
  30606=>"000000010",
  30607=>"111001111",
  30608=>"111111011",
  30609=>"110000000",
  30610=>"000111110",
  30611=>"001001110",
  30612=>"101011000",
  30613=>"101001110",
  30614=>"001100100",
  30615=>"000110100",
  30616=>"111100000",
  30617=>"100010010",
  30618=>"000110011",
  30619=>"101010100",
  30620=>"111011110",
  30621=>"110100110",
  30622=>"101110110",
  30623=>"110111001",
  30624=>"110100100",
  30625=>"110000101",
  30626=>"011001001",
  30627=>"011011111",
  30628=>"001000001",
  30629=>"101001011",
  30630=>"001110110",
  30631=>"111101011",
  30632=>"110111001",
  30633=>"011111110",
  30634=>"011011000",
  30635=>"111110111",
  30636=>"000001100",
  30637=>"111001010",
  30638=>"011001000",
  30639=>"011001000",
  30640=>"011001011",
  30641=>"010011000",
  30642=>"101000000",
  30643=>"001001111",
  30644=>"001101010",
  30645=>"000100011",
  30646=>"101100111",
  30647=>"011011110",
  30648=>"011001111",
  30649=>"010111010",
  30650=>"101011010",
  30651=>"110010100",
  30652=>"100100011",
  30653=>"100010001",
  30654=>"111011010",
  30655=>"001101100",
  30656=>"000000000",
  30657=>"000011000",
  30658=>"100111100",
  30659=>"110000000",
  30660=>"111110000",
  30661=>"100110011",
  30662=>"011001101",
  30663=>"000100011",
  30664=>"010010010",
  30665=>"101110101",
  30666=>"011010000",
  30667=>"110000110",
  30668=>"100100010",
  30669=>"110011011",
  30670=>"100011011",
  30671=>"111111101",
  30672=>"011000011",
  30673=>"001101001",
  30674=>"111101110",
  30675=>"001100001",
  30676=>"111101001",
  30677=>"111100000",
  30678=>"011110011",
  30679=>"010110110",
  30680=>"000100101",
  30681=>"101110101",
  30682=>"011100011",
  30683=>"011100100",
  30684=>"010111001",
  30685=>"100111101",
  30686=>"011010101",
  30687=>"001000001",
  30688=>"110001000",
  30689=>"011110010",
  30690=>"101000111",
  30691=>"000000101",
  30692=>"001010101",
  30693=>"010001011",
  30694=>"011101100",
  30695=>"100101101",
  30696=>"101000100",
  30697=>"010111110",
  30698=>"100101000",
  30699=>"110011111",
  30700=>"011100000",
  30701=>"100011010",
  30702=>"111110001",
  30703=>"011010110",
  30704=>"011011111",
  30705=>"100010110",
  30706=>"010100100",
  30707=>"001011000",
  30708=>"010110000",
  30709=>"110001001",
  30710=>"010010000",
  30711=>"010010111",
  30712=>"001001001",
  30713=>"000001111",
  30714=>"100100000",
  30715=>"001101100",
  30716=>"001100110",
  30717=>"110010110",
  30718=>"010111111",
  30719=>"110000111",
  30720=>"101001000",
  30721=>"000000111",
  30722=>"101000111",
  30723=>"100001101",
  30724=>"110011000",
  30725=>"001010011",
  30726=>"000011011",
  30727=>"001000100",
  30728=>"010100000",
  30729=>"100110110",
  30730=>"001010011",
  30731=>"000111010",
  30732=>"101101001",
  30733=>"001000011",
  30734=>"011000010",
  30735=>"101110111",
  30736=>"111101000",
  30737=>"111100000",
  30738=>"110100110",
  30739=>"010111010",
  30740=>"000011000",
  30741=>"010110010",
  30742=>"000110100",
  30743=>"010101010",
  30744=>"011001000",
  30745=>"101010111",
  30746=>"110100110",
  30747=>"010011000",
  30748=>"000000001",
  30749=>"011010110",
  30750=>"101001011",
  30751=>"011010100",
  30752=>"011101001",
  30753=>"100100101",
  30754=>"010000110",
  30755=>"000010000",
  30756=>"111011111",
  30757=>"100100100",
  30758=>"101100011",
  30759=>"010110001",
  30760=>"011011100",
  30761=>"100110111",
  30762=>"010000111",
  30763=>"101011010",
  30764=>"111001001",
  30765=>"100010110",
  30766=>"100110100",
  30767=>"000101000",
  30768=>"000101010",
  30769=>"001011000",
  30770=>"011001000",
  30771=>"111111010",
  30772=>"111001111",
  30773=>"101001001",
  30774=>"101000010",
  30775=>"010010110",
  30776=>"001101111",
  30777=>"010010010",
  30778=>"000000111",
  30779=>"111001111",
  30780=>"010000011",
  30781=>"101001110",
  30782=>"110101111",
  30783=>"001110101",
  30784=>"111001010",
  30785=>"001010010",
  30786=>"101111011",
  30787=>"011000001",
  30788=>"000000010",
  30789=>"101010101",
  30790=>"110000001",
  30791=>"011101000",
  30792=>"111101101",
  30793=>"000110000",
  30794=>"001101100",
  30795=>"111111111",
  30796=>"000011001",
  30797=>"101110010",
  30798=>"101011010",
  30799=>"100111000",
  30800=>"111000001",
  30801=>"010101101",
  30802=>"000001011",
  30803=>"001111101",
  30804=>"101110010",
  30805=>"000100001",
  30806=>"010100100",
  30807=>"001010010",
  30808=>"011110100",
  30809=>"010100010",
  30810=>"110000101",
  30811=>"100000110",
  30812=>"111011000",
  30813=>"000100010",
  30814=>"001010110",
  30815=>"100110010",
  30816=>"100011111",
  30817=>"010001000",
  30818=>"011111101",
  30819=>"011010010",
  30820=>"011011101",
  30821=>"110100101",
  30822=>"000010101",
  30823=>"110010100",
  30824=>"000010100",
  30825=>"010101000",
  30826=>"111010110",
  30827=>"110001010",
  30828=>"011111011",
  30829=>"101101100",
  30830=>"000000100",
  30831=>"110101111",
  30832=>"010010111",
  30833=>"000000011",
  30834=>"001111011",
  30835=>"110010001",
  30836=>"111011010",
  30837=>"100011001",
  30838=>"100001110",
  30839=>"100100001",
  30840=>"011011100",
  30841=>"011011000",
  30842=>"111010100",
  30843=>"011011101",
  30844=>"010101100",
  30845=>"011000011",
  30846=>"110010010",
  30847=>"000110110",
  30848=>"111010111",
  30849=>"010011000",
  30850=>"000011101",
  30851=>"110000110",
  30852=>"110010110",
  30853=>"000111100",
  30854=>"111010111",
  30855=>"100101010",
  30856=>"110100001",
  30857=>"101011110",
  30858=>"010001100",
  30859=>"110101001",
  30860=>"001001001",
  30861=>"101100101",
  30862=>"011110001",
  30863=>"011001001",
  30864=>"000100011",
  30865=>"011001010",
  30866=>"111011101",
  30867=>"101100011",
  30868=>"000110110",
  30869=>"111100100",
  30870=>"000100000",
  30871=>"101011110",
  30872=>"001111011",
  30873=>"100111000",
  30874=>"110001100",
  30875=>"010010010",
  30876=>"110011010",
  30877=>"010010110",
  30878=>"100111111",
  30879=>"010100100",
  30880=>"011011110",
  30881=>"110000010",
  30882=>"011001100",
  30883=>"011000011",
  30884=>"111010110",
  30885=>"100100110",
  30886=>"101000111",
  30887=>"111110001",
  30888=>"111011100",
  30889=>"101010101",
  30890=>"000000110",
  30891=>"010100010",
  30892=>"001000001",
  30893=>"101110010",
  30894=>"111100001",
  30895=>"010111101",
  30896=>"110001010",
  30897=>"101010111",
  30898=>"100111001",
  30899=>"100001110",
  30900=>"000010000",
  30901=>"000011010",
  30902=>"011001011",
  30903=>"001001111",
  30904=>"100010000",
  30905=>"101010101",
  30906=>"000011000",
  30907=>"011111011",
  30908=>"101100110",
  30909=>"110001010",
  30910=>"101100001",
  30911=>"001010100",
  30912=>"111011100",
  30913=>"000100110",
  30914=>"100111010",
  30915=>"111011111",
  30916=>"001100100",
  30917=>"000010000",
  30918=>"001110100",
  30919=>"111001000",
  30920=>"000111110",
  30921=>"001011011",
  30922=>"111101101",
  30923=>"000000100",
  30924=>"011010101",
  30925=>"111000100",
  30926=>"010101010",
  30927=>"000000010",
  30928=>"111110011",
  30929=>"011110011",
  30930=>"111001110",
  30931=>"000110000",
  30932=>"011110000",
  30933=>"100000101",
  30934=>"101001011",
  30935=>"010101110",
  30936=>"011000100",
  30937=>"110000001",
  30938=>"100100100",
  30939=>"010110111",
  30940=>"101001100",
  30941=>"011111000",
  30942=>"111100000",
  30943=>"011111111",
  30944=>"000001000",
  30945=>"011100001",
  30946=>"001000000",
  30947=>"111001100",
  30948=>"111011100",
  30949=>"000011001",
  30950=>"101101010",
  30951=>"000000000",
  30952=>"101110011",
  30953=>"010111101",
  30954=>"110111001",
  30955=>"100101100",
  30956=>"100110111",
  30957=>"001010011",
  30958=>"001010111",
  30959=>"000011000",
  30960=>"100000000",
  30961=>"011011010",
  30962=>"000000111",
  30963=>"100000000",
  30964=>"111100100",
  30965=>"100001101",
  30966=>"111100100",
  30967=>"010000000",
  30968=>"101010000",
  30969=>"010010100",
  30970=>"101001111",
  30971=>"000000100",
  30972=>"011011000",
  30973=>"010111110",
  30974=>"001000010",
  30975=>"111110110",
  30976=>"000100001",
  30977=>"010011110",
  30978=>"011010110",
  30979=>"101011000",
  30980=>"111110111",
  30981=>"011010010",
  30982=>"001000011",
  30983=>"000111011",
  30984=>"001010111",
  30985=>"001010011",
  30986=>"001011101",
  30987=>"000100011",
  30988=>"001000111",
  30989=>"000000110",
  30990=>"110111100",
  30991=>"011011010",
  30992=>"010001000",
  30993=>"111110000",
  30994=>"101010110",
  30995=>"111001111",
  30996=>"010010001",
  30997=>"110110011",
  30998=>"010010001",
  30999=>"010011000",
  31000=>"001000010",
  31001=>"111001110",
  31002=>"110110110",
  31003=>"100010001",
  31004=>"001100111",
  31005=>"000101011",
  31006=>"011011011",
  31007=>"011000110",
  31008=>"001101101",
  31009=>"100100001",
  31010=>"010101100",
  31011=>"110000111",
  31012=>"111111000",
  31013=>"011100101",
  31014=>"110010010",
  31015=>"110110100",
  31016=>"000110001",
  31017=>"101001100",
  31018=>"110100011",
  31019=>"000011100",
  31020=>"011100111",
  31021=>"101011010",
  31022=>"011000011",
  31023=>"101100111",
  31024=>"100011111",
  31025=>"100110111",
  31026=>"010000101",
  31027=>"001011111",
  31028=>"011101000",
  31029=>"111101100",
  31030=>"010100101",
  31031=>"000000100",
  31032=>"100110110",
  31033=>"110010010",
  31034=>"001011001",
  31035=>"011100001",
  31036=>"001010100",
  31037=>"111011111",
  31038=>"101110011",
  31039=>"011100010",
  31040=>"110111010",
  31041=>"010011100",
  31042=>"000100000",
  31043=>"110101000",
  31044=>"110010101",
  31045=>"010110011",
  31046=>"101011011",
  31047=>"100001111",
  31048=>"100110100",
  31049=>"100000000",
  31050=>"101100101",
  31051=>"100001111",
  31052=>"011110101",
  31053=>"111100101",
  31054=>"100110011",
  31055=>"001110000",
  31056=>"110011110",
  31057=>"000100110",
  31058=>"011110111",
  31059=>"110110011",
  31060=>"000111001",
  31061=>"100110111",
  31062=>"100100111",
  31063=>"101110010",
  31064=>"101110101",
  31065=>"111111001",
  31066=>"001011111",
  31067=>"010000000",
  31068=>"110111010",
  31069=>"111101001",
  31070=>"000110001",
  31071=>"111101011",
  31072=>"110010000",
  31073=>"011110001",
  31074=>"111000001",
  31075=>"111110011",
  31076=>"101000110",
  31077=>"111101111",
  31078=>"011010110",
  31079=>"010000000",
  31080=>"000101001",
  31081=>"100000111",
  31082=>"000010010",
  31083=>"001011100",
  31084=>"011011011",
  31085=>"100000100",
  31086=>"110010101",
  31087=>"101000101",
  31088=>"111001110",
  31089=>"101000010",
  31090=>"001111000",
  31091=>"110110000",
  31092=>"111110011",
  31093=>"110110010",
  31094=>"000000111",
  31095=>"111111111",
  31096=>"110110110",
  31097=>"111110000",
  31098=>"011001010",
  31099=>"111101010",
  31100=>"100100101",
  31101=>"000111001",
  31102=>"111001100",
  31103=>"010000110",
  31104=>"000101111",
  31105=>"001000100",
  31106=>"111100001",
  31107=>"010100010",
  31108=>"011110000",
  31109=>"110010010",
  31110=>"001000111",
  31111=>"101000010",
  31112=>"000010101",
  31113=>"100111101",
  31114=>"110011100",
  31115=>"000000010",
  31116=>"000000000",
  31117=>"110000010",
  31118=>"110010001",
  31119=>"010100110",
  31120=>"010110100",
  31121=>"000001000",
  31122=>"011000101",
  31123=>"101000110",
  31124=>"111011111",
  31125=>"000111100",
  31126=>"010011101",
  31127=>"001011101",
  31128=>"110001010",
  31129=>"001110010",
  31130=>"110110010",
  31131=>"011101011",
  31132=>"111010100",
  31133=>"111111111",
  31134=>"000101110",
  31135=>"101000111",
  31136=>"000000010",
  31137=>"111010011",
  31138=>"010100000",
  31139=>"001000010",
  31140=>"110011011",
  31141=>"000000010",
  31142=>"111000111",
  31143=>"110010011",
  31144=>"011111110",
  31145=>"101001100",
  31146=>"011111000",
  31147=>"001010101",
  31148=>"111100110",
  31149=>"110010100",
  31150=>"111111001",
  31151=>"001011010",
  31152=>"011100001",
  31153=>"110100110",
  31154=>"111101110",
  31155=>"011001110",
  31156=>"001100100",
  31157=>"010000100",
  31158=>"001101111",
  31159=>"011011010",
  31160=>"101111001",
  31161=>"000100001",
  31162=>"000010111",
  31163=>"100001100",
  31164=>"010011100",
  31165=>"000111010",
  31166=>"000000111",
  31167=>"010101000",
  31168=>"011010111",
  31169=>"000001010",
  31170=>"011111011",
  31171=>"001101111",
  31172=>"001111010",
  31173=>"011011001",
  31174=>"110000001",
  31175=>"111011100",
  31176=>"110010001",
  31177=>"100101011",
  31178=>"101001110",
  31179=>"010001101",
  31180=>"111000000",
  31181=>"000010001",
  31182=>"100011000",
  31183=>"000010101",
  31184=>"001000111",
  31185=>"010010111",
  31186=>"001111010",
  31187=>"100011000",
  31188=>"101101100",
  31189=>"000011100",
  31190=>"011100011",
  31191=>"100000011",
  31192=>"110010111",
  31193=>"010011001",
  31194=>"111110010",
  31195=>"111010010",
  31196=>"110011001",
  31197=>"010100001",
  31198=>"100110011",
  31199=>"101010000",
  31200=>"101000100",
  31201=>"011110001",
  31202=>"011010001",
  31203=>"111110101",
  31204=>"001101000",
  31205=>"101010111",
  31206=>"111100001",
  31207=>"100001001",
  31208=>"000110011",
  31209=>"000100010",
  31210=>"101010101",
  31211=>"000010001",
  31212=>"000001010",
  31213=>"110111011",
  31214=>"101110001",
  31215=>"011000100",
  31216=>"100001000",
  31217=>"110011010",
  31218=>"011110101",
  31219=>"001101100",
  31220=>"110110111",
  31221=>"111101101",
  31222=>"110010100",
  31223=>"011100001",
  31224=>"000100011",
  31225=>"011001000",
  31226=>"101011100",
  31227=>"001100110",
  31228=>"110001101",
  31229=>"000100001",
  31230=>"000010110",
  31231=>"001010000",
  31232=>"101110000",
  31233=>"011010001",
  31234=>"100100100",
  31235=>"011110011",
  31236=>"110011000",
  31237=>"001001001",
  31238=>"110010010",
  31239=>"000100100",
  31240=>"100011110",
  31241=>"100100001",
  31242=>"001010000",
  31243=>"001111100",
  31244=>"101111011",
  31245=>"010001100",
  31246=>"111111001",
  31247=>"101011111",
  31248=>"110111001",
  31249=>"011111011",
  31250=>"111110111",
  31251=>"111011000",
  31252=>"011010110",
  31253=>"111011011",
  31254=>"101010011",
  31255=>"100011101",
  31256=>"011111111",
  31257=>"000110011",
  31258=>"101010111",
  31259=>"100011000",
  31260=>"110010010",
  31261=>"110110001",
  31262=>"001000011",
  31263=>"010111111",
  31264=>"000010001",
  31265=>"001011101",
  31266=>"100100101",
  31267=>"110001100",
  31268=>"110001100",
  31269=>"110011000",
  31270=>"000000110",
  31271=>"001001101",
  31272=>"000110001",
  31273=>"100011100",
  31274=>"111010100",
  31275=>"011000001",
  31276=>"101000110",
  31277=>"100110111",
  31278=>"001101111",
  31279=>"100110101",
  31280=>"000000100",
  31281=>"011101100",
  31282=>"001011011",
  31283=>"101100011",
  31284=>"011110111",
  31285=>"010000000",
  31286=>"001101110",
  31287=>"110000010",
  31288=>"110111001",
  31289=>"000000100",
  31290=>"101001110",
  31291=>"000001011",
  31292=>"111101110",
  31293=>"110111111",
  31294=>"110110011",
  31295=>"101001111",
  31296=>"100111010",
  31297=>"010000101",
  31298=>"001100000",
  31299=>"001011010",
  31300=>"000110011",
  31301=>"101110000",
  31302=>"000101011",
  31303=>"100011011",
  31304=>"100011000",
  31305=>"010000011",
  31306=>"001110000",
  31307=>"000111001",
  31308=>"100000000",
  31309=>"110100010",
  31310=>"100000010",
  31311=>"001111101",
  31312=>"001111111",
  31313=>"000110110",
  31314=>"000100000",
  31315=>"000001011",
  31316=>"110000000",
  31317=>"000001110",
  31318=>"000101000",
  31319=>"110011111",
  31320=>"110010000",
  31321=>"100110001",
  31322=>"000011000",
  31323=>"000100001",
  31324=>"000101110",
  31325=>"100100110",
  31326=>"011011111",
  31327=>"111100111",
  31328=>"010011100",
  31329=>"001011011",
  31330=>"000010110",
  31331=>"001111001",
  31332=>"110110111",
  31333=>"011100100",
  31334=>"001100001",
  31335=>"001111111",
  31336=>"100100000",
  31337=>"000000011",
  31338=>"000101101",
  31339=>"111011000",
  31340=>"111101100",
  31341=>"000101001",
  31342=>"000111101",
  31343=>"011101000",
  31344=>"000101101",
  31345=>"001000000",
  31346=>"010110111",
  31347=>"111001110",
  31348=>"010101100",
  31349=>"110010111",
  31350=>"100010010",
  31351=>"011010110",
  31352=>"010110110",
  31353=>"101101001",
  31354=>"110011011",
  31355=>"101111001",
  31356=>"001111011",
  31357=>"000111010",
  31358=>"000001010",
  31359=>"000010010",
  31360=>"100100000",
  31361=>"011100100",
  31362=>"100111000",
  31363=>"001000100",
  31364=>"001010101",
  31365=>"011110011",
  31366=>"111000010",
  31367=>"000101010",
  31368=>"011110110",
  31369=>"011000011",
  31370=>"000001100",
  31371=>"111110101",
  31372=>"010000000",
  31373=>"101010100",
  31374=>"111000101",
  31375=>"100101000",
  31376=>"110100101",
  31377=>"101011111",
  31378=>"010010001",
  31379=>"011011101",
  31380=>"100010001",
  31381=>"101100001",
  31382=>"110011110",
  31383=>"011101011",
  31384=>"010010011",
  31385=>"011000011",
  31386=>"011110001",
  31387=>"110000110",
  31388=>"011101100",
  31389=>"011010100",
  31390=>"111101001",
  31391=>"101000000",
  31392=>"001100000",
  31393=>"100011110",
  31394=>"011001110",
  31395=>"010100001",
  31396=>"111110011",
  31397=>"000011010",
  31398=>"011001111",
  31399=>"010010101",
  31400=>"000101110",
  31401=>"110111111",
  31402=>"011001100",
  31403=>"100000110",
  31404=>"010001000",
  31405=>"000010010",
  31406=>"110100110",
  31407=>"010111100",
  31408=>"010001010",
  31409=>"011000101",
  31410=>"001110111",
  31411=>"001111011",
  31412=>"101110100",
  31413=>"001111101",
  31414=>"100111111",
  31415=>"010001110",
  31416=>"001010010",
  31417=>"100101111",
  31418=>"000101110",
  31419=>"100011000",
  31420=>"000000110",
  31421=>"110010101",
  31422=>"101101101",
  31423=>"000110101",
  31424=>"101110101",
  31425=>"010101111",
  31426=>"011000011",
  31427=>"110000111",
  31428=>"110111010",
  31429=>"100011011",
  31430=>"001111011",
  31431=>"011000000",
  31432=>"001001000",
  31433=>"000111110",
  31434=>"010010111",
  31435=>"010001111",
  31436=>"100011100",
  31437=>"001010110",
  31438=>"111111110",
  31439=>"011010011",
  31440=>"010101010",
  31441=>"110011110",
  31442=>"110101101",
  31443=>"110000010",
  31444=>"000001100",
  31445=>"000101001",
  31446=>"010110001",
  31447=>"111001010",
  31448=>"000011110",
  31449=>"010011110",
  31450=>"010100000",
  31451=>"111110001",
  31452=>"001001100",
  31453=>"000000101",
  31454=>"010001011",
  31455=>"001000110",
  31456=>"101000011",
  31457=>"010110110",
  31458=>"000000111",
  31459=>"011000001",
  31460=>"000010000",
  31461=>"011101101",
  31462=>"001100010",
  31463=>"100001001",
  31464=>"010101011",
  31465=>"100110001",
  31466=>"010100011",
  31467=>"010100010",
  31468=>"011010111",
  31469=>"111000111",
  31470=>"001001101",
  31471=>"110000011",
  31472=>"001010001",
  31473=>"111011001",
  31474=>"110111101",
  31475=>"001101011",
  31476=>"110001001",
  31477=>"000100110",
  31478=>"010011010",
  31479=>"101110100",
  31480=>"011100011",
  31481=>"110000111",
  31482=>"011011100",
  31483=>"000111011",
  31484=>"001111000",
  31485=>"000010111",
  31486=>"010101000",
  31487=>"111101111",
  31488=>"110101101",
  31489=>"111001101",
  31490=>"000100110",
  31491=>"010000010",
  31492=>"110100100",
  31493=>"000010101",
  31494=>"010000100",
  31495=>"110101000",
  31496=>"010000101",
  31497=>"000111001",
  31498=>"010100101",
  31499=>"000100010",
  31500=>"000011010",
  31501=>"011100011",
  31502=>"011101001",
  31503=>"100011000",
  31504=>"101001101",
  31505=>"000110011",
  31506=>"000101001",
  31507=>"011110110",
  31508=>"111010110",
  31509=>"000101001",
  31510=>"111101110",
  31511=>"110001011",
  31512=>"001111010",
  31513=>"010010110",
  31514=>"010100100",
  31515=>"100011011",
  31516=>"110000000",
  31517=>"101110110",
  31518=>"101001011",
  31519=>"010010110",
  31520=>"000011000",
  31521=>"000111001",
  31522=>"000110001",
  31523=>"101101000",
  31524=>"011100011",
  31525=>"111111011",
  31526=>"010000010",
  31527=>"000111011",
  31528=>"010010000",
  31529=>"110111101",
  31530=>"001101111",
  31531=>"000000100",
  31532=>"111111010",
  31533=>"110011101",
  31534=>"100011111",
  31535=>"000100010",
  31536=>"001010110",
  31537=>"011001101",
  31538=>"000010101",
  31539=>"001001010",
  31540=>"010111011",
  31541=>"100011100",
  31542=>"001000110",
  31543=>"011100010",
  31544=>"111110001",
  31545=>"101011000",
  31546=>"100101000",
  31547=>"101101011",
  31548=>"100010001",
  31549=>"010000011",
  31550=>"000010001",
  31551=>"011011101",
  31552=>"110011001",
  31553=>"111001010",
  31554=>"011101110",
  31555=>"101100111",
  31556=>"100011010",
  31557=>"101001101",
  31558=>"101010100",
  31559=>"011011001",
  31560=>"000011000",
  31561=>"000011110",
  31562=>"111011010",
  31563=>"110100110",
  31564=>"100100000",
  31565=>"001100001",
  31566=>"101001011",
  31567=>"111011011",
  31568=>"100101110",
  31569=>"101100000",
  31570=>"010010011",
  31571=>"001011111",
  31572=>"101100000",
  31573=>"011001101",
  31574=>"110110000",
  31575=>"110101100",
  31576=>"011101001",
  31577=>"011101101",
  31578=>"001101101",
  31579=>"110101110",
  31580=>"111000000",
  31581=>"111110001",
  31582=>"100110110",
  31583=>"101011101",
  31584=>"101000001",
  31585=>"001001011",
  31586=>"010111111",
  31587=>"001010101",
  31588=>"101101100",
  31589=>"111011100",
  31590=>"111000111",
  31591=>"001101000",
  31592=>"111011010",
  31593=>"111011001",
  31594=>"010001110",
  31595=>"101100111",
  31596=>"100011111",
  31597=>"011111011",
  31598=>"010011101",
  31599=>"010101001",
  31600=>"100101001",
  31601=>"001111001",
  31602=>"110001110",
  31603=>"001101010",
  31604=>"000001000",
  31605=>"100110100",
  31606=>"110000100",
  31607=>"100110011",
  31608=>"011000100",
  31609=>"000101010",
  31610=>"100010111",
  31611=>"101100101",
  31612=>"101110100",
  31613=>"101001001",
  31614=>"111011101",
  31615=>"010100101",
  31616=>"100111001",
  31617=>"000011101",
  31618=>"001000011",
  31619=>"111110100",
  31620=>"000000010",
  31621=>"100010001",
  31622=>"111100111",
  31623=>"111100101",
  31624=>"100101011",
  31625=>"101110000",
  31626=>"000101111",
  31627=>"111100001",
  31628=>"111101010",
  31629=>"001101111",
  31630=>"001011001",
  31631=>"101100011",
  31632=>"000101100",
  31633=>"001000110",
  31634=>"010011001",
  31635=>"000000101",
  31636=>"110011001",
  31637=>"110100000",
  31638=>"100001100",
  31639=>"010001011",
  31640=>"001001100",
  31641=>"111100000",
  31642=>"101101011",
  31643=>"001111101",
  31644=>"101000110",
  31645=>"001010010",
  31646=>"110000010",
  31647=>"011001010",
  31648=>"000100111",
  31649=>"111010000",
  31650=>"010101010",
  31651=>"111000011",
  31652=>"000010101",
  31653=>"000110110",
  31654=>"001100000",
  31655=>"100111010",
  31656=>"010001100",
  31657=>"010000011",
  31658=>"101011110",
  31659=>"001101001",
  31660=>"000100000",
  31661=>"110000011",
  31662=>"101100110",
  31663=>"000000011",
  31664=>"100010001",
  31665=>"000110110",
  31666=>"000110111",
  31667=>"001011011",
  31668=>"101101101",
  31669=>"110001101",
  31670=>"010101011",
  31671=>"011101010",
  31672=>"000000110",
  31673=>"000010100",
  31674=>"011101011",
  31675=>"001010011",
  31676=>"010110111",
  31677=>"010110110",
  31678=>"100100111",
  31679=>"101111000",
  31680=>"100001010",
  31681=>"111110111",
  31682=>"010110101",
  31683=>"010100100",
  31684=>"011101101",
  31685=>"101000101",
  31686=>"010011000",
  31687=>"010100111",
  31688=>"000000010",
  31689=>"001000111",
  31690=>"100110100",
  31691=>"000011011",
  31692=>"010100011",
  31693=>"101101111",
  31694=>"101011010",
  31695=>"000100110",
  31696=>"110111001",
  31697=>"110010101",
  31698=>"111011000",
  31699=>"100110011",
  31700=>"111111111",
  31701=>"011101101",
  31702=>"101011011",
  31703=>"000100110",
  31704=>"011010110",
  31705=>"101001001",
  31706=>"001001101",
  31707=>"010000101",
  31708=>"000111000",
  31709=>"000011110",
  31710=>"100110010",
  31711=>"000000110",
  31712=>"100101011",
  31713=>"110101000",
  31714=>"110111001",
  31715=>"111111000",
  31716=>"100001100",
  31717=>"100000010",
  31718=>"000010111",
  31719=>"110010100",
  31720=>"010110010",
  31721=>"110000000",
  31722=>"101000110",
  31723=>"100010011",
  31724=>"010110100",
  31725=>"011011010",
  31726=>"001000111",
  31727=>"111000011",
  31728=>"110011100",
  31729=>"100111100",
  31730=>"110111110",
  31731=>"001100100",
  31732=>"101011011",
  31733=>"010001000",
  31734=>"111111111",
  31735=>"010000010",
  31736=>"011100100",
  31737=>"111011100",
  31738=>"010011000",
  31739=>"101001111",
  31740=>"011111010",
  31741=>"101000001",
  31742=>"000010000",
  31743=>"110000011",
  31744=>"000010000",
  31745=>"011011001",
  31746=>"111001011",
  31747=>"101101011",
  31748=>"001101000",
  31749=>"111100000",
  31750=>"111100010",
  31751=>"101000001",
  31752=>"000001110",
  31753=>"010011000",
  31754=>"110111111",
  31755=>"111010110",
  31756=>"111111001",
  31757=>"011011101",
  31758=>"000100110",
  31759=>"111001010",
  31760=>"000101111",
  31761=>"000100100",
  31762=>"110011101",
  31763=>"101101011",
  31764=>"111111101",
  31765=>"011111111",
  31766=>"111001001",
  31767=>"011010101",
  31768=>"010010100",
  31769=>"001111000",
  31770=>"100101110",
  31771=>"111110110",
  31772=>"011000011",
  31773=>"101100011",
  31774=>"111110101",
  31775=>"111011111",
  31776=>"010111111",
  31777=>"111110001",
  31778=>"000011000",
  31779=>"110010101",
  31780=>"001110010",
  31781=>"010000110",
  31782=>"111010011",
  31783=>"000001100",
  31784=>"001111100",
  31785=>"001011010",
  31786=>"100000011",
  31787=>"111110110",
  31788=>"001111101",
  31789=>"111000011",
  31790=>"010011101",
  31791=>"000010010",
  31792=>"100101101",
  31793=>"101011011",
  31794=>"010110100",
  31795=>"001000000",
  31796=>"010010111",
  31797=>"001000100",
  31798=>"101101101",
  31799=>"010011110",
  31800=>"011011100",
  31801=>"111111001",
  31802=>"011101010",
  31803=>"010110000",
  31804=>"000001100",
  31805=>"000010011",
  31806=>"111000000",
  31807=>"100100011",
  31808=>"011000101",
  31809=>"000001000",
  31810=>"101100001",
  31811=>"100000010",
  31812=>"100111101",
  31813=>"110010001",
  31814=>"011011110",
  31815=>"111100000",
  31816=>"110011000",
  31817=>"101001001",
  31818=>"110000000",
  31819=>"010010001",
  31820=>"011110000",
  31821=>"101101000",
  31822=>"001111111",
  31823=>"100100100",
  31824=>"101001011",
  31825=>"110011000",
  31826=>"000101010",
  31827=>"110000110",
  31828=>"110010101",
  31829=>"011110110",
  31830=>"111110000",
  31831=>"100000000",
  31832=>"000010001",
  31833=>"111100010",
  31834=>"100111110",
  31835=>"000011101",
  31836=>"100110110",
  31837=>"010011100",
  31838=>"000000000",
  31839=>"001100110",
  31840=>"010100001",
  31841=>"111101100",
  31842=>"011110110",
  31843=>"100000110",
  31844=>"000011111",
  31845=>"111101010",
  31846=>"010110110",
  31847=>"010000101",
  31848=>"101110100",
  31849=>"000111110",
  31850=>"101001011",
  31851=>"000010101",
  31852=>"000001111",
  31853=>"010010011",
  31854=>"000111110",
  31855=>"010010001",
  31856=>"001110101",
  31857=>"000101101",
  31858=>"001100010",
  31859=>"101100000",
  31860=>"011000011",
  31861=>"010001110",
  31862=>"000100111",
  31863=>"101111011",
  31864=>"001110010",
  31865=>"100000000",
  31866=>"000010101",
  31867=>"010010011",
  31868=>"110110011",
  31869=>"000110110",
  31870=>"000111010",
  31871=>"000000011",
  31872=>"111001110",
  31873=>"111010010",
  31874=>"110001001",
  31875=>"001101011",
  31876=>"111111011",
  31877=>"000111111",
  31878=>"001100011",
  31879=>"101110000",
  31880=>"111000011",
  31881=>"011111111",
  31882=>"000010100",
  31883=>"011100111",
  31884=>"100100010",
  31885=>"011001100",
  31886=>"001011100",
  31887=>"011100000",
  31888=>"000001111",
  31889=>"110000011",
  31890=>"110111000",
  31891=>"100101011",
  31892=>"011000001",
  31893=>"010000001",
  31894=>"010001000",
  31895=>"001100101",
  31896=>"100011001",
  31897=>"001001011",
  31898=>"001001000",
  31899=>"110011010",
  31900=>"110101100",
  31901=>"111000000",
  31902=>"000000000",
  31903=>"001100101",
  31904=>"000111011",
  31905=>"110101001",
  31906=>"001110001",
  31907=>"101011001",
  31908=>"011010000",
  31909=>"000010000",
  31910=>"010001010",
  31911=>"101001110",
  31912=>"001010111",
  31913=>"000000111",
  31914=>"011011000",
  31915=>"010100000",
  31916=>"001100001",
  31917=>"010100011",
  31918=>"000110010",
  31919=>"110101101",
  31920=>"100100110",
  31921=>"100100111",
  31922=>"101101011",
  31923=>"111010000",
  31924=>"100100111",
  31925=>"000100000",
  31926=>"111001110",
  31927=>"000010001",
  31928=>"000001010",
  31929=>"011010010",
  31930=>"110010111",
  31931=>"000110011",
  31932=>"000000001",
  31933=>"000100101",
  31934=>"001001000",
  31935=>"100000010",
  31936=>"011000100",
  31937=>"101001010",
  31938=>"010010111",
  31939=>"001111011",
  31940=>"001111000",
  31941=>"000111000",
  31942=>"011001110",
  31943=>"001110101",
  31944=>"110101010",
  31945=>"111100110",
  31946=>"010110111",
  31947=>"110101010",
  31948=>"100010111",
  31949=>"000100100",
  31950=>"011111011",
  31951=>"011010001",
  31952=>"101000101",
  31953=>"000000001",
  31954=>"000000010",
  31955=>"000011111",
  31956=>"001111000",
  31957=>"110001100",
  31958=>"101101000",
  31959=>"101111100",
  31960=>"000000000",
  31961=>"111110011",
  31962=>"000011101",
  31963=>"100110001",
  31964=>"101001011",
  31965=>"100000011",
  31966=>"101110111",
  31967=>"001100100",
  31968=>"000000101",
  31969=>"011110101",
  31970=>"111000000",
  31971=>"111100110",
  31972=>"000110011",
  31973=>"000010101",
  31974=>"001001100",
  31975=>"000001111",
  31976=>"101001001",
  31977=>"110111010",
  31978=>"000001101",
  31979=>"001101110",
  31980=>"110111101",
  31981=>"000001111",
  31982=>"111101010",
  31983=>"010010101",
  31984=>"011000011",
  31985=>"010100010",
  31986=>"010001000",
  31987=>"010010100",
  31988=>"110110100",
  31989=>"011011001",
  31990=>"010101001",
  31991=>"110000110",
  31992=>"111110100",
  31993=>"110001100",
  31994=>"011000110",
  31995=>"000000110",
  31996=>"011000001",
  31997=>"001010001",
  31998=>"010100000",
  31999=>"011010110",
  32000=>"000110111",
  32001=>"110010110",
  32002=>"011110001",
  32003=>"010010011",
  32004=>"000011001",
  32005=>"011101011",
  32006=>"101011111",
  32007=>"110101101",
  32008=>"001011111",
  32009=>"111001011",
  32010=>"111101101",
  32011=>"001010000",
  32012=>"111101011",
  32013=>"001010101",
  32014=>"001000010",
  32015=>"010110001",
  32016=>"011011111",
  32017=>"110000001",
  32018=>"111110101",
  32019=>"110011010",
  32020=>"110100010",
  32021=>"111001100",
  32022=>"101101111",
  32023=>"011110001",
  32024=>"110110010",
  32025=>"001101011",
  32026=>"001010010",
  32027=>"101010001",
  32028=>"110111011",
  32029=>"000001111",
  32030=>"101111011",
  32031=>"000011101",
  32032=>"110000100",
  32033=>"110110011",
  32034=>"111101000",
  32035=>"101000111",
  32036=>"001000011",
  32037=>"100000110",
  32038=>"101101110",
  32039=>"001111111",
  32040=>"100110000",
  32041=>"010000100",
  32042=>"110101111",
  32043=>"111110101",
  32044=>"001101100",
  32045=>"100010000",
  32046=>"001110011",
  32047=>"001001100",
  32048=>"111111001",
  32049=>"111000110",
  32050=>"011110111",
  32051=>"111110010",
  32052=>"010010101",
  32053=>"000001011",
  32054=>"111011000",
  32055=>"110110011",
  32056=>"110110000",
  32057=>"010110100",
  32058=>"101110101",
  32059=>"100110110",
  32060=>"100000001",
  32061=>"111000101",
  32062=>"100011111",
  32063=>"001001100",
  32064=>"000000001",
  32065=>"011101001",
  32066=>"000101101",
  32067=>"000101101",
  32068=>"001101101",
  32069=>"111111001",
  32070=>"000110100",
  32071=>"000001001",
  32072=>"100011000",
  32073=>"110110110",
  32074=>"011001101",
  32075=>"001000110",
  32076=>"111010000",
  32077=>"100101010",
  32078=>"111111100",
  32079=>"001011101",
  32080=>"001000101",
  32081=>"010010111",
  32082=>"011111101",
  32083=>"111000010",
  32084=>"001111011",
  32085=>"011010110",
  32086=>"101101001",
  32087=>"000110000",
  32088=>"110001001",
  32089=>"101000111",
  32090=>"111000100",
  32091=>"011101101",
  32092=>"111000000",
  32093=>"000100111",
  32094=>"010001111",
  32095=>"000111111",
  32096=>"100100000",
  32097=>"011101101",
  32098=>"111000100",
  32099=>"110110101",
  32100=>"110111111",
  32101=>"111101011",
  32102=>"010001010",
  32103=>"000110010",
  32104=>"111001011",
  32105=>"010000000",
  32106=>"110100010",
  32107=>"101100000",
  32108=>"010010100",
  32109=>"001101101",
  32110=>"000000110",
  32111=>"000111011",
  32112=>"000110110",
  32113=>"100001101",
  32114=>"001110110",
  32115=>"111100100",
  32116=>"100111010",
  32117=>"111111101",
  32118=>"110101110",
  32119=>"100101010",
  32120=>"000001010",
  32121=>"001100101",
  32122=>"111111111",
  32123=>"011100000",
  32124=>"110110001",
  32125=>"101011010",
  32126=>"010000111",
  32127=>"110011000",
  32128=>"000010000",
  32129=>"110100010",
  32130=>"111000110",
  32131=>"110001011",
  32132=>"011001010",
  32133=>"001110111",
  32134=>"101010100",
  32135=>"101010000",
  32136=>"010001110",
  32137=>"001000001",
  32138=>"110111101",
  32139=>"001100111",
  32140=>"001110111",
  32141=>"100111111",
  32142=>"011010111",
  32143=>"111010111",
  32144=>"011101100",
  32145=>"010000100",
  32146=>"111100001",
  32147=>"101101010",
  32148=>"110000001",
  32149=>"000000010",
  32150=>"000011100",
  32151=>"001000101",
  32152=>"110111000",
  32153=>"100110010",
  32154=>"000011001",
  32155=>"010011111",
  32156=>"110001010",
  32157=>"100000101",
  32158=>"001111001",
  32159=>"000110001",
  32160=>"110010001",
  32161=>"010000000",
  32162=>"001101001",
  32163=>"111100011",
  32164=>"010010010",
  32165=>"100000101",
  32166=>"101110011",
  32167=>"010000111",
  32168=>"001111000",
  32169=>"111111111",
  32170=>"100111100",
  32171=>"001101111",
  32172=>"001111010",
  32173=>"000101110",
  32174=>"111011010",
  32175=>"100110110",
  32176=>"101100000",
  32177=>"100011001",
  32178=>"100001011",
  32179=>"000010010",
  32180=>"101111001",
  32181=>"101101001",
  32182=>"111011111",
  32183=>"001111111",
  32184=>"010110111",
  32185=>"101100010",
  32186=>"010000100",
  32187=>"111100110",
  32188=>"000101110",
  32189=>"000001000",
  32190=>"100100010",
  32191=>"110000100",
  32192=>"010010101",
  32193=>"111100011",
  32194=>"000100101",
  32195=>"010010101",
  32196=>"010000010",
  32197=>"000101001",
  32198=>"001100001",
  32199=>"000001010",
  32200=>"010100001",
  32201=>"000110000",
  32202=>"110110101",
  32203=>"111111110",
  32204=>"011111001",
  32205=>"110111101",
  32206=>"101011011",
  32207=>"001111010",
  32208=>"011100110",
  32209=>"010010001",
  32210=>"101110011",
  32211=>"010100000",
  32212=>"110100011",
  32213=>"001000101",
  32214=>"100100000",
  32215=>"000000100",
  32216=>"100111100",
  32217=>"100101010",
  32218=>"010010001",
  32219=>"100001011",
  32220=>"001100100",
  32221=>"001101011",
  32222=>"101010010",
  32223=>"000101111",
  32224=>"101000011",
  32225=>"101001001",
  32226=>"011111100",
  32227=>"001010011",
  32228=>"010001111",
  32229=>"100011011",
  32230=>"100001100",
  32231=>"001110010",
  32232=>"110101110",
  32233=>"110010011",
  32234=>"110001111",
  32235=>"011111011",
  32236=>"111000010",
  32237=>"110110000",
  32238=>"011111110",
  32239=>"011010101",
  32240=>"111110000",
  32241=>"110110000",
  32242=>"101101010",
  32243=>"110011010",
  32244=>"100111001",
  32245=>"010110110",
  32246=>"000110100",
  32247=>"100101100",
  32248=>"110001110",
  32249=>"110010101",
  32250=>"100011101",
  32251=>"101110000",
  32252=>"110011001",
  32253=>"011011101",
  32254=>"010001000",
  32255=>"000110100",
  32256=>"101010110",
  32257=>"100110110",
  32258=>"011101111",
  32259=>"010101010",
  32260=>"011010101",
  32261=>"101000111",
  32262=>"011000111",
  32263=>"111110101",
  32264=>"110000000",
  32265=>"110010100",
  32266=>"000111011",
  32267=>"000001010",
  32268=>"010100000",
  32269=>"010111111",
  32270=>"000010001",
  32271=>"110010110",
  32272=>"100100000",
  32273=>"010000000",
  32274=>"100101101",
  32275=>"111011111",
  32276=>"000000100",
  32277=>"011101000",
  32278=>"011011010",
  32279=>"111010100",
  32280=>"100101000",
  32281=>"010100100",
  32282=>"001000000",
  32283=>"000110111",
  32284=>"111001101",
  32285=>"110001011",
  32286=>"111101110",
  32287=>"111101100",
  32288=>"010110010",
  32289=>"111111100",
  32290=>"011010000",
  32291=>"011000010",
  32292=>"100110101",
  32293=>"001011000",
  32294=>"011111111",
  32295=>"001001110",
  32296=>"101111001",
  32297=>"101000100",
  32298=>"110011101",
  32299=>"001110011",
  32300=>"001111100",
  32301=>"101110010",
  32302=>"011011101",
  32303=>"110100100",
  32304=>"110001100",
  32305=>"000100010",
  32306=>"101001001",
  32307=>"011110001",
  32308=>"101010001",
  32309=>"100011101",
  32310=>"010000110",
  32311=>"000110111",
  32312=>"101110110",
  32313=>"010001000",
  32314=>"011100111",
  32315=>"011011101",
  32316=>"010000000",
  32317=>"010000010",
  32318=>"010100001",
  32319=>"011101101",
  32320=>"010111101",
  32321=>"000100000",
  32322=>"110010000",
  32323=>"000101110",
  32324=>"111010111",
  32325=>"000111001",
  32326=>"011110010",
  32327=>"010001111",
  32328=>"101011101",
  32329=>"010101101",
  32330=>"010110101",
  32331=>"100111010",
  32332=>"001111111",
  32333=>"000011101",
  32334=>"101011001",
  32335=>"010111000",
  32336=>"011000001",
  32337=>"110100011",
  32338=>"000101011",
  32339=>"110011110",
  32340=>"011100010",
  32341=>"000000111",
  32342=>"110101110",
  32343=>"101100100",
  32344=>"101011000",
  32345=>"110010011",
  32346=>"111010011",
  32347=>"101000111",
  32348=>"111101000",
  32349=>"010111100",
  32350=>"101001001",
  32351=>"000100101",
  32352=>"000100001",
  32353=>"001000010",
  32354=>"101111001",
  32355=>"011101000",
  32356=>"001001111",
  32357=>"011110111",
  32358=>"110111010",
  32359=>"000011011",
  32360=>"000000111",
  32361=>"010011011",
  32362=>"101101111",
  32363=>"010110011",
  32364=>"011011100",
  32365=>"010010110",
  32366=>"000010001",
  32367=>"111100100",
  32368=>"000110110",
  32369=>"111011010",
  32370=>"001010110",
  32371=>"001110101",
  32372=>"011000100",
  32373=>"110000100",
  32374=>"111111111",
  32375=>"010011100",
  32376=>"011110111",
  32377=>"111001110",
  32378=>"010101101",
  32379=>"110111111",
  32380=>"100001001",
  32381=>"111011011",
  32382=>"010001001",
  32383=>"010110100",
  32384=>"101001000",
  32385=>"100110010",
  32386=>"011111000",
  32387=>"100101110",
  32388=>"111001100",
  32389=>"101101100",
  32390=>"000011000",
  32391=>"111111110",
  32392=>"001011010",
  32393=>"010000101",
  32394=>"010011001",
  32395=>"011000010",
  32396=>"101100101",
  32397=>"001110111",
  32398=>"110011010",
  32399=>"001001000",
  32400=>"100101110",
  32401=>"011011000",
  32402=>"001011110",
  32403=>"110110011",
  32404=>"011000000",
  32405=>"110101000",
  32406=>"000100111",
  32407=>"001101111",
  32408=>"110111011",
  32409=>"110011001",
  32410=>"101010101",
  32411=>"011000000",
  32412=>"101110000",
  32413=>"110100111",
  32414=>"110111010",
  32415=>"110010110",
  32416=>"111110101",
  32417=>"110111101",
  32418=>"000100000",
  32419=>"101010100",
  32420=>"010110011",
  32421=>"100011110",
  32422=>"010011010",
  32423=>"111101011",
  32424=>"100010100",
  32425=>"111001010",
  32426=>"011101101",
  32427=>"001001011",
  32428=>"011011010",
  32429=>"011010010",
  32430=>"101111100",
  32431=>"110001001",
  32432=>"000100000",
  32433=>"001000101",
  32434=>"000110010",
  32435=>"101111001",
  32436=>"100100001",
  32437=>"010010110",
  32438=>"111111100",
  32439=>"111110100",
  32440=>"110101111",
  32441=>"000010011",
  32442=>"010110011",
  32443=>"000001110",
  32444=>"101010000",
  32445=>"000101111",
  32446=>"000010000",
  32447=>"110101110",
  32448=>"010010010",
  32449=>"011110111",
  32450=>"110100011",
  32451=>"110101111",
  32452=>"000010001",
  32453=>"000010011",
  32454=>"110000010",
  32455=>"010000101",
  32456=>"110000100",
  32457=>"010001000",
  32458=>"010101001",
  32459=>"000011001",
  32460=>"010001000",
  32461=>"001001101",
  32462=>"100110101",
  32463=>"010011000",
  32464=>"000110101",
  32465=>"111100110",
  32466=>"000011001",
  32467=>"011001101",
  32468=>"001111000",
  32469=>"101100100",
  32470=>"100100111",
  32471=>"000110000",
  32472=>"000010010",
  32473=>"111111000",
  32474=>"111100011",
  32475=>"100111011",
  32476=>"100011110",
  32477=>"010010111",
  32478=>"001101101",
  32479=>"000101100",
  32480=>"101001101",
  32481=>"010111010",
  32482=>"001100000",
  32483=>"111011011",
  32484=>"001101101",
  32485=>"110110001",
  32486=>"111011101",
  32487=>"000001100",
  32488=>"000110010",
  32489=>"101101100",
  32490=>"110011000",
  32491=>"011011010",
  32492=>"111100110",
  32493=>"100010011",
  32494=>"001001111",
  32495=>"010010011",
  32496=>"000101100",
  32497=>"110111000",
  32498=>"111001100",
  32499=>"101011100",
  32500=>"000100011",
  32501=>"100111101",
  32502=>"110010100",
  32503=>"111101101",
  32504=>"100101100",
  32505=>"111111111",
  32506=>"001100011",
  32507=>"111010000",
  32508=>"001100111",
  32509=>"010101111",
  32510=>"111010001",
  32511=>"100000100",
  32512=>"010101000",
  32513=>"001111101",
  32514=>"100101001",
  32515=>"101000001",
  32516=>"011010001",
  32517=>"101010110",
  32518=>"011101101",
  32519=>"011110001",
  32520=>"110100010",
  32521=>"001111001",
  32522=>"000101111",
  32523=>"001110000",
  32524=>"111100010",
  32525=>"100100100",
  32526=>"100000000",
  32527=>"001111111",
  32528=>"110111111",
  32529=>"100101000",
  32530=>"010101111",
  32531=>"110010100",
  32532=>"011010011",
  32533=>"010001111",
  32534=>"101010100",
  32535=>"111011000",
  32536=>"111011010",
  32537=>"100110000",
  32538=>"010110110",
  32539=>"010001011",
  32540=>"111001001",
  32541=>"101101000",
  32542=>"010011000",
  32543=>"001100000",
  32544=>"010100101",
  32545=>"001000010",
  32546=>"000111111",
  32547=>"111111110",
  32548=>"000101000",
  32549=>"010110000",
  32550=>"010010000",
  32551=>"101111000",
  32552=>"111000000",
  32553=>"101101000",
  32554=>"111111110",
  32555=>"010010001",
  32556=>"001100000",
  32557=>"111000000",
  32558=>"010100000",
  32559=>"011011011",
  32560=>"001110111",
  32561=>"110010110",
  32562=>"011100000",
  32563=>"101011111",
  32564=>"001000000",
  32565=>"011100011",
  32566=>"011000001",
  32567=>"000100000",
  32568=>"111100010",
  32569=>"110001011",
  32570=>"010001110",
  32571=>"011100010",
  32572=>"100111100",
  32573=>"101011011",
  32574=>"111011110",
  32575=>"100100110",
  32576=>"110101000",
  32577=>"110011011",
  32578=>"000001011",
  32579=>"101110100",
  32580=>"011000000",
  32581=>"001100000",
  32582=>"010100010",
  32583=>"111100001",
  32584=>"111111110",
  32585=>"100000000",
  32586=>"110010101",
  32587=>"001000000",
  32588=>"010001110",
  32589=>"101000001",
  32590=>"111110011",
  32591=>"110010111",
  32592=>"000100100",
  32593=>"011010101",
  32594=>"000000001",
  32595=>"101010001",
  32596=>"101001010",
  32597=>"011111000",
  32598=>"011001111",
  32599=>"111001011",
  32600=>"000001100",
  32601=>"101101100",
  32602=>"101001110",
  32603=>"110110000",
  32604=>"000001001",
  32605=>"010000101",
  32606=>"110110111",
  32607=>"110001111",
  32608=>"011100001",
  32609=>"001011000",
  32610=>"001000001",
  32611=>"010110110",
  32612=>"011100001",
  32613=>"010111001",
  32614=>"010110011",
  32615=>"111111010",
  32616=>"001011000",
  32617=>"111010100",
  32618=>"100111111",
  32619=>"110001000",
  32620=>"100001110",
  32621=>"000001010",
  32622=>"011110001",
  32623=>"101010011",
  32624=>"010110000",
  32625=>"111001101",
  32626=>"001101101",
  32627=>"111100010",
  32628=>"011010011",
  32629=>"110001000",
  32630=>"011111001",
  32631=>"111010100",
  32632=>"010101010",
  32633=>"110010111",
  32634=>"001000110",
  32635=>"000111001",
  32636=>"000000001",
  32637=>"101111010",
  32638=>"010001111",
  32639=>"000011001",
  32640=>"111101010",
  32641=>"010010100",
  32642=>"010000001",
  32643=>"101111001",
  32644=>"010110011",
  32645=>"110000001",
  32646=>"011010011",
  32647=>"100110111",
  32648=>"101110000",
  32649=>"010100101",
  32650=>"111110100",
  32651=>"111110010",
  32652=>"110011001",
  32653=>"001010010",
  32654=>"000100100",
  32655=>"111100100",
  32656=>"100100000",
  32657=>"110111110",
  32658=>"110111110",
  32659=>"100001111",
  32660=>"110001011",
  32661=>"010010111",
  32662=>"001000100",
  32663=>"000010110",
  32664=>"100001000",
  32665=>"000101101",
  32666=>"000110111",
  32667=>"101011010",
  32668=>"001000000",
  32669=>"011011000",
  32670=>"111100000",
  32671=>"010010001",
  32672=>"000111110",
  32673=>"101100101",
  32674=>"110000010",
  32675=>"110000111",
  32676=>"001110010",
  32677=>"111101111",
  32678=>"110011000",
  32679=>"011000000",
  32680=>"110101010",
  32681=>"000000100",
  32682=>"110100010",
  32683=>"011101100",
  32684=>"001000011",
  32685=>"000011110",
  32686=>"101000101",
  32687=>"110101010",
  32688=>"111000000",
  32689=>"101010001",
  32690=>"100101110",
  32691=>"000110010",
  32692=>"111111101",
  32693=>"111100110",
  32694=>"101010010",
  32695=>"001111101",
  32696=>"000100111",
  32697=>"111101111",
  32698=>"100010110",
  32699=>"100110111",
  32700=>"000100011",
  32701=>"010010010",
  32702=>"100101000",
  32703=>"111101101",
  32704=>"101010100",
  32705=>"001010011",
  32706=>"101101101",
  32707=>"001000011",
  32708=>"100100011",
  32709=>"110011111",
  32710=>"000110101",
  32711=>"010000101",
  32712=>"010000100",
  32713=>"011000001",
  32714=>"110001100",
  32715=>"110111011",
  32716=>"000101011",
  32717=>"001011001",
  32718=>"010110110",
  32719=>"001011000",
  32720=>"010000000",
  32721=>"011001000",
  32722=>"000101010",
  32723=>"001111111",
  32724=>"000000100",
  32725=>"010110011",
  32726=>"111100111",
  32727=>"011110010",
  32728=>"011000010",
  32729=>"111101011",
  32730=>"101101100",
  32731=>"100100110",
  32732=>"111111101",
  32733=>"001001001",
  32734=>"111110011",
  32735=>"000111011",
  32736=>"100100001",
  32737=>"111100001",
  32738=>"100010000",
  32739=>"001100000",
  32740=>"110101011",
  32741=>"101100010",
  32742=>"010001010",
  32743=>"100101010",
  32744=>"100010111",
  32745=>"110101011",
  32746=>"101100000",
  32747=>"111101111",
  32748=>"100000010",
  32749=>"111111111",
  32750=>"111100001",
  32751=>"100111111",
  32752=>"110010100",
  32753=>"111000001",
  32754=>"110101110",
  32755=>"111011110",
  32756=>"110000111",
  32757=>"101010000",
  32758=>"100110010",
  32759=>"010011111",
  32760=>"011111101",
  32761=>"110011101",
  32762=>"111011000",
  32763=>"110001011",
  32764=>"101000001",
  32765=>"110001101",
  32766=>"110010000",
  32767=>"000110101",
  32768=>"110010001",
  32769=>"010011010",
  32770=>"000001011",
  32771=>"001111110",
  32772=>"101000100",
  32773=>"000110010",
  32774=>"100001010",
  32775=>"010000000",
  32776=>"111100110",
  32777=>"001011001",
  32778=>"111010001",
  32779=>"101000100",
  32780=>"000000000",
  32781=>"111111010",
  32782=>"001000001",
  32783=>"100011001",
  32784=>"100011101",
  32785=>"001111100",
  32786=>"000001000",
  32787=>"000000110",
  32788=>"111100010",
  32789=>"010011000",
  32790=>"010010111",
  32791=>"010001111",
  32792=>"011010000",
  32793=>"111110111",
  32794=>"111010111",
  32795=>"010010000",
  32796=>"110101000",
  32797=>"110010101",
  32798=>"000110010",
  32799=>"100010011",
  32800=>"001111001",
  32801=>"010110011",
  32802=>"110011110",
  32803=>"011101110",
  32804=>"101001001",
  32805=>"110010101",
  32806=>"110110111",
  32807=>"111001110",
  32808=>"000010000",
  32809=>"100110000",
  32810=>"101000100",
  32811=>"100111011",
  32812=>"101001110",
  32813=>"011001110",
  32814=>"001110111",
  32815=>"101100110",
  32816=>"010111100",
  32817=>"111100110",
  32818=>"111100000",
  32819=>"010000101",
  32820=>"011001000",
  32821=>"100011000",
  32822=>"000000101",
  32823=>"011011000",
  32824=>"011111111",
  32825=>"000001100",
  32826=>"001111110",
  32827=>"111011000",
  32828=>"000010010",
  32829=>"011010111",
  32830=>"101011100",
  32831=>"011100101",
  32832=>"111010000",
  32833=>"000010100",
  32834=>"010101001",
  32835=>"100001110",
  32836=>"111101101",
  32837=>"101111011",
  32838=>"111110110",
  32839=>"011101001",
  32840=>"010010010",
  32841=>"111111100",
  32842=>"110101110",
  32843=>"100010111",
  32844=>"001101001",
  32845=>"111001001",
  32846=>"001011000",
  32847=>"000000011",
  32848=>"011010010",
  32849=>"101001111",
  32850=>"100010101",
  32851=>"010110000",
  32852=>"110011011",
  32853=>"011101011",
  32854=>"000001001",
  32855=>"100001010",
  32856=>"110111010",
  32857=>"001111010",
  32858=>"000101010",
  32859=>"011000000",
  32860=>"101011110",
  32861=>"110011011",
  32862=>"000000001",
  32863=>"001000111",
  32864=>"000100110",
  32865=>"000000110",
  32866=>"111101100",
  32867=>"110100011",
  32868=>"111011010",
  32869=>"001100011",
  32870=>"001111110",
  32871=>"001010101",
  32872=>"001010000",
  32873=>"011011001",
  32874=>"101101100",
  32875=>"011001101",
  32876=>"100011101",
  32877=>"100110010",
  32878=>"010000100",
  32879=>"101000000",
  32880=>"110000010",
  32881=>"000011111",
  32882=>"110001010",
  32883=>"111010101",
  32884=>"011111110",
  32885=>"100000111",
  32886=>"100111011",
  32887=>"011111110",
  32888=>"001000111",
  32889=>"000110000",
  32890=>"000111010",
  32891=>"001001010",
  32892=>"001010111",
  32893=>"111110111",
  32894=>"100100011",
  32895=>"000010000",
  32896=>"110000100",
  32897=>"011100101",
  32898=>"000111010",
  32899=>"010000000",
  32900=>"000000000",
  32901=>"011100011",
  32902=>"101011011",
  32903=>"100001010",
  32904=>"100010110",
  32905=>"100100000",
  32906=>"111101000",
  32907=>"110111110",
  32908=>"011000000",
  32909=>"110011100",
  32910=>"111000001",
  32911=>"001000001",
  32912=>"010111111",
  32913=>"110001111",
  32914=>"001001111",
  32915=>"010110001",
  32916=>"100010011",
  32917=>"010111111",
  32918=>"010110110",
  32919=>"000110000",
  32920=>"100001011",
  32921=>"111100010",
  32922=>"010010110",
  32923=>"010000000",
  32924=>"010010100",
  32925=>"100110110",
  32926=>"101101111",
  32927=>"000110011",
  32928=>"100110111",
  32929=>"011110010",
  32930=>"100101000",
  32931=>"010010010",
  32932=>"110101011",
  32933=>"000100001",
  32934=>"101110110",
  32935=>"010111101",
  32936=>"101011010",
  32937=>"100000000",
  32938=>"011101110",
  32939=>"111001101",
  32940=>"110001010",
  32941=>"110110110",
  32942=>"110111001",
  32943=>"000101001",
  32944=>"001001000",
  32945=>"000011011",
  32946=>"101100100",
  32947=>"011010010",
  32948=>"100001001",
  32949=>"100001111",
  32950=>"010101110",
  32951=>"100101111",
  32952=>"001100011",
  32953=>"100110110",
  32954=>"001000101",
  32955=>"000111110",
  32956=>"111000010",
  32957=>"001001010",
  32958=>"000001000",
  32959=>"010011110",
  32960=>"001011000",
  32961=>"111111000",
  32962=>"100011010",
  32963=>"010010100",
  32964=>"101100110",
  32965=>"100101111",
  32966=>"010011011",
  32967=>"000100010",
  32968=>"000010010",
  32969=>"110111001",
  32970=>"110010011",
  32971=>"111111110",
  32972=>"000111110",
  32973=>"110010100",
  32974=>"101110010",
  32975=>"101000100",
  32976=>"111100001",
  32977=>"101100110",
  32978=>"101110100",
  32979=>"011001001",
  32980=>"100101111",
  32981=>"101001110",
  32982=>"011111001",
  32983=>"110101010",
  32984=>"101000110",
  32985=>"000110100",
  32986=>"000000010",
  32987=>"000011000",
  32988=>"001110011",
  32989=>"000000100",
  32990=>"000000000",
  32991=>"010110010",
  32992=>"111001000",
  32993=>"101011101",
  32994=>"110001011",
  32995=>"000100110",
  32996=>"101101101",
  32997=>"001101001",
  32998=>"100001000",
  32999=>"110001101",
  33000=>"010010110",
  33001=>"010001111",
  33002=>"111101011",
  33003=>"101011011",
  33004=>"110000101",
  33005=>"000011010",
  33006=>"101100110",
  33007=>"000000000",
  33008=>"100001110",
  33009=>"101010011",
  33010=>"000110011",
  33011=>"001010101",
  33012=>"100100100",
  33013=>"001111110",
  33014=>"111010001",
  33015=>"000110000",
  33016=>"010101111",
  33017=>"100011101",
  33018=>"000110001",
  33019=>"000110000",
  33020=>"000100100",
  33021=>"100101100",
  33022=>"001011001",
  33023=>"110110001",
  33024=>"111011000",
  33025=>"000100001",
  33026=>"010111011",
  33027=>"111001100",
  33028=>"111111001",
  33029=>"100000101",
  33030=>"101011101",
  33031=>"000011111",
  33032=>"111110111",
  33033=>"111100100",
  33034=>"110110100",
  33035=>"100010000",
  33036=>"010011101",
  33037=>"011011101",
  33038=>"100010000",
  33039=>"000110011",
  33040=>"111110100",
  33041=>"111010010",
  33042=>"010101100",
  33043=>"001101010",
  33044=>"010011000",
  33045=>"000011110",
  33046=>"000000001",
  33047=>"110011011",
  33048=>"011100001",
  33049=>"101101000",
  33050=>"110011011",
  33051=>"000000000",
  33052=>"011001100",
  33053=>"100010001",
  33054=>"111111000",
  33055=>"100000111",
  33056=>"100110110",
  33057=>"100110010",
  33058=>"000111010",
  33059=>"011011111",
  33060=>"100011110",
  33061=>"110000010",
  33062=>"100011101",
  33063=>"111101010",
  33064=>"001101010",
  33065=>"110110100",
  33066=>"100011110",
  33067=>"001000011",
  33068=>"000000100",
  33069=>"000001111",
  33070=>"101101100",
  33071=>"010000111",
  33072=>"010011100",
  33073=>"101110010",
  33074=>"010001000",
  33075=>"011011101",
  33076=>"011010100",
  33077=>"011011101",
  33078=>"011101000",
  33079=>"000110110",
  33080=>"100110110",
  33081=>"001110000",
  33082=>"011001010",
  33083=>"110101001",
  33084=>"110000101",
  33085=>"010000110",
  33086=>"110101111",
  33087=>"001001001",
  33088=>"001001111",
  33089=>"010100100",
  33090=>"010000000",
  33091=>"111111110",
  33092=>"111011111",
  33093=>"100010011",
  33094=>"011111000",
  33095=>"011001001",
  33096=>"100010111",
  33097=>"101000101",
  33098=>"000110110",
  33099=>"010101111",
  33100=>"001111000",
  33101=>"101110101",
  33102=>"100000100",
  33103=>"101100100",
  33104=>"010100011",
  33105=>"000100011",
  33106=>"111110100",
  33107=>"110101100",
  33108=>"001010001",
  33109=>"110110101",
  33110=>"110101000",
  33111=>"100101010",
  33112=>"101001110",
  33113=>"000110111",
  33114=>"100011100",
  33115=>"001110100",
  33116=>"001100001",
  33117=>"111010001",
  33118=>"111001110",
  33119=>"101011010",
  33120=>"010010100",
  33121=>"000101111",
  33122=>"001100001",
  33123=>"000010111",
  33124=>"110111110",
  33125=>"011001110",
  33126=>"110101000",
  33127=>"010001101",
  33128=>"011000100",
  33129=>"001001111",
  33130=>"100011000",
  33131=>"010110010",
  33132=>"000001011",
  33133=>"111100111",
  33134=>"111111010",
  33135=>"010011101",
  33136=>"000000101",
  33137=>"010101101",
  33138=>"000101111",
  33139=>"101010100",
  33140=>"000100111",
  33141=>"110100101",
  33142=>"010111001",
  33143=>"101001110",
  33144=>"110111100",
  33145=>"010000101",
  33146=>"011011110",
  33147=>"100000011",
  33148=>"011011111",
  33149=>"111111010",
  33150=>"011011011",
  33151=>"101000010",
  33152=>"010111110",
  33153=>"011001100",
  33154=>"010011010",
  33155=>"001111100",
  33156=>"001001010",
  33157=>"001111000",
  33158=>"000110101",
  33159=>"011000011",
  33160=>"000101000",
  33161=>"100101100",
  33162=>"001100111",
  33163=>"100011111",
  33164=>"010000001",
  33165=>"100100010",
  33166=>"000001101",
  33167=>"010101010",
  33168=>"010000000",
  33169=>"000111011",
  33170=>"110110110",
  33171=>"001010011",
  33172=>"101001101",
  33173=>"001100111",
  33174=>"100001010",
  33175=>"000110011",
  33176=>"011000110",
  33177=>"100100101",
  33178=>"001111010",
  33179=>"100101000",
  33180=>"101001111",
  33181=>"100111011",
  33182=>"001111100",
  33183=>"111110001",
  33184=>"010111010",
  33185=>"010100010",
  33186=>"111001000",
  33187=>"000010001",
  33188=>"110010100",
  33189=>"011000010",
  33190=>"101000100",
  33191=>"111110100",
  33192=>"101000110",
  33193=>"011111000",
  33194=>"110111001",
  33195=>"101011010",
  33196=>"111111111",
  33197=>"100010000",
  33198=>"000100100",
  33199=>"110101111",
  33200=>"010100010",
  33201=>"110010111",
  33202=>"001101111",
  33203=>"110100110",
  33204=>"000011011",
  33205=>"101011011",
  33206=>"111011110",
  33207=>"110011010",
  33208=>"001010100",
  33209=>"001000001",
  33210=>"001100000",
  33211=>"111000000",
  33212=>"000100101",
  33213=>"000011101",
  33214=>"100100001",
  33215=>"100010011",
  33216=>"011001000",
  33217=>"011110000",
  33218=>"100011001",
  33219=>"010100100",
  33220=>"010100101",
  33221=>"101010100",
  33222=>"000001101",
  33223=>"010000100",
  33224=>"010110110",
  33225=>"011001110",
  33226=>"010010110",
  33227=>"111010000",
  33228=>"000111010",
  33229=>"101110000",
  33230=>"011110110",
  33231=>"101101110",
  33232=>"110111100",
  33233=>"000010000",
  33234=>"111010111",
  33235=>"000100001",
  33236=>"110101111",
  33237=>"110110110",
  33238=>"101010111",
  33239=>"111000100",
  33240=>"010000101",
  33241=>"011000010",
  33242=>"001111000",
  33243=>"110011010",
  33244=>"011000111",
  33245=>"010111010",
  33246=>"011000000",
  33247=>"010111011",
  33248=>"110001111",
  33249=>"010101000",
  33250=>"100111111",
  33251=>"010000010",
  33252=>"011101111",
  33253=>"100111111",
  33254=>"000110001",
  33255=>"100000000",
  33256=>"001100001",
  33257=>"111001101",
  33258=>"000001100",
  33259=>"010010010",
  33260=>"011000010",
  33261=>"001011000",
  33262=>"011110101",
  33263=>"101000001",
  33264=>"110010110",
  33265=>"100111001",
  33266=>"111110001",
  33267=>"011001001",
  33268=>"110100100",
  33269=>"110100111",
  33270=>"110001000",
  33271=>"110000001",
  33272=>"010011101",
  33273=>"111000011",
  33274=>"010011100",
  33275=>"110111110",
  33276=>"001010101",
  33277=>"010010001",
  33278=>"111111010",
  33279=>"101010111",
  33280=>"010111010",
  33281=>"001010010",
  33282=>"111011010",
  33283=>"000010111",
  33284=>"011101001",
  33285=>"001111000",
  33286=>"110000111",
  33287=>"101100110",
  33288=>"100111001",
  33289=>"010001110",
  33290=>"111101101",
  33291=>"111101010",
  33292=>"001000010",
  33293=>"010011101",
  33294=>"011000001",
  33295=>"111000010",
  33296=>"010011000",
  33297=>"111000011",
  33298=>"111111000",
  33299=>"001101110",
  33300=>"001100011",
  33301=>"001011000",
  33302=>"111011100",
  33303=>"001110000",
  33304=>"101111101",
  33305=>"001111100",
  33306=>"111101010",
  33307=>"001000011",
  33308=>"101010010",
  33309=>"100101111",
  33310=>"001100010",
  33311=>"010011001",
  33312=>"010000010",
  33313=>"000010101",
  33314=>"100010011",
  33315=>"010111111",
  33316=>"011010111",
  33317=>"011100011",
  33318=>"001000010",
  33319=>"111111001",
  33320=>"000001100",
  33321=>"000100000",
  33322=>"110110000",
  33323=>"010111010",
  33324=>"010110111",
  33325=>"000010101",
  33326=>"011011101",
  33327=>"010010110",
  33328=>"111011101",
  33329=>"100100001",
  33330=>"111000100",
  33331=>"101011000",
  33332=>"100010100",
  33333=>"111001011",
  33334=>"000101101",
  33335=>"000100110",
  33336=>"000100010",
  33337=>"010000110",
  33338=>"001011010",
  33339=>"011110001",
  33340=>"010100100",
  33341=>"011100001",
  33342=>"001011110",
  33343=>"001001101",
  33344=>"101101111",
  33345=>"000100100",
  33346=>"000110111",
  33347=>"001011110",
  33348=>"110010000",
  33349=>"101011000",
  33350=>"010100100",
  33351=>"000111001",
  33352=>"001000111",
  33353=>"110000110",
  33354=>"011101101",
  33355=>"101011111",
  33356=>"011100011",
  33357=>"111110010",
  33358=>"111001011",
  33359=>"000111011",
  33360=>"110001010",
  33361=>"000110010",
  33362=>"111100001",
  33363=>"000101111",
  33364=>"111110011",
  33365=>"011101001",
  33366=>"100001011",
  33367=>"010011111",
  33368=>"010110011",
  33369=>"111100111",
  33370=>"111000000",
  33371=>"001100010",
  33372=>"000110010",
  33373=>"110001101",
  33374=>"110010110",
  33375=>"010000100",
  33376=>"110011001",
  33377=>"011000011",
  33378=>"000000000",
  33379=>"101101010",
  33380=>"000100010",
  33381=>"111100111",
  33382=>"000000110",
  33383=>"011111111",
  33384=>"001001011",
  33385=>"010011001",
  33386=>"100110100",
  33387=>"001101110",
  33388=>"001001101",
  33389=>"001010011",
  33390=>"101110111",
  33391=>"110101101",
  33392=>"001010010",
  33393=>"000100010",
  33394=>"111001111",
  33395=>"010101100",
  33396=>"001000000",
  33397=>"001011011",
  33398=>"111110101",
  33399=>"001000111",
  33400=>"110110111",
  33401=>"001000110",
  33402=>"001111010",
  33403=>"110010111",
  33404=>"111101001",
  33405=>"110001110",
  33406=>"100001011",
  33407=>"000001111",
  33408=>"101001111",
  33409=>"101010010",
  33410=>"101010010",
  33411=>"011000011",
  33412=>"111100111",
  33413=>"111111001",
  33414=>"110100001",
  33415=>"101000011",
  33416=>"011000110",
  33417=>"000111011",
  33418=>"001010000",
  33419=>"100110011",
  33420=>"100110111",
  33421=>"100111100",
  33422=>"110111101",
  33423=>"111111110",
  33424=>"100100000",
  33425=>"110111101",
  33426=>"100100001",
  33427=>"110111100",
  33428=>"010001100",
  33429=>"111010010",
  33430=>"010000001",
  33431=>"010000011",
  33432=>"101011100",
  33433=>"010011100",
  33434=>"100110010",
  33435=>"011010111",
  33436=>"000011001",
  33437=>"011010111",
  33438=>"110001100",
  33439=>"100110011",
  33440=>"110011000",
  33441=>"011011111",
  33442=>"110110110",
  33443=>"011001011",
  33444=>"101011010",
  33445=>"011001000",
  33446=>"111110010",
  33447=>"000101100",
  33448=>"011011010",
  33449=>"000011111",
  33450=>"000101001",
  33451=>"110100111",
  33452=>"101111011",
  33453=>"011111000",
  33454=>"111111000",
  33455=>"010001000",
  33456=>"000101101",
  33457=>"000100101",
  33458=>"000111100",
  33459=>"000000001",
  33460=>"011000010",
  33461=>"110000110",
  33462=>"110110111",
  33463=>"001100110",
  33464=>"110101010",
  33465=>"111100111",
  33466=>"011110111",
  33467=>"100000001",
  33468=>"001100011",
  33469=>"111110111",
  33470=>"100010001",
  33471=>"101010100",
  33472=>"000101011",
  33473=>"011001111",
  33474=>"110001111",
  33475=>"011011001",
  33476=>"011000101",
  33477=>"001111010",
  33478=>"011100100",
  33479=>"001011011",
  33480=>"000100101",
  33481=>"001111101",
  33482=>"110011100",
  33483=>"001000001",
  33484=>"000111100",
  33485=>"111010011",
  33486=>"011000011",
  33487=>"001110111",
  33488=>"010101001",
  33489=>"101001000",
  33490=>"000010010",
  33491=>"000101011",
  33492=>"000110100",
  33493=>"011000101",
  33494=>"000001001",
  33495=>"101101101",
  33496=>"010001000",
  33497=>"000000011",
  33498=>"001000111",
  33499=>"111111001",
  33500=>"110110011",
  33501=>"000000110",
  33502=>"010111111",
  33503=>"011100101",
  33504=>"011111011",
  33505=>"010101111",
  33506=>"110111010",
  33507=>"110111011",
  33508=>"011001111",
  33509=>"111010100",
  33510=>"010001001",
  33511=>"000000100",
  33512=>"100111101",
  33513=>"110011111",
  33514=>"000011110",
  33515=>"111011001",
  33516=>"001100010",
  33517=>"100011100",
  33518=>"110011010",
  33519=>"001100101",
  33520=>"001100101",
  33521=>"101111100",
  33522=>"100000100",
  33523=>"110100001",
  33524=>"100010000",
  33525=>"100010001",
  33526=>"111011010",
  33527=>"000000011",
  33528=>"110110000",
  33529=>"110000001",
  33530=>"001011010",
  33531=>"101011110",
  33532=>"111000011",
  33533=>"011000101",
  33534=>"001100001",
  33535=>"001010001",
  33536=>"101011001",
  33537=>"101010000",
  33538=>"001001111",
  33539=>"101010001",
  33540=>"110000001",
  33541=>"010000001",
  33542=>"101011000",
  33543=>"001010000",
  33544=>"101001101",
  33545=>"011110010",
  33546=>"100010010",
  33547=>"000010001",
  33548=>"111010010",
  33549=>"000100101",
  33550=>"010000110",
  33551=>"011000010",
  33552=>"010100110",
  33553=>"111011101",
  33554=>"011101101",
  33555=>"000010101",
  33556=>"101010100",
  33557=>"101100110",
  33558=>"011101000",
  33559=>"100010111",
  33560=>"010110111",
  33561=>"001101001",
  33562=>"110001011",
  33563=>"000010001",
  33564=>"101111000",
  33565=>"010100000",
  33566=>"101010100",
  33567=>"010100001",
  33568=>"010011110",
  33569=>"111010111",
  33570=>"001100101",
  33571=>"010011001",
  33572=>"000000101",
  33573=>"100001000",
  33574=>"101101101",
  33575=>"111010100",
  33576=>"001111011",
  33577=>"011101000",
  33578=>"100000001",
  33579=>"100000101",
  33580=>"101001010",
  33581=>"111011111",
  33582=>"000011010",
  33583=>"110110011",
  33584=>"101101010",
  33585=>"111101011",
  33586=>"101101010",
  33587=>"000010000",
  33588=>"101100111",
  33589=>"101000010",
  33590=>"110000011",
  33591=>"001100000",
  33592=>"011101011",
  33593=>"001101000",
  33594=>"100011000",
  33595=>"011001110",
  33596=>"101100100",
  33597=>"000111101",
  33598=>"001110001",
  33599=>"101110110",
  33600=>"100010000",
  33601=>"001111011",
  33602=>"011111011",
  33603=>"110111011",
  33604=>"101000011",
  33605=>"000011001",
  33606=>"011100001",
  33607=>"001101101",
  33608=>"110000101",
  33609=>"100000100",
  33610=>"011011101",
  33611=>"101011001",
  33612=>"111100111",
  33613=>"111011110",
  33614=>"110100110",
  33615=>"011111111",
  33616=>"001010110",
  33617=>"110101010",
  33618=>"100010111",
  33619=>"000010011",
  33620=>"010100010",
  33621=>"100101100",
  33622=>"101000100",
  33623=>"101111110",
  33624=>"010100110",
  33625=>"110111100",
  33626=>"000011010",
  33627=>"011011011",
  33628=>"001011111",
  33629=>"111110001",
  33630=>"001111011",
  33631=>"100100111",
  33632=>"011100100",
  33633=>"010101110",
  33634=>"001001010",
  33635=>"110101100",
  33636=>"010011010",
  33637=>"000010110",
  33638=>"100010000",
  33639=>"100100000",
  33640=>"111000001",
  33641=>"001111010",
  33642=>"001110100",
  33643=>"011011111",
  33644=>"000000101",
  33645=>"101010000",
  33646=>"001001000",
  33647=>"000001101",
  33648=>"100110101",
  33649=>"100000111",
  33650=>"000010001",
  33651=>"010111111",
  33652=>"001001000",
  33653=>"110101110",
  33654=>"001001001",
  33655=>"100001011",
  33656=>"000000010",
  33657=>"101010010",
  33658=>"001101000",
  33659=>"111110000",
  33660=>"001000000",
  33661=>"011000000",
  33662=>"011000010",
  33663=>"010001001",
  33664=>"101111100",
  33665=>"001010110",
  33666=>"010101010",
  33667=>"100011011",
  33668=>"111110111",
  33669=>"110010011",
  33670=>"000100101",
  33671=>"111000000",
  33672=>"011110010",
  33673=>"000100111",
  33674=>"111100011",
  33675=>"110101100",
  33676=>"000110101",
  33677=>"000101000",
  33678=>"110110100",
  33679=>"100010001",
  33680=>"100111001",
  33681=>"111111111",
  33682=>"000001100",
  33683=>"011000000",
  33684=>"100000001",
  33685=>"110010100",
  33686=>"001000100",
  33687=>"100001001",
  33688=>"110101001",
  33689=>"100010010",
  33690=>"111011101",
  33691=>"010010001",
  33692=>"010111010",
  33693=>"000000100",
  33694=>"000100101",
  33695=>"010110011",
  33696=>"111000000",
  33697=>"101101110",
  33698=>"100100010",
  33699=>"011110010",
  33700=>"001111110",
  33701=>"101100001",
  33702=>"100110111",
  33703=>"000100100",
  33704=>"100111111",
  33705=>"000001110",
  33706=>"101101000",
  33707=>"111000010",
  33708=>"000000111",
  33709=>"010111000",
  33710=>"000111110",
  33711=>"100111111",
  33712=>"011110001",
  33713=>"111110101",
  33714=>"111011011",
  33715=>"111110001",
  33716=>"010101101",
  33717=>"100101101",
  33718=>"000101010",
  33719=>"001011111",
  33720=>"000100110",
  33721=>"100010110",
  33722=>"000110011",
  33723=>"000110000",
  33724=>"100101000",
  33725=>"101101000",
  33726=>"000011000",
  33727=>"011100100",
  33728=>"111001110",
  33729=>"010101011",
  33730=>"000110100",
  33731=>"100111010",
  33732=>"011101000",
  33733=>"111010111",
  33734=>"101111011",
  33735=>"011000011",
  33736=>"101010000",
  33737=>"010000000",
  33738=>"111011001",
  33739=>"000000100",
  33740=>"100011010",
  33741=>"110110000",
  33742=>"000011111",
  33743=>"011000110",
  33744=>"101111111",
  33745=>"000111000",
  33746=>"111111000",
  33747=>"111101100",
  33748=>"100000010",
  33749=>"010010001",
  33750=>"101101100",
  33751=>"010111101",
  33752=>"111111110",
  33753=>"100111111",
  33754=>"100101000",
  33755=>"010000001",
  33756=>"101101011",
  33757=>"011001010",
  33758=>"010101011",
  33759=>"010001000",
  33760=>"010111011",
  33761=>"011010011",
  33762=>"000011000",
  33763=>"011010001",
  33764=>"010110000",
  33765=>"101100111",
  33766=>"111100011",
  33767=>"010010011",
  33768=>"101000101",
  33769=>"000010111",
  33770=>"010101001",
  33771=>"010011011",
  33772=>"010011000",
  33773=>"101001110",
  33774=>"101001101",
  33775=>"100010101",
  33776=>"011011011",
  33777=>"001111000",
  33778=>"010001011",
  33779=>"001100111",
  33780=>"101110100",
  33781=>"000110000",
  33782=>"100101001",
  33783=>"101111000",
  33784=>"000100101",
  33785=>"100010101",
  33786=>"010000100",
  33787=>"111011110",
  33788=>"100000010",
  33789=>"111111111",
  33790=>"010101111",
  33791=>"000111000",
  33792=>"011000000",
  33793=>"100111100",
  33794=>"011100000",
  33795=>"101100101",
  33796=>"000000111",
  33797=>"001111111",
  33798=>"110100010",
  33799=>"111110100",
  33800=>"010111100",
  33801=>"011000101",
  33802=>"010001011",
  33803=>"011110011",
  33804=>"110000111",
  33805=>"001100011",
  33806=>"011100000",
  33807=>"000000000",
  33808=>"011100111",
  33809=>"000100011",
  33810=>"101000110",
  33811=>"110000000",
  33812=>"010110010",
  33813=>"000000111",
  33814=>"000000110",
  33815=>"111011110",
  33816=>"110100001",
  33817=>"000101011",
  33818=>"000100010",
  33819=>"101111111",
  33820=>"111111110",
  33821=>"111100011",
  33822=>"000101010",
  33823=>"101000000",
  33824=>"000010110",
  33825=>"100010100",
  33826=>"000100010",
  33827=>"111110110",
  33828=>"111010001",
  33829=>"101100010",
  33830=>"001110100",
  33831=>"100101101",
  33832=>"101011010",
  33833=>"011100010",
  33834=>"111001011",
  33835=>"001110101",
  33836=>"101010000",
  33837=>"000001010",
  33838=>"111110010",
  33839=>"010001101",
  33840=>"001100001",
  33841=>"010010000",
  33842=>"011110010",
  33843=>"011111110",
  33844=>"100100110",
  33845=>"010011101",
  33846=>"001000000",
  33847=>"010110001",
  33848=>"001000101",
  33849=>"100100011",
  33850=>"100111011",
  33851=>"001010110",
  33852=>"011011000",
  33853=>"111000000",
  33854=>"000110011",
  33855=>"011111100",
  33856=>"001011000",
  33857=>"000011001",
  33858=>"111000000",
  33859=>"110000000",
  33860=>"111010101",
  33861=>"100010001",
  33862=>"000101111",
  33863=>"010111100",
  33864=>"011110010",
  33865=>"100010100",
  33866=>"010011001",
  33867=>"100001000",
  33868=>"010100010",
  33869=>"000011110",
  33870=>"111110110",
  33871=>"001110011",
  33872=>"011100010",
  33873=>"011111001",
  33874=>"111001100",
  33875=>"001111101",
  33876=>"101110101",
  33877=>"111000001",
  33878=>"101001110",
  33879=>"001100001",
  33880=>"101000011",
  33881=>"110010010",
  33882=>"010101011",
  33883=>"100001101",
  33884=>"001000011",
  33885=>"011011010",
  33886=>"010001001",
  33887=>"000111011",
  33888=>"000000011",
  33889=>"100010110",
  33890=>"111100111",
  33891=>"101001110",
  33892=>"100110101",
  33893=>"100010001",
  33894=>"010111011",
  33895=>"011011001",
  33896=>"100100001",
  33897=>"101001000",
  33898=>"111110001",
  33899=>"001101111",
  33900=>"000101110",
  33901=>"110010100",
  33902=>"100101001",
  33903=>"011011111",
  33904=>"010000011",
  33905=>"010010001",
  33906=>"101110010",
  33907=>"100111001",
  33908=>"100010011",
  33909=>"101000101",
  33910=>"001000110",
  33911=>"100100111",
  33912=>"010111110",
  33913=>"000001111",
  33914=>"001001010",
  33915=>"010110111",
  33916=>"000101011",
  33917=>"111101111",
  33918=>"010101001",
  33919=>"010101101",
  33920=>"000101111",
  33921=>"011110011",
  33922=>"011100001",
  33923=>"011000000",
  33924=>"000001111",
  33925=>"011110001",
  33926=>"111011100",
  33927=>"111010001",
  33928=>"011110001",
  33929=>"110101100",
  33930=>"010011011",
  33931=>"001001000",
  33932=>"011010000",
  33933=>"010000001",
  33934=>"111000001",
  33935=>"110001001",
  33936=>"010111000",
  33937=>"010011000",
  33938=>"000101111",
  33939=>"110000011",
  33940=>"011000100",
  33941=>"001100100",
  33942=>"111101111",
  33943=>"110000100",
  33944=>"011100111",
  33945=>"011101100",
  33946=>"011110000",
  33947=>"011111001",
  33948=>"111101010",
  33949=>"100010100",
  33950=>"011101110",
  33951=>"001011001",
  33952=>"111101000",
  33953=>"000011110",
  33954=>"001100110",
  33955=>"010001000",
  33956=>"010110111",
  33957=>"110100101",
  33958=>"100000011",
  33959=>"001100100",
  33960=>"000011000",
  33961=>"001001100",
  33962=>"111111010",
  33963=>"110000000",
  33964=>"011000010",
  33965=>"100101111",
  33966=>"001011111",
  33967=>"001000010",
  33968=>"011000101",
  33969=>"010000010",
  33970=>"110001001",
  33971=>"011110101",
  33972=>"110110000",
  33973=>"110100110",
  33974=>"101110000",
  33975=>"100001110",
  33976=>"110100010",
  33977=>"011010101",
  33978=>"000000010",
  33979=>"100111010",
  33980=>"110100111",
  33981=>"011110000",
  33982=>"100010011",
  33983=>"011100101",
  33984=>"111010011",
  33985=>"001110111",
  33986=>"011010110",
  33987=>"110100111",
  33988=>"111101101",
  33989=>"101100011",
  33990=>"000001110",
  33991=>"110000000",
  33992=>"010011100",
  33993=>"110010111",
  33994=>"101000010",
  33995=>"000110011",
  33996=>"110111010",
  33997=>"010001101",
  33998=>"010111000",
  33999=>"111011111",
  34000=>"011100101",
  34001=>"000011101",
  34002=>"000111110",
  34003=>"011011001",
  34004=>"101010011",
  34005=>"011000011",
  34006=>"001100110",
  34007=>"111101100",
  34008=>"110001000",
  34009=>"101010000",
  34010=>"001011001",
  34011=>"110010110",
  34012=>"101001011",
  34013=>"111100111",
  34014=>"000010001",
  34015=>"110000111",
  34016=>"111001000",
  34017=>"010000000",
  34018=>"010010111",
  34019=>"100011000",
  34020=>"000010010",
  34021=>"101110011",
  34022=>"001110010",
  34023=>"000000101",
  34024=>"111101000",
  34025=>"100110010",
  34026=>"011011001",
  34027=>"110001000",
  34028=>"110011000",
  34029=>"011011011",
  34030=>"011011001",
  34031=>"010110110",
  34032=>"101010100",
  34033=>"110111111",
  34034=>"011101010",
  34035=>"010101100",
  34036=>"000111111",
  34037=>"010010110",
  34038=>"011100001",
  34039=>"101001011",
  34040=>"010010000",
  34041=>"000100101",
  34042=>"011101100",
  34043=>"010001001",
  34044=>"000100000",
  34045=>"011100111",
  34046=>"001100100",
  34047=>"111011111",
  34048=>"111011101",
  34049=>"110000011",
  34050=>"111010000",
  34051=>"111000001",
  34052=>"100001101",
  34053=>"011001100",
  34054=>"000011100",
  34055=>"100110100",
  34056=>"101010000",
  34057=>"111010000",
  34058=>"000010111",
  34059=>"001000011",
  34060=>"110011001",
  34061=>"011011101",
  34062=>"001100111",
  34063=>"110110011",
  34064=>"001010000",
  34065=>"011010100",
  34066=>"010001100",
  34067=>"111101111",
  34068=>"011100100",
  34069=>"101100000",
  34070=>"111010000",
  34071=>"100000110",
  34072=>"001011010",
  34073=>"010010100",
  34074=>"100001001",
  34075=>"101011011",
  34076=>"011001111",
  34077=>"010111101",
  34078=>"110011100",
  34079=>"100100111",
  34080=>"111100110",
  34081=>"100111001",
  34082=>"001001110",
  34083=>"011101111",
  34084=>"000010010",
  34085=>"010111101",
  34086=>"101100101",
  34087=>"010110110",
  34088=>"000000000",
  34089=>"110110101",
  34090=>"011010010",
  34091=>"100001000",
  34092=>"111101001",
  34093=>"110100000",
  34094=>"100001110",
  34095=>"000001000",
  34096=>"000000110",
  34097=>"000100111",
  34098=>"001110100",
  34099=>"101110101",
  34100=>"011011101",
  34101=>"000001000",
  34102=>"001010001",
  34103=>"000101010",
  34104=>"110001110",
  34105=>"110000100",
  34106=>"110101110",
  34107=>"111100010",
  34108=>"011001101",
  34109=>"011010110",
  34110=>"110101000",
  34111=>"111110100",
  34112=>"011001101",
  34113=>"100011010",
  34114=>"000010001",
  34115=>"100011000",
  34116=>"110011010",
  34117=>"000000100",
  34118=>"110101111",
  34119=>"111100000",
  34120=>"101010010",
  34121=>"011100001",
  34122=>"110010001",
  34123=>"110001000",
  34124=>"000100111",
  34125=>"011011100",
  34126=>"001010001",
  34127=>"011100000",
  34128=>"010010001",
  34129=>"110000010",
  34130=>"111010101",
  34131=>"011101111",
  34132=>"111001111",
  34133=>"111101000",
  34134=>"101000010",
  34135=>"111000010",
  34136=>"000000000",
  34137=>"011111010",
  34138=>"101001011",
  34139=>"011100000",
  34140=>"001110001",
  34141=>"011110110",
  34142=>"011100101",
  34143=>"110011101",
  34144=>"010011000",
  34145=>"010010010",
  34146=>"111100001",
  34147=>"100111111",
  34148=>"110110000",
  34149=>"011100000",
  34150=>"101000111",
  34151=>"101010110",
  34152=>"110101110",
  34153=>"000011000",
  34154=>"101011101",
  34155=>"110110010",
  34156=>"000110010",
  34157=>"001010101",
  34158=>"111100100",
  34159=>"000001110",
  34160=>"110011000",
  34161=>"000001110",
  34162=>"110011000",
  34163=>"111001011",
  34164=>"001100010",
  34165=>"111000100",
  34166=>"000001100",
  34167=>"100010011",
  34168=>"010011010",
  34169=>"100101101",
  34170=>"100111101",
  34171=>"100110011",
  34172=>"000010010",
  34173=>"011101010",
  34174=>"110001100",
  34175=>"100000000",
  34176=>"111111111",
  34177=>"100111000",
  34178=>"110100111",
  34179=>"000011011",
  34180=>"100010110",
  34181=>"011110001",
  34182=>"100000010",
  34183=>"011110010",
  34184=>"101011100",
  34185=>"001110000",
  34186=>"110111110",
  34187=>"111111101",
  34188=>"101000100",
  34189=>"101010011",
  34190=>"000010011",
  34191=>"000010010",
  34192=>"110010100",
  34193=>"000111100",
  34194=>"100101111",
  34195=>"101011000",
  34196=>"111110101",
  34197=>"011011010",
  34198=>"001100101",
  34199=>"011101000",
  34200=>"000110101",
  34201=>"000101101",
  34202=>"010000011",
  34203=>"000001100",
  34204=>"111001101",
  34205=>"010000110",
  34206=>"101100010",
  34207=>"101110011",
  34208=>"010011001",
  34209=>"011111000",
  34210=>"001111011",
  34211=>"100101101",
  34212=>"111100011",
  34213=>"010000101",
  34214=>"110001101",
  34215=>"010100010",
  34216=>"101101000",
  34217=>"100011010",
  34218=>"100111110",
  34219=>"010010100",
  34220=>"000111100",
  34221=>"100101111",
  34222=>"111011010",
  34223=>"011011001",
  34224=>"001010010",
  34225=>"110010111",
  34226=>"111001110",
  34227=>"010010010",
  34228=>"110101010",
  34229=>"000101101",
  34230=>"111101010",
  34231=>"111001001",
  34232=>"001101111",
  34233=>"101110001",
  34234=>"101110111",
  34235=>"001011110",
  34236=>"101101100",
  34237=>"001101111",
  34238=>"111101010",
  34239=>"011100001",
  34240=>"011011010",
  34241=>"001111001",
  34242=>"010001011",
  34243=>"010101011",
  34244=>"111000011",
  34245=>"100000100",
  34246=>"110101011",
  34247=>"001110010",
  34248=>"111101111",
  34249=>"100010000",
  34250=>"011000101",
  34251=>"011001111",
  34252=>"011110010",
  34253=>"001011011",
  34254=>"000000001",
  34255=>"111101100",
  34256=>"100010100",
  34257=>"011101110",
  34258=>"010010101",
  34259=>"101110110",
  34260=>"010010010",
  34261=>"010011110",
  34262=>"011101111",
  34263=>"111110000",
  34264=>"010111100",
  34265=>"010101111",
  34266=>"011000000",
  34267=>"101010100",
  34268=>"010100010",
  34269=>"000111110",
  34270=>"000010111",
  34271=>"110111111",
  34272=>"111111011",
  34273=>"111011110",
  34274=>"110101110",
  34275=>"100010011",
  34276=>"011110001",
  34277=>"011111111",
  34278=>"100110001",
  34279=>"001011100",
  34280=>"001001110",
  34281=>"110001000",
  34282=>"000010000",
  34283=>"111010110",
  34284=>"010110101",
  34285=>"110111100",
  34286=>"100010010",
  34287=>"011110010",
  34288=>"011000001",
  34289=>"110111100",
  34290=>"100111101",
  34291=>"000010010",
  34292=>"000010011",
  34293=>"110001100",
  34294=>"011111101",
  34295=>"111101110",
  34296=>"110111111",
  34297=>"011001000",
  34298=>"111001000",
  34299=>"111000001",
  34300=>"111100111",
  34301=>"011110100",
  34302=>"111110111",
  34303=>"111111111",
  34304=>"011100001",
  34305=>"101010010",
  34306=>"010010101",
  34307=>"100000101",
  34308=>"011101101",
  34309=>"000010010",
  34310=>"111100111",
  34311=>"001010111",
  34312=>"101100011",
  34313=>"101100011",
  34314=>"110011000",
  34315=>"001110101",
  34316=>"000001111",
  34317=>"111010010",
  34318=>"010100100",
  34319=>"111000110",
  34320=>"010000101",
  34321=>"110110011",
  34322=>"001101010",
  34323=>"001010110",
  34324=>"101000000",
  34325=>"100011001",
  34326=>"101101100",
  34327=>"010100111",
  34328=>"111010110",
  34329=>"100110010",
  34330=>"000011000",
  34331=>"101011000",
  34332=>"001001100",
  34333=>"000000110",
  34334=>"101111101",
  34335=>"001110001",
  34336=>"001000111",
  34337=>"000001001",
  34338=>"011110101",
  34339=>"010010001",
  34340=>"001000110",
  34341=>"001100011",
  34342=>"111111100",
  34343=>"001011111",
  34344=>"101011110",
  34345=>"000111111",
  34346=>"011111111",
  34347=>"010001011",
  34348=>"110111110",
  34349=>"110001001",
  34350=>"010111100",
  34351=>"001010111",
  34352=>"011110101",
  34353=>"001100000",
  34354=>"010010000",
  34355=>"010110011",
  34356=>"111100011",
  34357=>"000100110",
  34358=>"000001111",
  34359=>"101110010",
  34360=>"000100001",
  34361=>"000100111",
  34362=>"100100000",
  34363=>"111100111",
  34364=>"001111000",
  34365=>"111010100",
  34366=>"111101111",
  34367=>"110010000",
  34368=>"101000101",
  34369=>"010001001",
  34370=>"101000111",
  34371=>"110111111",
  34372=>"011010000",
  34373=>"011001100",
  34374=>"000100000",
  34375=>"101000000",
  34376=>"101110010",
  34377=>"110001110",
  34378=>"010000011",
  34379=>"100111110",
  34380=>"000000111",
  34381=>"010011100",
  34382=>"000010010",
  34383=>"111110010",
  34384=>"000111101",
  34385=>"110010000",
  34386=>"101101111",
  34387=>"111010000",
  34388=>"001000000",
  34389=>"010011001",
  34390=>"100110011",
  34391=>"111011110",
  34392=>"010100010",
  34393=>"111101100",
  34394=>"111111000",
  34395=>"010001110",
  34396=>"010011100",
  34397=>"000000110",
  34398=>"100100000",
  34399=>"100000100",
  34400=>"000111110",
  34401=>"100000010",
  34402=>"111011001",
  34403=>"010000101",
  34404=>"111010010",
  34405=>"000010110",
  34406=>"100011000",
  34407=>"000011011",
  34408=>"110000100",
  34409=>"111110101",
  34410=>"111101011",
  34411=>"110000010",
  34412=>"100111111",
  34413=>"111010001",
  34414=>"000100011",
  34415=>"011101101",
  34416=>"101110001",
  34417=>"010111100",
  34418=>"010101110",
  34419=>"010000010",
  34420=>"000000001",
  34421=>"010000110",
  34422=>"011001111",
  34423=>"110111000",
  34424=>"110010100",
  34425=>"110101101",
  34426=>"000011111",
  34427=>"000111110",
  34428=>"000000110",
  34429=>"011001111",
  34430=>"100111100",
  34431=>"100101011",
  34432=>"001110001",
  34433=>"110110001",
  34434=>"100110001",
  34435=>"111111111",
  34436=>"011111100",
  34437=>"111101100",
  34438=>"001100010",
  34439=>"111111010",
  34440=>"101000000",
  34441=>"001101000",
  34442=>"000000001",
  34443=>"110011110",
  34444=>"010010100",
  34445=>"101110000",
  34446=>"110000111",
  34447=>"001100010",
  34448=>"011110111",
  34449=>"110001010",
  34450=>"010101110",
  34451=>"011001000",
  34452=>"011011010",
  34453=>"010101101",
  34454=>"111101111",
  34455=>"011111111",
  34456=>"100100000",
  34457=>"111100111",
  34458=>"000011111",
  34459=>"101111010",
  34460=>"010110111",
  34461=>"000100100",
  34462=>"101000010",
  34463=>"011000101",
  34464=>"001111111",
  34465=>"010001111",
  34466=>"010010011",
  34467=>"001011101",
  34468=>"000001111",
  34469=>"010000100",
  34470=>"011100011",
  34471=>"010101111",
  34472=>"101001111",
  34473=>"000001011",
  34474=>"100101011",
  34475=>"010100010",
  34476=>"110011111",
  34477=>"011011000",
  34478=>"000111000",
  34479=>"110111101",
  34480=>"011001100",
  34481=>"111010010",
  34482=>"011111111",
  34483=>"110101001",
  34484=>"011110010",
  34485=>"101101011",
  34486=>"110100110",
  34487=>"010000011",
  34488=>"101111111",
  34489=>"011100010",
  34490=>"011011111",
  34491=>"111110000",
  34492=>"001000101",
  34493=>"111110101",
  34494=>"011111110",
  34495=>"111111110",
  34496=>"001100101",
  34497=>"111111011",
  34498=>"001010000",
  34499=>"101100101",
  34500=>"011000010",
  34501=>"000101010",
  34502=>"001110110",
  34503=>"000111000",
  34504=>"110011000",
  34505=>"001000011",
  34506=>"011110010",
  34507=>"000101101",
  34508=>"001000111",
  34509=>"000110010",
  34510=>"011000110",
  34511=>"100010000",
  34512=>"010101010",
  34513=>"010000011",
  34514=>"100101100",
  34515=>"000110000",
  34516=>"011101011",
  34517=>"000111111",
  34518=>"010000000",
  34519=>"011110111",
  34520=>"000110010",
  34521=>"001111000",
  34522=>"000010011",
  34523=>"100001101",
  34524=>"110011111",
  34525=>"011000110",
  34526=>"101110000",
  34527=>"011111010",
  34528=>"010111110",
  34529=>"100000100",
  34530=>"100000001",
  34531=>"111010000",
  34532=>"000111100",
  34533=>"000010001",
  34534=>"001001100",
  34535=>"111111001",
  34536=>"101001001",
  34537=>"000001011",
  34538=>"100111111",
  34539=>"011010111",
  34540=>"000001010",
  34541=>"011100100",
  34542=>"111001001",
  34543=>"001111000",
  34544=>"111010100",
  34545=>"100010100",
  34546=>"000000100",
  34547=>"100101101",
  34548=>"101000100",
  34549=>"110110010",
  34550=>"111100011",
  34551=>"000000000",
  34552=>"011010000",
  34553=>"111110111",
  34554=>"111111100",
  34555=>"100000110",
  34556=>"001011000",
  34557=>"001011110",
  34558=>"100111000",
  34559=>"010101000",
  34560=>"001011011",
  34561=>"100010110",
  34562=>"110100010",
  34563=>"101001011",
  34564=>"111100010",
  34565=>"000000100",
  34566=>"110110010",
  34567=>"111011000",
  34568=>"001010100",
  34569=>"010011100",
  34570=>"011101000",
  34571=>"011011001",
  34572=>"001101110",
  34573=>"110111100",
  34574=>"010001001",
  34575=>"111110010",
  34576=>"010100101",
  34577=>"000100010",
  34578=>"011111100",
  34579=>"110000101",
  34580=>"101011110",
  34581=>"110010110",
  34582=>"001011001",
  34583=>"000100001",
  34584=>"000111100",
  34585=>"001010110",
  34586=>"100101101",
  34587=>"110000110",
  34588=>"000000011",
  34589=>"111111100",
  34590=>"110010000",
  34591=>"011100110",
  34592=>"110100111",
  34593=>"011001101",
  34594=>"111011011",
  34595=>"000101001",
  34596=>"011110111",
  34597=>"100000100",
  34598=>"011001100",
  34599=>"100001000",
  34600=>"100010111",
  34601=>"010001011",
  34602=>"111010010",
  34603=>"101011111",
  34604=>"111010001",
  34605=>"100101100",
  34606=>"111011110",
  34607=>"100011101",
  34608=>"001100100",
  34609=>"101010101",
  34610=>"000111100",
  34611=>"100001001",
  34612=>"000100100",
  34613=>"100011101",
  34614=>"001001110",
  34615=>"100111111",
  34616=>"101110001",
  34617=>"110001010",
  34618=>"011100111",
  34619=>"000100110",
  34620=>"100100010",
  34621=>"010000000",
  34622=>"100010000",
  34623=>"000001101",
  34624=>"000110000",
  34625=>"100010010",
  34626=>"101010100",
  34627=>"101110111",
  34628=>"001100101",
  34629=>"011000111",
  34630=>"111000101",
  34631=>"000101101",
  34632=>"100101110",
  34633=>"110110111",
  34634=>"001001000",
  34635=>"001000011",
  34636=>"010011100",
  34637=>"111110001",
  34638=>"000010110",
  34639=>"110011000",
  34640=>"000010100",
  34641=>"010111100",
  34642=>"000010100",
  34643=>"010101000",
  34644=>"101100100",
  34645=>"110011000",
  34646=>"000110010",
  34647=>"100101100",
  34648=>"110000110",
  34649=>"011000110",
  34650=>"011001100",
  34651=>"100111010",
  34652=>"101000110",
  34653=>"110111000",
  34654=>"011001111",
  34655=>"011111010",
  34656=>"100011011",
  34657=>"011100000",
  34658=>"111101010",
  34659=>"001100111",
  34660=>"011110011",
  34661=>"111011101",
  34662=>"001110111",
  34663=>"110101101",
  34664=>"000100111",
  34665=>"010001001",
  34666=>"100000000",
  34667=>"010110001",
  34668=>"001010001",
  34669=>"001110100",
  34670=>"100001101",
  34671=>"110001100",
  34672=>"010110010",
  34673=>"111110001",
  34674=>"110011101",
  34675=>"000101100",
  34676=>"010000101",
  34677=>"101011100",
  34678=>"001001010",
  34679=>"110110110",
  34680=>"110111101",
  34681=>"011100001",
  34682=>"111100011",
  34683=>"111101110",
  34684=>"100010000",
  34685=>"101110011",
  34686=>"111010010",
  34687=>"100011100",
  34688=>"011111001",
  34689=>"110100011",
  34690=>"000100111",
  34691=>"001001010",
  34692=>"011110011",
  34693=>"001000110",
  34694=>"111011000",
  34695=>"111001100",
  34696=>"000010110",
  34697=>"110001011",
  34698=>"111011111",
  34699=>"011000001",
  34700=>"101101111",
  34701=>"101000000",
  34702=>"100000110",
  34703=>"001010000",
  34704=>"101110001",
  34705=>"100001111",
  34706=>"000011110",
  34707=>"101011011",
  34708=>"001000000",
  34709=>"111110011",
  34710=>"011011011",
  34711=>"111111010",
  34712=>"111111110",
  34713=>"111001011",
  34714=>"111101010",
  34715=>"101011011",
  34716=>"110100100",
  34717=>"001000111",
  34718=>"101110100",
  34719=>"100011010",
  34720=>"101100110",
  34721=>"011001011",
  34722=>"101111011",
  34723=>"000010110",
  34724=>"100011010",
  34725=>"011111100",
  34726=>"111001011",
  34727=>"010100000",
  34728=>"011101010",
  34729=>"101110101",
  34730=>"100010011",
  34731=>"111101001",
  34732=>"010101001",
  34733=>"010100001",
  34734=>"110010011",
  34735=>"110100010",
  34736=>"000110111",
  34737=>"011011111",
  34738=>"001010010",
  34739=>"011110011",
  34740=>"110100111",
  34741=>"101111011",
  34742=>"000010011",
  34743=>"101011101",
  34744=>"100101111",
  34745=>"111100101",
  34746=>"101101110",
  34747=>"010001101",
  34748=>"101000010",
  34749=>"010100001",
  34750=>"000000111",
  34751=>"001000100",
  34752=>"011010011",
  34753=>"100000101",
  34754=>"100011011",
  34755=>"010011000",
  34756=>"100110110",
  34757=>"101001101",
  34758=>"111010100",
  34759=>"111001110",
  34760=>"000100001",
  34761=>"100111000",
  34762=>"101110001",
  34763=>"110001011",
  34764=>"101010001",
  34765=>"011100001",
  34766=>"110110111",
  34767=>"010110110",
  34768=>"111111010",
  34769=>"000001110",
  34770=>"101111010",
  34771=>"000011001",
  34772=>"010100010",
  34773=>"001000001",
  34774=>"100000010",
  34775=>"111000001",
  34776=>"111011001",
  34777=>"011011111",
  34778=>"010010001",
  34779=>"100000111",
  34780=>"011001001",
  34781=>"011000101",
  34782=>"010010001",
  34783=>"101000010",
  34784=>"100100011",
  34785=>"100001100",
  34786=>"011001110",
  34787=>"100011011",
  34788=>"110011000",
  34789=>"111001000",
  34790=>"001111111",
  34791=>"000000011",
  34792=>"101011111",
  34793=>"111111101",
  34794=>"111010001",
  34795=>"000001101",
  34796=>"000100100",
  34797=>"111000000",
  34798=>"111101011",
  34799=>"110000111",
  34800=>"001000011",
  34801=>"100011110",
  34802=>"110100110",
  34803=>"100101010",
  34804=>"100110101",
  34805=>"110111100",
  34806=>"100001000",
  34807=>"111001001",
  34808=>"111101011",
  34809=>"100000111",
  34810=>"111110101",
  34811=>"111100101",
  34812=>"100100001",
  34813=>"010001101",
  34814=>"011001001",
  34815=>"110010110",
  34816=>"010100101",
  34817=>"100011010",
  34818=>"100100111",
  34819=>"111110000",
  34820=>"001111001",
  34821=>"110101000",
  34822=>"110111011",
  34823=>"010101011",
  34824=>"001110011",
  34825=>"101101110",
  34826=>"110000100",
  34827=>"110000000",
  34828=>"111010110",
  34829=>"101011010",
  34830=>"100100000",
  34831=>"111110011",
  34832=>"110101100",
  34833=>"000111111",
  34834=>"111000110",
  34835=>"001101011",
  34836=>"111001010",
  34837=>"111111110",
  34838=>"100111101",
  34839=>"001010010",
  34840=>"000000010",
  34841=>"111101101",
  34842=>"001001101",
  34843=>"111000101",
  34844=>"000000010",
  34845=>"111101001",
  34846=>"010010000",
  34847=>"011111010",
  34848=>"010111111",
  34849=>"010001100",
  34850=>"100011100",
  34851=>"110100100",
  34852=>"111101101",
  34853=>"000111000",
  34854=>"001111011",
  34855=>"010101111",
  34856=>"000010010",
  34857=>"110011111",
  34858=>"110111010",
  34859=>"000011010",
  34860=>"000101100",
  34861=>"001110000",
  34862=>"011001001",
  34863=>"010111001",
  34864=>"010100010",
  34865=>"100000100",
  34866=>"111010100",
  34867=>"011010110",
  34868=>"000000100",
  34869=>"000110001",
  34870=>"010001011",
  34871=>"111111110",
  34872=>"100010110",
  34873=>"100010101",
  34874=>"011000111",
  34875=>"100101011",
  34876=>"001111011",
  34877=>"100111001",
  34878=>"100011100",
  34879=>"001011011",
  34880=>"100011001",
  34881=>"101001101",
  34882=>"101110110",
  34883=>"101011101",
  34884=>"000001001",
  34885=>"000110111",
  34886=>"101011101",
  34887=>"101010010",
  34888=>"100100100",
  34889=>"011110000",
  34890=>"110000101",
  34891=>"101011110",
  34892=>"000000001",
  34893=>"101110001",
  34894=>"011010000",
  34895=>"101001010",
  34896=>"101101011",
  34897=>"111111111",
  34898=>"111111000",
  34899=>"010100011",
  34900=>"000000101",
  34901=>"111111111",
  34902=>"110101010",
  34903=>"100111011",
  34904=>"000010011",
  34905=>"000000110",
  34906=>"110001000",
  34907=>"111100101",
  34908=>"011110000",
  34909=>"000110110",
  34910=>"101110010",
  34911=>"111011011",
  34912=>"010000111",
  34913=>"011101111",
  34914=>"001110101",
  34915=>"100000110",
  34916=>"100111110",
  34917=>"001010111",
  34918=>"111111010",
  34919=>"101111111",
  34920=>"000001010",
  34921=>"001000100",
  34922=>"101111111",
  34923=>"000000011",
  34924=>"011010001",
  34925=>"100111110",
  34926=>"001111110",
  34927=>"111101000",
  34928=>"101111111",
  34929=>"001101101",
  34930=>"000001101",
  34931=>"101001111",
  34932=>"110110000",
  34933=>"001000011",
  34934=>"010000101",
  34935=>"000011011",
  34936=>"000100101",
  34937=>"101100100",
  34938=>"001111011",
  34939=>"000100001",
  34940=>"110010010",
  34941=>"011100011",
  34942=>"101001010",
  34943=>"101110111",
  34944=>"110001001",
  34945=>"001001011",
  34946=>"101011101",
  34947=>"001110101",
  34948=>"100111010",
  34949=>"001101001",
  34950=>"001100011",
  34951=>"010111001",
  34952=>"000001111",
  34953=>"111011010",
  34954=>"010000111",
  34955=>"001100100",
  34956=>"001111110",
  34957=>"100100010",
  34958=>"000000100",
  34959=>"101001000",
  34960=>"010000110",
  34961=>"011101100",
  34962=>"011011001",
  34963=>"111111110",
  34964=>"101000001",
  34965=>"111001110",
  34966=>"111000100",
  34967=>"001101000",
  34968=>"110000110",
  34969=>"011100111",
  34970=>"010010110",
  34971=>"111010111",
  34972=>"110001010",
  34973=>"000011011",
  34974=>"110001110",
  34975=>"000101011",
  34976=>"011000110",
  34977=>"101000001",
  34978=>"101101000",
  34979=>"101100111",
  34980=>"001111000",
  34981=>"110101110",
  34982=>"100110010",
  34983=>"011110000",
  34984=>"010001111",
  34985=>"111101101",
  34986=>"011010010",
  34987=>"100001110",
  34988=>"011011001",
  34989=>"000001111",
  34990=>"110100011",
  34991=>"001011000",
  34992=>"000011011",
  34993=>"010100101",
  34994=>"000001111",
  34995=>"110111101",
  34996=>"011010010",
  34997=>"101011110",
  34998=>"011011110",
  34999=>"000001011",
  35000=>"001111100",
  35001=>"010100011",
  35002=>"100110101",
  35003=>"000101100",
  35004=>"010001100",
  35005=>"001001011",
  35006=>"011011111",
  35007=>"000001111",
  35008=>"110111100",
  35009=>"110001101",
  35010=>"110101111",
  35011=>"101000110",
  35012=>"110111110",
  35013=>"000000110",
  35014=>"001010100",
  35015=>"010001101",
  35016=>"010001101",
  35017=>"111011101",
  35018=>"011011001",
  35019=>"110101010",
  35020=>"100100000",
  35021=>"101000000",
  35022=>"100000001",
  35023=>"000010001",
  35024=>"111110010",
  35025=>"111000111",
  35026=>"001010010",
  35027=>"111001000",
  35028=>"111001110",
  35029=>"000011011",
  35030=>"010010001",
  35031=>"110101100",
  35032=>"001000111",
  35033=>"010010101",
  35034=>"000111101",
  35035=>"111111100",
  35036=>"111001110",
  35037=>"101101101",
  35038=>"111010011",
  35039=>"000111110",
  35040=>"101000100",
  35041=>"011111010",
  35042=>"101001110",
  35043=>"000101000",
  35044=>"100000000",
  35045=>"101111100",
  35046=>"010100010",
  35047=>"000010011",
  35048=>"000100001",
  35049=>"111101101",
  35050=>"001001011",
  35051=>"011110111",
  35052=>"110110111",
  35053=>"011100001",
  35054=>"000101000",
  35055=>"110110001",
  35056=>"010110110",
  35057=>"000100011",
  35058=>"101111111",
  35059=>"101000100",
  35060=>"100110110",
  35061=>"010111110",
  35062=>"100000101",
  35063=>"000100100",
  35064=>"001110101",
  35065=>"011100100",
  35066=>"001011100",
  35067=>"001000011",
  35068=>"110011011",
  35069=>"010101010",
  35070=>"000100010",
  35071=>"110001001",
  35072=>"010100010",
  35073=>"101101010",
  35074=>"101011001",
  35075=>"100011111",
  35076=>"101011110",
  35077=>"111101000",
  35078=>"111000100",
  35079=>"000000101",
  35080=>"100110111",
  35081=>"011110100",
  35082=>"100010010",
  35083=>"011001000",
  35084=>"111110010",
  35085=>"110101000",
  35086=>"001011110",
  35087=>"100010100",
  35088=>"001100111",
  35089=>"000011010",
  35090=>"111011111",
  35091=>"110110000",
  35092=>"100100111",
  35093=>"111110011",
  35094=>"001100110",
  35095=>"001101110",
  35096=>"011101100",
  35097=>"010011101",
  35098=>"001111101",
  35099=>"001101001",
  35100=>"110011111",
  35101=>"011010011",
  35102=>"101110100",
  35103=>"000000010",
  35104=>"111101111",
  35105=>"110000000",
  35106=>"110101000",
  35107=>"100111111",
  35108=>"011000010",
  35109=>"101111010",
  35110=>"100110110",
  35111=>"000011110",
  35112=>"000111111",
  35113=>"110111100",
  35114=>"111111001",
  35115=>"100000100",
  35116=>"010100011",
  35117=>"110000111",
  35118=>"010011100",
  35119=>"010010010",
  35120=>"100010000",
  35121=>"100000010",
  35122=>"010010110",
  35123=>"101001101",
  35124=>"110010001",
  35125=>"001000111",
  35126=>"101000100",
  35127=>"101100000",
  35128=>"100001111",
  35129=>"111001100",
  35130=>"001001101",
  35131=>"001010100",
  35132=>"110101010",
  35133=>"011010100",
  35134=>"011001111",
  35135=>"101001110",
  35136=>"011101100",
  35137=>"110000100",
  35138=>"101100111",
  35139=>"000010110",
  35140=>"110110110",
  35141=>"110011010",
  35142=>"101000001",
  35143=>"001110011",
  35144=>"101111011",
  35145=>"100000110",
  35146=>"110110000",
  35147=>"010010000",
  35148=>"000100101",
  35149=>"000100111",
  35150=>"010001010",
  35151=>"110110101",
  35152=>"101100100",
  35153=>"001101000",
  35154=>"101110010",
  35155=>"111010101",
  35156=>"100100100",
  35157=>"110110110",
  35158=>"101010001",
  35159=>"111001000",
  35160=>"100011010",
  35161=>"010010110",
  35162=>"001000010",
  35163=>"001011111",
  35164=>"101001110",
  35165=>"110010111",
  35166=>"010011100",
  35167=>"101001111",
  35168=>"100101001",
  35169=>"010100001",
  35170=>"001110011",
  35171=>"011000100",
  35172=>"001101011",
  35173=>"000000000",
  35174=>"011011111",
  35175=>"100011110",
  35176=>"001101100",
  35177=>"010011101",
  35178=>"011000001",
  35179=>"001000000",
  35180=>"011010010",
  35181=>"010000101",
  35182=>"100100101",
  35183=>"101001011",
  35184=>"101110001",
  35185=>"110010100",
  35186=>"001111010",
  35187=>"011100001",
  35188=>"101011100",
  35189=>"111110011",
  35190=>"001111000",
  35191=>"111111011",
  35192=>"011101101",
  35193=>"110101110",
  35194=>"001111100",
  35195=>"110011010",
  35196=>"100010100",
  35197=>"110100111",
  35198=>"011001111",
  35199=>"000000110",
  35200=>"100100001",
  35201=>"010100110",
  35202=>"000111110",
  35203=>"001010111",
  35204=>"111001101",
  35205=>"110010111",
  35206=>"011011001",
  35207=>"110010001",
  35208=>"110111101",
  35209=>"011110000",
  35210=>"100001111",
  35211=>"011011100",
  35212=>"010000101",
  35213=>"000000111",
  35214=>"011000101",
  35215=>"011001101",
  35216=>"101100111",
  35217=>"100011010",
  35218=>"100110100",
  35219=>"011011011",
  35220=>"000000000",
  35221=>"001000110",
  35222=>"100010000",
  35223=>"101010010",
  35224=>"101111111",
  35225=>"111100010",
  35226=>"000110010",
  35227=>"110110111",
  35228=>"101000001",
  35229=>"100110100",
  35230=>"100100000",
  35231=>"010000011",
  35232=>"000011010",
  35233=>"111100110",
  35234=>"010100100",
  35235=>"110100110",
  35236=>"011000100",
  35237=>"000011100",
  35238=>"101010001",
  35239=>"110101100",
  35240=>"101010001",
  35241=>"010000110",
  35242=>"000110010",
  35243=>"101000001",
  35244=>"101001010",
  35245=>"101101001",
  35246=>"000101111",
  35247=>"001001101",
  35248=>"010100001",
  35249=>"001100110",
  35250=>"000110001",
  35251=>"110101110",
  35252=>"010110110",
  35253=>"110111111",
  35254=>"010110001",
  35255=>"100001001",
  35256=>"010101001",
  35257=>"110001010",
  35258=>"001110111",
  35259=>"101001100",
  35260=>"001100100",
  35261=>"110010000",
  35262=>"100010001",
  35263=>"110001100",
  35264=>"001100100",
  35265=>"011000111",
  35266=>"000110100",
  35267=>"011100100",
  35268=>"011110011",
  35269=>"010111111",
  35270=>"101111011",
  35271=>"000010000",
  35272=>"001000111",
  35273=>"011111011",
  35274=>"001111000",
  35275=>"111110110",
  35276=>"010011101",
  35277=>"011010110",
  35278=>"101010110",
  35279=>"010011010",
  35280=>"111100100",
  35281=>"000010110",
  35282=>"110111111",
  35283=>"101100010",
  35284=>"111111010",
  35285=>"010010010",
  35286=>"000100010",
  35287=>"100110011",
  35288=>"111100011",
  35289=>"000010110",
  35290=>"001101001",
  35291=>"010100000",
  35292=>"100111010",
  35293=>"010110011",
  35294=>"110011110",
  35295=>"100001011",
  35296=>"100011001",
  35297=>"001010010",
  35298=>"001011111",
  35299=>"101010111",
  35300=>"001100111",
  35301=>"001001011",
  35302=>"111110101",
  35303=>"111011010",
  35304=>"001001010",
  35305=>"110110110",
  35306=>"100110101",
  35307=>"001110011",
  35308=>"010110111",
  35309=>"010000000",
  35310=>"110010001",
  35311=>"011101111",
  35312=>"111100100",
  35313=>"000110101",
  35314=>"101100110",
  35315=>"110011010",
  35316=>"000110000",
  35317=>"010010111",
  35318=>"001100110",
  35319=>"111110010",
  35320=>"100110011",
  35321=>"111010100",
  35322=>"111111110",
  35323=>"010000000",
  35324=>"100101000",
  35325=>"111101010",
  35326=>"110011011",
  35327=>"111001000",
  35328=>"010001111",
  35329=>"100000001",
  35330=>"011110111",
  35331=>"100011010",
  35332=>"101100000",
  35333=>"011011010",
  35334=>"111000111",
  35335=>"000101100",
  35336=>"111111100",
  35337=>"010001010",
  35338=>"110000110",
  35339=>"011010100",
  35340=>"001100101",
  35341=>"111000011",
  35342=>"000000011",
  35343=>"111000101",
  35344=>"000011100",
  35345=>"001111011",
  35346=>"010110101",
  35347=>"011000000",
  35348=>"000000110",
  35349=>"111001101",
  35350=>"011101101",
  35351=>"100000000",
  35352=>"100101010",
  35353=>"010111110",
  35354=>"110000001",
  35355=>"010000101",
  35356=>"111100101",
  35357=>"111100101",
  35358=>"000110001",
  35359=>"100111000",
  35360=>"010011100",
  35361=>"010001101",
  35362=>"000111100",
  35363=>"101011000",
  35364=>"000000101",
  35365=>"101101001",
  35366=>"101000000",
  35367=>"110000111",
  35368=>"000110001",
  35369=>"010100011",
  35370=>"111111111",
  35371=>"000100100",
  35372=>"111010001",
  35373=>"101001010",
  35374=>"110111110",
  35375=>"010001110",
  35376=>"010111111",
  35377=>"010110100",
  35378=>"100101000",
  35379=>"001000100",
  35380=>"011101111",
  35381=>"110000000",
  35382=>"001001010",
  35383=>"100110100",
  35384=>"010011010",
  35385=>"010110001",
  35386=>"011001011",
  35387=>"100010111",
  35388=>"010000110",
  35389=>"011010100",
  35390=>"110011011",
  35391=>"000100000",
  35392=>"110010010",
  35393=>"000110101",
  35394=>"001101000",
  35395=>"110010001",
  35396=>"101110000",
  35397=>"010100011",
  35398=>"000100011",
  35399=>"100110101",
  35400=>"010111111",
  35401=>"001001000",
  35402=>"011001000",
  35403=>"010101110",
  35404=>"001010110",
  35405=>"101101100",
  35406=>"100011001",
  35407=>"111000010",
  35408=>"000110110",
  35409=>"001010100",
  35410=>"100000001",
  35411=>"100100000",
  35412=>"011100001",
  35413=>"000000110",
  35414=>"001111111",
  35415=>"011101011",
  35416=>"111111001",
  35417=>"101000101",
  35418=>"101000010",
  35419=>"100001110",
  35420=>"000011001",
  35421=>"001010100",
  35422=>"010100011",
  35423=>"111010110",
  35424=>"100100110",
  35425=>"100001001",
  35426=>"100100001",
  35427=>"111111100",
  35428=>"100111010",
  35429=>"100100011",
  35430=>"001011100",
  35431=>"101111011",
  35432=>"001001011",
  35433=>"110001111",
  35434=>"111010000",
  35435=>"111110000",
  35436=>"101101010",
  35437=>"011110110",
  35438=>"111110100",
  35439=>"100001111",
  35440=>"101010111",
  35441=>"101100001",
  35442=>"111111111",
  35443=>"011010111",
  35444=>"010111001",
  35445=>"101011001",
  35446=>"100110110",
  35447=>"110101010",
  35448=>"100111010",
  35449=>"111011110",
  35450=>"000000000",
  35451=>"001000111",
  35452=>"001100010",
  35453=>"001110010",
  35454=>"001000010",
  35455=>"010010111",
  35456=>"100011110",
  35457=>"010101001",
  35458=>"011111111",
  35459=>"111110010",
  35460=>"101001001",
  35461=>"000110100",
  35462=>"011000010",
  35463=>"011010011",
  35464=>"101100101",
  35465=>"000000000",
  35466=>"110010101",
  35467=>"001010001",
  35468=>"001000000",
  35469=>"111100000",
  35470=>"000000010",
  35471=>"011101111",
  35472=>"100011011",
  35473=>"110100001",
  35474=>"111111111",
  35475=>"101111111",
  35476=>"111001111",
  35477=>"111110010",
  35478=>"101101111",
  35479=>"100011101",
  35480=>"001000010",
  35481=>"101001111",
  35482=>"000111101",
  35483=>"110110010",
  35484=>"100010111",
  35485=>"000011000",
  35486=>"011100110",
  35487=>"111011001",
  35488=>"011100000",
  35489=>"111110010",
  35490=>"111001001",
  35491=>"111111111",
  35492=>"110111101",
  35493=>"011110011",
  35494=>"010111110",
  35495=>"000001000",
  35496=>"111111000",
  35497=>"110011111",
  35498=>"001111111",
  35499=>"110011011",
  35500=>"100111100",
  35501=>"110101001",
  35502=>"110110111",
  35503=>"111111001",
  35504=>"100010110",
  35505=>"011110111",
  35506=>"111111001",
  35507=>"000100110",
  35508=>"001000110",
  35509=>"111100001",
  35510=>"001110000",
  35511=>"001110010",
  35512=>"110101000",
  35513=>"111010011",
  35514=>"000111100",
  35515=>"111000101",
  35516=>"110110110",
  35517=>"110000101",
  35518=>"010011000",
  35519=>"110100110",
  35520=>"010000101",
  35521=>"111011100",
  35522=>"001000010",
  35523=>"110111001",
  35524=>"001101010",
  35525=>"101010100",
  35526=>"111001001",
  35527=>"101110010",
  35528=>"100011100",
  35529=>"111010010",
  35530=>"101011100",
  35531=>"101101111",
  35532=>"111111011",
  35533=>"011111011",
  35534=>"110111111",
  35535=>"111101110",
  35536=>"101011000",
  35537=>"101100100",
  35538=>"011110000",
  35539=>"101110111",
  35540=>"100000110",
  35541=>"010000001",
  35542=>"010100101",
  35543=>"111101110",
  35544=>"101001101",
  35545=>"100110000",
  35546=>"111110100",
  35547=>"111011101",
  35548=>"010111011",
  35549=>"010110101",
  35550=>"010000011",
  35551=>"100101001",
  35552=>"000100111",
  35553=>"011110000",
  35554=>"000001001",
  35555=>"001101100",
  35556=>"010111111",
  35557=>"110000101",
  35558=>"001101000",
  35559=>"000000000",
  35560=>"011001011",
  35561=>"110010001",
  35562=>"110000011",
  35563=>"100000111",
  35564=>"000000011",
  35565=>"100110110",
  35566=>"000110001",
  35567=>"001000100",
  35568=>"110101101",
  35569=>"000001111",
  35570=>"000111110",
  35571=>"101101111",
  35572=>"010111111",
  35573=>"001101000",
  35574=>"110010100",
  35575=>"110111010",
  35576=>"100001001",
  35577=>"110010011",
  35578=>"100011011",
  35579=>"101001100",
  35580=>"111110100",
  35581=>"111100000",
  35582=>"010100010",
  35583=>"011101111",
  35584=>"111010100",
  35585=>"011010001",
  35586=>"100001100",
  35587=>"111011010",
  35588=>"011110000",
  35589=>"101001100",
  35590=>"100110111",
  35591=>"010100010",
  35592=>"101100010",
  35593=>"000000110",
  35594=>"110100011",
  35595=>"000111011",
  35596=>"101101100",
  35597=>"000111101",
  35598=>"111001111",
  35599=>"011011111",
  35600=>"001111101",
  35601=>"110011011",
  35602=>"101001101",
  35603=>"110001100",
  35604=>"111001101",
  35605=>"000000111",
  35606=>"010011010",
  35607=>"110000010",
  35608=>"000100000",
  35609=>"111101111",
  35610=>"010110000",
  35611=>"110000011",
  35612=>"100010101",
  35613=>"110001100",
  35614=>"110010110",
  35615=>"110100100",
  35616=>"001110111",
  35617=>"011110000",
  35618=>"011100100",
  35619=>"001001101",
  35620=>"010100011",
  35621=>"000011011",
  35622=>"101010011",
  35623=>"111110111",
  35624=>"111111000",
  35625=>"111000011",
  35626=>"011110000",
  35627=>"101001110",
  35628=>"011011100",
  35629=>"001110011",
  35630=>"100010100",
  35631=>"100010110",
  35632=>"111110001",
  35633=>"011001111",
  35634=>"011100001",
  35635=>"101010101",
  35636=>"110000011",
  35637=>"110110010",
  35638=>"011001100",
  35639=>"001001010",
  35640=>"111111100",
  35641=>"101110000",
  35642=>"001101101",
  35643=>"011000010",
  35644=>"110001100",
  35645=>"011000010",
  35646=>"011011100",
  35647=>"001001001",
  35648=>"100011001",
  35649=>"001100001",
  35650=>"000000100",
  35651=>"111011101",
  35652=>"011000011",
  35653=>"000001011",
  35654=>"110011101",
  35655=>"001101001",
  35656=>"001011000",
  35657=>"111100100",
  35658=>"110100100",
  35659=>"001000101",
  35660=>"100001101",
  35661=>"000110010",
  35662=>"001010110",
  35663=>"100101100",
  35664=>"111100010",
  35665=>"111000101",
  35666=>"110110011",
  35667=>"010001010",
  35668=>"101011101",
  35669=>"110110111",
  35670=>"010110000",
  35671=>"001000000",
  35672=>"111100111",
  35673=>"100110011",
  35674=>"000101101",
  35675=>"010010111",
  35676=>"100001000",
  35677=>"111111110",
  35678=>"011111011",
  35679=>"000001000",
  35680=>"110011011",
  35681=>"010011110",
  35682=>"110001100",
  35683=>"111011010",
  35684=>"100000110",
  35685=>"000100001",
  35686=>"101000000",
  35687=>"110010001",
  35688=>"110100000",
  35689=>"111000010",
  35690=>"101100001",
  35691=>"001101001",
  35692=>"010101100",
  35693=>"100000100",
  35694=>"100111101",
  35695=>"100011011",
  35696=>"001011110",
  35697=>"000000100",
  35698=>"111010110",
  35699=>"101001111",
  35700=>"000111000",
  35701=>"100110101",
  35702=>"000010111",
  35703=>"011001100",
  35704=>"001110110",
  35705=>"001111011",
  35706=>"101000101",
  35707=>"011101101",
  35708=>"100101000",
  35709=>"001110001",
  35710=>"101011100",
  35711=>"110110101",
  35712=>"101111101",
  35713=>"110100101",
  35714=>"000100010",
  35715=>"111000001",
  35716=>"101111101",
  35717=>"000111111",
  35718=>"111110011",
  35719=>"011110101",
  35720=>"000000000",
  35721=>"001101001",
  35722=>"001010110",
  35723=>"101000000",
  35724=>"110100011",
  35725=>"000101100",
  35726=>"000101011",
  35727=>"000100000",
  35728=>"111011011",
  35729=>"100010101",
  35730=>"010010111",
  35731=>"011001110",
  35732=>"110111100",
  35733=>"010100000",
  35734=>"100000011",
  35735=>"010110111",
  35736=>"001010011",
  35737=>"110100011",
  35738=>"101101111",
  35739=>"100111100",
  35740=>"000101000",
  35741=>"111011001",
  35742=>"001110011",
  35743=>"101100100",
  35744=>"101110100",
  35745=>"101111111",
  35746=>"001001110",
  35747=>"010110001",
  35748=>"001110011",
  35749=>"010111101",
  35750=>"111110001",
  35751=>"000010000",
  35752=>"001000000",
  35753=>"010110110",
  35754=>"010101101",
  35755=>"000101010",
  35756=>"100001101",
  35757=>"110111011",
  35758=>"000111101",
  35759=>"110110110",
  35760=>"101000000",
  35761=>"001000100",
  35762=>"101001110",
  35763=>"010111001",
  35764=>"110001000",
  35765=>"000111101",
  35766=>"111010010",
  35767=>"010011011",
  35768=>"110100000",
  35769=>"000010110",
  35770=>"101101000",
  35771=>"100000111",
  35772=>"011000101",
  35773=>"000001001",
  35774=>"100011001",
  35775=>"100000011",
  35776=>"001000110",
  35777=>"000010001",
  35778=>"110000111",
  35779=>"100000011",
  35780=>"011001001",
  35781=>"111100011",
  35782=>"101001000",
  35783=>"110101110",
  35784=>"001010111",
  35785=>"010101001",
  35786=>"101010010",
  35787=>"001011111",
  35788=>"001111001",
  35789=>"001001000",
  35790=>"000110111",
  35791=>"110111010",
  35792=>"101101001",
  35793=>"110000000",
  35794=>"110101011",
  35795=>"011011101",
  35796=>"100100101",
  35797=>"011010000",
  35798=>"011011111",
  35799=>"011110110",
  35800=>"111110111",
  35801=>"100011001",
  35802=>"000010000",
  35803=>"000101000",
  35804=>"000000000",
  35805=>"011011100",
  35806=>"111001011",
  35807=>"010000110",
  35808=>"001110010",
  35809=>"101001101",
  35810=>"011001010",
  35811=>"101111000",
  35812=>"010011001",
  35813=>"101101100",
  35814=>"101100100",
  35815=>"111011000",
  35816=>"001101111",
  35817=>"111100110",
  35818=>"110100101",
  35819=>"011111011",
  35820=>"011110101",
  35821=>"111010110",
  35822=>"101100000",
  35823=>"001011010",
  35824=>"100010100",
  35825=>"111011100",
  35826=>"100011010",
  35827=>"100110010",
  35828=>"010100010",
  35829=>"000001100",
  35830=>"100011010",
  35831=>"111100111",
  35832=>"100000011",
  35833=>"001111111",
  35834=>"000011010",
  35835=>"100100100",
  35836=>"001010101",
  35837=>"111001111",
  35838=>"110111101",
  35839=>"000001010",
  35840=>"000000010",
  35841=>"111101100",
  35842=>"100100111",
  35843=>"011001000",
  35844=>"011100100",
  35845=>"001111000",
  35846=>"111011001",
  35847=>"010000011",
  35848=>"111111100",
  35849=>"001010000",
  35850=>"000010110",
  35851=>"100111010",
  35852=>"001110000",
  35853=>"111100011",
  35854=>"001001111",
  35855=>"000100000",
  35856=>"111101111",
  35857=>"011001100",
  35858=>"110100111",
  35859=>"101010010",
  35860=>"010010110",
  35861=>"001100111",
  35862=>"000100000",
  35863=>"011110101",
  35864=>"110001110",
  35865=>"010111000",
  35866=>"010100100",
  35867=>"110111010",
  35868=>"011001110",
  35869=>"001010101",
  35870=>"111011101",
  35871=>"000000010",
  35872=>"100010111",
  35873=>"011110011",
  35874=>"001110001",
  35875=>"100101111",
  35876=>"000101110",
  35877=>"001001011",
  35878=>"010101000",
  35879=>"111001101",
  35880=>"010101001",
  35881=>"000010100",
  35882=>"111101000",
  35883=>"111011111",
  35884=>"010000001",
  35885=>"110101100",
  35886=>"001100011",
  35887=>"001111111",
  35888=>"010011011",
  35889=>"001000100",
  35890=>"100100000",
  35891=>"101000101",
  35892=>"011111100",
  35893=>"010110101",
  35894=>"001001000",
  35895=>"011000110",
  35896=>"111010111",
  35897=>"101000000",
  35898=>"011001101",
  35899=>"111011010",
  35900=>"001110110",
  35901=>"101101001",
  35902=>"001101010",
  35903=>"111010011",
  35904=>"001111110",
  35905=>"010111000",
  35906=>"011110110",
  35907=>"100111000",
  35908=>"001011101",
  35909=>"100010101",
  35910=>"011000011",
  35911=>"100000111",
  35912=>"100000001",
  35913=>"101101000",
  35914=>"011011001",
  35915=>"101111100",
  35916=>"010100010",
  35917=>"101111001",
  35918=>"111101001",
  35919=>"011010111",
  35920=>"000111010",
  35921=>"001010111",
  35922=>"111001000",
  35923=>"000100010",
  35924=>"000110011",
  35925=>"011100011",
  35926=>"100010000",
  35927=>"110010001",
  35928=>"001011101",
  35929=>"011001010",
  35930=>"101100001",
  35931=>"001010111",
  35932=>"001010011",
  35933=>"001011101",
  35934=>"010111100",
  35935=>"001101110",
  35936=>"010000110",
  35937=>"101110110",
  35938=>"000000001",
  35939=>"101001001",
  35940=>"000011100",
  35941=>"001000100",
  35942=>"010011111",
  35943=>"111011100",
  35944=>"001111101",
  35945=>"010000000",
  35946=>"001100010",
  35947=>"100110110",
  35948=>"000010110",
  35949=>"001001000",
  35950=>"000011011",
  35951=>"100111000",
  35952=>"001111000",
  35953=>"110000000",
  35954=>"010101001",
  35955=>"101110100",
  35956=>"000000010",
  35957=>"101000001",
  35958=>"100011000",
  35959=>"010111000",
  35960=>"001001100",
  35961=>"010101011",
  35962=>"001111001",
  35963=>"101000110",
  35964=>"111101011",
  35965=>"110001011",
  35966=>"111010011",
  35967=>"011111111",
  35968=>"100111001",
  35969=>"000100010",
  35970=>"011111010",
  35971=>"000000110",
  35972=>"000001100",
  35973=>"101100110",
  35974=>"101010110",
  35975=>"110101000",
  35976=>"000001100",
  35977=>"011010001",
  35978=>"011100100",
  35979=>"101100000",
  35980=>"000000001",
  35981=>"101100001",
  35982=>"101010011",
  35983=>"011000100",
  35984=>"010110001",
  35985=>"111100011",
  35986=>"110001001",
  35987=>"000110101",
  35988=>"010011100",
  35989=>"111101101",
  35990=>"000010100",
  35991=>"100110111",
  35992=>"110111101",
  35993=>"010101110",
  35994=>"100101010",
  35995=>"111110111",
  35996=>"001000010",
  35997=>"100110000",
  35998=>"110001110",
  35999=>"010110100",
  36000=>"000101110",
  36001=>"001101101",
  36002=>"001110101",
  36003=>"001000100",
  36004=>"100001111",
  36005=>"000010111",
  36006=>"100110111",
  36007=>"110001000",
  36008=>"101010011",
  36009=>"110111110",
  36010=>"001110000",
  36011=>"001000111",
  36012=>"011110000",
  36013=>"011011100",
  36014=>"111010000",
  36015=>"011010111",
  36016=>"011011101",
  36017=>"000000101",
  36018=>"100011111",
  36019=>"101011011",
  36020=>"101100100",
  36021=>"111110100",
  36022=>"111110101",
  36023=>"001100110",
  36024=>"110000100",
  36025=>"100000111",
  36026=>"001010000",
  36027=>"100101000",
  36028=>"111111111",
  36029=>"111001011",
  36030=>"110100010",
  36031=>"111101000",
  36032=>"110010111",
  36033=>"111110010",
  36034=>"110111001",
  36035=>"001110111",
  36036=>"011000110",
  36037=>"111001000",
  36038=>"001101011",
  36039=>"110110110",
  36040=>"000000001",
  36041=>"100000101",
  36042=>"110001101",
  36043=>"111011001",
  36044=>"101000100",
  36045=>"001100100",
  36046=>"001001110",
  36047=>"101011000",
  36048=>"111010110",
  36049=>"101111011",
  36050=>"100110000",
  36051=>"110000100",
  36052=>"101001111",
  36053=>"001101001",
  36054=>"100001010",
  36055=>"101001111",
  36056=>"101001101",
  36057=>"110101110",
  36058=>"101010111",
  36059=>"110110011",
  36060=>"110110100",
  36061=>"100110111",
  36062=>"111101110",
  36063=>"111111010",
  36064=>"011101101",
  36065=>"111100010",
  36066=>"000000101",
  36067=>"101000111",
  36068=>"011100011",
  36069=>"001101100",
  36070=>"100100001",
  36071=>"110011111",
  36072=>"011001110",
  36073=>"111101111",
  36074=>"101011100",
  36075=>"000001110",
  36076=>"101010100",
  36077=>"100001111",
  36078=>"001011110",
  36079=>"110111110",
  36080=>"101000110",
  36081=>"000101110",
  36082=>"100001000",
  36083=>"110011000",
  36084=>"011100001",
  36085=>"111110010",
  36086=>"101101111",
  36087=>"000110010",
  36088=>"110010111",
  36089=>"101100010",
  36090=>"011110000",
  36091=>"011101101",
  36092=>"000011110",
  36093=>"100001111",
  36094=>"011001010",
  36095=>"010110010",
  36096=>"010010111",
  36097=>"010110100",
  36098=>"111101011",
  36099=>"100000011",
  36100=>"001100100",
  36101=>"011110000",
  36102=>"000110000",
  36103=>"001001100",
  36104=>"000000111",
  36105=>"101000010",
  36106=>"010000011",
  36107=>"101000010",
  36108=>"110010111",
  36109=>"110110000",
  36110=>"101100011",
  36111=>"000110011",
  36112=>"000110010",
  36113=>"000111100",
  36114=>"110100000",
  36115=>"101011110",
  36116=>"010000101",
  36117=>"010011000",
  36118=>"011101010",
  36119=>"111010011",
  36120=>"111111110",
  36121=>"011000000",
  36122=>"110011010",
  36123=>"100011000",
  36124=>"101111000",
  36125=>"111000001",
  36126=>"100011000",
  36127=>"001111111",
  36128=>"101111110",
  36129=>"100001101",
  36130=>"011010010",
  36131=>"001111011",
  36132=>"001010110",
  36133=>"000101011",
  36134=>"101001011",
  36135=>"000010110",
  36136=>"110111011",
  36137=>"011101110",
  36138=>"011100001",
  36139=>"010010000",
  36140=>"011110010",
  36141=>"000001001",
  36142=>"100000101",
  36143=>"011010110",
  36144=>"100000010",
  36145=>"011001000",
  36146=>"000011110",
  36147=>"001000010",
  36148=>"100011100",
  36149=>"001010100",
  36150=>"111111100",
  36151=>"110001010",
  36152=>"000101111",
  36153=>"101110110",
  36154=>"010010110",
  36155=>"001000100",
  36156=>"000101101",
  36157=>"101010000",
  36158=>"110010101",
  36159=>"111010111",
  36160=>"001000101",
  36161=>"010001001",
  36162=>"001001101",
  36163=>"100001011",
  36164=>"101101111",
  36165=>"111101001",
  36166=>"110010000",
  36167=>"011100111",
  36168=>"000101101",
  36169=>"010001110",
  36170=>"000011010",
  36171=>"001110010",
  36172=>"011101110",
  36173=>"100011000",
  36174=>"100101000",
  36175=>"100001100",
  36176=>"101110001",
  36177=>"111010010",
  36178=>"111111111",
  36179=>"100100010",
  36180=>"100011011",
  36181=>"000100110",
  36182=>"110101001",
  36183=>"101001001",
  36184=>"011111000",
  36185=>"011101010",
  36186=>"000101111",
  36187=>"110001001",
  36188=>"000111111",
  36189=>"011010010",
  36190=>"011101011",
  36191=>"010101010",
  36192=>"011001101",
  36193=>"100001100",
  36194=>"101101100",
  36195=>"011011111",
  36196=>"101100000",
  36197=>"101011100",
  36198=>"100101110",
  36199=>"011010110",
  36200=>"111011111",
  36201=>"111110000",
  36202=>"100011110",
  36203=>"010010101",
  36204=>"001110110",
  36205=>"101000001",
  36206=>"101000001",
  36207=>"101110001",
  36208=>"111111111",
  36209=>"100000111",
  36210=>"010111101",
  36211=>"000100101",
  36212=>"001100110",
  36213=>"011011010",
  36214=>"100101100",
  36215=>"100111110",
  36216=>"001110111",
  36217=>"010110001",
  36218=>"000000010",
  36219=>"101010110",
  36220=>"001111010",
  36221=>"111010010",
  36222=>"000100100",
  36223=>"111010110",
  36224=>"101011010",
  36225=>"010000000",
  36226=>"111110110",
  36227=>"010000110",
  36228=>"000011100",
  36229=>"000101010",
  36230=>"110011000",
  36231=>"110111101",
  36232=>"101011001",
  36233=>"011100010",
  36234=>"011000101",
  36235=>"010010011",
  36236=>"100101100",
  36237=>"111011111",
  36238=>"100110111",
  36239=>"111101110",
  36240=>"111111110",
  36241=>"000101100",
  36242=>"110010000",
  36243=>"100010011",
  36244=>"111000000",
  36245=>"001001010",
  36246=>"110010010",
  36247=>"000001100",
  36248=>"010111000",
  36249=>"001000100",
  36250=>"101010010",
  36251=>"110010110",
  36252=>"000101011",
  36253=>"100101111",
  36254=>"110100110",
  36255=>"001001010",
  36256=>"101110100",
  36257=>"011000111",
  36258=>"111011110",
  36259=>"100110111",
  36260=>"100011011",
  36261=>"111100100",
  36262=>"000110110",
  36263=>"011010000",
  36264=>"100111111",
  36265=>"000111101",
  36266=>"000101100",
  36267=>"100000001",
  36268=>"110110101",
  36269=>"110011110",
  36270=>"001100001",
  36271=>"001101111",
  36272=>"010000101",
  36273=>"000010001",
  36274=>"010101111",
  36275=>"111100100",
  36276=>"010000001",
  36277=>"010010110",
  36278=>"111101001",
  36279=>"010100010",
  36280=>"101001110",
  36281=>"101110100",
  36282=>"101011110",
  36283=>"001010101",
  36284=>"111010100",
  36285=>"011101111",
  36286=>"010011000",
  36287=>"010100101",
  36288=>"101011000",
  36289=>"010101011",
  36290=>"111110010",
  36291=>"101000001",
  36292=>"010001100",
  36293=>"100010110",
  36294=>"101010000",
  36295=>"000011001",
  36296=>"011000111",
  36297=>"101000010",
  36298=>"000011010",
  36299=>"101100111",
  36300=>"100100000",
  36301=>"110110001",
  36302=>"100001100",
  36303=>"010101010",
  36304=>"001110011",
  36305=>"010011100",
  36306=>"110100000",
  36307=>"001011101",
  36308=>"000011010",
  36309=>"011011101",
  36310=>"100010011",
  36311=>"010101001",
  36312=>"100000011",
  36313=>"100010110",
  36314=>"000001010",
  36315=>"010110000",
  36316=>"111111100",
  36317=>"010000000",
  36318=>"000010010",
  36319=>"011011100",
  36320=>"110000000",
  36321=>"010111001",
  36322=>"110111111",
  36323=>"101111011",
  36324=>"000001101",
  36325=>"100111100",
  36326=>"001000101",
  36327=>"111011100",
  36328=>"011101010",
  36329=>"101011111",
  36330=>"010000100",
  36331=>"111000111",
  36332=>"110111110",
  36333=>"010011100",
  36334=>"110110010",
  36335=>"010000001",
  36336=>"111001001",
  36337=>"111011111",
  36338=>"110010110",
  36339=>"110010010",
  36340=>"111111011",
  36341=>"111111111",
  36342=>"100000111",
  36343=>"111011100",
  36344=>"110011101",
  36345=>"111010110",
  36346=>"101000100",
  36347=>"111110111",
  36348=>"011011100",
  36349=>"110101111",
  36350=>"110101011",
  36351=>"000000001",
  36352=>"100011110",
  36353=>"000000000",
  36354=>"100110101",
  36355=>"100110100",
  36356=>"110010011",
  36357=>"011100100",
  36358=>"000100110",
  36359=>"010111111",
  36360=>"001110100",
  36361=>"010001111",
  36362=>"011011100",
  36363=>"010000010",
  36364=>"010010000",
  36365=>"010101101",
  36366=>"001111011",
  36367=>"101101100",
  36368=>"011110110",
  36369=>"011111110",
  36370=>"111100010",
  36371=>"011011101",
  36372=>"011110010",
  36373=>"010011000",
  36374=>"011110100",
  36375=>"100101111",
  36376=>"101001010",
  36377=>"011001101",
  36378=>"001011111",
  36379=>"101101001",
  36380=>"111010110",
  36381=>"010110100",
  36382=>"110101011",
  36383=>"001000010",
  36384=>"101010110",
  36385=>"110001011",
  36386=>"100000000",
  36387=>"110101110",
  36388=>"011000001",
  36389=>"010011101",
  36390=>"110011000",
  36391=>"000100110",
  36392=>"001101011",
  36393=>"100111000",
  36394=>"111010111",
  36395=>"100001000",
  36396=>"110111000",
  36397=>"001100011",
  36398=>"011010001",
  36399=>"010111100",
  36400=>"011110011",
  36401=>"001010011",
  36402=>"000001100",
  36403=>"001100100",
  36404=>"101001110",
  36405=>"010100100",
  36406=>"100001100",
  36407=>"110111100",
  36408=>"001101111",
  36409=>"000000001",
  36410=>"111101000",
  36411=>"110000010",
  36412=>"110101111",
  36413=>"010100100",
  36414=>"111111011",
  36415=>"010110100",
  36416=>"000000101",
  36417=>"101010111",
  36418=>"010100011",
  36419=>"010000111",
  36420=>"000000000",
  36421=>"101010111",
  36422=>"010010010",
  36423=>"110011011",
  36424=>"000011001",
  36425=>"101000100",
  36426=>"101010001",
  36427=>"101111001",
  36428=>"101101010",
  36429=>"100101001",
  36430=>"100110000",
  36431=>"010111100",
  36432=>"101100010",
  36433=>"000001011",
  36434=>"100111010",
  36435=>"100011111",
  36436=>"000001001",
  36437=>"011100101",
  36438=>"000000000",
  36439=>"101100110",
  36440=>"001001011",
  36441=>"111010110",
  36442=>"110000101",
  36443=>"110000001",
  36444=>"100001001",
  36445=>"010110010",
  36446=>"101101111",
  36447=>"000111011",
  36448=>"000011111",
  36449=>"010001010",
  36450=>"110110110",
  36451=>"010011011",
  36452=>"100001010",
  36453=>"010011001",
  36454=>"100100000",
  36455=>"000001111",
  36456=>"011100100",
  36457=>"111111001",
  36458=>"010111111",
  36459=>"000000100",
  36460=>"001011010",
  36461=>"111101010",
  36462=>"101111000",
  36463=>"101001000",
  36464=>"100000111",
  36465=>"111010000",
  36466=>"111001110",
  36467=>"110001001",
  36468=>"101011100",
  36469=>"100000100",
  36470=>"001010111",
  36471=>"000110010",
  36472=>"101101011",
  36473=>"000100010",
  36474=>"100000101",
  36475=>"000101010",
  36476=>"101101010",
  36477=>"000001010",
  36478=>"000011101",
  36479=>"111111100",
  36480=>"110111001",
  36481=>"100111010",
  36482=>"001000001",
  36483=>"111101001",
  36484=>"101111010",
  36485=>"100001111",
  36486=>"111001001",
  36487=>"100000110",
  36488=>"111001010",
  36489=>"011001010",
  36490=>"100110100",
  36491=>"010011011",
  36492=>"101011010",
  36493=>"100100010",
  36494=>"010110101",
  36495=>"101011101",
  36496=>"111001001",
  36497=>"010010101",
  36498=>"101101111",
  36499=>"000001100",
  36500=>"011100010",
  36501=>"011010010",
  36502=>"001010010",
  36503=>"001100001",
  36504=>"101110111",
  36505=>"100000101",
  36506=>"011001010",
  36507=>"101011100",
  36508=>"000110011",
  36509=>"011011100",
  36510=>"001000101",
  36511=>"000100100",
  36512=>"000110110",
  36513=>"010001001",
  36514=>"110000101",
  36515=>"111100111",
  36516=>"001010001",
  36517=>"011001011",
  36518=>"101011000",
  36519=>"000101110",
  36520=>"011100100",
  36521=>"011000001",
  36522=>"011000110",
  36523=>"001111011",
  36524=>"010101000",
  36525=>"111000010",
  36526=>"000111000",
  36527=>"000011100",
  36528=>"001011001",
  36529=>"101010100",
  36530=>"010111010",
  36531=>"000010100",
  36532=>"001000001",
  36533=>"100100101",
  36534=>"001000001",
  36535=>"110011001",
  36536=>"000010000",
  36537=>"100001010",
  36538=>"101000010",
  36539=>"100010001",
  36540=>"010110011",
  36541=>"001001011",
  36542=>"100111101",
  36543=>"101110001",
  36544=>"011011101",
  36545=>"000010000",
  36546=>"000111110",
  36547=>"011001100",
  36548=>"010100100",
  36549=>"111011011",
  36550=>"101010011",
  36551=>"111011011",
  36552=>"100011011",
  36553=>"001100101",
  36554=>"110111011",
  36555=>"010111000",
  36556=>"000101101",
  36557=>"010010101",
  36558=>"010110011",
  36559=>"100000001",
  36560=>"100100000",
  36561=>"011001110",
  36562=>"110110110",
  36563=>"001000010",
  36564=>"110101110",
  36565=>"001001111",
  36566=>"010111011",
  36567=>"001011101",
  36568=>"010011100",
  36569=>"001000100",
  36570=>"010010101",
  36571=>"110100111",
  36572=>"101111110",
  36573=>"000110110",
  36574=>"010100010",
  36575=>"010010100",
  36576=>"001100001",
  36577=>"010110111",
  36578=>"100010011",
  36579=>"111100110",
  36580=>"101110001",
  36581=>"000101010",
  36582=>"010101100",
  36583=>"110011000",
  36584=>"111000010",
  36585=>"001001001",
  36586=>"001001010",
  36587=>"111000101",
  36588=>"110010101",
  36589=>"000010111",
  36590=>"100110100",
  36591=>"011011101",
  36592=>"001000101",
  36593=>"011001011",
  36594=>"001101000",
  36595=>"010001011",
  36596=>"010001100",
  36597=>"111010010",
  36598=>"100000111",
  36599=>"011000100",
  36600=>"110101111",
  36601=>"010001011",
  36602=>"000100011",
  36603=>"001011001",
  36604=>"010110011",
  36605=>"000000001",
  36606=>"101001000",
  36607=>"110010001",
  36608=>"011101100",
  36609=>"010010110",
  36610=>"011111000",
  36611=>"000011101",
  36612=>"110101100",
  36613=>"010001010",
  36614=>"111011010",
  36615=>"010110000",
  36616=>"100000010",
  36617=>"001110000",
  36618=>"011111110",
  36619=>"011011110",
  36620=>"110110000",
  36621=>"011110101",
  36622=>"001101000",
  36623=>"111111100",
  36624=>"001000110",
  36625=>"000000101",
  36626=>"000111100",
  36627=>"011110101",
  36628=>"101001000",
  36629=>"101010010",
  36630=>"001110111",
  36631=>"010110000",
  36632=>"011110000",
  36633=>"101110010",
  36634=>"100011000",
  36635=>"101010110",
  36636=>"100101110",
  36637=>"100011000",
  36638=>"110000100",
  36639=>"000001001",
  36640=>"111010011",
  36641=>"100001100",
  36642=>"110011111",
  36643=>"001011001",
  36644=>"000001001",
  36645=>"111001110",
  36646=>"000010100",
  36647=>"111010011",
  36648=>"010110001",
  36649=>"101010010",
  36650=>"111010111",
  36651=>"101000110",
  36652=>"100101101",
  36653=>"011011010",
  36654=>"000110011",
  36655=>"100001100",
  36656=>"011000000",
  36657=>"111011111",
  36658=>"100100010",
  36659=>"010000110",
  36660=>"011111000",
  36661=>"010111001",
  36662=>"110110011",
  36663=>"111001001",
  36664=>"000010100",
  36665=>"000010111",
  36666=>"101101010",
  36667=>"110011110",
  36668=>"001011111",
  36669=>"100000010",
  36670=>"111111111",
  36671=>"010110101",
  36672=>"011010000",
  36673=>"001101111",
  36674=>"000111001",
  36675=>"011001000",
  36676=>"001110101",
  36677=>"110001000",
  36678=>"011110100",
  36679=>"010101000",
  36680=>"111111111",
  36681=>"011100110",
  36682=>"000010100",
  36683=>"000100111",
  36684=>"000010000",
  36685=>"010011100",
  36686=>"100111010",
  36687=>"000111010",
  36688=>"010101111",
  36689=>"000000111",
  36690=>"010101110",
  36691=>"010100110",
  36692=>"110111101",
  36693=>"010110001",
  36694=>"001110101",
  36695=>"010101011",
  36696=>"111011110",
  36697=>"000101011",
  36698=>"111101010",
  36699=>"010111111",
  36700=>"010110011",
  36701=>"001111111",
  36702=>"011111111",
  36703=>"000001011",
  36704=>"100000010",
  36705=>"101010000",
  36706=>"111101000",
  36707=>"011111010",
  36708=>"001110000",
  36709=>"001011110",
  36710=>"001001010",
  36711=>"110100101",
  36712=>"010010010",
  36713=>"110100010",
  36714=>"100110000",
  36715=>"100100111",
  36716=>"010000010",
  36717=>"000010010",
  36718=>"001111010",
  36719=>"001101011",
  36720=>"001111111",
  36721=>"000000000",
  36722=>"000111101",
  36723=>"011001110",
  36724=>"100010100",
  36725=>"001110111",
  36726=>"100111011",
  36727=>"111001010",
  36728=>"100111001",
  36729=>"011110111",
  36730=>"110111101",
  36731=>"111010001",
  36732=>"000001001",
  36733=>"010100011",
  36734=>"110111111",
  36735=>"011111011",
  36736=>"100101100",
  36737=>"010011010",
  36738=>"001100000",
  36739=>"000100011",
  36740=>"100001010",
  36741=>"110110011",
  36742=>"011101111",
  36743=>"001100000",
  36744=>"101001101",
  36745=>"010111110",
  36746=>"011000000",
  36747=>"000001000",
  36748=>"110001011",
  36749=>"000010000",
  36750=>"110101011",
  36751=>"110010000",
  36752=>"010011000",
  36753=>"011100110",
  36754=>"010010001",
  36755=>"110111111",
  36756=>"011101111",
  36757=>"011001101",
  36758=>"011000001",
  36759=>"000110100",
  36760=>"100000010",
  36761=>"001110000",
  36762=>"010000001",
  36763=>"110000110",
  36764=>"101101011",
  36765=>"100011000",
  36766=>"110011000",
  36767=>"010100001",
  36768=>"001010000",
  36769=>"010000001",
  36770=>"011101011",
  36771=>"000000111",
  36772=>"111010000",
  36773=>"011100110",
  36774=>"111101010",
  36775=>"100010010",
  36776=>"010011101",
  36777=>"001000011",
  36778=>"100001101",
  36779=>"110111101",
  36780=>"100100001",
  36781=>"001001011",
  36782=>"000101111",
  36783=>"110110010",
  36784=>"111000100",
  36785=>"000011010",
  36786=>"111001001",
  36787=>"000110100",
  36788=>"110011101",
  36789=>"110101010",
  36790=>"010101101",
  36791=>"001011100",
  36792=>"011000001",
  36793=>"010000001",
  36794=>"001101101",
  36795=>"011001011",
  36796=>"000001000",
  36797=>"110000000",
  36798=>"011111100",
  36799=>"001111100",
  36800=>"100100011",
  36801=>"011000010",
  36802=>"010101011",
  36803=>"011000100",
  36804=>"000011101",
  36805=>"011001111",
  36806=>"010100100",
  36807=>"101010001",
  36808=>"000100010",
  36809=>"000110010",
  36810=>"010101010",
  36811=>"010000011",
  36812=>"011110011",
  36813=>"111000011",
  36814=>"101110010",
  36815=>"110100011",
  36816=>"011001001",
  36817=>"101101010",
  36818=>"110100000",
  36819=>"001011001",
  36820=>"100101011",
  36821=>"011100100",
  36822=>"111101101",
  36823=>"011000110",
  36824=>"100001000",
  36825=>"001110010",
  36826=>"010101110",
  36827=>"111000010",
  36828=>"001001000",
  36829=>"000010011",
  36830=>"110111110",
  36831=>"111000100",
  36832=>"111100100",
  36833=>"100001000",
  36834=>"000000000",
  36835=>"000111111",
  36836=>"000100100",
  36837=>"111110000",
  36838=>"010000000",
  36839=>"011000000",
  36840=>"000011010",
  36841=>"011110010",
  36842=>"000001010",
  36843=>"010011110",
  36844=>"111101110",
  36845=>"110000011",
  36846=>"000100100",
  36847=>"011101101",
  36848=>"011101101",
  36849=>"011100111",
  36850=>"011010111",
  36851=>"101101000",
  36852=>"111110111",
  36853=>"100001001",
  36854=>"100001001",
  36855=>"111011111",
  36856=>"111110111",
  36857=>"010000110",
  36858=>"000000000",
  36859=>"111111001",
  36860=>"011001111",
  36861=>"000110110",
  36862=>"111110100",
  36863=>"100000011",
  36864=>"100001000",
  36865=>"100011110",
  36866=>"011011111",
  36867=>"111110101",
  36868=>"100010010",
  36869=>"110101110",
  36870=>"100010001",
  36871=>"111011011",
  36872=>"110110000",
  36873=>"111001111",
  36874=>"111101010",
  36875=>"001111010",
  36876=>"010010001",
  36877=>"000110101",
  36878=>"110010010",
  36879=>"110010001",
  36880=>"100010110",
  36881=>"001101001",
  36882=>"110001001",
  36883=>"011010111",
  36884=>"110011111",
  36885=>"010100101",
  36886=>"110000011",
  36887=>"100000101",
  36888=>"000000000",
  36889=>"101111101",
  36890=>"111001011",
  36891=>"010000111",
  36892=>"111101111",
  36893=>"010000101",
  36894=>"000000000",
  36895=>"111011000",
  36896=>"000101010",
  36897=>"000011001",
  36898=>"110000011",
  36899=>"110010011",
  36900=>"000110000",
  36901=>"110111111",
  36902=>"000100000",
  36903=>"011111100",
  36904=>"001001010",
  36905=>"110101001",
  36906=>"000111001",
  36907=>"000011000",
  36908=>"100000100",
  36909=>"000001010",
  36910=>"000101011",
  36911=>"110111110",
  36912=>"110011001",
  36913=>"001011101",
  36914=>"111001100",
  36915=>"110111011",
  36916=>"101100001",
  36917=>"101100101",
  36918=>"011001100",
  36919=>"100101011",
  36920=>"110110010",
  36921=>"000110000",
  36922=>"110011101",
  36923=>"100100010",
  36924=>"010000101",
  36925=>"101001110",
  36926=>"000001111",
  36927=>"001111101",
  36928=>"001000001",
  36929=>"100010001",
  36930=>"011001111",
  36931=>"010010000",
  36932=>"000001100",
  36933=>"000100010",
  36934=>"000110100",
  36935=>"100010100",
  36936=>"010011110",
  36937=>"110011111",
  36938=>"100101101",
  36939=>"111011100",
  36940=>"010111111",
  36941=>"000111011",
  36942=>"100100110",
  36943=>"001011110",
  36944=>"100010100",
  36945=>"010000010",
  36946=>"100100010",
  36947=>"101111101",
  36948=>"010101101",
  36949=>"110000101",
  36950=>"011001111",
  36951=>"111101110",
  36952=>"001100010",
  36953=>"111111010",
  36954=>"000101111",
  36955=>"101101000",
  36956=>"111110000",
  36957=>"001011111",
  36958=>"111101010",
  36959=>"001000001",
  36960=>"001110100",
  36961=>"011111001",
  36962=>"111100110",
  36963=>"110011000",
  36964=>"111101000",
  36965=>"010001010",
  36966=>"001110101",
  36967=>"000100100",
  36968=>"000000110",
  36969=>"010001100",
  36970=>"111010100",
  36971=>"010101001",
  36972=>"101011110",
  36973=>"010101110",
  36974=>"101110010",
  36975=>"101110001",
  36976=>"011001001",
  36977=>"010111110",
  36978=>"101001001",
  36979=>"010111110",
  36980=>"100100111",
  36981=>"010010011",
  36982=>"001101100",
  36983=>"110010110",
  36984=>"110111101",
  36985=>"100110001",
  36986=>"100001101",
  36987=>"110011001",
  36988=>"000101110",
  36989=>"001101110",
  36990=>"100010101",
  36991=>"101000001",
  36992=>"110101100",
  36993=>"001011101",
  36994=>"001111100",
  36995=>"100100011",
  36996=>"011001011",
  36997=>"110111001",
  36998=>"011110101",
  36999=>"010110100",
  37000=>"001000001",
  37001=>"110000110",
  37002=>"010100001",
  37003=>"011001001",
  37004=>"100110010",
  37005=>"010010010",
  37006=>"010010100",
  37007=>"101111111",
  37008=>"010100010",
  37009=>"011110110",
  37010=>"110010111",
  37011=>"010111011",
  37012=>"110101011",
  37013=>"100100001",
  37014=>"100000000",
  37015=>"011001001",
  37016=>"110011111",
  37017=>"110100101",
  37018=>"110111010",
  37019=>"001110011",
  37020=>"100110001",
  37021=>"110011001",
  37022=>"010001010",
  37023=>"001011000",
  37024=>"111100100",
  37025=>"110000110",
  37026=>"010101000",
  37027=>"001100001",
  37028=>"010111000",
  37029=>"111101011",
  37030=>"001111000",
  37031=>"100010001",
  37032=>"011001001",
  37033=>"101000101",
  37034=>"010011011",
  37035=>"000010101",
  37036=>"101111011",
  37037=>"111011001",
  37038=>"010101000",
  37039=>"000011101",
  37040=>"111100011",
  37041=>"010111111",
  37042=>"010100000",
  37043=>"001101001",
  37044=>"111101110",
  37045=>"110100111",
  37046=>"001001001",
  37047=>"110100010",
  37048=>"100111100",
  37049=>"110111000",
  37050=>"000001110",
  37051=>"001101100",
  37052=>"100100001",
  37053=>"110101011",
  37054=>"100001010",
  37055=>"111110100",
  37056=>"100001010",
  37057=>"111010110",
  37058=>"100110111",
  37059=>"100010000",
  37060=>"010010101",
  37061=>"001100001",
  37062=>"111011111",
  37063=>"111011101",
  37064=>"101000010",
  37065=>"010000111",
  37066=>"110010000",
  37067=>"010101111",
  37068=>"000100011",
  37069=>"010100010",
  37070=>"000110110",
  37071=>"010010101",
  37072=>"000001001",
  37073=>"011111100",
  37074=>"001010000",
  37075=>"101001001",
  37076=>"110111011",
  37077=>"001001010",
  37078=>"101101001",
  37079=>"110101011",
  37080=>"100001011",
  37081=>"011101001",
  37082=>"010001001",
  37083=>"001111001",
  37084=>"000101100",
  37085=>"111110110",
  37086=>"010010111",
  37087=>"100000111",
  37088=>"111110001",
  37089=>"000000010",
  37090=>"100100111",
  37091=>"010111110",
  37092=>"101101011",
  37093=>"001100110",
  37094=>"001100000",
  37095=>"110110001",
  37096=>"100111011",
  37097=>"010010011",
  37098=>"110011001",
  37099=>"011100011",
  37100=>"110011001",
  37101=>"011100001",
  37102=>"011111110",
  37103=>"110100110",
  37104=>"110110010",
  37105=>"111101110",
  37106=>"101000001",
  37107=>"111111111",
  37108=>"100010000",
  37109=>"000101111",
  37110=>"111001011",
  37111=>"011001110",
  37112=>"001110000",
  37113=>"111111100",
  37114=>"001110101",
  37115=>"101001100",
  37116=>"011111110",
  37117=>"001000001",
  37118=>"000000000",
  37119=>"111011011",
  37120=>"110001101",
  37121=>"000010001",
  37122=>"001000010",
  37123=>"111101111",
  37124=>"000011110",
  37125=>"111110101",
  37126=>"100101110",
  37127=>"011101011",
  37128=>"100001011",
  37129=>"001000000",
  37130=>"010011110",
  37131=>"111001011",
  37132=>"011110100",
  37133=>"111000110",
  37134=>"101100001",
  37135=>"010100011",
  37136=>"100000110",
  37137=>"000010010",
  37138=>"000000110",
  37139=>"110111001",
  37140=>"001100110",
  37141=>"011111011",
  37142=>"011010010",
  37143=>"110000001",
  37144=>"100100101",
  37145=>"001000101",
  37146=>"110110100",
  37147=>"010100010",
  37148=>"000010111",
  37149=>"010011111",
  37150=>"111110011",
  37151=>"000001010",
  37152=>"110110110",
  37153=>"101101101",
  37154=>"100100010",
  37155=>"001111001",
  37156=>"010001000",
  37157=>"110111101",
  37158=>"000000010",
  37159=>"110010101",
  37160=>"101101111",
  37161=>"111000000",
  37162=>"010000110",
  37163=>"101011010",
  37164=>"001100101",
  37165=>"001000101",
  37166=>"010101011",
  37167=>"000001000",
  37168=>"010010000",
  37169=>"101111000",
  37170=>"001001101",
  37171=>"111101111",
  37172=>"001110111",
  37173=>"000010011",
  37174=>"100110000",
  37175=>"000110111",
  37176=>"000111000",
  37177=>"100000110",
  37178=>"110001001",
  37179=>"011001101",
  37180=>"100010001",
  37181=>"111110010",
  37182=>"010100000",
  37183=>"010110111",
  37184=>"011101000",
  37185=>"001101101",
  37186=>"101111110",
  37187=>"110100110",
  37188=>"000111000",
  37189=>"110010001",
  37190=>"001000100",
  37191=>"110010100",
  37192=>"110110111",
  37193=>"100001011",
  37194=>"001100010",
  37195=>"101010011",
  37196=>"001011000",
  37197=>"101110010",
  37198=>"011100100",
  37199=>"101110111",
  37200=>"100111111",
  37201=>"100110111",
  37202=>"101101100",
  37203=>"111011111",
  37204=>"010011110",
  37205=>"110101100",
  37206=>"110101110",
  37207=>"110111101",
  37208=>"010111000",
  37209=>"100000001",
  37210=>"010001110",
  37211=>"011110011",
  37212=>"111011111",
  37213=>"101111010",
  37214=>"001011000",
  37215=>"000001001",
  37216=>"100000011",
  37217=>"111100111",
  37218=>"011100100",
  37219=>"111100111",
  37220=>"010000100",
  37221=>"111000000",
  37222=>"111011111",
  37223=>"010000101",
  37224=>"100100110",
  37225=>"100110111",
  37226=>"111110100",
  37227=>"111011001",
  37228=>"001101110",
  37229=>"010111101",
  37230=>"100101101",
  37231=>"010010110",
  37232=>"001111111",
  37233=>"010010011",
  37234=>"001111111",
  37235=>"000000010",
  37236=>"011011000",
  37237=>"101000011",
  37238=>"110011000",
  37239=>"100010110",
  37240=>"001111101",
  37241=>"100100101",
  37242=>"010110101",
  37243=>"001111011",
  37244=>"001100000",
  37245=>"011111111",
  37246=>"100110010",
  37247=>"101000001",
  37248=>"111111111",
  37249=>"000101011",
  37250=>"101001111",
  37251=>"010010001",
  37252=>"100011101",
  37253=>"001000110",
  37254=>"101110110",
  37255=>"011011000",
  37256=>"011101010",
  37257=>"111100101",
  37258=>"011011010",
  37259=>"111111100",
  37260=>"111100001",
  37261=>"111111011",
  37262=>"110001000",
  37263=>"000011100",
  37264=>"000001111",
  37265=>"011011111",
  37266=>"010110101",
  37267=>"101000010",
  37268=>"101011000",
  37269=>"011011011",
  37270=>"001000100",
  37271=>"010000000",
  37272=>"011110110",
  37273=>"001011010",
  37274=>"001110111",
  37275=>"000000011",
  37276=>"011011110",
  37277=>"110001110",
  37278=>"110011100",
  37279=>"000101001",
  37280=>"010000000",
  37281=>"001011000",
  37282=>"000000001",
  37283=>"110100011",
  37284=>"011010000",
  37285=>"110111011",
  37286=>"001010111",
  37287=>"110010000",
  37288=>"010000101",
  37289=>"001110101",
  37290=>"000010000",
  37291=>"110100011",
  37292=>"001010110",
  37293=>"100110010",
  37294=>"101100011",
  37295=>"000100000",
  37296=>"100101000",
  37297=>"011001010",
  37298=>"100010000",
  37299=>"111110100",
  37300=>"010011110",
  37301=>"010110101",
  37302=>"110110010",
  37303=>"111100000",
  37304=>"011001110",
  37305=>"111100000",
  37306=>"101011010",
  37307=>"100110100",
  37308=>"010111111",
  37309=>"111000011",
  37310=>"111101011",
  37311=>"001100000",
  37312=>"011100011",
  37313=>"011011111",
  37314=>"110001110",
  37315=>"010000011",
  37316=>"111010010",
  37317=>"111010111",
  37318=>"111101010",
  37319=>"010001010",
  37320=>"101111100",
  37321=>"001111011",
  37322=>"111000111",
  37323=>"011111111",
  37324=>"001010101",
  37325=>"101000100",
  37326=>"011101010",
  37327=>"000100101",
  37328=>"001000110",
  37329=>"111011011",
  37330=>"100001000",
  37331=>"001000100",
  37332=>"000101011",
  37333=>"111001111",
  37334=>"111100101",
  37335=>"000001011",
  37336=>"011010111",
  37337=>"100000010",
  37338=>"110000100",
  37339=>"011001100",
  37340=>"000111011",
  37341=>"001001110",
  37342=>"010000010",
  37343=>"011111001",
  37344=>"101111010",
  37345=>"000010101",
  37346=>"000011001",
  37347=>"110001000",
  37348=>"111010000",
  37349=>"100011000",
  37350=>"001011011",
  37351=>"100111001",
  37352=>"110101000",
  37353=>"011101100",
  37354=>"010010010",
  37355=>"001010111",
  37356=>"100001100",
  37357=>"110101101",
  37358=>"110011001",
  37359=>"101001000",
  37360=>"011000110",
  37361=>"111111011",
  37362=>"101111010",
  37363=>"100100110",
  37364=>"010001000",
  37365=>"111011101",
  37366=>"100100110",
  37367=>"101001011",
  37368=>"100111100",
  37369=>"011111100",
  37370=>"001110111",
  37371=>"001011001",
  37372=>"001101000",
  37373=>"001101010",
  37374=>"000001100",
  37375=>"111111011",
  37376=>"110000101",
  37377=>"010000010",
  37378=>"001011001",
  37379=>"000100010",
  37380=>"101011010",
  37381=>"011100110",
  37382=>"010011001",
  37383=>"010001111",
  37384=>"110011000",
  37385=>"001000000",
  37386=>"011111001",
  37387=>"100000101",
  37388=>"100111010",
  37389=>"101000000",
  37390=>"100100110",
  37391=>"100101010",
  37392=>"000010001",
  37393=>"001110011",
  37394=>"110111001",
  37395=>"100011001",
  37396=>"101110101",
  37397=>"101010101",
  37398=>"110100010",
  37399=>"101101011",
  37400=>"100101010",
  37401=>"110101110",
  37402=>"100100000",
  37403=>"011110100",
  37404=>"000101100",
  37405=>"000100101",
  37406=>"100110101",
  37407=>"100000101",
  37408=>"110001010",
  37409=>"101100100",
  37410=>"001001010",
  37411=>"100010010",
  37412=>"100101010",
  37413=>"111011111",
  37414=>"100010110",
  37415=>"110010011",
  37416=>"110000000",
  37417=>"001101101",
  37418=>"000100101",
  37419=>"100001100",
  37420=>"111110100",
  37421=>"100011001",
  37422=>"010111111",
  37423=>"100000110",
  37424=>"001000000",
  37425=>"100111111",
  37426=>"010001101",
  37427=>"100001111",
  37428=>"010010100",
  37429=>"001100011",
  37430=>"000001101",
  37431=>"100001011",
  37432=>"000000011",
  37433=>"110100110",
  37434=>"101011100",
  37435=>"011011001",
  37436=>"000111011",
  37437=>"100000110",
  37438=>"100111111",
  37439=>"111001001",
  37440=>"100111110",
  37441=>"011110101",
  37442=>"100110010",
  37443=>"001011111",
  37444=>"110100111",
  37445=>"010110001",
  37446=>"111111001",
  37447=>"111000100",
  37448=>"100011000",
  37449=>"111101101",
  37450=>"111100011",
  37451=>"000101110",
  37452=>"011110110",
  37453=>"110011100",
  37454=>"001111111",
  37455=>"110100111",
  37456=>"000000100",
  37457=>"111011110",
  37458=>"111110001",
  37459=>"010011001",
  37460=>"001001100",
  37461=>"100110101",
  37462=>"000110110",
  37463=>"101011010",
  37464=>"100010010",
  37465=>"001001101",
  37466=>"111111000",
  37467=>"101000000",
  37468=>"110111101",
  37469=>"011001010",
  37470=>"111111110",
  37471=>"100000010",
  37472=>"100111111",
  37473=>"001110100",
  37474=>"010010110",
  37475=>"110011000",
  37476=>"010000100",
  37477=>"000110101",
  37478=>"001001100",
  37479=>"011110010",
  37480=>"010001111",
  37481=>"110010000",
  37482=>"111010111",
  37483=>"001001101",
  37484=>"101101110",
  37485=>"000100001",
  37486=>"101101010",
  37487=>"011010010",
  37488=>"110010000",
  37489=>"000011010",
  37490=>"101101111",
  37491=>"100011011",
  37492=>"000111011",
  37493=>"111100101",
  37494=>"110010100",
  37495=>"110101011",
  37496=>"110010001",
  37497=>"001001101",
  37498=>"000111101",
  37499=>"100000001",
  37500=>"110110101",
  37501=>"001000011",
  37502=>"010101001",
  37503=>"010110000",
  37504=>"010100101",
  37505=>"111111111",
  37506=>"100000001",
  37507=>"101011011",
  37508=>"110011101",
  37509=>"001001111",
  37510=>"101100111",
  37511=>"111100111",
  37512=>"101111110",
  37513=>"010101000",
  37514=>"011010101",
  37515=>"010110110",
  37516=>"100011100",
  37517=>"000111110",
  37518=>"010110011",
  37519=>"010110111",
  37520=>"001110111",
  37521=>"101110100",
  37522=>"010101010",
  37523=>"001010101",
  37524=>"111101010",
  37525=>"111010010",
  37526=>"011100101",
  37527=>"100001111",
  37528=>"101000000",
  37529=>"011101111",
  37530=>"100110000",
  37531=>"000110001",
  37532=>"101101101",
  37533=>"000100000",
  37534=>"010010000",
  37535=>"110001010",
  37536=>"100100000",
  37537=>"001010111",
  37538=>"101010000",
  37539=>"100100001",
  37540=>"100001110",
  37541=>"110010010",
  37542=>"010111000",
  37543=>"100000100",
  37544=>"101110101",
  37545=>"100001000",
  37546=>"001010000",
  37547=>"000101110",
  37548=>"110000011",
  37549=>"000001000",
  37550=>"001010111",
  37551=>"000101111",
  37552=>"000001011",
  37553=>"101000010",
  37554=>"111010000",
  37555=>"010000111",
  37556=>"110111011",
  37557=>"101110110",
  37558=>"101010110",
  37559=>"100010000",
  37560=>"011101001",
  37561=>"010101010",
  37562=>"111101101",
  37563=>"011011011",
  37564=>"111111001",
  37565=>"000101011",
  37566=>"100001001",
  37567=>"010010101",
  37568=>"101100000",
  37569=>"000101000",
  37570=>"110111010",
  37571=>"111100111",
  37572=>"110111010",
  37573=>"010011000",
  37574=>"010101100",
  37575=>"100100101",
  37576=>"001000010",
  37577=>"100010001",
  37578=>"011011101",
  37579=>"101100011",
  37580=>"100001100",
  37581=>"011111110",
  37582=>"001001000",
  37583=>"010110010",
  37584=>"011110010",
  37585=>"001110101",
  37586=>"100101001",
  37587=>"110100111",
  37588=>"000010010",
  37589=>"001011111",
  37590=>"011001000",
  37591=>"101000000",
  37592=>"101011001",
  37593=>"010000001",
  37594=>"000010000",
  37595=>"101100111",
  37596=>"010011110",
  37597=>"010000110",
  37598=>"110011101",
  37599=>"011101011",
  37600=>"001011111",
  37601=>"100110001",
  37602=>"111011111",
  37603=>"100101100",
  37604=>"110001101",
  37605=>"111001011",
  37606=>"100010111",
  37607=>"011100111",
  37608=>"010101011",
  37609=>"010001111",
  37610=>"101000001",
  37611=>"101000100",
  37612=>"100100101",
  37613=>"100001000",
  37614=>"001001110",
  37615=>"101001011",
  37616=>"011100010",
  37617=>"110001101",
  37618=>"010111111",
  37619=>"000010010",
  37620=>"010010110",
  37621=>"111111110",
  37622=>"010010111",
  37623=>"100000111",
  37624=>"111010001",
  37625=>"110000001",
  37626=>"001001111",
  37627=>"101000011",
  37628=>"110000001",
  37629=>"010010100",
  37630=>"000001111",
  37631=>"001110001",
  37632=>"100001001",
  37633=>"111000001",
  37634=>"101101101",
  37635=>"101000111",
  37636=>"001010100",
  37637=>"011001001",
  37638=>"000111100",
  37639=>"011001011",
  37640=>"000100101",
  37641=>"001001101",
  37642=>"010011000",
  37643=>"001110011",
  37644=>"001010000",
  37645=>"111100100",
  37646=>"010110110",
  37647=>"110000000",
  37648=>"111011111",
  37649=>"111000011",
  37650=>"011100100",
  37651=>"001100001",
  37652=>"010011111",
  37653=>"101000111",
  37654=>"101100000",
  37655=>"100011011",
  37656=>"000011100",
  37657=>"010100001",
  37658=>"001010101",
  37659=>"110011110",
  37660=>"010110011",
  37661=>"110100010",
  37662=>"100111011",
  37663=>"001000100",
  37664=>"101111101",
  37665=>"010010110",
  37666=>"001001111",
  37667=>"000000110",
  37668=>"010110100",
  37669=>"010001011",
  37670=>"100101111",
  37671=>"100111011",
  37672=>"111101100",
  37673=>"111101100",
  37674=>"011010111",
  37675=>"111011000",
  37676=>"111101001",
  37677=>"011001110",
  37678=>"110101111",
  37679=>"010000001",
  37680=>"001001110",
  37681=>"000100111",
  37682=>"110110101",
  37683=>"111001001",
  37684=>"101111111",
  37685=>"101000100",
  37686=>"010000110",
  37687=>"010011100",
  37688=>"011101100",
  37689=>"000011010",
  37690=>"101111110",
  37691=>"001101000",
  37692=>"111111011",
  37693=>"101000001",
  37694=>"100100010",
  37695=>"001100000",
  37696=>"100001001",
  37697=>"000000001",
  37698=>"010101011",
  37699=>"110110001",
  37700=>"000010001",
  37701=>"001110010",
  37702=>"000011111",
  37703=>"110101101",
  37704=>"011100100",
  37705=>"011100101",
  37706=>"111010000",
  37707=>"000000000",
  37708=>"010000010",
  37709=>"110000101",
  37710=>"000110011",
  37711=>"000000110",
  37712=>"000110100",
  37713=>"110111011",
  37714=>"111111100",
  37715=>"101100100",
  37716=>"101010011",
  37717=>"000110011",
  37718=>"000100001",
  37719=>"110010110",
  37720=>"001111001",
  37721=>"001001010",
  37722=>"011001010",
  37723=>"001101001",
  37724=>"001011110",
  37725=>"101011100",
  37726=>"000111000",
  37727=>"010101010",
  37728=>"100101100",
  37729=>"000011111",
  37730=>"101101101",
  37731=>"111010100",
  37732=>"011100001",
  37733=>"110001000",
  37734=>"100100011",
  37735=>"101011111",
  37736=>"100101010",
  37737=>"111010010",
  37738=>"100011111",
  37739=>"010011001",
  37740=>"011101001",
  37741=>"100100000",
  37742=>"110000001",
  37743=>"001000100",
  37744=>"001110011",
  37745=>"110010000",
  37746=>"001010111",
  37747=>"001011001",
  37748=>"110100101",
  37749=>"011111011",
  37750=>"000100000",
  37751=>"011011110",
  37752=>"110110101",
  37753=>"000101001",
  37754=>"100111100",
  37755=>"010011111",
  37756=>"000101000",
  37757=>"100110111",
  37758=>"000011111",
  37759=>"000001111",
  37760=>"011000100",
  37761=>"111100111",
  37762=>"110100111",
  37763=>"000101011",
  37764=>"110111110",
  37765=>"110001000",
  37766=>"110111110",
  37767=>"000010010",
  37768=>"001000110",
  37769=>"100111000",
  37770=>"000000001",
  37771=>"110101010",
  37772=>"000000010",
  37773=>"000100111",
  37774=>"100100110",
  37775=>"101111011",
  37776=>"111110100",
  37777=>"010111101",
  37778=>"011010011",
  37779=>"101100000",
  37780=>"011110001",
  37781=>"100100010",
  37782=>"101101111",
  37783=>"100001100",
  37784=>"011011100",
  37785=>"111011101",
  37786=>"011111010",
  37787=>"111001110",
  37788=>"001010001",
  37789=>"010001110",
  37790=>"001111001",
  37791=>"010000010",
  37792=>"100000100",
  37793=>"000100100",
  37794=>"110010101",
  37795=>"100110001",
  37796=>"010100011",
  37797=>"011110101",
  37798=>"101001010",
  37799=>"101110101",
  37800=>"100001101",
  37801=>"101110000",
  37802=>"010110001",
  37803=>"101011010",
  37804=>"010001011",
  37805=>"001101111",
  37806=>"011111011",
  37807=>"100000010",
  37808=>"010100010",
  37809=>"000000001",
  37810=>"100000101",
  37811=>"110010110",
  37812=>"001100101",
  37813=>"000101111",
  37814=>"010110000",
  37815=>"011011110",
  37816=>"011000000",
  37817=>"000001011",
  37818=>"111010000",
  37819=>"010001101",
  37820=>"110010010",
  37821=>"010110011",
  37822=>"111011010",
  37823=>"111100100",
  37824=>"010011000",
  37825=>"110111001",
  37826=>"101100101",
  37827=>"101101010",
  37828=>"101011111",
  37829=>"010001010",
  37830=>"110000011",
  37831=>"100011111",
  37832=>"011001010",
  37833=>"001011111",
  37834=>"001111011",
  37835=>"010010000",
  37836=>"110001010",
  37837=>"110110010",
  37838=>"111001101",
  37839=>"101001100",
  37840=>"011001000",
  37841=>"011000011",
  37842=>"001100111",
  37843=>"000000000",
  37844=>"000010001",
  37845=>"100000000",
  37846=>"111000010",
  37847=>"110010001",
  37848=>"110111100",
  37849=>"110011110",
  37850=>"100001000",
  37851=>"011001001",
  37852=>"001111110",
  37853=>"010110000",
  37854=>"111000000",
  37855=>"111001011",
  37856=>"011011000",
  37857=>"100011101",
  37858=>"000010101",
  37859=>"110011100",
  37860=>"000101001",
  37861=>"011011101",
  37862=>"100011001",
  37863=>"010001100",
  37864=>"100101101",
  37865=>"011101101",
  37866=>"111001111",
  37867=>"110110110",
  37868=>"101100101",
  37869=>"000010110",
  37870=>"110110111",
  37871=>"100001010",
  37872=>"000010010",
  37873=>"010001011",
  37874=>"000101001",
  37875=>"001011001",
  37876=>"111000001",
  37877=>"010101101",
  37878=>"000011111",
  37879=>"001000101",
  37880=>"110011100",
  37881=>"100111000",
  37882=>"111001001",
  37883=>"100001110",
  37884=>"011000000",
  37885=>"000000011",
  37886=>"100100010",
  37887=>"111000011",
  37888=>"101101101",
  37889=>"101001101",
  37890=>"100000010",
  37891=>"100010100",
  37892=>"100110001",
  37893=>"001100001",
  37894=>"000111010",
  37895=>"011011100",
  37896=>"010010100",
  37897=>"010001001",
  37898=>"000100111",
  37899=>"001110011",
  37900=>"011110010",
  37901=>"101001100",
  37902=>"011000101",
  37903=>"100001001",
  37904=>"000011111",
  37905=>"100101111",
  37906=>"101000000",
  37907=>"011101001",
  37908=>"010110111",
  37909=>"001100110",
  37910=>"111001111",
  37911=>"001100111",
  37912=>"010001110",
  37913=>"000000001",
  37914=>"010001011",
  37915=>"001110010",
  37916=>"010111001",
  37917=>"001001111",
  37918=>"111010010",
  37919=>"100001101",
  37920=>"001010111",
  37921=>"110000100",
  37922=>"011000001",
  37923=>"011111100",
  37924=>"100110000",
  37925=>"001001001",
  37926=>"010010111",
  37927=>"100000110",
  37928=>"111101110",
  37929=>"000010100",
  37930=>"000111100",
  37931=>"001001100",
  37932=>"101110001",
  37933=>"110101010",
  37934=>"111100110",
  37935=>"000100110",
  37936=>"000010110",
  37937=>"010110100",
  37938=>"111100000",
  37939=>"111010011",
  37940=>"010100101",
  37941=>"011001000",
  37942=>"010010011",
  37943=>"011000110",
  37944=>"110101100",
  37945=>"100101010",
  37946=>"010100001",
  37947=>"010110000",
  37948=>"101011010",
  37949=>"010010100",
  37950=>"101011110",
  37951=>"010010110",
  37952=>"101000000",
  37953=>"111110101",
  37954=>"010110101",
  37955=>"000111101",
  37956=>"001010110",
  37957=>"100100000",
  37958=>"101111001",
  37959=>"101101001",
  37960=>"101101010",
  37961=>"101010111",
  37962=>"010100011",
  37963=>"101011110",
  37964=>"101000101",
  37965=>"010100011",
  37966=>"101011101",
  37967=>"101111111",
  37968=>"110111010",
  37969=>"000010110",
  37970=>"011011110",
  37971=>"100000100",
  37972=>"100100101",
  37973=>"111001100",
  37974=>"111010110",
  37975=>"001100110",
  37976=>"001010111",
  37977=>"011110010",
  37978=>"000100101",
  37979=>"100100010",
  37980=>"001111011",
  37981=>"101110111",
  37982=>"111001000",
  37983=>"110101010",
  37984=>"101000001",
  37985=>"010101111",
  37986=>"010101110",
  37987=>"011000110",
  37988=>"110000111",
  37989=>"000101011",
  37990=>"111100111",
  37991=>"000010101",
  37992=>"110101100",
  37993=>"100110010",
  37994=>"111011111",
  37995=>"010101001",
  37996=>"111011001",
  37997=>"111001101",
  37998=>"010000111",
  37999=>"011011010",
  38000=>"111100000",
  38001=>"001111011",
  38002=>"010111000",
  38003=>"101001111",
  38004=>"111101111",
  38005=>"111100110",
  38006=>"000100000",
  38007=>"010000100",
  38008=>"010110110",
  38009=>"000010110",
  38010=>"000100110",
  38011=>"001100101",
  38012=>"001000010",
  38013=>"101111000",
  38014=>"001110000",
  38015=>"101001001",
  38016=>"011000101",
  38017=>"110000011",
  38018=>"000100010",
  38019=>"110010001",
  38020=>"110111010",
  38021=>"011000011",
  38022=>"011111101",
  38023=>"001111110",
  38024=>"110000000",
  38025=>"110110101",
  38026=>"000101110",
  38027=>"010001110",
  38028=>"010000110",
  38029=>"111111110",
  38030=>"111111010",
  38031=>"011011101",
  38032=>"001011111",
  38033=>"111100111",
  38034=>"001100000",
  38035=>"001001011",
  38036=>"110001101",
  38037=>"111101011",
  38038=>"100110111",
  38039=>"110111010",
  38040=>"110011100",
  38041=>"000110001",
  38042=>"100010000",
  38043=>"001001000",
  38044=>"010001100",
  38045=>"100100100",
  38046=>"110011001",
  38047=>"111001010",
  38048=>"100110110",
  38049=>"101100110",
  38050=>"011100100",
  38051=>"110100100",
  38052=>"001000110",
  38053=>"001111100",
  38054=>"100010011",
  38055=>"100111001",
  38056=>"100111110",
  38057=>"101011101",
  38058=>"010011001",
  38059=>"111000101",
  38060=>"110101111",
  38061=>"001011100",
  38062=>"100110101",
  38063=>"111110101",
  38064=>"010101111",
  38065=>"011000000",
  38066=>"111011100",
  38067=>"011101011",
  38068=>"111110001",
  38069=>"010110101",
  38070=>"011111011",
  38071=>"111110100",
  38072=>"000000101",
  38073=>"111001001",
  38074=>"100100001",
  38075=>"011110100",
  38076=>"001111101",
  38077=>"011100000",
  38078=>"011001001",
  38079=>"001101001",
  38080=>"110111100",
  38081=>"011110101",
  38082=>"001100111",
  38083=>"101100100",
  38084=>"011110010",
  38085=>"100010001",
  38086=>"111000110",
  38087=>"000010110",
  38088=>"001101010",
  38089=>"101110011",
  38090=>"010110001",
  38091=>"000011000",
  38092=>"111001110",
  38093=>"000110100",
  38094=>"111011100",
  38095=>"101100000",
  38096=>"100110101",
  38097=>"110111010",
  38098=>"000100010",
  38099=>"101100011",
  38100=>"001011110",
  38101=>"011110111",
  38102=>"010101101",
  38103=>"110001110",
  38104=>"000001001",
  38105=>"100000100",
  38106=>"101110100",
  38107=>"001100111",
  38108=>"101111100",
  38109=>"111011001",
  38110=>"101011110",
  38111=>"010110011",
  38112=>"000010001",
  38113=>"101110011",
  38114=>"010111100",
  38115=>"011110100",
  38116=>"000101110",
  38117=>"110101011",
  38118=>"110010111",
  38119=>"010011001",
  38120=>"110010001",
  38121=>"100100001",
  38122=>"000000001",
  38123=>"110110111",
  38124=>"010011111",
  38125=>"110110011",
  38126=>"000000011",
  38127=>"011011101",
  38128=>"000000010",
  38129=>"101110111",
  38130=>"110100011",
  38131=>"010001101",
  38132=>"111111100",
  38133=>"000100101",
  38134=>"001100011",
  38135=>"100101101",
  38136=>"011001110",
  38137=>"011011111",
  38138=>"011111110",
  38139=>"100010000",
  38140=>"101000100",
  38141=>"001001110",
  38142=>"110111100",
  38143=>"110010111",
  38144=>"001001100",
  38145=>"100010001",
  38146=>"100001100",
  38147=>"110000010",
  38148=>"011000101",
  38149=>"100000110",
  38150=>"101101111",
  38151=>"000101000",
  38152=>"110001110",
  38153=>"101000110",
  38154=>"011001010",
  38155=>"000011100",
  38156=>"010000011",
  38157=>"011101001",
  38158=>"100010010",
  38159=>"000110100",
  38160=>"101011001",
  38161=>"101000100",
  38162=>"000101110",
  38163=>"100111101",
  38164=>"001010000",
  38165=>"100111100",
  38166=>"010111011",
  38167=>"100001000",
  38168=>"011100011",
  38169=>"110001011",
  38170=>"111010100",
  38171=>"010101110",
  38172=>"100011000",
  38173=>"111001101",
  38174=>"110101011",
  38175=>"001001011",
  38176=>"111000100",
  38177=>"100011010",
  38178=>"010111111",
  38179=>"010010010",
  38180=>"010010011",
  38181=>"000000001",
  38182=>"101111011",
  38183=>"010100101",
  38184=>"001000101",
  38185=>"101000100",
  38186=>"000111001",
  38187=>"001011110",
  38188=>"100010001",
  38189=>"100100000",
  38190=>"101000011",
  38191=>"100100010",
  38192=>"101011010",
  38193=>"111111111",
  38194=>"110010111",
  38195=>"101111010",
  38196=>"100011010",
  38197=>"000100110",
  38198=>"011001011",
  38199=>"000110111",
  38200=>"111010001",
  38201=>"101001011",
  38202=>"110001100",
  38203=>"110111110",
  38204=>"111011111",
  38205=>"011011101",
  38206=>"001101010",
  38207=>"100011100",
  38208=>"011001100",
  38209=>"000100100",
  38210=>"100100010",
  38211=>"100000011",
  38212=>"100000101",
  38213=>"101010011",
  38214=>"111110011",
  38215=>"000001011",
  38216=>"001110001",
  38217=>"101001010",
  38218=>"001111011",
  38219=>"111000010",
  38220=>"000010011",
  38221=>"111001110",
  38222=>"001101101",
  38223=>"111101111",
  38224=>"001101101",
  38225=>"011111001",
  38226=>"000110110",
  38227=>"011011111",
  38228=>"000001111",
  38229=>"100100010",
  38230=>"001010110",
  38231=>"000110101",
  38232=>"011110101",
  38233=>"011000111",
  38234=>"000000111",
  38235=>"001101100",
  38236=>"011100001",
  38237=>"101111110",
  38238=>"000001001",
  38239=>"000100100",
  38240=>"110100000",
  38241=>"100110011",
  38242=>"101101100",
  38243=>"000001010",
  38244=>"100011000",
  38245=>"110010100",
  38246=>"100110010",
  38247=>"001111110",
  38248=>"011101110",
  38249=>"101000001",
  38250=>"000110001",
  38251=>"111001010",
  38252=>"111110010",
  38253=>"010101100",
  38254=>"010000110",
  38255=>"111100001",
  38256=>"000110000",
  38257=>"101000101",
  38258=>"001000111",
  38259=>"101110111",
  38260=>"011100111",
  38261=>"110101001",
  38262=>"110111110",
  38263=>"101011001",
  38264=>"111111011",
  38265=>"111011100",
  38266=>"011100111",
  38267=>"111101100",
  38268=>"000101111",
  38269=>"000011110",
  38270=>"011101101",
  38271=>"110010010",
  38272=>"010101100",
  38273=>"100001111",
  38274=>"110100100",
  38275=>"001101001",
  38276=>"100000000",
  38277=>"000010000",
  38278=>"001010011",
  38279=>"111100110",
  38280=>"110110100",
  38281=>"101010100",
  38282=>"111111000",
  38283=>"101110000",
  38284=>"011010010",
  38285=>"111110101",
  38286=>"010000000",
  38287=>"001110000",
  38288=>"001000111",
  38289=>"110101000",
  38290=>"100010110",
  38291=>"010011001",
  38292=>"111110111",
  38293=>"011011110",
  38294=>"001010000",
  38295=>"100110000",
  38296=>"101011000",
  38297=>"010111110",
  38298=>"001101111",
  38299=>"011010111",
  38300=>"111011011",
  38301=>"101011111",
  38302=>"011110110",
  38303=>"110110111",
  38304=>"010011100",
  38305=>"010001101",
  38306=>"111011000",
  38307=>"101001100",
  38308=>"001101100",
  38309=>"100111000",
  38310=>"111101000",
  38311=>"001101000",
  38312=>"100101110",
  38313=>"100011100",
  38314=>"101000111",
  38315=>"110101011",
  38316=>"101111011",
  38317=>"010010010",
  38318=>"100001110",
  38319=>"001010110",
  38320=>"101001000",
  38321=>"001101111",
  38322=>"100100000",
  38323=>"110100101",
  38324=>"011111001",
  38325=>"111001100",
  38326=>"011100110",
  38327=>"100010100",
  38328=>"011111010",
  38329=>"010111111",
  38330=>"101000111",
  38331=>"101010000",
  38332=>"011011101",
  38333=>"011010110",
  38334=>"110001000",
  38335=>"011011101",
  38336=>"011110001",
  38337=>"111110101",
  38338=>"011110010",
  38339=>"110110111",
  38340=>"111101100",
  38341=>"100001000",
  38342=>"111110000",
  38343=>"111011010",
  38344=>"100010110",
  38345=>"010111111",
  38346=>"011000010",
  38347=>"011011001",
  38348=>"111100111",
  38349=>"110000011",
  38350=>"100100111",
  38351=>"111101001",
  38352=>"110010101",
  38353=>"001011110",
  38354=>"111101010",
  38355=>"110000010",
  38356=>"010101001",
  38357=>"000001001",
  38358=>"011001111",
  38359=>"100100000",
  38360=>"110010100",
  38361=>"110011000",
  38362=>"111011111",
  38363=>"110011101",
  38364=>"110101011",
  38365=>"000000100",
  38366=>"001001000",
  38367=>"100110100",
  38368=>"110111110",
  38369=>"111011011",
  38370=>"000110010",
  38371=>"010100111",
  38372=>"110100000",
  38373=>"101001101",
  38374=>"001010101",
  38375=>"100011101",
  38376=>"110101100",
  38377=>"110100001",
  38378=>"111000101",
  38379=>"100111111",
  38380=>"100101101",
  38381=>"100000110",
  38382=>"111101111",
  38383=>"100011110",
  38384=>"001100101",
  38385=>"110001011",
  38386=>"110000110",
  38387=>"110010011",
  38388=>"101001011",
  38389=>"011011000",
  38390=>"111011010",
  38391=>"100110000",
  38392=>"110100101",
  38393=>"101101110",
  38394=>"011011101",
  38395=>"110011111",
  38396=>"110001111",
  38397=>"000000010",
  38398=>"111011001",
  38399=>"001010000",
  38400=>"111110111",
  38401=>"101011010",
  38402=>"101101011",
  38403=>"011001001",
  38404=>"011000001",
  38405=>"100010011",
  38406=>"010100001",
  38407=>"101100100",
  38408=>"100000110",
  38409=>"001001111",
  38410=>"111010001",
  38411=>"001010001",
  38412=>"101011111",
  38413=>"001001100",
  38414=>"101110110",
  38415=>"101101100",
  38416=>"000011011",
  38417=>"110011000",
  38418=>"010010100",
  38419=>"010100011",
  38420=>"110100100",
  38421=>"111010011",
  38422=>"000110011",
  38423=>"110010000",
  38424=>"000001000",
  38425=>"000011011",
  38426=>"110000001",
  38427=>"010011001",
  38428=>"110001100",
  38429=>"000111111",
  38430=>"011000101",
  38431=>"100001110",
  38432=>"111001111",
  38433=>"010011101",
  38434=>"110110001",
  38435=>"101001001",
  38436=>"011111111",
  38437=>"000000011",
  38438=>"100001000",
  38439=>"010101101",
  38440=>"000111010",
  38441=>"000000000",
  38442=>"110010010",
  38443=>"001100001",
  38444=>"011011011",
  38445=>"110011010",
  38446=>"001000001",
  38447=>"011010101",
  38448=>"010000010",
  38449=>"000001010",
  38450=>"000110111",
  38451=>"110111001",
  38452=>"010110101",
  38453=>"000011010",
  38454=>"101100111",
  38455=>"011100010",
  38456=>"110011100",
  38457=>"001100111",
  38458=>"100010010",
  38459=>"010101101",
  38460=>"001011001",
  38461=>"000110000",
  38462=>"001110100",
  38463=>"100001010",
  38464=>"010001001",
  38465=>"101000111",
  38466=>"110000101",
  38467=>"000000100",
  38468=>"010110011",
  38469=>"001010111",
  38470=>"000001001",
  38471=>"100100001",
  38472=>"101000000",
  38473=>"100011001",
  38474=>"010000001",
  38475=>"101110000",
  38476=>"101000000",
  38477=>"000011111",
  38478=>"101110101",
  38479=>"110001001",
  38480=>"010101110",
  38481=>"001000111",
  38482=>"101100011",
  38483=>"101110101",
  38484=>"010101101",
  38485=>"111010010",
  38486=>"110100001",
  38487=>"011101011",
  38488=>"101101011",
  38489=>"000110101",
  38490=>"111111011",
  38491=>"011100101",
  38492=>"001111001",
  38493=>"011010100",
  38494=>"111011100",
  38495=>"000001001",
  38496=>"111001000",
  38497=>"101110111",
  38498=>"010010101",
  38499=>"110010010",
  38500=>"111000110",
  38501=>"101111000",
  38502=>"110111010",
  38503=>"000110000",
  38504=>"110110010",
  38505=>"010010101",
  38506=>"001111001",
  38507=>"101001111",
  38508=>"000100110",
  38509=>"101111001",
  38510=>"010011001",
  38511=>"101110000",
  38512=>"111010101",
  38513=>"000010010",
  38514=>"110110001",
  38515=>"111101100",
  38516=>"000110111",
  38517=>"001000010",
  38518=>"001010111",
  38519=>"111110001",
  38520=>"101011111",
  38521=>"001001100",
  38522=>"010101000",
  38523=>"111001000",
  38524=>"001000001",
  38525=>"000101101",
  38526=>"111011010",
  38527=>"101101000",
  38528=>"111000001",
  38529=>"101011000",
  38530=>"100001001",
  38531=>"100011110",
  38532=>"111011001",
  38533=>"001101010",
  38534=>"111011111",
  38535=>"000100010",
  38536=>"000101010",
  38537=>"001110000",
  38538=>"111000101",
  38539=>"000001101",
  38540=>"001010001",
  38541=>"100001110",
  38542=>"110111011",
  38543=>"101110110",
  38544=>"101110111",
  38545=>"111001111",
  38546=>"010001001",
  38547=>"000010000",
  38548=>"000100000",
  38549=>"010110001",
  38550=>"100110000",
  38551=>"101100100",
  38552=>"111010010",
  38553=>"111011001",
  38554=>"111100111",
  38555=>"100001011",
  38556=>"110110010",
  38557=>"001110110",
  38558=>"001101101",
  38559=>"100000111",
  38560=>"010011110",
  38561=>"110010010",
  38562=>"001100010",
  38563=>"001111111",
  38564=>"011111111",
  38565=>"010001000",
  38566=>"001111110",
  38567=>"111010001",
  38568=>"000000011",
  38569=>"010101000",
  38570=>"110100110",
  38571=>"010000101",
  38572=>"011101010",
  38573=>"000001111",
  38574=>"011110010",
  38575=>"001000101",
  38576=>"110101111",
  38577=>"111010011",
  38578=>"001100001",
  38579=>"100101010",
  38580=>"110101010",
  38581=>"000000011",
  38582=>"100101111",
  38583=>"110110111",
  38584=>"010100101",
  38585=>"011100110",
  38586=>"001111001",
  38587=>"011101001",
  38588=>"000000010",
  38589=>"010010011",
  38590=>"000110101",
  38591=>"001111000",
  38592=>"000011100",
  38593=>"101110001",
  38594=>"011110011",
  38595=>"010000000",
  38596=>"000000011",
  38597=>"010001011",
  38598=>"011010000",
  38599=>"110110110",
  38600=>"010001000",
  38601=>"001111010",
  38602=>"110000000",
  38603=>"011100101",
  38604=>"111111101",
  38605=>"010100001",
  38606=>"111001111",
  38607=>"011100101",
  38608=>"100001011",
  38609=>"100111110",
  38610=>"011011010",
  38611=>"000001000",
  38612=>"111110111",
  38613=>"100110100",
  38614=>"101110010",
  38615=>"100111111",
  38616=>"101100001",
  38617=>"000010011",
  38618=>"011101001",
  38619=>"010111000",
  38620=>"000001111",
  38621=>"100101000",
  38622=>"011111100",
  38623=>"111100001",
  38624=>"010011100",
  38625=>"110011110",
  38626=>"010000100",
  38627=>"011101001",
  38628=>"100011011",
  38629=>"100010100",
  38630=>"100000010",
  38631=>"101110011",
  38632=>"001000111",
  38633=>"101111001",
  38634=>"101111101",
  38635=>"111101100",
  38636=>"101001010",
  38637=>"001011011",
  38638=>"100000000",
  38639=>"110011101",
  38640=>"011101111",
  38641=>"010010101",
  38642=>"110100101",
  38643=>"010000101",
  38644=>"110000111",
  38645=>"101110100",
  38646=>"100110110",
  38647=>"010001110",
  38648=>"111011001",
  38649=>"000000111",
  38650=>"111110101",
  38651=>"010000001",
  38652=>"010100110",
  38653=>"010011110",
  38654=>"111110001",
  38655=>"010001010",
  38656=>"110001001",
  38657=>"111010101",
  38658=>"010110010",
  38659=>"100010000",
  38660=>"101101011",
  38661=>"001000100",
  38662=>"110010100",
  38663=>"110001011",
  38664=>"100011110",
  38665=>"011010111",
  38666=>"110101010",
  38667=>"110100001",
  38668=>"001010000",
  38669=>"011110011",
  38670=>"111010001",
  38671=>"110011010",
  38672=>"011000001",
  38673=>"100100000",
  38674=>"100111101",
  38675=>"000110010",
  38676=>"001100010",
  38677=>"001111111",
  38678=>"101111101",
  38679=>"001111000",
  38680=>"001000000",
  38681=>"101001010",
  38682=>"000011100",
  38683=>"111110101",
  38684=>"100100000",
  38685=>"011000101",
  38686=>"100111101",
  38687=>"110001000",
  38688=>"101110101",
  38689=>"011110011",
  38690=>"101100111",
  38691=>"111110110",
  38692=>"001001101",
  38693=>"101100000",
  38694=>"001011110",
  38695=>"110110001",
  38696=>"011010100",
  38697=>"001110110",
  38698=>"010101111",
  38699=>"011101100",
  38700=>"101000001",
  38701=>"011110110",
  38702=>"000010010",
  38703=>"100001000",
  38704=>"000011011",
  38705=>"101110011",
  38706=>"011111011",
  38707=>"010001111",
  38708=>"011000101",
  38709=>"001010100",
  38710=>"000011100",
  38711=>"011101111",
  38712=>"111111010",
  38713=>"101011000",
  38714=>"011111001",
  38715=>"111110000",
  38716=>"010101101",
  38717=>"000111101",
  38718=>"101101010",
  38719=>"101101111",
  38720=>"111111011",
  38721=>"001000010",
  38722=>"100111011",
  38723=>"110100000",
  38724=>"001101011",
  38725=>"001000010",
  38726=>"101011001",
  38727=>"011010011",
  38728=>"001011110",
  38729=>"001011001",
  38730=>"100110000",
  38731=>"101010010",
  38732=>"011010010",
  38733=>"100111101",
  38734=>"011010101",
  38735=>"000000011",
  38736=>"011001000",
  38737=>"101001001",
  38738=>"101000001",
  38739=>"001010101",
  38740=>"001001001",
  38741=>"110100110",
  38742=>"001110011",
  38743=>"010100010",
  38744=>"010010001",
  38745=>"110010111",
  38746=>"111101100",
  38747=>"001110100",
  38748=>"000100000",
  38749=>"011011010",
  38750=>"110011011",
  38751=>"000010100",
  38752=>"000010000",
  38753=>"001010010",
  38754=>"011100011",
  38755=>"110111011",
  38756=>"011111001",
  38757=>"111110000",
  38758=>"000111010",
  38759=>"111101111",
  38760=>"001011100",
  38761=>"101011000",
  38762=>"110010100",
  38763=>"100000000",
  38764=>"100011100",
  38765=>"000001111",
  38766=>"111011010",
  38767=>"101001101",
  38768=>"001000001",
  38769=>"101010011",
  38770=>"100001101",
  38771=>"110000001",
  38772=>"111101011",
  38773=>"010110001",
  38774=>"110111000",
  38775=>"001100101",
  38776=>"111001100",
  38777=>"100000001",
  38778=>"000101100",
  38779=>"001000100",
  38780=>"000001111",
  38781=>"101110000",
  38782=>"100000100",
  38783=>"001111101",
  38784=>"110110111",
  38785=>"110011001",
  38786=>"100000011",
  38787=>"101001110",
  38788=>"101110001",
  38789=>"100100101",
  38790=>"100101111",
  38791=>"001000000",
  38792=>"110111101",
  38793=>"011110000",
  38794=>"111100011",
  38795=>"011010101",
  38796=>"111111010",
  38797=>"110110000",
  38798=>"101011111",
  38799=>"001101110",
  38800=>"001001100",
  38801=>"010001011",
  38802=>"100001011",
  38803=>"100110111",
  38804=>"111010101",
  38805=>"000101011",
  38806=>"111110111",
  38807=>"001000101",
  38808=>"011010110",
  38809=>"001111101",
  38810=>"000111011",
  38811=>"111010000",
  38812=>"010100000",
  38813=>"110111000",
  38814=>"111100011",
  38815=>"101000001",
  38816=>"111001001",
  38817=>"111110101",
  38818=>"110111110",
  38819=>"011100101",
  38820=>"000111010",
  38821=>"011000101",
  38822=>"010110011",
  38823=>"000111010",
  38824=>"110000101",
  38825=>"010101011",
  38826=>"111110111",
  38827=>"010110000",
  38828=>"110010110",
  38829=>"101010100",
  38830=>"100111101",
  38831=>"111011101",
  38832=>"100010100",
  38833=>"000101110",
  38834=>"110011000",
  38835=>"100000100",
  38836=>"010011110",
  38837=>"111001011",
  38838=>"001000111",
  38839=>"100110000",
  38840=>"001010010",
  38841=>"101100111",
  38842=>"001000000",
  38843=>"110110010",
  38844=>"010111011",
  38845=>"000001110",
  38846=>"111010110",
  38847=>"001101001",
  38848=>"000010011",
  38849=>"011011111",
  38850=>"101010111",
  38851=>"110100100",
  38852=>"000100100",
  38853=>"011010011",
  38854=>"110001000",
  38855=>"111011010",
  38856=>"100110011",
  38857=>"010000111",
  38858=>"001100100",
  38859=>"110101110",
  38860=>"101111000",
  38861=>"010100001",
  38862=>"111000011",
  38863=>"010111101",
  38864=>"010111100",
  38865=>"000101100",
  38866=>"001111110",
  38867=>"101000000",
  38868=>"001000100",
  38869=>"010010100",
  38870=>"001101010",
  38871=>"000100101",
  38872=>"100111101",
  38873=>"010001011",
  38874=>"111011010",
  38875=>"101111010",
  38876=>"011111001",
  38877=>"111100110",
  38878=>"011011111",
  38879=>"111111111",
  38880=>"010000011",
  38881=>"010011001",
  38882=>"000110011",
  38883=>"001100110",
  38884=>"011000010",
  38885=>"000011000",
  38886=>"010011110",
  38887=>"111000111",
  38888=>"000101001",
  38889=>"011101001",
  38890=>"111110111",
  38891=>"010110011",
  38892=>"110111110",
  38893=>"110000100",
  38894=>"010111111",
  38895=>"010110000",
  38896=>"111000111",
  38897=>"100010000",
  38898=>"001001100",
  38899=>"101101100",
  38900=>"011010000",
  38901=>"111101100",
  38902=>"010011010",
  38903=>"111110110",
  38904=>"000010100",
  38905=>"101101000",
  38906=>"000101100",
  38907=>"001101011",
  38908=>"011100001",
  38909=>"111001000",
  38910=>"011011100",
  38911=>"101011001",
  38912=>"011100011",
  38913=>"000000000",
  38914=>"101010101",
  38915=>"000111100",
  38916=>"101000110",
  38917=>"100111010",
  38918=>"011001000",
  38919=>"001001011",
  38920=>"010011101",
  38921=>"010000110",
  38922=>"101000111",
  38923=>"110010100",
  38924=>"111111111",
  38925=>"011101010",
  38926=>"011110011",
  38927=>"001011000",
  38928=>"101110001",
  38929=>"000010101",
  38930=>"101110110",
  38931=>"011110001",
  38932=>"110011100",
  38933=>"101101011",
  38934=>"000110101",
  38935=>"101100100",
  38936=>"101001001",
  38937=>"111000011",
  38938=>"100001001",
  38939=>"111011111",
  38940=>"000011110",
  38941=>"101110110",
  38942=>"111111111",
  38943=>"101001010",
  38944=>"010000001",
  38945=>"000110101",
  38946=>"010101111",
  38947=>"011100011",
  38948=>"011000101",
  38949=>"010011000",
  38950=>"110100101",
  38951=>"111111011",
  38952=>"011010100",
  38953=>"001111011",
  38954=>"100011101",
  38955=>"010110101",
  38956=>"110011100",
  38957=>"010001111",
  38958=>"001100001",
  38959=>"111111100",
  38960=>"111100001",
  38961=>"000011110",
  38962=>"010100110",
  38963=>"110010010",
  38964=>"101001010",
  38965=>"011010110",
  38966=>"001001100",
  38967=>"111000010",
  38968=>"001000011",
  38969=>"000111011",
  38970=>"111111100",
  38971=>"101111110",
  38972=>"100101000",
  38973=>"100111111",
  38974=>"111100000",
  38975=>"011111101",
  38976=>"001010000",
  38977=>"001000111",
  38978=>"001110001",
  38979=>"111111001",
  38980=>"111100100",
  38981=>"000101010",
  38982=>"000110100",
  38983=>"010010001",
  38984=>"011000111",
  38985=>"111101111",
  38986=>"001001100",
  38987=>"000000110",
  38988=>"100001001",
  38989=>"101000110",
  38990=>"001000100",
  38991=>"111010100",
  38992=>"000010010",
  38993=>"011100101",
  38994=>"001001000",
  38995=>"010110100",
  38996=>"100010010",
  38997=>"001001111",
  38998=>"010101101",
  38999=>"000110000",
  39000=>"001001100",
  39001=>"001010000",
  39002=>"101111101",
  39003=>"001001010",
  39004=>"001110011",
  39005=>"010110011",
  39006=>"110100011",
  39007=>"101111101",
  39008=>"000010001",
  39009=>"100101100",
  39010=>"111010111",
  39011=>"000011100",
  39012=>"111100011",
  39013=>"011110010",
  39014=>"111001111",
  39015=>"011110101",
  39016=>"011100001",
  39017=>"011100001",
  39018=>"010010001",
  39019=>"100111011",
  39020=>"100000010",
  39021=>"101111011",
  39022=>"101010000",
  39023=>"011001111",
  39024=>"101111000",
  39025=>"110001000",
  39026=>"110010111",
  39027=>"101011011",
  39028=>"110001111",
  39029=>"110001111",
  39030=>"011001011",
  39031=>"111100111",
  39032=>"000001000",
  39033=>"010101101",
  39034=>"101000111",
  39035=>"110110101",
  39036=>"001000001",
  39037=>"011100100",
  39038=>"111001101",
  39039=>"100010011",
  39040=>"000001001",
  39041=>"010101001",
  39042=>"010010001",
  39043=>"001001111",
  39044=>"011111101",
  39045=>"101101110",
  39046=>"000001101",
  39047=>"110111010",
  39048=>"011101000",
  39049=>"001100000",
  39050=>"011110011",
  39051=>"100100000",
  39052=>"101011010",
  39053=>"010110111",
  39054=>"011100111",
  39055=>"101000001",
  39056=>"011001111",
  39057=>"010011110",
  39058=>"000010010",
  39059=>"011010100",
  39060=>"010001000",
  39061=>"001100111",
  39062=>"111000111",
  39063=>"101101111",
  39064=>"100110100",
  39065=>"110110010",
  39066=>"001000100",
  39067=>"101111111",
  39068=>"001000100",
  39069=>"101010000",
  39070=>"001111001",
  39071=>"010111010",
  39072=>"111101111",
  39073=>"011001001",
  39074=>"100001101",
  39075=>"101001101",
  39076=>"101001011",
  39077=>"010011100",
  39078=>"100110000",
  39079=>"001010000",
  39080=>"001001000",
  39081=>"111111011",
  39082=>"001101101",
  39083=>"101010111",
  39084=>"000100010",
  39085=>"001110011",
  39086=>"010111110",
  39087=>"110000100",
  39088=>"111011011",
  39089=>"000001001",
  39090=>"010011110",
  39091=>"100001100",
  39092=>"001011000",
  39093=>"111011101",
  39094=>"010011011",
  39095=>"110001001",
  39096=>"011101001",
  39097=>"001100110",
  39098=>"010001111",
  39099=>"100100110",
  39100=>"000111100",
  39101=>"000010101",
  39102=>"001001111",
  39103=>"111110111",
  39104=>"001110110",
  39105=>"001111110",
  39106=>"001010011",
  39107=>"010111100",
  39108=>"110111000",
  39109=>"101101111",
  39110=>"011010000",
  39111=>"101000011",
  39112=>"100010101",
  39113=>"000110100",
  39114=>"011101001",
  39115=>"001000111",
  39116=>"001000101",
  39117=>"010111000",
  39118=>"000011100",
  39119=>"101111100",
  39120=>"110100011",
  39121=>"000001100",
  39122=>"001101111",
  39123=>"110001101",
  39124=>"101000101",
  39125=>"001111010",
  39126=>"011001001",
  39127=>"111101010",
  39128=>"000000000",
  39129=>"100001111",
  39130=>"010011101",
  39131=>"101111000",
  39132=>"000101000",
  39133=>"101001111",
  39134=>"110010110",
  39135=>"100100000",
  39136=>"100011001",
  39137=>"000101110",
  39138=>"011110000",
  39139=>"110100000",
  39140=>"111111010",
  39141=>"011101100",
  39142=>"000110001",
  39143=>"010110110",
  39144=>"000001000",
  39145=>"000000101",
  39146=>"101111100",
  39147=>"111010001",
  39148=>"111010011",
  39149=>"001001110",
  39150=>"111001011",
  39151=>"111010011",
  39152=>"111000001",
  39153=>"111111111",
  39154=>"100111111",
  39155=>"101110000",
  39156=>"000100010",
  39157=>"111110101",
  39158=>"001101111",
  39159=>"011101011",
  39160=>"010110101",
  39161=>"110000111",
  39162=>"000011100",
  39163=>"011001101",
  39164=>"010001000",
  39165=>"110000000",
  39166=>"011101111",
  39167=>"001001000",
  39168=>"011010010",
  39169=>"101110001",
  39170=>"111101100",
  39171=>"010111001",
  39172=>"000110010",
  39173=>"110101111",
  39174=>"010111100",
  39175=>"100111011",
  39176=>"010011100",
  39177=>"011100101",
  39178=>"011100001",
  39179=>"101011000",
  39180=>"000010000",
  39181=>"100000101",
  39182=>"100101011",
  39183=>"100100010",
  39184=>"011101001",
  39185=>"000100100",
  39186=>"011000000",
  39187=>"001110101",
  39188=>"100100101",
  39189=>"100011011",
  39190=>"010010100",
  39191=>"001001100",
  39192=>"110100100",
  39193=>"100100111",
  39194=>"110010001",
  39195=>"011110010",
  39196=>"110100011",
  39197=>"001000010",
  39198=>"101000010",
  39199=>"000000100",
  39200=>"001100100",
  39201=>"100000101",
  39202=>"011111100",
  39203=>"100100101",
  39204=>"011000010",
  39205=>"101011001",
  39206=>"100110100",
  39207=>"000101010",
  39208=>"110001010",
  39209=>"110110110",
  39210=>"101010101",
  39211=>"010010010",
  39212=>"110010001",
  39213=>"110111100",
  39214=>"100000001",
  39215=>"011100001",
  39216=>"011011011",
  39217=>"101100000",
  39218=>"010011110",
  39219=>"110110110",
  39220=>"010111011",
  39221=>"010100000",
  39222=>"111111000",
  39223=>"110101011",
  39224=>"000010110",
  39225=>"111011000",
  39226=>"001010010",
  39227=>"000011100",
  39228=>"110011010",
  39229=>"100000110",
  39230=>"101010011",
  39231=>"001000110",
  39232=>"100011001",
  39233=>"011001010",
  39234=>"010011100",
  39235=>"100010110",
  39236=>"100100011",
  39237=>"111010110",
  39238=>"111111011",
  39239=>"111111010",
  39240=>"111010110",
  39241=>"010100001",
  39242=>"101111010",
  39243=>"001001110",
  39244=>"011010000",
  39245=>"100101100",
  39246=>"001011010",
  39247=>"010101000",
  39248=>"101110000",
  39249=>"100101110",
  39250=>"110000010",
  39251=>"000011111",
  39252=>"100010110",
  39253=>"011111111",
  39254=>"011010110",
  39255=>"111111111",
  39256=>"000100100",
  39257=>"100101010",
  39258=>"110101110",
  39259=>"111011110",
  39260=>"110000011",
  39261=>"111101010",
  39262=>"010100101",
  39263=>"111000100",
  39264=>"101100100",
  39265=>"110001001",
  39266=>"000011110",
  39267=>"010100001",
  39268=>"101110011",
  39269=>"011001000",
  39270=>"000001100",
  39271=>"011011100",
  39272=>"010110010",
  39273=>"000001100",
  39274=>"010100001",
  39275=>"010011011",
  39276=>"001001110",
  39277=>"001100101",
  39278=>"101111001",
  39279=>"100111111",
  39280=>"001111010",
  39281=>"100010010",
  39282=>"110110001",
  39283=>"111100011",
  39284=>"101111010",
  39285=>"001001110",
  39286=>"000110010",
  39287=>"100110110",
  39288=>"110000010",
  39289=>"101110001",
  39290=>"010100010",
  39291=>"111111101",
  39292=>"111001011",
  39293=>"111011110",
  39294=>"010110011",
  39295=>"100001001",
  39296=>"001111110",
  39297=>"000100100",
  39298=>"110000001",
  39299=>"001100111",
  39300=>"011111110",
  39301=>"000100111",
  39302=>"001101011",
  39303=>"101010100",
  39304=>"110111001",
  39305=>"001101010",
  39306=>"100110000",
  39307=>"101110111",
  39308=>"001010110",
  39309=>"110111011",
  39310=>"100000110",
  39311=>"001110110",
  39312=>"111011111",
  39313=>"111010011",
  39314=>"000110001",
  39315=>"011111101",
  39316=>"010100101",
  39317=>"100010001",
  39318=>"000011011",
  39319=>"101111101",
  39320=>"101001010",
  39321=>"011000111",
  39322=>"000001010",
  39323=>"111000100",
  39324=>"111001101",
  39325=>"111100011",
  39326=>"011110100",
  39327=>"111110111",
  39328=>"011010011",
  39329=>"100000000",
  39330=>"010000101",
  39331=>"011101111",
  39332=>"001111000",
  39333=>"100101000",
  39334=>"000110111",
  39335=>"000001100",
  39336=>"011100101",
  39337=>"100000000",
  39338=>"000011100",
  39339=>"010100111",
  39340=>"010111110",
  39341=>"001011001",
  39342=>"011001101",
  39343=>"001100000",
  39344=>"101111000",
  39345=>"100010001",
  39346=>"000000001",
  39347=>"100100101",
  39348=>"110011110",
  39349=>"010010000",
  39350=>"001010010",
  39351=>"010000010",
  39352=>"110011001",
  39353=>"000110010",
  39354=>"100110011",
  39355=>"000100101",
  39356=>"100011000",
  39357=>"000110001",
  39358=>"001111011",
  39359=>"010000010",
  39360=>"101001010",
  39361=>"111110010",
  39362=>"000001010",
  39363=>"011101001",
  39364=>"111010101",
  39365=>"010110100",
  39366=>"101111111",
  39367=>"011011010",
  39368=>"111001010",
  39369=>"110101110",
  39370=>"000100101",
  39371=>"111011001",
  39372=>"111001101",
  39373=>"010110101",
  39374=>"110100111",
  39375=>"000011011",
  39376=>"101001101",
  39377=>"010010011",
  39378=>"001011100",
  39379=>"000001000",
  39380=>"100010110",
  39381=>"011001111",
  39382=>"001100011",
  39383=>"011010100",
  39384=>"010010110",
  39385=>"101110111",
  39386=>"100000001",
  39387=>"101001000",
  39388=>"000001011",
  39389=>"110011111",
  39390=>"111000000",
  39391=>"101010100",
  39392=>"010101010",
  39393=>"110011011",
  39394=>"111110001",
  39395=>"110011010",
  39396=>"001011101",
  39397=>"000000100",
  39398=>"010000000",
  39399=>"011001010",
  39400=>"001110011",
  39401=>"111011101",
  39402=>"000110000",
  39403=>"001010101",
  39404=>"111101011",
  39405=>"101111001",
  39406=>"011001000",
  39407=>"000001110",
  39408=>"101010111",
  39409=>"110011100",
  39410=>"100000000",
  39411=>"000100110",
  39412=>"101111101",
  39413=>"001111100",
  39414=>"010101101",
  39415=>"000000011",
  39416=>"110000100",
  39417=>"100100001",
  39418=>"000100000",
  39419=>"010000000",
  39420=>"000110001",
  39421=>"110111111",
  39422=>"110001001",
  39423=>"110101000",
  39424=>"100111100",
  39425=>"011101111",
  39426=>"101111110",
  39427=>"010011001",
  39428=>"100101100",
  39429=>"001111111",
  39430=>"111011101",
  39431=>"101010010",
  39432=>"011011111",
  39433=>"000110100",
  39434=>"101111001",
  39435=>"010010011",
  39436=>"011001010",
  39437=>"111110111",
  39438=>"100001101",
  39439=>"111110010",
  39440=>"000000011",
  39441=>"011001110",
  39442=>"000001101",
  39443=>"011101110",
  39444=>"010111100",
  39445=>"111100000",
  39446=>"111100001",
  39447=>"000001001",
  39448=>"001010111",
  39449=>"111001011",
  39450=>"010010001",
  39451=>"010110010",
  39452=>"111010111",
  39453=>"010110100",
  39454=>"011111001",
  39455=>"011111010",
  39456=>"001111000",
  39457=>"001000101",
  39458=>"000011000",
  39459=>"111010111",
  39460=>"001010100",
  39461=>"011011001",
  39462=>"100010110",
  39463=>"011110000",
  39464=>"100000100",
  39465=>"000000000",
  39466=>"100001101",
  39467=>"011001100",
  39468=>"011001000",
  39469=>"111000010",
  39470=>"010110100",
  39471=>"101101000",
  39472=>"001101110",
  39473=>"101001101",
  39474=>"011001110",
  39475=>"101110001",
  39476=>"111010111",
  39477=>"001011100",
  39478=>"111000111",
  39479=>"100100001",
  39480=>"000011111",
  39481=>"111100101",
  39482=>"001101010",
  39483=>"010100001",
  39484=>"000100011",
  39485=>"110011011",
  39486=>"010010011",
  39487=>"000001011",
  39488=>"100010100",
  39489=>"001101000",
  39490=>"110011111",
  39491=>"011101111",
  39492=>"100010001",
  39493=>"110111101",
  39494=>"011000100",
  39495=>"110010111",
  39496=>"110110011",
  39497=>"100101110",
  39498=>"010101111",
  39499=>"100100111",
  39500=>"010010010",
  39501=>"000001001",
  39502=>"111110111",
  39503=>"110110100",
  39504=>"001001110",
  39505=>"010111111",
  39506=>"101001010",
  39507=>"101111110",
  39508=>"010011010",
  39509=>"111110111",
  39510=>"001011100",
  39511=>"100110110",
  39512=>"101111111",
  39513=>"111011011",
  39514=>"110000010",
  39515=>"010000000",
  39516=>"010011001",
  39517=>"001110100",
  39518=>"011100011",
  39519=>"001100111",
  39520=>"111000010",
  39521=>"010010110",
  39522=>"001111010",
  39523=>"101001011",
  39524=>"001010100",
  39525=>"111001000",
  39526=>"101010001",
  39527=>"111101111",
  39528=>"000010011",
  39529=>"111110001",
  39530=>"100100010",
  39531=>"100000111",
  39532=>"100100001",
  39533=>"100111110",
  39534=>"111011001",
  39535=>"011011101",
  39536=>"011101011",
  39537=>"000001000",
  39538=>"111100011",
  39539=>"100011010",
  39540=>"000011000",
  39541=>"011101011",
  39542=>"010011001",
  39543=>"001011111",
  39544=>"001010100",
  39545=>"010000101",
  39546=>"110110001",
  39547=>"011100101",
  39548=>"100011001",
  39549=>"000011111",
  39550=>"110111010",
  39551=>"101011101",
  39552=>"001010101",
  39553=>"110010000",
  39554=>"011000110",
  39555=>"100011001",
  39556=>"010000111",
  39557=>"011000001",
  39558=>"000001010",
  39559=>"001111101",
  39560=>"000010010",
  39561=>"101000010",
  39562=>"100001111",
  39563=>"000100010",
  39564=>"110000000",
  39565=>"010100010",
  39566=>"101000000",
  39567=>"010011111",
  39568=>"111000010",
  39569=>"111111100",
  39570=>"111011010",
  39571=>"100011000",
  39572=>"111001111",
  39573=>"111000101",
  39574=>"011111111",
  39575=>"001100100",
  39576=>"110011111",
  39577=>"100011000",
  39578=>"110100101",
  39579=>"111001000",
  39580=>"010111000",
  39581=>"101100101",
  39582=>"011111111",
  39583=>"100000000",
  39584=>"100001100",
  39585=>"000101101",
  39586=>"000010110",
  39587=>"100101001",
  39588=>"111111010",
  39589=>"000110101",
  39590=>"011010100",
  39591=>"010000100",
  39592=>"011010100",
  39593=>"101101100",
  39594=>"101100001",
  39595=>"100111010",
  39596=>"001100001",
  39597=>"111001000",
  39598=>"001010011",
  39599=>"110011000",
  39600=>"010010010",
  39601=>"111000111",
  39602=>"010010100",
  39603=>"101110010",
  39604=>"010011000",
  39605=>"011110000",
  39606=>"000000010",
  39607=>"010000010",
  39608=>"111110011",
  39609=>"111101011",
  39610=>"111001101",
  39611=>"110000101",
  39612=>"111101100",
  39613=>"011001110",
  39614=>"000011100",
  39615=>"110101101",
  39616=>"010111101",
  39617=>"010010000",
  39618=>"010010111",
  39619=>"011011101",
  39620=>"011111000",
  39621=>"010100010",
  39622=>"000011001",
  39623=>"110111001",
  39624=>"011000110",
  39625=>"000001110",
  39626=>"011010001",
  39627=>"011000000",
  39628=>"000011000",
  39629=>"101011110",
  39630=>"001010100",
  39631=>"000111011",
  39632=>"101101111",
  39633=>"001001011",
  39634=>"110110100",
  39635=>"110100110",
  39636=>"111101100",
  39637=>"001000110",
  39638=>"110101011",
  39639=>"001100100",
  39640=>"010011011",
  39641=>"101101100",
  39642=>"001000001",
  39643=>"010110000",
  39644=>"000101100",
  39645=>"000010001",
  39646=>"001110000",
  39647=>"010010010",
  39648=>"110110011",
  39649=>"000000000",
  39650=>"100100011",
  39651=>"100111110",
  39652=>"010010011",
  39653=>"100101000",
  39654=>"001011011",
  39655=>"010111100",
  39656=>"101001111",
  39657=>"111100100",
  39658=>"111000100",
  39659=>"100001101",
  39660=>"000011010",
  39661=>"011100011",
  39662=>"010101000",
  39663=>"111011101",
  39664=>"100111000",
  39665=>"110001110",
  39666=>"010111001",
  39667=>"001110101",
  39668=>"110100010",
  39669=>"101001111",
  39670=>"101001111",
  39671=>"011100001",
  39672=>"110100100",
  39673=>"100011001",
  39674=>"101001000",
  39675=>"100001010",
  39676=>"111000110",
  39677=>"000000110",
  39678=>"000001011",
  39679=>"111111111",
  39680=>"000011000",
  39681=>"000110010",
  39682=>"011111110",
  39683=>"001100001",
  39684=>"010001000",
  39685=>"001001000",
  39686=>"011010011",
  39687=>"100000100",
  39688=>"010101001",
  39689=>"100101111",
  39690=>"101111001",
  39691=>"000101001",
  39692=>"111101101",
  39693=>"101001001",
  39694=>"100100011",
  39695=>"000011110",
  39696=>"011100011",
  39697=>"010011011",
  39698=>"011001001",
  39699=>"110011111",
  39700=>"010110111",
  39701=>"001001001",
  39702=>"101001001",
  39703=>"001100010",
  39704=>"010010110",
  39705=>"001000011",
  39706=>"000100111",
  39707=>"110100100",
  39708=>"101010001",
  39709=>"101100101",
  39710=>"110111011",
  39711=>"010110110",
  39712=>"000001110",
  39713=>"101000110",
  39714=>"011000111",
  39715=>"100001111",
  39716=>"001100011",
  39717=>"000110000",
  39718=>"000001110",
  39719=>"001010100",
  39720=>"010001100",
  39721=>"111101101",
  39722=>"011100001",
  39723=>"000101110",
  39724=>"110111001",
  39725=>"000010000",
  39726=>"011010010",
  39727=>"011010110",
  39728=>"001001111",
  39729=>"010101001",
  39730=>"010111010",
  39731=>"000010011",
  39732=>"100110111",
  39733=>"001110110",
  39734=>"010100011",
  39735=>"111000001",
  39736=>"010000110",
  39737=>"010000001",
  39738=>"101111010",
  39739=>"000110011",
  39740=>"111111001",
  39741=>"111101001",
  39742=>"111100001",
  39743=>"101011110",
  39744=>"011100001",
  39745=>"100000111",
  39746=>"111111011",
  39747=>"110001001",
  39748=>"111000100",
  39749=>"100000001",
  39750=>"111111111",
  39751=>"101010100",
  39752=>"011110100",
  39753=>"000100111",
  39754=>"001111010",
  39755=>"110000010",
  39756=>"010111011",
  39757=>"000111001",
  39758=>"010110111",
  39759=>"011000110",
  39760=>"110011110",
  39761=>"110001100",
  39762=>"000111101",
  39763=>"101010010",
  39764=>"111101001",
  39765=>"111110110",
  39766=>"010010110",
  39767=>"010011111",
  39768=>"010010010",
  39769=>"101111010",
  39770=>"010110101",
  39771=>"010010101",
  39772=>"111111100",
  39773=>"001110000",
  39774=>"010001000",
  39775=>"001011110",
  39776=>"101011111",
  39777=>"111011010",
  39778=>"101111100",
  39779=>"000110110",
  39780=>"101000001",
  39781=>"000001011",
  39782=>"011111001",
  39783=>"001010100",
  39784=>"010111001",
  39785=>"101010111",
  39786=>"000010100",
  39787=>"001010110",
  39788=>"000001100",
  39789=>"101111011",
  39790=>"100001110",
  39791=>"001011100",
  39792=>"001001100",
  39793=>"101110011",
  39794=>"111000111",
  39795=>"101100000",
  39796=>"000001010",
  39797=>"110111010",
  39798=>"010100111",
  39799=>"000001001",
  39800=>"011110110",
  39801=>"110101000",
  39802=>"101000110",
  39803=>"001111000",
  39804=>"111101011",
  39805=>"100111101",
  39806=>"101010011",
  39807=>"110011110",
  39808=>"011110100",
  39809=>"111001010",
  39810=>"011001010",
  39811=>"011001010",
  39812=>"011011100",
  39813=>"101110100",
  39814=>"001110011",
  39815=>"000011001",
  39816=>"110011000",
  39817=>"100101010",
  39818=>"110011100",
  39819=>"100000101",
  39820=>"000000111",
  39821=>"111110010",
  39822=>"110111101",
  39823=>"010001111",
  39824=>"000100011",
  39825=>"111111011",
  39826=>"010000110",
  39827=>"010111010",
  39828=>"100010011",
  39829=>"111100111",
  39830=>"101101000",
  39831=>"111000100",
  39832=>"001111001",
  39833=>"010010101",
  39834=>"001100000",
  39835=>"001101001",
  39836=>"111101100",
  39837=>"001100111",
  39838=>"000001101",
  39839=>"100111110",
  39840=>"010101101",
  39841=>"011111000",
  39842=>"100110101",
  39843=>"011101011",
  39844=>"100001001",
  39845=>"111101111",
  39846=>"000001100",
  39847=>"101110101",
  39848=>"000110111",
  39849=>"010011000",
  39850=>"000010000",
  39851=>"010001001",
  39852=>"010001101",
  39853=>"001101111",
  39854=>"010000000",
  39855=>"011101101",
  39856=>"101100101",
  39857=>"111011011",
  39858=>"001100000",
  39859=>"101110111",
  39860=>"001000110",
  39861=>"000011000",
  39862=>"110110100",
  39863=>"000100001",
  39864=>"111001100",
  39865=>"001110010",
  39866=>"000100101",
  39867=>"001101110",
  39868=>"110011110",
  39869=>"001010111",
  39870=>"000000001",
  39871=>"001001000",
  39872=>"001000000",
  39873=>"000001000",
  39874=>"010001101",
  39875=>"001101110",
  39876=>"111101001",
  39877=>"100100100",
  39878=>"011101110",
  39879=>"100110110",
  39880=>"011111000",
  39881=>"010011011",
  39882=>"101110111",
  39883=>"100010111",
  39884=>"001010100",
  39885=>"100100000",
  39886=>"111000101",
  39887=>"100011000",
  39888=>"001100111",
  39889=>"101000100",
  39890=>"100111100",
  39891=>"010111101",
  39892=>"010111110",
  39893=>"011011111",
  39894=>"001111110",
  39895=>"001100000",
  39896=>"011010101",
  39897=>"010111110",
  39898=>"111010100",
  39899=>"011010010",
  39900=>"010111111",
  39901=>"011100011",
  39902=>"110000111",
  39903=>"011000010",
  39904=>"111001110",
  39905=>"101110010",
  39906=>"010000111",
  39907=>"100110100",
  39908=>"011011000",
  39909=>"111101101",
  39910=>"011110011",
  39911=>"001111001",
  39912=>"010010110",
  39913=>"001101100",
  39914=>"100011000",
  39915=>"001111001",
  39916=>"110010101",
  39917=>"100010000",
  39918=>"000111001",
  39919=>"011101101",
  39920=>"001011000",
  39921=>"111110101",
  39922=>"110101101",
  39923=>"001100001",
  39924=>"110001110",
  39925=>"010110100",
  39926=>"000000111",
  39927=>"010101001",
  39928=>"101110001",
  39929=>"010100100",
  39930=>"000001001",
  39931=>"000110001",
  39932=>"111011001",
  39933=>"001111011",
  39934=>"000100001",
  39935=>"110001100",
  39936=>"101010111",
  39937=>"100001000",
  39938=>"110110110",
  39939=>"011101100",
  39940=>"111100011",
  39941=>"000010101",
  39942=>"100000100",
  39943=>"101000101",
  39944=>"000011001",
  39945=>"000010111",
  39946=>"110111011",
  39947=>"011000100",
  39948=>"010000110",
  39949=>"110111111",
  39950=>"011001111",
  39951=>"001011101",
  39952=>"111111101",
  39953=>"101010011",
  39954=>"110001000",
  39955=>"110000001",
  39956=>"000101010",
  39957=>"110100010",
  39958=>"111000011",
  39959=>"100000000",
  39960=>"100001100",
  39961=>"101000101",
  39962=>"111101101",
  39963=>"011110111",
  39964=>"001110111",
  39965=>"000110010",
  39966=>"011010101",
  39967=>"011110101",
  39968=>"100000111",
  39969=>"101110011",
  39970=>"011010010",
  39971=>"101001101",
  39972=>"001011011",
  39973=>"110001011",
  39974=>"111101010",
  39975=>"101011101",
  39976=>"110110110",
  39977=>"100011110",
  39978=>"111100011",
  39979=>"010101111",
  39980=>"000100110",
  39981=>"001010001",
  39982=>"011010111",
  39983=>"110011011",
  39984=>"101011101",
  39985=>"000011111",
  39986=>"100011010",
  39987=>"001101101",
  39988=>"001001010",
  39989=>"100101011",
  39990=>"010101110",
  39991=>"100010011",
  39992=>"110010011",
  39993=>"111001111",
  39994=>"110101010",
  39995=>"100010000",
  39996=>"100000010",
  39997=>"011000101",
  39998=>"111101101",
  39999=>"110011011",
  40000=>"001000000",
  40001=>"111000000",
  40002=>"011000011",
  40003=>"111001001",
  40004=>"000111100",
  40005=>"111110011",
  40006=>"110110100",
  40007=>"100101101",
  40008=>"000101010",
  40009=>"101011110",
  40010=>"100110011",
  40011=>"001110010",
  40012=>"000111100",
  40013=>"111111000",
  40014=>"100011001",
  40015=>"000100000",
  40016=>"110001100",
  40017=>"001111000",
  40018=>"001110111",
  40019=>"110110001",
  40020=>"110001101",
  40021=>"101000000",
  40022=>"011011111",
  40023=>"001101001",
  40024=>"100001111",
  40025=>"010011011",
  40026=>"000000101",
  40027=>"100001110",
  40028=>"010010001",
  40029=>"010100101",
  40030=>"001011101",
  40031=>"100110010",
  40032=>"101000010",
  40033=>"111011000",
  40034=>"110100010",
  40035=>"001001010",
  40036=>"100111101",
  40037=>"001001011",
  40038=>"010000011",
  40039=>"011001010",
  40040=>"001111011",
  40041=>"110011101",
  40042=>"001100111",
  40043=>"000100001",
  40044=>"010001011",
  40045=>"001010101",
  40046=>"000000001",
  40047=>"101111000",
  40048=>"001110111",
  40049=>"100001100",
  40050=>"010011101",
  40051=>"101000001",
  40052=>"110110011",
  40053=>"100100011",
  40054=>"101000010",
  40055=>"011011001",
  40056=>"101100111",
  40057=>"000100110",
  40058=>"001001010",
  40059=>"111010000",
  40060=>"000000100",
  40061=>"111111111",
  40062=>"010110101",
  40063=>"001010100",
  40064=>"110000000",
  40065=>"011111100",
  40066=>"111101011",
  40067=>"101011110",
  40068=>"100000101",
  40069=>"110110001",
  40070=>"000010001",
  40071=>"111011010",
  40072=>"010000100",
  40073=>"011101001",
  40074=>"011100000",
  40075=>"110100011",
  40076=>"010011100",
  40077=>"101001000",
  40078=>"001101100",
  40079=>"000010001",
  40080=>"111010111",
  40081=>"111111001",
  40082=>"110001110",
  40083=>"000110101",
  40084=>"101101001",
  40085=>"011111011",
  40086=>"100001000",
  40087=>"111101001",
  40088=>"110111010",
  40089=>"011000100",
  40090=>"111111101",
  40091=>"101010101",
  40092=>"111110101",
  40093=>"110000101",
  40094=>"011100111",
  40095=>"100110010",
  40096=>"000001110",
  40097=>"110110110",
  40098=>"100110100",
  40099=>"110110011",
  40100=>"111000010",
  40101=>"001101111",
  40102=>"000101101",
  40103=>"110111010",
  40104=>"101110000",
  40105=>"110001000",
  40106=>"001010110",
  40107=>"011001010",
  40108=>"001101111",
  40109=>"100110101",
  40110=>"110010101",
  40111=>"100011010",
  40112=>"001000011",
  40113=>"000011110",
  40114=>"100101000",
  40115=>"111100001",
  40116=>"100111110",
  40117=>"011100000",
  40118=>"100110110",
  40119=>"000100010",
  40120=>"011010011",
  40121=>"010010100",
  40122=>"101110000",
  40123=>"001010000",
  40124=>"110100101",
  40125=>"000011110",
  40126=>"111010000",
  40127=>"111010011",
  40128=>"111000010",
  40129=>"101101000",
  40130=>"001100111",
  40131=>"010101100",
  40132=>"111110010",
  40133=>"001110010",
  40134=>"000110001",
  40135=>"111001000",
  40136=>"011100010",
  40137=>"101111000",
  40138=>"000000100",
  40139=>"111101111",
  40140=>"101111110",
  40141=>"010000100",
  40142=>"101101001",
  40143=>"110011010",
  40144=>"110000011",
  40145=>"100111011",
  40146=>"101011001",
  40147=>"011110011",
  40148=>"000001110",
  40149=>"010010010",
  40150=>"001111110",
  40151=>"110111110",
  40152=>"101101110",
  40153=>"111010101",
  40154=>"101111000",
  40155=>"001011010",
  40156=>"101100001",
  40157=>"100111111",
  40158=>"010010000",
  40159=>"100010111",
  40160=>"000101001",
  40161=>"110000000",
  40162=>"110010010",
  40163=>"101000000",
  40164=>"111110110",
  40165=>"101100001",
  40166=>"011101110",
  40167=>"111010101",
  40168=>"001101010",
  40169=>"110001010",
  40170=>"100010001",
  40171=>"110011101",
  40172=>"101110001",
  40173=>"101001011",
  40174=>"001011100",
  40175=>"011100010",
  40176=>"010111010",
  40177=>"000101010",
  40178=>"101110011",
  40179=>"000100100",
  40180=>"000110011",
  40181=>"111010001",
  40182=>"111000110",
  40183=>"001010011",
  40184=>"111010101",
  40185=>"100111101",
  40186=>"111010110",
  40187=>"111100001",
  40188=>"001000001",
  40189=>"011000110",
  40190=>"000100011",
  40191=>"000011001",
  40192=>"110001100",
  40193=>"011110000",
  40194=>"000110100",
  40195=>"110111111",
  40196=>"010100101",
  40197=>"110100100",
  40198=>"000111000",
  40199=>"111110001",
  40200=>"011000001",
  40201=>"101110011",
  40202=>"010010111",
  40203=>"110001000",
  40204=>"011000100",
  40205=>"000111011",
  40206=>"110001010",
  40207=>"010001000",
  40208=>"110011011",
  40209=>"111110100",
  40210=>"100000111",
  40211=>"001000001",
  40212=>"000101011",
  40213=>"011110110",
  40214=>"100000010",
  40215=>"011101011",
  40216=>"110001001",
  40217=>"010110111",
  40218=>"011100000",
  40219=>"100010100",
  40220=>"000010001",
  40221=>"101100011",
  40222=>"101111011",
  40223=>"001110101",
  40224=>"010000101",
  40225=>"111111010",
  40226=>"010111101",
  40227=>"101100100",
  40228=>"000101000",
  40229=>"110011111",
  40230=>"001010000",
  40231=>"111100010",
  40232=>"101011001",
  40233=>"010010100",
  40234=>"001011010",
  40235=>"110010110",
  40236=>"000011011",
  40237=>"001011101",
  40238=>"100100000",
  40239=>"001110110",
  40240=>"011000100",
  40241=>"111101100",
  40242=>"100111100",
  40243=>"001001011",
  40244=>"000101000",
  40245=>"010011110",
  40246=>"111101100",
  40247=>"001111010",
  40248=>"011010010",
  40249=>"100001111",
  40250=>"000010010",
  40251=>"111111111",
  40252=>"000101101",
  40253=>"110001001",
  40254=>"100110101",
  40255=>"101010100",
  40256=>"011001001",
  40257=>"110100100",
  40258=>"011010110",
  40259=>"010010101",
  40260=>"101001011",
  40261=>"110011010",
  40262=>"010001000",
  40263=>"101001001",
  40264=>"001001000",
  40265=>"100010000",
  40266=>"010101010",
  40267=>"001000110",
  40268=>"111010101",
  40269=>"100011100",
  40270=>"000110111",
  40271=>"111101010",
  40272=>"100001001",
  40273=>"001111100",
  40274=>"110110001",
  40275=>"110100010",
  40276=>"001001110",
  40277=>"001101011",
  40278=>"101011011",
  40279=>"110101011",
  40280=>"001010010",
  40281=>"100010011",
  40282=>"101011101",
  40283=>"010001011",
  40284=>"010111110",
  40285=>"000110111",
  40286=>"000110000",
  40287=>"001101101",
  40288=>"010111111",
  40289=>"101110101",
  40290=>"101000111",
  40291=>"101000010",
  40292=>"100001010",
  40293=>"011011010",
  40294=>"001111000",
  40295=>"101010110",
  40296=>"001000101",
  40297=>"110101111",
  40298=>"001000011",
  40299=>"000000001",
  40300=>"100010100",
  40301=>"101100011",
  40302=>"110000110",
  40303=>"011000111",
  40304=>"111111100",
  40305=>"011101010",
  40306=>"111101111",
  40307=>"001011111",
  40308=>"000000001",
  40309=>"101111101",
  40310=>"000000001",
  40311=>"110010001",
  40312=>"001101001",
  40313=>"011010000",
  40314=>"101000000",
  40315=>"111101101",
  40316=>"000111101",
  40317=>"101010111",
  40318=>"000101011",
  40319=>"100111110",
  40320=>"100001000",
  40321=>"010001011",
  40322=>"011101101",
  40323=>"010100010",
  40324=>"101011011",
  40325=>"100101100",
  40326=>"000010001",
  40327=>"100110010",
  40328=>"100000001",
  40329=>"011001010",
  40330=>"010100000",
  40331=>"110101100",
  40332=>"110010011",
  40333=>"100100000",
  40334=>"101010011",
  40335=>"001001111",
  40336=>"111011011",
  40337=>"010110010",
  40338=>"100100111",
  40339=>"111001110",
  40340=>"000011110",
  40341=>"101010011",
  40342=>"101110001",
  40343=>"010101111",
  40344=>"000000001",
  40345=>"100001111",
  40346=>"000101110",
  40347=>"001101101",
  40348=>"010101011",
  40349=>"011111110",
  40350=>"111010111",
  40351=>"111111111",
  40352=>"011000110",
  40353=>"110111010",
  40354=>"110001101",
  40355=>"010000110",
  40356=>"010001001",
  40357=>"011100001",
  40358=>"011101110",
  40359=>"001000011",
  40360=>"011000100",
  40361=>"100100101",
  40362=>"101100000",
  40363=>"110011011",
  40364=>"010110001",
  40365=>"001001010",
  40366=>"101010001",
  40367=>"001010000",
  40368=>"100010001",
  40369=>"111000001",
  40370=>"110101000",
  40371=>"011000101",
  40372=>"000000101",
  40373=>"011101001",
  40374=>"111010110",
  40375=>"001111010",
  40376=>"110010111",
  40377=>"111010011",
  40378=>"010110001",
  40379=>"010100011",
  40380=>"110001001",
  40381=>"000011000",
  40382=>"001100001",
  40383=>"000111010",
  40384=>"010001000",
  40385=>"111111110",
  40386=>"010101000",
  40387=>"000000110",
  40388=>"000011011",
  40389=>"111011011",
  40390=>"011001100",
  40391=>"011100100",
  40392=>"100101001",
  40393=>"110110100",
  40394=>"111111111",
  40395=>"110011001",
  40396=>"011111001",
  40397=>"101111001",
  40398=>"110110111",
  40399=>"000101110",
  40400=>"001011101",
  40401=>"010011101",
  40402=>"010110011",
  40403=>"111101100",
  40404=>"010100101",
  40405=>"100001101",
  40406=>"001100000",
  40407=>"110100010",
  40408=>"110001011",
  40409=>"010010101",
  40410=>"010110010",
  40411=>"011011110",
  40412=>"100011111",
  40413=>"011101110",
  40414=>"100110111",
  40415=>"111100111",
  40416=>"101001001",
  40417=>"110111011",
  40418=>"111100101",
  40419=>"100011000",
  40420=>"000100011",
  40421=>"100100011",
  40422=>"001001111",
  40423=>"101001001",
  40424=>"101000010",
  40425=>"010101010",
  40426=>"010110011",
  40427=>"001100110",
  40428=>"111011000",
  40429=>"010111101",
  40430=>"011010010",
  40431=>"001001000",
  40432=>"111011000",
  40433=>"001101100",
  40434=>"111110110",
  40435=>"001100100",
  40436=>"110011011",
  40437=>"101011010",
  40438=>"001110010",
  40439=>"110101110",
  40440=>"110011110",
  40441=>"011010010",
  40442=>"001011100",
  40443=>"001110011",
  40444=>"111101001",
  40445=>"011001010",
  40446=>"111000101",
  40447=>"000000010",
  40448=>"001011100",
  40449=>"110001101",
  40450=>"101000001",
  40451=>"010000000",
  40452=>"110001000",
  40453=>"111110101",
  40454=>"110010100",
  40455=>"001000100",
  40456=>"100100000",
  40457=>"010010001",
  40458=>"111101110",
  40459=>"111001000",
  40460=>"010100010",
  40461=>"110000100",
  40462=>"110100001",
  40463=>"001011101",
  40464=>"011101101",
  40465=>"011111000",
  40466=>"111111100",
  40467=>"000110000",
  40468=>"101101100",
  40469=>"011010110",
  40470=>"001000101",
  40471=>"110010100",
  40472=>"011000110",
  40473=>"000011111",
  40474=>"001100010",
  40475=>"000010100",
  40476=>"010111100",
  40477=>"001101101",
  40478=>"001001111",
  40479=>"101010010",
  40480=>"111111111",
  40481=>"010110001",
  40482=>"010111011",
  40483=>"100011111",
  40484=>"101000000",
  40485=>"000010010",
  40486=>"101110100",
  40487=>"111101010",
  40488=>"110101011",
  40489=>"111111100",
  40490=>"111100101",
  40491=>"000001111",
  40492=>"101111111",
  40493=>"000111011",
  40494=>"101010000",
  40495=>"010100100",
  40496=>"011001001",
  40497=>"101111000",
  40498=>"100110011",
  40499=>"001011110",
  40500=>"110010100",
  40501=>"010111011",
  40502=>"101110011",
  40503=>"110110111",
  40504=>"001010101",
  40505=>"111010001",
  40506=>"001101100",
  40507=>"101100011",
  40508=>"110000000",
  40509=>"101000010",
  40510=>"010010001",
  40511=>"011110100",
  40512=>"011101010",
  40513=>"110111111",
  40514=>"110110011",
  40515=>"001110011",
  40516=>"000011010",
  40517=>"010011001",
  40518=>"000011100",
  40519=>"011101000",
  40520=>"010101101",
  40521=>"011001000",
  40522=>"001001011",
  40523=>"000100100",
  40524=>"000000110",
  40525=>"010010101",
  40526=>"001001011",
  40527=>"110110111",
  40528=>"110010101",
  40529=>"010000000",
  40530=>"110101100",
  40531=>"010110000",
  40532=>"010100010",
  40533=>"111001000",
  40534=>"010110010",
  40535=>"010110111",
  40536=>"110011010",
  40537=>"110000010",
  40538=>"001111001",
  40539=>"100001100",
  40540=>"100100011",
  40541=>"001111100",
  40542=>"011000110",
  40543=>"001000011",
  40544=>"101011000",
  40545=>"111001000",
  40546=>"110011111",
  40547=>"011001111",
  40548=>"111011101",
  40549=>"111000000",
  40550=>"001110100",
  40551=>"011110111",
  40552=>"011100011",
  40553=>"100001000",
  40554=>"110000001",
  40555=>"010011010",
  40556=>"101110100",
  40557=>"011101001",
  40558=>"000011101",
  40559=>"000101010",
  40560=>"010111111",
  40561=>"110111011",
  40562=>"101100011",
  40563=>"000111001",
  40564=>"110110111",
  40565=>"011110001",
  40566=>"111001010",
  40567=>"001001011",
  40568=>"000000010",
  40569=>"001011111",
  40570=>"010101111",
  40571=>"111000110",
  40572=>"000100111",
  40573=>"001010011",
  40574=>"001111000",
  40575=>"111100000",
  40576=>"000010110",
  40577=>"001100110",
  40578=>"100110111",
  40579=>"100010101",
  40580=>"111110101",
  40581=>"100011000",
  40582=>"101000000",
  40583=>"111110000",
  40584=>"111010011",
  40585=>"100110100",
  40586=>"111110001",
  40587=>"001011111",
  40588=>"000000100",
  40589=>"111100011",
  40590=>"011100100",
  40591=>"111110110",
  40592=>"000110010",
  40593=>"101001001",
  40594=>"110101010",
  40595=>"011110100",
  40596=>"111001010",
  40597=>"101111000",
  40598=>"110000000",
  40599=>"001000001",
  40600=>"010101010",
  40601=>"011010000",
  40602=>"000100111",
  40603=>"110011100",
  40604=>"010100001",
  40605=>"110010111",
  40606=>"000100000",
  40607=>"001011101",
  40608=>"111110000",
  40609=>"110110111",
  40610=>"001000010",
  40611=>"111001010",
  40612=>"100000001",
  40613=>"101001010",
  40614=>"011000111",
  40615=>"010110011",
  40616=>"111001001",
  40617=>"110110101",
  40618=>"001011110",
  40619=>"010101111",
  40620=>"010011111",
  40621=>"010000100",
  40622=>"001100111",
  40623=>"100010101",
  40624=>"000000010",
  40625=>"100100010",
  40626=>"110011011",
  40627=>"001111010",
  40628=>"000001111",
  40629=>"001111110",
  40630=>"110001100",
  40631=>"101011001",
  40632=>"011011100",
  40633=>"101111011",
  40634=>"101000101",
  40635=>"011011110",
  40636=>"001001000",
  40637=>"000101001",
  40638=>"010001000",
  40639=>"100011100",
  40640=>"100001001",
  40641=>"100111100",
  40642=>"001101100",
  40643=>"000101111",
  40644=>"110011011",
  40645=>"001110000",
  40646=>"100010001",
  40647=>"110101111",
  40648=>"110000110",
  40649=>"110001000",
  40650=>"010111111",
  40651=>"110000000",
  40652=>"101101000",
  40653=>"011111010",
  40654=>"110100011",
  40655=>"011110100",
  40656=>"011000010",
  40657=>"111110110",
  40658=>"111001110",
  40659=>"100010100",
  40660=>"000000011",
  40661=>"000100100",
  40662=>"001000100",
  40663=>"011000101",
  40664=>"000100000",
  40665=>"111111011",
  40666=>"110010100",
  40667=>"010010000",
  40668=>"110100111",
  40669=>"011010111",
  40670=>"111101010",
  40671=>"111000011",
  40672=>"000010101",
  40673=>"011011101",
  40674=>"110100000",
  40675=>"111000101",
  40676=>"100101111",
  40677=>"010001111",
  40678=>"110111101",
  40679=>"010011001",
  40680=>"111110100",
  40681=>"001001101",
  40682=>"001100000",
  40683=>"110100000",
  40684=>"000001000",
  40685=>"100010001",
  40686=>"110001111",
  40687=>"011010001",
  40688=>"001000011",
  40689=>"110001011",
  40690=>"111110110",
  40691=>"100001101",
  40692=>"011110111",
  40693=>"100100001",
  40694=>"010010111",
  40695=>"110010011",
  40696=>"111000100",
  40697=>"100010101",
  40698=>"001010100",
  40699=>"100111000",
  40700=>"010101110",
  40701=>"111001100",
  40702=>"001111111",
  40703=>"111001111",
  40704=>"001100010",
  40705=>"101011111",
  40706=>"110010010",
  40707=>"001000011",
  40708=>"001111101",
  40709=>"011000111",
  40710=>"010101111",
  40711=>"111001001",
  40712=>"101111101",
  40713=>"101111001",
  40714=>"111111001",
  40715=>"000001101",
  40716=>"011010011",
  40717=>"110110001",
  40718=>"010101000",
  40719=>"101101010",
  40720=>"010010001",
  40721=>"000000100",
  40722=>"111011100",
  40723=>"100010010",
  40724=>"001111001",
  40725=>"001011110",
  40726=>"111110111",
  40727=>"111011110",
  40728=>"100000000",
  40729=>"111000111",
  40730=>"100111001",
  40731=>"011111111",
  40732=>"001110010",
  40733=>"011010000",
  40734=>"100111101",
  40735=>"111110100",
  40736=>"110111110",
  40737=>"100101010",
  40738=>"110111111",
  40739=>"100111111",
  40740=>"111011101",
  40741=>"000000110",
  40742=>"110000100",
  40743=>"100001100",
  40744=>"011000101",
  40745=>"001101110",
  40746=>"000110100",
  40747=>"011001001",
  40748=>"010100111",
  40749=>"000000000",
  40750=>"100010100",
  40751=>"000101101",
  40752=>"011111101",
  40753=>"011100111",
  40754=>"101010111",
  40755=>"101111011",
  40756=>"011101011",
  40757=>"000001001",
  40758=>"000101111",
  40759=>"010000110",
  40760=>"000001111",
  40761=>"000111001",
  40762=>"100110001",
  40763=>"110100001",
  40764=>"101101000",
  40765=>"100100010",
  40766=>"000110101",
  40767=>"110010101",
  40768=>"111000000",
  40769=>"001101000",
  40770=>"111010001",
  40771=>"111010111",
  40772=>"011001100",
  40773=>"100011100",
  40774=>"111000100",
  40775=>"101001101",
  40776=>"000101111",
  40777=>"101010100",
  40778=>"011111010",
  40779=>"101100110",
  40780=>"011110110",
  40781=>"110011100",
  40782=>"110100101",
  40783=>"000100111",
  40784=>"101110000",
  40785=>"111011010",
  40786=>"100110010",
  40787=>"101001001",
  40788=>"101101101",
  40789=>"011010101",
  40790=>"001010000",
  40791=>"110000000",
  40792=>"111000001",
  40793=>"100010010",
  40794=>"011010100",
  40795=>"001100010",
  40796=>"111100111",
  40797=>"010110000",
  40798=>"111001110",
  40799=>"000011000",
  40800=>"011001010",
  40801=>"000001101",
  40802=>"010110101",
  40803=>"000010010",
  40804=>"100111111",
  40805=>"110000111",
  40806=>"001010011",
  40807=>"101111000",
  40808=>"110101110",
  40809=>"111100101",
  40810=>"111101011",
  40811=>"100110110",
  40812=>"110110100",
  40813=>"001010000",
  40814=>"110110100",
  40815=>"111000011",
  40816=>"000000100",
  40817=>"011000111",
  40818=>"101001001",
  40819=>"011010000",
  40820=>"101110001",
  40821=>"111000000",
  40822=>"011000000",
  40823=>"111100101",
  40824=>"011100011",
  40825=>"000110000",
  40826=>"001110011",
  40827=>"001010001",
  40828=>"010001011",
  40829=>"101111001",
  40830=>"010010101",
  40831=>"010101111",
  40832=>"111111001",
  40833=>"010101101",
  40834=>"100001111",
  40835=>"111011101",
  40836=>"110110011",
  40837=>"001110100",
  40838=>"110000111",
  40839=>"000001101",
  40840=>"101111111",
  40841=>"111111001",
  40842=>"000011011",
  40843=>"001110011",
  40844=>"110101011",
  40845=>"011010011",
  40846=>"100101001",
  40847=>"100101101",
  40848=>"000000100",
  40849=>"100111011",
  40850=>"110000100",
  40851=>"001011110",
  40852=>"001100011",
  40853=>"100110101",
  40854=>"001000011",
  40855=>"011000011",
  40856=>"000010110",
  40857=>"001011010",
  40858=>"101000111",
  40859=>"111000100",
  40860=>"111111110",
  40861=>"011001000",
  40862=>"011000000",
  40863=>"111011011",
  40864=>"100101110",
  40865=>"110100101",
  40866=>"110010000",
  40867=>"001101110",
  40868=>"111001101",
  40869=>"100100011",
  40870=>"101110110",
  40871=>"000111010",
  40872=>"000111010",
  40873=>"011100111",
  40874=>"100001000",
  40875=>"011011011",
  40876=>"110110110",
  40877=>"110111111",
  40878=>"001000100",
  40879=>"001001100",
  40880=>"110001000",
  40881=>"111111100",
  40882=>"010001110",
  40883=>"000110111",
  40884=>"101111111",
  40885=>"101100101",
  40886=>"100000001",
  40887=>"011101111",
  40888=>"001111001",
  40889=>"101100001",
  40890=>"011000111",
  40891=>"111111111",
  40892=>"110011010",
  40893=>"010110000",
  40894=>"101011111",
  40895=>"100110001",
  40896=>"001010100",
  40897=>"110000110",
  40898=>"111110100",
  40899=>"100101000",
  40900=>"001110101",
  40901=>"111010101",
  40902=>"011011100",
  40903=>"011111011",
  40904=>"100101000",
  40905=>"000000111",
  40906=>"101100000",
  40907=>"101101101",
  40908=>"110100001",
  40909=>"100010000",
  40910=>"110010010",
  40911=>"010111010",
  40912=>"010111010",
  40913=>"101000111",
  40914=>"101001100",
  40915=>"000100111",
  40916=>"111110111",
  40917=>"010100111",
  40918=>"001111100",
  40919=>"001110110",
  40920=>"100001000",
  40921=>"100000111",
  40922=>"000110110",
  40923=>"011001010",
  40924=>"011111110",
  40925=>"101101100",
  40926=>"100101010",
  40927=>"101101110",
  40928=>"001010010",
  40929=>"100100101",
  40930=>"111111101",
  40931=>"010010010",
  40932=>"101010100",
  40933=>"100110010",
  40934=>"100010001",
  40935=>"111011011",
  40936=>"010110101",
  40937=>"111000001",
  40938=>"111001010",
  40939=>"110011100",
  40940=>"111110110",
  40941=>"111110111",
  40942=>"010110101",
  40943=>"110010011",
  40944=>"001100001",
  40945=>"010100011",
  40946=>"111000100",
  40947=>"111010100",
  40948=>"000110010",
  40949=>"010100111",
  40950=>"000111011",
  40951=>"011110001",
  40952=>"000001101",
  40953=>"001001001",
  40954=>"001111101",
  40955=>"101110000",
  40956=>"111100101",
  40957=>"111011111",
  40958=>"100101011",
  40959=>"100001011",
  40960=>"000101111",
  40961=>"000001011",
  40962=>"001011010",
  40963=>"011010000",
  40964=>"101111110",
  40965=>"111101100",
  40966=>"010011001",
  40967=>"101011010",
  40968=>"110101110",
  40969=>"110000111",
  40970=>"011010100",
  40971=>"001110110",
  40972=>"101001100",
  40973=>"011011010",
  40974=>"100110000",
  40975=>"011100110",
  40976=>"011100011",
  40977=>"001010001",
  40978=>"111111011",
  40979=>"000010101",
  40980=>"010011100",
  40981=>"110010011",
  40982=>"001110111",
  40983=>"010111000",
  40984=>"101111100",
  40985=>"110100110",
  40986=>"111110110",
  40987=>"111000100",
  40988=>"111010110",
  40989=>"011011001",
  40990=>"100101100",
  40991=>"000000100",
  40992=>"100111110",
  40993=>"101010010",
  40994=>"011011101",
  40995=>"110110111",
  40996=>"101100101",
  40997=>"100001101",
  40998=>"001011110",
  40999=>"011100111",
  41000=>"110100001",
  41001=>"000110111",
  41002=>"111010110",
  41003=>"111011110",
  41004=>"101001000",
  41005=>"010010110",
  41006=>"001101111",
  41007=>"111011101",
  41008=>"010111000",
  41009=>"010000010",
  41010=>"101000100",
  41011=>"000000001",
  41012=>"001001000",
  41013=>"101010000",
  41014=>"101101000",
  41015=>"010010001",
  41016=>"001001100",
  41017=>"111111001",
  41018=>"000100110",
  41019=>"011011111",
  41020=>"000100010",
  41021=>"101100100",
  41022=>"010100001",
  41023=>"011011010",
  41024=>"011100000",
  41025=>"011000110",
  41026=>"001100000",
  41027=>"011001000",
  41028=>"111110110",
  41029=>"110010101",
  41030=>"010110100",
  41031=>"000010000",
  41032=>"010111110",
  41033=>"011011010",
  41034=>"110101010",
  41035=>"011111100",
  41036=>"000100000",
  41037=>"001011101",
  41038=>"000111101",
  41039=>"100011110",
  41040=>"100000111",
  41041=>"110110111",
  41042=>"110100000",
  41043=>"111011010",
  41044=>"111111111",
  41045=>"110111100",
  41046=>"001001111",
  41047=>"000000000",
  41048=>"001000010",
  41049=>"111000001",
  41050=>"101110110",
  41051=>"101000010",
  41052=>"000000010",
  41053=>"101101011",
  41054=>"000100111",
  41055=>"100001000",
  41056=>"110110000",
  41057=>"111100110",
  41058=>"100100000",
  41059=>"010000001",
  41060=>"000001010",
  41061=>"111000010",
  41062=>"101001101",
  41063=>"000000010",
  41064=>"000001001",
  41065=>"001101101",
  41066=>"100000000",
  41067=>"110111111",
  41068=>"011000000",
  41069=>"110101000",
  41070=>"111000011",
  41071=>"010100101",
  41072=>"001000001",
  41073=>"000000101",
  41074=>"010010010",
  41075=>"111000111",
  41076=>"011010110",
  41077=>"100000000",
  41078=>"110010101",
  41079=>"110000101",
  41080=>"011100100",
  41081=>"000010110",
  41082=>"010101101",
  41083=>"000001101",
  41084=>"100010100",
  41085=>"110111001",
  41086=>"101101110",
  41087=>"101000101",
  41088=>"000001001",
  41089=>"100000011",
  41090=>"110101010",
  41091=>"111110110",
  41092=>"100011000",
  41093=>"100101000",
  41094=>"010001011",
  41095=>"000101100",
  41096=>"110111101",
  41097=>"001100111",
  41098=>"001000100",
  41099=>"111001110",
  41100=>"000011000",
  41101=>"100100111",
  41102=>"110000111",
  41103=>"001000100",
  41104=>"100110111",
  41105=>"100110010",
  41106=>"110101011",
  41107=>"100100110",
  41108=>"111101001",
  41109=>"001100010",
  41110=>"100010100",
  41111=>"011000100",
  41112=>"100111011",
  41113=>"111110100",
  41114=>"011010111",
  41115=>"011000111",
  41116=>"100110010",
  41117=>"011101110",
  41118=>"101111110",
  41119=>"110010110",
  41120=>"001000110",
  41121=>"101111110",
  41122=>"110100011",
  41123=>"101101000",
  41124=>"001110101",
  41125=>"101010100",
  41126=>"101111010",
  41127=>"111101100",
  41128=>"100110001",
  41129=>"110111001",
  41130=>"110100100",
  41131=>"001011011",
  41132=>"001000101",
  41133=>"110010111",
  41134=>"001011011",
  41135=>"111101000",
  41136=>"000001000",
  41137=>"110100010",
  41138=>"010010111",
  41139=>"110110100",
  41140=>"101100101",
  41141=>"110010110",
  41142=>"011101111",
  41143=>"001100100",
  41144=>"100001001",
  41145=>"110110100",
  41146=>"001100010",
  41147=>"001000110",
  41148=>"111100001",
  41149=>"000010001",
  41150=>"110101011",
  41151=>"000100111",
  41152=>"111110101",
  41153=>"001110111",
  41154=>"010010001",
  41155=>"011000000",
  41156=>"100001000",
  41157=>"011100000",
  41158=>"011101100",
  41159=>"000010101",
  41160=>"111010111",
  41161=>"000101000",
  41162=>"111111001",
  41163=>"001011110",
  41164=>"010000000",
  41165=>"010110110",
  41166=>"000100101",
  41167=>"010110110",
  41168=>"000001011",
  41169=>"010001110",
  41170=>"100111101",
  41171=>"110101110",
  41172=>"011001000",
  41173=>"000001110",
  41174=>"000100000",
  41175=>"000000011",
  41176=>"101001110",
  41177=>"101101100",
  41178=>"010000111",
  41179=>"010110001",
  41180=>"000001010",
  41181=>"010010011",
  41182=>"000000010",
  41183=>"001100010",
  41184=>"000000110",
  41185=>"110101110",
  41186=>"011010000",
  41187=>"000100100",
  41188=>"110111000",
  41189=>"001000111",
  41190=>"100100110",
  41191=>"011100110",
  41192=>"000101101",
  41193=>"101111010",
  41194=>"100101010",
  41195=>"001011110",
  41196=>"101101011",
  41197=>"100100010",
  41198=>"100111101",
  41199=>"110110000",
  41200=>"011101001",
  41201=>"001110011",
  41202=>"100000101",
  41203=>"010111011",
  41204=>"110010010",
  41205=>"110011010",
  41206=>"100010000",
  41207=>"100100111",
  41208=>"000010010",
  41209=>"101010110",
  41210=>"100000011",
  41211=>"010010000",
  41212=>"100100100",
  41213=>"010010100",
  41214=>"000110100",
  41215=>"110001111",
  41216=>"111001011",
  41217=>"101100110",
  41218=>"010000010",
  41219=>"100000001",
  41220=>"000110011",
  41221=>"111111111",
  41222=>"100000011",
  41223=>"111110010",
  41224=>"011100110",
  41225=>"100011111",
  41226=>"000111011",
  41227=>"000111001",
  41228=>"100000110",
  41229=>"101000101",
  41230=>"110101111",
  41231=>"000101001",
  41232=>"010010001",
  41233=>"110000110",
  41234=>"000100000",
  41235=>"111111110",
  41236=>"101010011",
  41237=>"100011110",
  41238=>"010111011",
  41239=>"100110111",
  41240=>"001000010",
  41241=>"011011000",
  41242=>"010100001",
  41243=>"011100100",
  41244=>"110111010",
  41245=>"011111110",
  41246=>"110010011",
  41247=>"001010011",
  41248=>"001000110",
  41249=>"000011101",
  41250=>"100000010",
  41251=>"001000000",
  41252=>"111100110",
  41253=>"111011110",
  41254=>"011100110",
  41255=>"111101101",
  41256=>"011010111",
  41257=>"111111111",
  41258=>"100011110",
  41259=>"010010101",
  41260=>"001011010",
  41261=>"110111111",
  41262=>"000000011",
  41263=>"011000100",
  41264=>"100101010",
  41265=>"101100101",
  41266=>"000010000",
  41267=>"010111111",
  41268=>"000011011",
  41269=>"101110110",
  41270=>"110010101",
  41271=>"011011100",
  41272=>"001011101",
  41273=>"010001000",
  41274=>"100111111",
  41275=>"100111110",
  41276=>"101010000",
  41277=>"111101101",
  41278=>"110101100",
  41279=>"001110010",
  41280=>"110111101",
  41281=>"110011000",
  41282=>"010000010",
  41283=>"101100100",
  41284=>"010001000",
  41285=>"010011110",
  41286=>"100011101",
  41287=>"111100101",
  41288=>"011011110",
  41289=>"000000000",
  41290=>"101111010",
  41291=>"001100111",
  41292=>"011000111",
  41293=>"100001010",
  41294=>"100010000",
  41295=>"001011001",
  41296=>"011101011",
  41297=>"111010011",
  41298=>"000011100",
  41299=>"111010111",
  41300=>"111100000",
  41301=>"000011011",
  41302=>"101110011",
  41303=>"110101010",
  41304=>"100011011",
  41305=>"110001000",
  41306=>"100000111",
  41307=>"110110111",
  41308=>"101001110",
  41309=>"100011101",
  41310=>"101110001",
  41311=>"101001110",
  41312=>"111000001",
  41313=>"110000101",
  41314=>"100101110",
  41315=>"011111011",
  41316=>"000001000",
  41317=>"000001111",
  41318=>"001011001",
  41319=>"011101010",
  41320=>"011001010",
  41321=>"100111110",
  41322=>"101000000",
  41323=>"001001110",
  41324=>"101110111",
  41325=>"011101010",
  41326=>"010111110",
  41327=>"111111111",
  41328=>"000011101",
  41329=>"111110001",
  41330=>"111100110",
  41331=>"011100100",
  41332=>"101000111",
  41333=>"001011100",
  41334=>"100111101",
  41335=>"110000110",
  41336=>"011001000",
  41337=>"011001000",
  41338=>"110110011",
  41339=>"111001101",
  41340=>"011011010",
  41341=>"000010101",
  41342=>"110101101",
  41343=>"110011101",
  41344=>"010111000",
  41345=>"010010010",
  41346=>"001011111",
  41347=>"111000100",
  41348=>"100110010",
  41349=>"101100111",
  41350=>"001111110",
  41351=>"010100100",
  41352=>"001010010",
  41353=>"010111010",
  41354=>"001100110",
  41355=>"001011011",
  41356=>"110100111",
  41357=>"000001000",
  41358=>"100111010",
  41359=>"011011111",
  41360=>"111001011",
  41361=>"110000000",
  41362=>"110100101",
  41363=>"010100011",
  41364=>"110110101",
  41365=>"110101101",
  41366=>"110111111",
  41367=>"011111101",
  41368=>"001010001",
  41369=>"101010001",
  41370=>"010010111",
  41371=>"101011110",
  41372=>"001101010",
  41373=>"100100101",
  41374=>"110001100",
  41375=>"111101111",
  41376=>"110100111",
  41377=>"111000100",
  41378=>"101010001",
  41379=>"000000011",
  41380=>"111001111",
  41381=>"010010110",
  41382=>"001001000",
  41383=>"001100001",
  41384=>"001100010",
  41385=>"111010111",
  41386=>"110110111",
  41387=>"001000100",
  41388=>"110101110",
  41389=>"101100100",
  41390=>"000110110",
  41391=>"110000010",
  41392=>"101000010",
  41393=>"110111110",
  41394=>"010110010",
  41395=>"000100000",
  41396=>"100001000",
  41397=>"010011110",
  41398=>"010100110",
  41399=>"110011011",
  41400=>"100010011",
  41401=>"011010011",
  41402=>"101110101",
  41403=>"101010001",
  41404=>"111101011",
  41405=>"100010000",
  41406=>"110110100",
  41407=>"110101000",
  41408=>"101001000",
  41409=>"000100010",
  41410=>"110111000",
  41411=>"100001011",
  41412=>"101100110",
  41413=>"000011000",
  41414=>"010101010",
  41415=>"010010100",
  41416=>"110000000",
  41417=>"011110111",
  41418=>"010100001",
  41419=>"001001101",
  41420=>"110000111",
  41421=>"000111001",
  41422=>"000101001",
  41423=>"001110011",
  41424=>"110010010",
  41425=>"000000100",
  41426=>"100000001",
  41427=>"001110110",
  41428=>"001101001",
  41429=>"111111100",
  41430=>"000011100",
  41431=>"000110111",
  41432=>"010111000",
  41433=>"101111100",
  41434=>"001110000",
  41435=>"100000101",
  41436=>"010101011",
  41437=>"100111100",
  41438=>"000000001",
  41439=>"101111011",
  41440=>"000010110",
  41441=>"100001011",
  41442=>"100110110",
  41443=>"011101110",
  41444=>"000000110",
  41445=>"010111001",
  41446=>"111110111",
  41447=>"100011000",
  41448=>"011011110",
  41449=>"111101000",
  41450=>"101111110",
  41451=>"000101011",
  41452=>"110011100",
  41453=>"111100100",
  41454=>"010001000",
  41455=>"001000110",
  41456=>"010000111",
  41457=>"101101010",
  41458=>"101100100",
  41459=>"010001001",
  41460=>"101101110",
  41461=>"000110010",
  41462=>"001101001",
  41463=>"110111001",
  41464=>"011101101",
  41465=>"100010100",
  41466=>"110111111",
  41467=>"111111011",
  41468=>"110100110",
  41469=>"100110011",
  41470=>"001110000",
  41471=>"100100111",
  41472=>"000000110",
  41473=>"101000110",
  41474=>"000101101",
  41475=>"010100110",
  41476=>"100100100",
  41477=>"100111111",
  41478=>"111111100",
  41479=>"100111011",
  41480=>"001100001",
  41481=>"101100111",
  41482=>"000100000",
  41483=>"001011000",
  41484=>"010010011",
  41485=>"001010001",
  41486=>"000100111",
  41487=>"010001110",
  41488=>"010000100",
  41489=>"001111010",
  41490=>"110001010",
  41491=>"010101000",
  41492=>"010110100",
  41493=>"000010110",
  41494=>"100111111",
  41495=>"100110111",
  41496=>"100100000",
  41497=>"011110101",
  41498=>"100010101",
  41499=>"110110010",
  41500=>"010011000",
  41501=>"000100100",
  41502=>"111110000",
  41503=>"111111101",
  41504=>"000100101",
  41505=>"000010010",
  41506=>"010001001",
  41507=>"011000001",
  41508=>"000111000",
  41509=>"000101011",
  41510=>"100110110",
  41511=>"100111111",
  41512=>"000111110",
  41513=>"110011010",
  41514=>"100101010",
  41515=>"111110010",
  41516=>"100110010",
  41517=>"001111001",
  41518=>"111000110",
  41519=>"010001101",
  41520=>"111100100",
  41521=>"001001100",
  41522=>"111001100",
  41523=>"111010011",
  41524=>"001111011",
  41525=>"101101111",
  41526=>"100010000",
  41527=>"011001100",
  41528=>"000011010",
  41529=>"111110110",
  41530=>"011111011",
  41531=>"001011011",
  41532=>"011010110",
  41533=>"111001010",
  41534=>"101101110",
  41535=>"100001001",
  41536=>"100100100",
  41537=>"011011001",
  41538=>"100011011",
  41539=>"000110100",
  41540=>"101010111",
  41541=>"000011101",
  41542=>"101101110",
  41543=>"010111010",
  41544=>"010000000",
  41545=>"110101111",
  41546=>"111011100",
  41547=>"100111111",
  41548=>"001001100",
  41549=>"110001110",
  41550=>"000111110",
  41551=>"011010000",
  41552=>"100110010",
  41553=>"101010100",
  41554=>"000010010",
  41555=>"001010111",
  41556=>"000011001",
  41557=>"111100101",
  41558=>"000001011",
  41559=>"110100110",
  41560=>"001000001",
  41561=>"111111100",
  41562=>"010101011",
  41563=>"000100011",
  41564=>"101010010",
  41565=>"111001110",
  41566=>"001010101",
  41567=>"100000110",
  41568=>"010111001",
  41569=>"000000000",
  41570=>"010110001",
  41571=>"111001001",
  41572=>"111000000",
  41573=>"101111011",
  41574=>"000010001",
  41575=>"101001111",
  41576=>"011000000",
  41577=>"110010101",
  41578=>"011100111",
  41579=>"100110111",
  41580=>"101110000",
  41581=>"011010000",
  41582=>"001001100",
  41583=>"100011000",
  41584=>"000100011",
  41585=>"010000001",
  41586=>"001100011",
  41587=>"101100001",
  41588=>"010001101",
  41589=>"001000001",
  41590=>"111011110",
  41591=>"001110111",
  41592=>"101110000",
  41593=>"100110110",
  41594=>"101101000",
  41595=>"001010001",
  41596=>"111000011",
  41597=>"111000001",
  41598=>"110100101",
  41599=>"010110111",
  41600=>"101100110",
  41601=>"110110110",
  41602=>"110101100",
  41603=>"110000000",
  41604=>"100101010",
  41605=>"000100010",
  41606=>"100000011",
  41607=>"001011010",
  41608=>"111010000",
  41609=>"000110111",
  41610=>"111111010",
  41611=>"010011011",
  41612=>"000010011",
  41613=>"000101101",
  41614=>"011110100",
  41615=>"100110111",
  41616=>"000001010",
  41617=>"000101011",
  41618=>"111110111",
  41619=>"011101100",
  41620=>"011011100",
  41621=>"011001010",
  41622=>"010011110",
  41623=>"000101100",
  41624=>"110100110",
  41625=>"000110101",
  41626=>"111110001",
  41627=>"001111100",
  41628=>"100001110",
  41629=>"110111010",
  41630=>"001101110",
  41631=>"110110100",
  41632=>"110000110",
  41633=>"110100001",
  41634=>"110001100",
  41635=>"111000100",
  41636=>"000100100",
  41637=>"111101100",
  41638=>"111111000",
  41639=>"110100001",
  41640=>"010000000",
  41641=>"100100000",
  41642=>"110100010",
  41643=>"111000111",
  41644=>"100001011",
  41645=>"110111101",
  41646=>"010100011",
  41647=>"001001101",
  41648=>"001101100",
  41649=>"101100111",
  41650=>"111001010",
  41651=>"000101100",
  41652=>"011001001",
  41653=>"011010101",
  41654=>"111101001",
  41655=>"101101110",
  41656=>"110100011",
  41657=>"100001100",
  41658=>"100001001",
  41659=>"000111111",
  41660=>"110111100",
  41661=>"010110100",
  41662=>"110111111",
  41663=>"111000101",
  41664=>"100101011",
  41665=>"011010111",
  41666=>"111101010",
  41667=>"000100001",
  41668=>"001000010",
  41669=>"111110101",
  41670=>"110101001",
  41671=>"110010111",
  41672=>"110000110",
  41673=>"001010011",
  41674=>"100111110",
  41675=>"000100000",
  41676=>"100110011",
  41677=>"011001000",
  41678=>"101000011",
  41679=>"001111101",
  41680=>"100111111",
  41681=>"001110110",
  41682=>"100011100",
  41683=>"110000000",
  41684=>"110110111",
  41685=>"111001111",
  41686=>"011011011",
  41687=>"100110101",
  41688=>"100100001",
  41689=>"010010001",
  41690=>"110001010",
  41691=>"000111101",
  41692=>"110110110",
  41693=>"110111111",
  41694=>"011011101",
  41695=>"000011000",
  41696=>"001110100",
  41697=>"010000001",
  41698=>"110100110",
  41699=>"011111001",
  41700=>"101111101",
  41701=>"000100111",
  41702=>"001011100",
  41703=>"100001010",
  41704=>"010111001",
  41705=>"000111110",
  41706=>"010101000",
  41707=>"010110011",
  41708=>"010000110",
  41709=>"100111010",
  41710=>"001001110",
  41711=>"100101001",
  41712=>"111001011",
  41713=>"011100100",
  41714=>"010011111",
  41715=>"111111010",
  41716=>"000100010",
  41717=>"110110101",
  41718=>"011001010",
  41719=>"110000001",
  41720=>"001000011",
  41721=>"011000101",
  41722=>"001100101",
  41723=>"011110000",
  41724=>"100010000",
  41725=>"101110001",
  41726=>"000001100",
  41727=>"110010101",
  41728=>"110000101",
  41729=>"100010010",
  41730=>"000000011",
  41731=>"010101010",
  41732=>"000001010",
  41733=>"110111000",
  41734=>"011010010",
  41735=>"110000101",
  41736=>"010110110",
  41737=>"111100001",
  41738=>"011110110",
  41739=>"001110000",
  41740=>"011001011",
  41741=>"000011001",
  41742=>"100000100",
  41743=>"000010011",
  41744=>"101111011",
  41745=>"100101110",
  41746=>"000100001",
  41747=>"111010001",
  41748=>"010110000",
  41749=>"001010000",
  41750=>"100011000",
  41751=>"000001110",
  41752=>"000100000",
  41753=>"000001001",
  41754=>"011101100",
  41755=>"010000100",
  41756=>"011011111",
  41757=>"101000111",
  41758=>"100100111",
  41759=>"111111001",
  41760=>"101111111",
  41761=>"000000111",
  41762=>"001010110",
  41763=>"100110110",
  41764=>"011100100",
  41765=>"110110010",
  41766=>"001000001",
  41767=>"110011110",
  41768=>"110000011",
  41769=>"001001000",
  41770=>"110011100",
  41771=>"110111100",
  41772=>"010010111",
  41773=>"111111111",
  41774=>"100100101",
  41775=>"101100111",
  41776=>"011000010",
  41777=>"001100101",
  41778=>"011110000",
  41779=>"010111001",
  41780=>"100110110",
  41781=>"010100101",
  41782=>"110001000",
  41783=>"101101011",
  41784=>"000000000",
  41785=>"110100110",
  41786=>"100011111",
  41787=>"110011100",
  41788=>"010101011",
  41789=>"010111111",
  41790=>"001000100",
  41791=>"101101101",
  41792=>"101011100",
  41793=>"101011001",
  41794=>"100011001",
  41795=>"101111100",
  41796=>"111111110",
  41797=>"100101010",
  41798=>"100110110",
  41799=>"010111100",
  41800=>"010111000",
  41801=>"011110000",
  41802=>"011110000",
  41803=>"000110100",
  41804=>"101101100",
  41805=>"110100101",
  41806=>"100000111",
  41807=>"011000101",
  41808=>"111110100",
  41809=>"110111101",
  41810=>"110110010",
  41811=>"000010101",
  41812=>"100000010",
  41813=>"100011111",
  41814=>"101000010",
  41815=>"000001101",
  41816=>"010011010",
  41817=>"000100011",
  41818=>"110101001",
  41819=>"010110000",
  41820=>"100100101",
  41821=>"110000001",
  41822=>"011010100",
  41823=>"110101110",
  41824=>"111000010",
  41825=>"100110111",
  41826=>"010001000",
  41827=>"000011100",
  41828=>"110011100",
  41829=>"110010101",
  41830=>"110010000",
  41831=>"010000111",
  41832=>"000000111",
  41833=>"010000001",
  41834=>"111011100",
  41835=>"101110111",
  41836=>"110111000",
  41837=>"000000010",
  41838=>"100000010",
  41839=>"011011011",
  41840=>"011000010",
  41841=>"010010101",
  41842=>"101101010",
  41843=>"001101010",
  41844=>"010100110",
  41845=>"011001101",
  41846=>"010100111",
  41847=>"111101110",
  41848=>"011101001",
  41849=>"100110110",
  41850=>"111101000",
  41851=>"010001011",
  41852=>"100000000",
  41853=>"101110001",
  41854=>"111100111",
  41855=>"111111100",
  41856=>"011000000",
  41857=>"111011001",
  41858=>"010000111",
  41859=>"000111100",
  41860=>"000100111",
  41861=>"011101011",
  41862=>"101110001",
  41863=>"011000110",
  41864=>"101100001",
  41865=>"100111000",
  41866=>"011101000",
  41867=>"101010000",
  41868=>"000101001",
  41869=>"100001001",
  41870=>"000101111",
  41871=>"101110010",
  41872=>"100011100",
  41873=>"111000110",
  41874=>"100010110",
  41875=>"101010100",
  41876=>"100011010",
  41877=>"110100110",
  41878=>"101101101",
  41879=>"100101001",
  41880=>"011010001",
  41881=>"110111110",
  41882=>"101100100",
  41883=>"001000011",
  41884=>"110110101",
  41885=>"110001101",
  41886=>"100001101",
  41887=>"100000100",
  41888=>"000000000",
  41889=>"100000000",
  41890=>"101000111",
  41891=>"010111001",
  41892=>"110000010",
  41893=>"111110100",
  41894=>"010111100",
  41895=>"001100100",
  41896=>"001101100",
  41897=>"110100010",
  41898=>"100010101",
  41899=>"001001010",
  41900=>"111000000",
  41901=>"101110011",
  41902=>"110010000",
  41903=>"100101110",
  41904=>"011111110",
  41905=>"111100111",
  41906=>"011111111",
  41907=>"101010001",
  41908=>"111010101",
  41909=>"100000010",
  41910=>"011011010",
  41911=>"001101010",
  41912=>"101010101",
  41913=>"011110111",
  41914=>"000001011",
  41915=>"000100010",
  41916=>"000010001",
  41917=>"111010100",
  41918=>"111111101",
  41919=>"010101100",
  41920=>"011100111",
  41921=>"010001001",
  41922=>"110001101",
  41923=>"100101001",
  41924=>"001000011",
  41925=>"010110100",
  41926=>"001001001",
  41927=>"010110010",
  41928=>"000001001",
  41929=>"110011011",
  41930=>"000011111",
  41931=>"110110101",
  41932=>"111101110",
  41933=>"100000010",
  41934=>"001111010",
  41935=>"111010001",
  41936=>"110100011",
  41937=>"100001001",
  41938=>"110011100",
  41939=>"101010011",
  41940=>"000010101",
  41941=>"000100001",
  41942=>"101011101",
  41943=>"001111011",
  41944=>"111111001",
  41945=>"000000001",
  41946=>"101100000",
  41947=>"110000111",
  41948=>"110101100",
  41949=>"101001000",
  41950=>"001001010",
  41951=>"111101100",
  41952=>"010000000",
  41953=>"011110001",
  41954=>"000010001",
  41955=>"001000110",
  41956=>"100110000",
  41957=>"111010110",
  41958=>"101101100",
  41959=>"001100110",
  41960=>"101100100",
  41961=>"000010110",
  41962=>"001110100",
  41963=>"100000101",
  41964=>"010001100",
  41965=>"100011000",
  41966=>"010011011",
  41967=>"111011101",
  41968=>"010110111",
  41969=>"110110110",
  41970=>"000111101",
  41971=>"100110101",
  41972=>"110101000",
  41973=>"000000001",
  41974=>"100101110",
  41975=>"110000111",
  41976=>"011111111",
  41977=>"101110000",
  41978=>"100101000",
  41979=>"111110000",
  41980=>"111110111",
  41981=>"001010010",
  41982=>"011011010",
  41983=>"001000010",
  41984=>"000000101",
  41985=>"111100100",
  41986=>"000100110",
  41987=>"010001000",
  41988=>"110101010",
  41989=>"010100111",
  41990=>"110011111",
  41991=>"001111000",
  41992=>"110111011",
  41993=>"000101101",
  41994=>"110100010",
  41995=>"011010011",
  41996=>"110000101",
  41997=>"101111100",
  41998=>"010010101",
  41999=>"100100011",
  42000=>"111001001",
  42001=>"001111111",
  42002=>"111110011",
  42003=>"111010110",
  42004=>"111000111",
  42005=>"110010110",
  42006=>"001111000",
  42007=>"001111001",
  42008=>"001011010",
  42009=>"110110010",
  42010=>"101001001",
  42011=>"111101100",
  42012=>"010001111",
  42013=>"000000001",
  42014=>"010101110",
  42015=>"000011010",
  42016=>"000000101",
  42017=>"000011000",
  42018=>"100111110",
  42019=>"001110111",
  42020=>"000001100",
  42021=>"111111011",
  42022=>"110111111",
  42023=>"010111101",
  42024=>"001100101",
  42025=>"100011100",
  42026=>"100001011",
  42027=>"111000010",
  42028=>"000000001",
  42029=>"000011011",
  42030=>"101011001",
  42031=>"001000101",
  42032=>"001000100",
  42033=>"010000110",
  42034=>"100111000",
  42035=>"110100101",
  42036=>"101101110",
  42037=>"001000011",
  42038=>"000010110",
  42039=>"100010011",
  42040=>"110011100",
  42041=>"111010111",
  42042=>"001101101",
  42043=>"000000000",
  42044=>"000000010",
  42045=>"011011111",
  42046=>"110011000",
  42047=>"011000110",
  42048=>"010001101",
  42049=>"010000110",
  42050=>"011000110",
  42051=>"010110110",
  42052=>"110100011",
  42053=>"100110111",
  42054=>"111110111",
  42055=>"101101100",
  42056=>"101010111",
  42057=>"011001110",
  42058=>"101111100",
  42059=>"010001010",
  42060=>"000110000",
  42061=>"100001100",
  42062=>"111000100",
  42063=>"000111001",
  42064=>"011100111",
  42065=>"011011010",
  42066=>"101110001",
  42067=>"110100011",
  42068=>"111001000",
  42069=>"111000101",
  42070=>"000001011",
  42071=>"101001011",
  42072=>"110101111",
  42073=>"010110011",
  42074=>"011101100",
  42075=>"011100100",
  42076=>"000100100",
  42077=>"000000000",
  42078=>"010001100",
  42079=>"110110001",
  42080=>"000000010",
  42081=>"011111101",
  42082=>"101101010",
  42083=>"000001111",
  42084=>"111010100",
  42085=>"000010111",
  42086=>"111111110",
  42087=>"010111000",
  42088=>"001111111",
  42089=>"010000101",
  42090=>"111100001",
  42091=>"100010111",
  42092=>"100010010",
  42093=>"001011111",
  42094=>"001000000",
  42095=>"001111011",
  42096=>"001010010",
  42097=>"110110111",
  42098=>"101100010",
  42099=>"011100001",
  42100=>"111000000",
  42101=>"010011101",
  42102=>"010011001",
  42103=>"000111110",
  42104=>"001111010",
  42105=>"111011011",
  42106=>"010000000",
  42107=>"011100010",
  42108=>"011100010",
  42109=>"010110110",
  42110=>"100100111",
  42111=>"000011111",
  42112=>"011110101",
  42113=>"001011111",
  42114=>"101011011",
  42115=>"001110011",
  42116=>"000010110",
  42117=>"111000101",
  42118=>"110010110",
  42119=>"110111100",
  42120=>"000011110",
  42121=>"010100111",
  42122=>"010001101",
  42123=>"100000111",
  42124=>"010010101",
  42125=>"100101010",
  42126=>"110100111",
  42127=>"101001111",
  42128=>"101000110",
  42129=>"011010111",
  42130=>"010101010",
  42131=>"011100110",
  42132=>"100100110",
  42133=>"000000100",
  42134=>"111111110",
  42135=>"111000001",
  42136=>"101111110",
  42137=>"111111011",
  42138=>"001011110",
  42139=>"000110001",
  42140=>"101111001",
  42141=>"011111010",
  42142=>"011011101",
  42143=>"001000111",
  42144=>"001000101",
  42145=>"001010011",
  42146=>"010101101",
  42147=>"110000111",
  42148=>"011110011",
  42149=>"111110110",
  42150=>"001110011",
  42151=>"111100101",
  42152=>"111001110",
  42153=>"011111111",
  42154=>"101111011",
  42155=>"011110111",
  42156=>"101010101",
  42157=>"101001011",
  42158=>"110000100",
  42159=>"000101110",
  42160=>"000100010",
  42161=>"001010010",
  42162=>"111001001",
  42163=>"111100011",
  42164=>"001100010",
  42165=>"001011011",
  42166=>"111101001",
  42167=>"011100000",
  42168=>"101101101",
  42169=>"110000011",
  42170=>"110001011",
  42171=>"010111001",
  42172=>"010100001",
  42173=>"011100110",
  42174=>"111101011",
  42175=>"111100111",
  42176=>"000001101",
  42177=>"101111111",
  42178=>"110110000",
  42179=>"110000101",
  42180=>"100110010",
  42181=>"111111100",
  42182=>"000100010",
  42183=>"100100101",
  42184=>"011101010",
  42185=>"111011001",
  42186=>"110001001",
  42187=>"001100111",
  42188=>"011110011",
  42189=>"100110011",
  42190=>"011010110",
  42191=>"101011001",
  42192=>"000001110",
  42193=>"110011011",
  42194=>"100100111",
  42195=>"010111000",
  42196=>"101011001",
  42197=>"111100001",
  42198=>"010001001",
  42199=>"000010011",
  42200=>"000101111",
  42201=>"011101111",
  42202=>"101000010",
  42203=>"000000000",
  42204=>"001001010",
  42205=>"111101110",
  42206=>"111100101",
  42207=>"101011001",
  42208=>"101001111",
  42209=>"000000010",
  42210=>"010011111",
  42211=>"111111000",
  42212=>"111100001",
  42213=>"011000101",
  42214=>"101111001",
  42215=>"011011011",
  42216=>"110100111",
  42217=>"000001011",
  42218=>"100001010",
  42219=>"100010000",
  42220=>"000111010",
  42221=>"101010000",
  42222=>"010101011",
  42223=>"111100001",
  42224=>"111100100",
  42225=>"111010011",
  42226=>"011100111",
  42227=>"000011011",
  42228=>"011000110",
  42229=>"000110011",
  42230=>"110111000",
  42231=>"100111111",
  42232=>"011010111",
  42233=>"001100100",
  42234=>"000111100",
  42235=>"001011110",
  42236=>"110101111",
  42237=>"101110001",
  42238=>"110101110",
  42239=>"000101001",
  42240=>"111100100",
  42241=>"100110010",
  42242=>"111000101",
  42243=>"001000111",
  42244=>"101111001",
  42245=>"011101111",
  42246=>"111010000",
  42247=>"110001000",
  42248=>"001000101",
  42249=>"111000001",
  42250=>"100001000",
  42251=>"100000111",
  42252=>"001101100",
  42253=>"110111111",
  42254=>"101110011",
  42255=>"000010010",
  42256=>"101010000",
  42257=>"111101001",
  42258=>"111011101",
  42259=>"101001101",
  42260=>"010011101",
  42261=>"100000100",
  42262=>"100001000",
  42263=>"101101010",
  42264=>"110101111",
  42265=>"010000100",
  42266=>"100000111",
  42267=>"100111000",
  42268=>"000011100",
  42269=>"101111111",
  42270=>"111101100",
  42271=>"110001010",
  42272=>"000000100",
  42273=>"010110001",
  42274=>"001111101",
  42275=>"011010101",
  42276=>"001100001",
  42277=>"011111101",
  42278=>"110011100",
  42279=>"100001111",
  42280=>"000101110",
  42281=>"111110110",
  42282=>"000000011",
  42283=>"111111101",
  42284=>"111011111",
  42285=>"100010000",
  42286=>"100000111",
  42287=>"110010010",
  42288=>"000000000",
  42289=>"010000110",
  42290=>"110000110",
  42291=>"011110001",
  42292=>"111111010",
  42293=>"111000001",
  42294=>"110100111",
  42295=>"011101111",
  42296=>"001000000",
  42297=>"111110110",
  42298=>"111111100",
  42299=>"111000000",
  42300=>"101110011",
  42301=>"100111010",
  42302=>"001110111",
  42303=>"011100100",
  42304=>"011101111",
  42305=>"010101101",
  42306=>"111100001",
  42307=>"110101111",
  42308=>"001111011",
  42309=>"011111101",
  42310=>"010101100",
  42311=>"110101110",
  42312=>"001101101",
  42313=>"011011010",
  42314=>"011001111",
  42315=>"000100001",
  42316=>"011111110",
  42317=>"111110000",
  42318=>"110101010",
  42319=>"100001000",
  42320=>"110001111",
  42321=>"101001111",
  42322=>"011001110",
  42323=>"110010001",
  42324=>"011111101",
  42325=>"010001100",
  42326=>"000111100",
  42327=>"001101100",
  42328=>"000100000",
  42329=>"011101101",
  42330=>"011000101",
  42331=>"011111110",
  42332=>"111011100",
  42333=>"110100101",
  42334=>"111000011",
  42335=>"110010111",
  42336=>"100111000",
  42337=>"010110111",
  42338=>"010011010",
  42339=>"111101101",
  42340=>"100101100",
  42341=>"010101100",
  42342=>"000110001",
  42343=>"001111111",
  42344=>"101110101",
  42345=>"100010010",
  42346=>"111010111",
  42347=>"000011010",
  42348=>"111010110",
  42349=>"101010010",
  42350=>"000010000",
  42351=>"010101110",
  42352=>"101000100",
  42353=>"100111110",
  42354=>"010100010",
  42355=>"001101101",
  42356=>"100011010",
  42357=>"000010100",
  42358=>"111000110",
  42359=>"100111010",
  42360=>"101010010",
  42361=>"110100110",
  42362=>"100101011",
  42363=>"100001000",
  42364=>"000011111",
  42365=>"100101000",
  42366=>"000100010",
  42367=>"111001001",
  42368=>"000000110",
  42369=>"101010011",
  42370=>"000101001",
  42371=>"000111011",
  42372=>"111010111",
  42373=>"110011001",
  42374=>"010111011",
  42375=>"111101011",
  42376=>"010100000",
  42377=>"111110110",
  42378=>"011011011",
  42379=>"101000110",
  42380=>"110000001",
  42381=>"110110101",
  42382=>"101101111",
  42383=>"101001100",
  42384=>"111100000",
  42385=>"000110000",
  42386=>"101111010",
  42387=>"111010111",
  42388=>"110100111",
  42389=>"000000010",
  42390=>"000001100",
  42391=>"001110101",
  42392=>"101100110",
  42393=>"010110111",
  42394=>"110110110",
  42395=>"000001000",
  42396=>"101011111",
  42397=>"000011010",
  42398=>"111110000",
  42399=>"011010111",
  42400=>"001111011",
  42401=>"100011011",
  42402=>"101001000",
  42403=>"000101000",
  42404=>"000000010",
  42405=>"000100101",
  42406=>"001101101",
  42407=>"011100000",
  42408=>"110110010",
  42409=>"001110000",
  42410=>"101110101",
  42411=>"101010010",
  42412=>"111000010",
  42413=>"001111010",
  42414=>"101000000",
  42415=>"110111100",
  42416=>"001010100",
  42417=>"111100011",
  42418=>"111110100",
  42419=>"100100100",
  42420=>"110001110",
  42421=>"001011110",
  42422=>"011001001",
  42423=>"110110010",
  42424=>"010000100",
  42425=>"101100001",
  42426=>"101001101",
  42427=>"111110111",
  42428=>"011000100",
  42429=>"000101111",
  42430=>"000011110",
  42431=>"010110111",
  42432=>"111110100",
  42433=>"101010111",
  42434=>"000001100",
  42435=>"110001010",
  42436=>"011110001",
  42437=>"010011100",
  42438=>"000101000",
  42439=>"010000000",
  42440=>"111011110",
  42441=>"001101001",
  42442=>"010010100",
  42443=>"111001110",
  42444=>"001111010",
  42445=>"010010100",
  42446=>"110001100",
  42447=>"101101011",
  42448=>"100101000",
  42449=>"101110000",
  42450=>"010010101",
  42451=>"110010001",
  42452=>"010000100",
  42453=>"000000101",
  42454=>"010101010",
  42455=>"101000001",
  42456=>"111110010",
  42457=>"011000000",
  42458=>"000110010",
  42459=>"000101100",
  42460=>"110011111",
  42461=>"000111110",
  42462=>"110000100",
  42463=>"111110011",
  42464=>"101000000",
  42465=>"010010111",
  42466=>"001010110",
  42467=>"011101110",
  42468=>"100000111",
  42469=>"100101000",
  42470=>"000101000",
  42471=>"001010001",
  42472=>"011111000",
  42473=>"101110111",
  42474=>"110100110",
  42475=>"010011110",
  42476=>"111100100",
  42477=>"101110111",
  42478=>"010001001",
  42479=>"010100011",
  42480=>"110110100",
  42481=>"100101101",
  42482=>"101111111",
  42483=>"001110111",
  42484=>"010010010",
  42485=>"001100100",
  42486=>"111010111",
  42487=>"110110100",
  42488=>"111010010",
  42489=>"001110000",
  42490=>"100001111",
  42491=>"011000011",
  42492=>"010000010",
  42493=>"111001011",
  42494=>"011110001",
  42495=>"000010111",
  42496=>"110011111",
  42497=>"001000110",
  42498=>"101010100",
  42499=>"111000111",
  42500=>"011011110",
  42501=>"000001000",
  42502=>"100101000",
  42503=>"111100001",
  42504=>"000101110",
  42505=>"011101100",
  42506=>"100100110",
  42507=>"001111000",
  42508=>"001001111",
  42509=>"111100000",
  42510=>"100001100",
  42511=>"111111100",
  42512=>"011111110",
  42513=>"001110011",
  42514=>"111100000",
  42515=>"000000001",
  42516=>"000101111",
  42517=>"001010001",
  42518=>"011110101",
  42519=>"010011101",
  42520=>"111001101",
  42521=>"000111111",
  42522=>"101110011",
  42523=>"101010000",
  42524=>"101101111",
  42525=>"100010111",
  42526=>"011001110",
  42527=>"001001010",
  42528=>"100010100",
  42529=>"110100001",
  42530=>"011111001",
  42531=>"100001111",
  42532=>"111011011",
  42533=>"000000111",
  42534=>"100000100",
  42535=>"111000000",
  42536=>"110100100",
  42537=>"001010000",
  42538=>"000111001",
  42539=>"100010000",
  42540=>"000001010",
  42541=>"011001110",
  42542=>"001001000",
  42543=>"001111000",
  42544=>"010111010",
  42545=>"101110000",
  42546=>"111100110",
  42547=>"100000010",
  42548=>"110101101",
  42549=>"001001001",
  42550=>"010001100",
  42551=>"001111100",
  42552=>"100101111",
  42553=>"111001110",
  42554=>"101110101",
  42555=>"101110101",
  42556=>"110100111",
  42557=>"000001100",
  42558=>"011101111",
  42559=>"111001010",
  42560=>"011010100",
  42561=>"100100010",
  42562=>"100101111",
  42563=>"011000110",
  42564=>"100000000",
  42565=>"010110101",
  42566=>"010011000",
  42567=>"111111110",
  42568=>"100111100",
  42569=>"111100010",
  42570=>"010001111",
  42571=>"001011111",
  42572=>"110000100",
  42573=>"101101011",
  42574=>"101101011",
  42575=>"001011011",
  42576=>"010010011",
  42577=>"110100001",
  42578=>"000011011",
  42579=>"110110101",
  42580=>"000001000",
  42581=>"100110100",
  42582=>"000101011",
  42583=>"111010001",
  42584=>"111001010",
  42585=>"111001001",
  42586=>"011101101",
  42587=>"001101100",
  42588=>"101000101",
  42589=>"111100000",
  42590=>"111011000",
  42591=>"100101110",
  42592=>"011001011",
  42593=>"000010110",
  42594=>"100110011",
  42595=>"100101011",
  42596=>"110000010",
  42597=>"000100110",
  42598=>"011111100",
  42599=>"110011111",
  42600=>"000010001",
  42601=>"100101011",
  42602=>"010110101",
  42603=>"000011010",
  42604=>"101011111",
  42605=>"001010101",
  42606=>"100011111",
  42607=>"101111000",
  42608=>"100111000",
  42609=>"110001110",
  42610=>"000001111",
  42611=>"011110000",
  42612=>"100001100",
  42613=>"101000000",
  42614=>"010100101",
  42615=>"101101101",
  42616=>"000101111",
  42617=>"010101000",
  42618=>"010000000",
  42619=>"011010111",
  42620=>"101110101",
  42621=>"101110100",
  42622=>"000100001",
  42623=>"010011100",
  42624=>"101000101",
  42625=>"001001110",
  42626=>"101100000",
  42627=>"100111100",
  42628=>"100001011",
  42629=>"101001010",
  42630=>"000011110",
  42631=>"111001111",
  42632=>"000000111",
  42633=>"111101011",
  42634=>"111011110",
  42635=>"001110011",
  42636=>"111000110",
  42637=>"100011110",
  42638=>"110110010",
  42639=>"011000110",
  42640=>"101001101",
  42641=>"011100100",
  42642=>"001011010",
  42643=>"000001011",
  42644=>"000001100",
  42645=>"011011001",
  42646=>"001000110",
  42647=>"010100101",
  42648=>"110011101",
  42649=>"100011101",
  42650=>"110010010",
  42651=>"010101111",
  42652=>"100011110",
  42653=>"010000001",
  42654=>"000000000",
  42655=>"001001001",
  42656=>"111000000",
  42657=>"000001001",
  42658=>"000111011",
  42659=>"000110110",
  42660=>"101000010",
  42661=>"101010101",
  42662=>"111111111",
  42663=>"011100110",
  42664=>"010110100",
  42665=>"000111100",
  42666=>"011101110",
  42667=>"100011111",
  42668=>"011010011",
  42669=>"000111010",
  42670=>"000100100",
  42671=>"110001011",
  42672=>"010001010",
  42673=>"001000000",
  42674=>"110000000",
  42675=>"011111011",
  42676=>"011001000",
  42677=>"110110000",
  42678=>"111110110",
  42679=>"101101011",
  42680=>"010000101",
  42681=>"000110110",
  42682=>"111101110",
  42683=>"001001010",
  42684=>"110010000",
  42685=>"111010010",
  42686=>"000010111",
  42687=>"111111100",
  42688=>"100110000",
  42689=>"101001111",
  42690=>"010101111",
  42691=>"001100101",
  42692=>"010010011",
  42693=>"111000101",
  42694=>"100110000",
  42695=>"111100100",
  42696=>"011000111",
  42697=>"010111100",
  42698=>"000111111",
  42699=>"110010011",
  42700=>"111000110",
  42701=>"011001001",
  42702=>"110011010",
  42703=>"110100000",
  42704=>"000111000",
  42705=>"000101010",
  42706=>"001110110",
  42707=>"110000000",
  42708=>"000011010",
  42709=>"000100110",
  42710=>"011111111",
  42711=>"011010101",
  42712=>"111000111",
  42713=>"100100101",
  42714=>"010110010",
  42715=>"100110000",
  42716=>"110001100",
  42717=>"100100001",
  42718=>"011011101",
  42719=>"101000000",
  42720=>"001001110",
  42721=>"011001000",
  42722=>"011110110",
  42723=>"111011110",
  42724=>"001111101",
  42725=>"000000001",
  42726=>"011110111",
  42727=>"101101111",
  42728=>"111010001",
  42729=>"111111000",
  42730=>"101110010",
  42731=>"100011011",
  42732=>"000111111",
  42733=>"111011001",
  42734=>"000101010",
  42735=>"001101101",
  42736=>"110110111",
  42737=>"010001010",
  42738=>"001000110",
  42739=>"010000001",
  42740=>"110100101",
  42741=>"010010000",
  42742=>"010101010",
  42743=>"011101011",
  42744=>"000111110",
  42745=>"001111101",
  42746=>"100010111",
  42747=>"000010011",
  42748=>"001110001",
  42749=>"100101000",
  42750=>"010000111",
  42751=>"100100101",
  42752=>"000000000",
  42753=>"101101011",
  42754=>"011011101",
  42755=>"110101110",
  42756=>"110000101",
  42757=>"011000111",
  42758=>"111001001",
  42759=>"000010011",
  42760=>"000010100",
  42761=>"100011000",
  42762=>"110110111",
  42763=>"101010110",
  42764=>"111101101",
  42765=>"100101000",
  42766=>"100000001",
  42767=>"011001100",
  42768=>"100100111",
  42769=>"010100110",
  42770=>"010010101",
  42771=>"001100110",
  42772=>"110010111",
  42773=>"010111111",
  42774=>"000110101",
  42775=>"000111111",
  42776=>"100011000",
  42777=>"000000010",
  42778=>"110011100",
  42779=>"010001111",
  42780=>"010010110",
  42781=>"110010101",
  42782=>"011101101",
  42783=>"010001010",
  42784=>"000100101",
  42785=>"011110101",
  42786=>"000000111",
  42787=>"011010110",
  42788=>"110011001",
  42789=>"000010000",
  42790=>"001111111",
  42791=>"100111101",
  42792=>"100111011",
  42793=>"001101110",
  42794=>"001010011",
  42795=>"001100110",
  42796=>"110000001",
  42797=>"101011111",
  42798=>"010101101",
  42799=>"101001011",
  42800=>"010110010",
  42801=>"011111011",
  42802=>"011011111",
  42803=>"000001001",
  42804=>"110110010",
  42805=>"010001111",
  42806=>"100010011",
  42807=>"000101001",
  42808=>"111011010",
  42809=>"111010011",
  42810=>"001100010",
  42811=>"101110000",
  42812=>"110010110",
  42813=>"101100100",
  42814=>"100000010",
  42815=>"110110011",
  42816=>"000000001",
  42817=>"111110010",
  42818=>"011001100",
  42819=>"111000111",
  42820=>"000110111",
  42821=>"110011100",
  42822=>"010010000",
  42823=>"101001101",
  42824=>"100111100",
  42825=>"111001111",
  42826=>"010110000",
  42827=>"011101010",
  42828=>"111011010",
  42829=>"011101110",
  42830=>"000011010",
  42831=>"111111101",
  42832=>"000000010",
  42833=>"100001000",
  42834=>"000001001",
  42835=>"011110011",
  42836=>"010100110",
  42837=>"000101110",
  42838=>"000101101",
  42839=>"110111100",
  42840=>"111110000",
  42841=>"110001001",
  42842=>"010111000",
  42843=>"100010010",
  42844=>"010010111",
  42845=>"001001010",
  42846=>"000011001",
  42847=>"000001110",
  42848=>"000111011",
  42849=>"111001111",
  42850=>"010001101",
  42851=>"001101000",
  42852=>"111010110",
  42853=>"001111101",
  42854=>"010000011",
  42855=>"010101010",
  42856=>"001110110",
  42857=>"100001010",
  42858=>"101101110",
  42859=>"001101001",
  42860=>"001111101",
  42861=>"010000100",
  42862=>"000000000",
  42863=>"111001011",
  42864=>"001010000",
  42865=>"110011011",
  42866=>"101101111",
  42867=>"110011101",
  42868=>"110110111",
  42869=>"001010011",
  42870=>"100011110",
  42871=>"000110010",
  42872=>"010010100",
  42873=>"001110000",
  42874=>"111100000",
  42875=>"001100100",
  42876=>"000001001",
  42877=>"111101111",
  42878=>"001001110",
  42879=>"011111100",
  42880=>"110001100",
  42881=>"110010000",
  42882=>"100111101",
  42883=>"010001110",
  42884=>"110110100",
  42885=>"110011000",
  42886=>"110000101",
  42887=>"000111001",
  42888=>"101101000",
  42889=>"111001011",
  42890=>"001110100",
  42891=>"001000000",
  42892=>"101000101",
  42893=>"010011110",
  42894=>"011110100",
  42895=>"101111110",
  42896=>"011101011",
  42897=>"100011100",
  42898=>"001111001",
  42899=>"111011111",
  42900=>"011010011",
  42901=>"110000010",
  42902=>"011110111",
  42903=>"100011011",
  42904=>"101111011",
  42905=>"111111111",
  42906=>"111111101",
  42907=>"100101011",
  42908=>"101111101",
  42909=>"011110001",
  42910=>"000110001",
  42911=>"111111000",
  42912=>"011111010",
  42913=>"000101101",
  42914=>"010011100",
  42915=>"101111001",
  42916=>"101001111",
  42917=>"000011111",
  42918=>"001101111",
  42919=>"110011111",
  42920=>"000110000",
  42921=>"011001010",
  42922=>"011101101",
  42923=>"110111011",
  42924=>"100101011",
  42925=>"011110001",
  42926=>"000100011",
  42927=>"001001001",
  42928=>"110110001",
  42929=>"110011111",
  42930=>"101101001",
  42931=>"000100010",
  42932=>"010010100",
  42933=>"011101010",
  42934=>"011001000",
  42935=>"101011100",
  42936=>"110111110",
  42937=>"001111001",
  42938=>"011010110",
  42939=>"001111011",
  42940=>"100111101",
  42941=>"001000100",
  42942=>"001110010",
  42943=>"111011111",
  42944=>"101010011",
  42945=>"111101111",
  42946=>"000000111",
  42947=>"110101100",
  42948=>"110101000",
  42949=>"001100001",
  42950=>"000001111",
  42951=>"100001010",
  42952=>"000000001",
  42953=>"000110110",
  42954=>"111101001",
  42955=>"011011110",
  42956=>"000000000",
  42957=>"001110010",
  42958=>"010110011",
  42959=>"011001000",
  42960=>"100000000",
  42961=>"011000111",
  42962=>"101100111",
  42963=>"101110001",
  42964=>"010101000",
  42965=>"010111100",
  42966=>"001011110",
  42967=>"001110010",
  42968=>"001101100",
  42969=>"001011011",
  42970=>"110000110",
  42971=>"001100011",
  42972=>"100010100",
  42973=>"100000100",
  42974=>"101100010",
  42975=>"111000101",
  42976=>"010010000",
  42977=>"001000011",
  42978=>"101100010",
  42979=>"101110111",
  42980=>"100010101",
  42981=>"111011100",
  42982=>"111100000",
  42983=>"111110010",
  42984=>"111001110",
  42985=>"110110111",
  42986=>"111101110",
  42987=>"000000100",
  42988=>"101100010",
  42989=>"000011110",
  42990=>"000110011",
  42991=>"011101100",
  42992=>"100010010",
  42993=>"010101101",
  42994=>"001100010",
  42995=>"101101011",
  42996=>"101010000",
  42997=>"100101011",
  42998=>"001100000",
  42999=>"000111010",
  43000=>"111111001",
  43001=>"101100100",
  43002=>"111011111",
  43003=>"000000101",
  43004=>"011011100",
  43005=>"110001011",
  43006=>"110011010",
  43007=>"111010111",
  43008=>"011000111",
  43009=>"110011101",
  43010=>"000111011",
  43011=>"011010101",
  43012=>"111111110",
  43013=>"100111001",
  43014=>"011111111",
  43015=>"010010101",
  43016=>"110001011",
  43017=>"000101001",
  43018=>"001000000",
  43019=>"010111001",
  43020=>"011111010",
  43021=>"100000101",
  43022=>"011011111",
  43023=>"011100000",
  43024=>"001011100",
  43025=>"000101111",
  43026=>"100111000",
  43027=>"100100011",
  43028=>"011011000",
  43029=>"011100101",
  43030=>"110101110",
  43031=>"101000001",
  43032=>"110111100",
  43033=>"010001101",
  43034=>"011011101",
  43035=>"010101111",
  43036=>"110110011",
  43037=>"101100011",
  43038=>"101100000",
  43039=>"000101011",
  43040=>"010111101",
  43041=>"110111100",
  43042=>"010111001",
  43043=>"101111000",
  43044=>"111110001",
  43045=>"110110011",
  43046=>"010011001",
  43047=>"100011010",
  43048=>"111110110",
  43049=>"101100001",
  43050=>"010110100",
  43051=>"101111000",
  43052=>"101101101",
  43053=>"101100010",
  43054=>"110100100",
  43055=>"011000000",
  43056=>"110111011",
  43057=>"111100101",
  43058=>"011000011",
  43059=>"010000101",
  43060=>"001000001",
  43061=>"100011000",
  43062=>"101111100",
  43063=>"000111111",
  43064=>"000001110",
  43065=>"010111010",
  43066=>"101101000",
  43067=>"101000110",
  43068=>"001111101",
  43069=>"110001100",
  43070=>"111100111",
  43071=>"010011011",
  43072=>"111000101",
  43073=>"010100001",
  43074=>"000000100",
  43075=>"001100110",
  43076=>"011011111",
  43077=>"110000100",
  43078=>"111100000",
  43079=>"100000110",
  43080=>"001011100",
  43081=>"111111111",
  43082=>"100010001",
  43083=>"011001011",
  43084=>"010001000",
  43085=>"100110100",
  43086=>"010010100",
  43087=>"001111010",
  43088=>"011111101",
  43089=>"000000010",
  43090=>"010111110",
  43091=>"110110111",
  43092=>"010010011",
  43093=>"101110100",
  43094=>"110011001",
  43095=>"110100101",
  43096=>"001011100",
  43097=>"100010011",
  43098=>"001110011",
  43099=>"111011110",
  43100=>"011001100",
  43101=>"010110110",
  43102=>"000111110",
  43103=>"000111000",
  43104=>"011111011",
  43105=>"000101100",
  43106=>"100011111",
  43107=>"001101101",
  43108=>"101011000",
  43109=>"101010010",
  43110=>"000110101",
  43111=>"001010111",
  43112=>"100001001",
  43113=>"001100101",
  43114=>"010101111",
  43115=>"111100001",
  43116=>"010110000",
  43117=>"001000011",
  43118=>"010100100",
  43119=>"000101101",
  43120=>"111011111",
  43121=>"001110011",
  43122=>"000001010",
  43123=>"110011110",
  43124=>"110111110",
  43125=>"100111111",
  43126=>"101110101",
  43127=>"000110111",
  43128=>"001001110",
  43129=>"010100010",
  43130=>"110110110",
  43131=>"001101001",
  43132=>"011001111",
  43133=>"111100010",
  43134=>"101101110",
  43135=>"001000010",
  43136=>"110001100",
  43137=>"011010011",
  43138=>"101011110",
  43139=>"010101010",
  43140=>"011001001",
  43141=>"111101010",
  43142=>"110010011",
  43143=>"001011111",
  43144=>"100011100",
  43145=>"101000110",
  43146=>"111100001",
  43147=>"101011101",
  43148=>"001010000",
  43149=>"010011000",
  43150=>"101001110",
  43151=>"101011011",
  43152=>"010101111",
  43153=>"100110101",
  43154=>"010110100",
  43155=>"101111100",
  43156=>"001001011",
  43157=>"011110010",
  43158=>"111101110",
  43159=>"101111101",
  43160=>"101000000",
  43161=>"100011111",
  43162=>"001110110",
  43163=>"000010001",
  43164=>"100010001",
  43165=>"111101100",
  43166=>"110100010",
  43167=>"011011111",
  43168=>"010111110",
  43169=>"110100000",
  43170=>"001011100",
  43171=>"110110111",
  43172=>"001110010",
  43173=>"001011010",
  43174=>"000110101",
  43175=>"110100110",
  43176=>"110000101",
  43177=>"000101000",
  43178=>"011011010",
  43179=>"110001010",
  43180=>"111111010",
  43181=>"000100110",
  43182=>"001100101",
  43183=>"101111011",
  43184=>"011001110",
  43185=>"101110100",
  43186=>"011101101",
  43187=>"110010010",
  43188=>"101010001",
  43189=>"010011110",
  43190=>"000111001",
  43191=>"000101000",
  43192=>"101010100",
  43193=>"010100000",
  43194=>"010010110",
  43195=>"011111001",
  43196=>"111001000",
  43197=>"110100100",
  43198=>"010110100",
  43199=>"110101000",
  43200=>"110110000",
  43201=>"100100011",
  43202=>"110111110",
  43203=>"101111010",
  43204=>"110100011",
  43205=>"010001010",
  43206=>"010001000",
  43207=>"100111001",
  43208=>"000110010",
  43209=>"110001110",
  43210=>"110010100",
  43211=>"100011110",
  43212=>"110011110",
  43213=>"001000111",
  43214=>"100010110",
  43215=>"001100101",
  43216=>"101111110",
  43217=>"111100100",
  43218=>"000001100",
  43219=>"111101101",
  43220=>"010111000",
  43221=>"101001100",
  43222=>"101101000",
  43223=>"010100001",
  43224=>"110010111",
  43225=>"010101000",
  43226=>"010000011",
  43227=>"011010010",
  43228=>"110101000",
  43229=>"100111011",
  43230=>"001100010",
  43231=>"001000011",
  43232=>"011010001",
  43233=>"000010111",
  43234=>"001010000",
  43235=>"001001100",
  43236=>"111000101",
  43237=>"001010101",
  43238=>"001010001",
  43239=>"110011101",
  43240=>"100000010",
  43241=>"110011010",
  43242=>"111111000",
  43243=>"111011100",
  43244=>"111000000",
  43245=>"011001111",
  43246=>"011101110",
  43247=>"000100100",
  43248=>"011010000",
  43249=>"100110111",
  43250=>"001011110",
  43251=>"010010101",
  43252=>"100000010",
  43253=>"101011001",
  43254=>"110100001",
  43255=>"010010000",
  43256=>"011000111",
  43257=>"111011101",
  43258=>"111101110",
  43259=>"001100010",
  43260=>"000101100",
  43261=>"001100101",
  43262=>"001001100",
  43263=>"101010010",
  43264=>"001010011",
  43265=>"101011110",
  43266=>"110101111",
  43267=>"110000000",
  43268=>"001111000",
  43269=>"110000001",
  43270=>"010010100",
  43271=>"101101011",
  43272=>"101011001",
  43273=>"110010111",
  43274=>"011010110",
  43275=>"110000010",
  43276=>"100101100",
  43277=>"001110110",
  43278=>"111000011",
  43279=>"001001101",
  43280=>"101001010",
  43281=>"010111000",
  43282=>"100111111",
  43283=>"111011101",
  43284=>"101000000",
  43285=>"010100000",
  43286=>"001010100",
  43287=>"010010111",
  43288=>"000011000",
  43289=>"100011011",
  43290=>"011011010",
  43291=>"011011010",
  43292=>"001001101",
  43293=>"111010001",
  43294=>"101110000",
  43295=>"011110000",
  43296=>"000110001",
  43297=>"010000000",
  43298=>"111100111",
  43299=>"100100001",
  43300=>"100111010",
  43301=>"101011101",
  43302=>"001010010",
  43303=>"000011100",
  43304=>"010000010",
  43305=>"110111111",
  43306=>"100000010",
  43307=>"000001010",
  43308=>"100110011",
  43309=>"001101000",
  43310=>"111111000",
  43311=>"011110101",
  43312=>"111111001",
  43313=>"001010110",
  43314=>"110111100",
  43315=>"110111000",
  43316=>"111011001",
  43317=>"010011001",
  43318=>"001111000",
  43319=>"011101011",
  43320=>"001001000",
  43321=>"001001101",
  43322=>"000101111",
  43323=>"001000011",
  43324=>"001001000",
  43325=>"000111101",
  43326=>"001010101",
  43327=>"000100011",
  43328=>"110101010",
  43329=>"111110010",
  43330=>"000000001",
  43331=>"011101001",
  43332=>"000111000",
  43333=>"111100101",
  43334=>"010001110",
  43335=>"101011101",
  43336=>"011001001",
  43337=>"010000110",
  43338=>"100111001",
  43339=>"111011001",
  43340=>"100110000",
  43341=>"011100010",
  43342=>"110010010",
  43343=>"110111110",
  43344=>"011010011",
  43345=>"010010001",
  43346=>"111011110",
  43347=>"011101010",
  43348=>"110000100",
  43349=>"010010111",
  43350=>"110111110",
  43351=>"000110000",
  43352=>"001001100",
  43353=>"110101101",
  43354=>"100010000",
  43355=>"000111111",
  43356=>"011011100",
  43357=>"100111100",
  43358=>"001010010",
  43359=>"100101110",
  43360=>"010100010",
  43361=>"110011111",
  43362=>"010010011",
  43363=>"100100000",
  43364=>"100111001",
  43365=>"110000000",
  43366=>"111001000",
  43367=>"010100010",
  43368=>"110110011",
  43369=>"001000001",
  43370=>"100010011",
  43371=>"111111111",
  43372=>"100010001",
  43373=>"110111110",
  43374=>"011100100",
  43375=>"010111001",
  43376=>"000001010",
  43377=>"111001000",
  43378=>"011000101",
  43379=>"111010010",
  43380=>"011101111",
  43381=>"010001110",
  43382=>"001000000",
  43383=>"011101111",
  43384=>"001000010",
  43385=>"001110110",
  43386=>"011000000",
  43387=>"110100111",
  43388=>"000011000",
  43389=>"110110101",
  43390=>"101001011",
  43391=>"000100011",
  43392=>"110001011",
  43393=>"000010100",
  43394=>"111000101",
  43395=>"001010011",
  43396=>"000011011",
  43397=>"001100100",
  43398=>"101011111",
  43399=>"011101001",
  43400=>"110100000",
  43401=>"111101010",
  43402=>"000110100",
  43403=>"110011100",
  43404=>"110110100",
  43405=>"111110011",
  43406=>"010000101",
  43407=>"110100100",
  43408=>"011000000",
  43409=>"100101011",
  43410=>"010000101",
  43411=>"001000101",
  43412=>"011111000",
  43413=>"101110111",
  43414=>"100010010",
  43415=>"110001001",
  43416=>"001000011",
  43417=>"111111101",
  43418=>"000100111",
  43419=>"111111000",
  43420=>"101101111",
  43421=>"010100100",
  43422=>"011111001",
  43423=>"001011000",
  43424=>"111011100",
  43425=>"100100111",
  43426=>"101000111",
  43427=>"110100101",
  43428=>"100110011",
  43429=>"010001101",
  43430=>"011111001",
  43431=>"010011000",
  43432=>"101010111",
  43433=>"001001100",
  43434=>"010010001",
  43435=>"100001110",
  43436=>"111100101",
  43437=>"000110010",
  43438=>"100111010",
  43439=>"011100100",
  43440=>"011100011",
  43441=>"000000010",
  43442=>"010010100",
  43443=>"001100001",
  43444=>"101011011",
  43445=>"101000000",
  43446=>"101001100",
  43447=>"011101000",
  43448=>"111101000",
  43449=>"110100111",
  43450=>"000000101",
  43451=>"101100011",
  43452=>"100100111",
  43453=>"000010001",
  43454=>"101110010",
  43455=>"101111101",
  43456=>"001110110",
  43457=>"010011000",
  43458=>"000100010",
  43459=>"010010110",
  43460=>"111001110",
  43461=>"110101100",
  43462=>"010011101",
  43463=>"000001000",
  43464=>"111100011",
  43465=>"000111111",
  43466=>"001101000",
  43467=>"001010111",
  43468=>"001010001",
  43469=>"111100001",
  43470=>"001010101",
  43471=>"001000111",
  43472=>"011111001",
  43473=>"001011011",
  43474=>"011001100",
  43475=>"101100101",
  43476=>"001110111",
  43477=>"011001101",
  43478=>"000000011",
  43479=>"001111111",
  43480=>"000110110",
  43481=>"011101101",
  43482=>"010111011",
  43483=>"010110011",
  43484=>"001110000",
  43485=>"000101001",
  43486=>"011110000",
  43487=>"001010011",
  43488=>"000101100",
  43489=>"101011111",
  43490=>"010010101",
  43491=>"100110001",
  43492=>"101000001",
  43493=>"100000000",
  43494=>"110111110",
  43495=>"011110100",
  43496=>"111100010",
  43497=>"010010100",
  43498=>"011001001",
  43499=>"111011001",
  43500=>"010010100",
  43501=>"010010010",
  43502=>"000110101",
  43503=>"000100011",
  43504=>"010011110",
  43505=>"000100000",
  43506=>"010011000",
  43507=>"001011000",
  43508=>"010000111",
  43509=>"101001000",
  43510=>"011001010",
  43511=>"101000000",
  43512=>"110010000",
  43513=>"111110101",
  43514=>"000100001",
  43515=>"010000111",
  43516=>"110001001",
  43517=>"101101101",
  43518=>"110011010",
  43519=>"001001000",
  43520=>"101001110",
  43521=>"100111100",
  43522=>"101100100",
  43523=>"001100000",
  43524=>"001010110",
  43525=>"000010101",
  43526=>"011100001",
  43527=>"111110010",
  43528=>"001011110",
  43529=>"000110011",
  43530=>"101010000",
  43531=>"010000011",
  43532=>"111110111",
  43533=>"100111000",
  43534=>"001111111",
  43535=>"011100100",
  43536=>"111111001",
  43537=>"011110110",
  43538=>"011011111",
  43539=>"010100011",
  43540=>"101000010",
  43541=>"100011111",
  43542=>"110110101",
  43543=>"100101011",
  43544=>"010111111",
  43545=>"111000010",
  43546=>"100001110",
  43547=>"001001110",
  43548=>"111000001",
  43549=>"110101010",
  43550=>"001000000",
  43551=>"010101111",
  43552=>"111110101",
  43553=>"010011001",
  43554=>"010011001",
  43555=>"010101010",
  43556=>"010001011",
  43557=>"000010000",
  43558=>"111110111",
  43559=>"011000101",
  43560=>"001010110",
  43561=>"010011101",
  43562=>"000000110",
  43563=>"011000110",
  43564=>"101101010",
  43565=>"111110111",
  43566=>"011110010",
  43567=>"111110111",
  43568=>"110001001",
  43569=>"011100110",
  43570=>"101010011",
  43571=>"000101000",
  43572=>"010010110",
  43573=>"000110000",
  43574=>"101001101",
  43575=>"110111011",
  43576=>"111000000",
  43577=>"100110001",
  43578=>"011001100",
  43579=>"000000100",
  43580=>"101000011",
  43581=>"001101111",
  43582=>"001110000",
  43583=>"001101100",
  43584=>"000000001",
  43585=>"001110101",
  43586=>"001011011",
  43587=>"111000010",
  43588=>"111011010",
  43589=>"011001110",
  43590=>"110111111",
  43591=>"110010010",
  43592=>"100001001",
  43593=>"111000101",
  43594=>"010000011",
  43595=>"111110000",
  43596=>"111110011",
  43597=>"101010111",
  43598=>"100110111",
  43599=>"111010001",
  43600=>"111001111",
  43601=>"100110010",
  43602=>"000101111",
  43603=>"010000001",
  43604=>"100000010",
  43605=>"110000011",
  43606=>"011000011",
  43607=>"110110110",
  43608=>"001001001",
  43609=>"001111111",
  43610=>"001110001",
  43611=>"001001111",
  43612=>"000001000",
  43613=>"111110011",
  43614=>"010010011",
  43615=>"011001000",
  43616=>"110000010",
  43617=>"001110000",
  43618=>"101101010",
  43619=>"010011010",
  43620=>"111111011",
  43621=>"011110001",
  43622=>"000001111",
  43623=>"000101111",
  43624=>"001001110",
  43625=>"000101100",
  43626=>"101010000",
  43627=>"111110111",
  43628=>"000011111",
  43629=>"100100110",
  43630=>"101110111",
  43631=>"010101001",
  43632=>"110111101",
  43633=>"000010110",
  43634=>"010000001",
  43635=>"000100100",
  43636=>"101011111",
  43637=>"010000010",
  43638=>"010101000",
  43639=>"110100000",
  43640=>"101000101",
  43641=>"100011000",
  43642=>"000000001",
  43643=>"000100010",
  43644=>"100011010",
  43645=>"001000010",
  43646=>"111001000",
  43647=>"011101011",
  43648=>"101001110",
  43649=>"000101000",
  43650=>"001010101",
  43651=>"110000101",
  43652=>"111010000",
  43653=>"010011101",
  43654=>"010101110",
  43655=>"001001100",
  43656=>"110011001",
  43657=>"000000111",
  43658=>"010101111",
  43659=>"000100100",
  43660=>"110010101",
  43661=>"010000110",
  43662=>"110010011",
  43663=>"100111001",
  43664=>"101111011",
  43665=>"000011001",
  43666=>"100011011",
  43667=>"001101110",
  43668=>"000101001",
  43669=>"101001011",
  43670=>"011101100",
  43671=>"001100101",
  43672=>"001110000",
  43673=>"011011111",
  43674=>"000110000",
  43675=>"100011010",
  43676=>"001011000",
  43677=>"100111100",
  43678=>"111001011",
  43679=>"111001010",
  43680=>"111111101",
  43681=>"000010011",
  43682=>"101100010",
  43683=>"110010001",
  43684=>"000100011",
  43685=>"010111001",
  43686=>"100000110",
  43687=>"111010001",
  43688=>"011011110",
  43689=>"001010101",
  43690=>"011000100",
  43691=>"111000000",
  43692=>"101011111",
  43693=>"111010100",
  43694=>"000011100",
  43695=>"010001010",
  43696=>"000101110",
  43697=>"011111111",
  43698=>"011110001",
  43699=>"100101001",
  43700=>"000101011",
  43701=>"000110100",
  43702=>"010001000",
  43703=>"001111010",
  43704=>"001110000",
  43705=>"001000101",
  43706=>"001100100",
  43707=>"101100110",
  43708=>"101111101",
  43709=>"111010000",
  43710=>"000011111",
  43711=>"111110011",
  43712=>"101101101",
  43713=>"101011100",
  43714=>"001001101",
  43715=>"011001000",
  43716=>"000001000",
  43717=>"011100000",
  43718=>"110101100",
  43719=>"100100110",
  43720=>"101101111",
  43721=>"100010110",
  43722=>"100111010",
  43723=>"011100111",
  43724=>"000110010",
  43725=>"000011101",
  43726=>"100111111",
  43727=>"100001100",
  43728=>"001011100",
  43729=>"001110111",
  43730=>"100001111",
  43731=>"001001110",
  43732=>"101001101",
  43733=>"000000111",
  43734=>"000110100",
  43735=>"001111110",
  43736=>"111011011",
  43737=>"100011001",
  43738=>"111101101",
  43739=>"100000100",
  43740=>"100110100",
  43741=>"000010110",
  43742=>"101010110",
  43743=>"010001100",
  43744=>"010011001",
  43745=>"110111001",
  43746=>"010100010",
  43747=>"101110010",
  43748=>"000110011",
  43749=>"111001001",
  43750=>"000111010",
  43751=>"100100100",
  43752=>"001101100",
  43753=>"010010100",
  43754=>"111000000",
  43755=>"100101011",
  43756=>"010011001",
  43757=>"100110100",
  43758=>"101001111",
  43759=>"001100010",
  43760=>"011101000",
  43761=>"001101001",
  43762=>"011110110",
  43763=>"000101100",
  43764=>"111011111",
  43765=>"010001011",
  43766=>"111011100",
  43767=>"000111101",
  43768=>"110010100",
  43769=>"010000011",
  43770=>"100011110",
  43771=>"000000001",
  43772=>"111100011",
  43773=>"001001000",
  43774=>"111100001",
  43775=>"111001100",
  43776=>"010000101",
  43777=>"011100101",
  43778=>"100110111",
  43779=>"010000100",
  43780=>"011110010",
  43781=>"100000110",
  43782=>"101010100",
  43783=>"101000110",
  43784=>"101101010",
  43785=>"111000011",
  43786=>"101001100",
  43787=>"110110111",
  43788=>"000000001",
  43789=>"000011011",
  43790=>"001001000",
  43791=>"100011100",
  43792=>"000001011",
  43793=>"111110101",
  43794=>"111000011",
  43795=>"100011111",
  43796=>"100010111",
  43797=>"000111010",
  43798=>"101000001",
  43799=>"001011101",
  43800=>"100100100",
  43801=>"110111101",
  43802=>"010000110",
  43803=>"001101010",
  43804=>"110101001",
  43805=>"100001100",
  43806=>"110001101",
  43807=>"101101110",
  43808=>"110010111",
  43809=>"101101001",
  43810=>"101110000",
  43811=>"110000011",
  43812=>"101011101",
  43813=>"000100111",
  43814=>"001101110",
  43815=>"011000101",
  43816=>"000000101",
  43817=>"000000101",
  43818=>"101101111",
  43819=>"100100110",
  43820=>"011101010",
  43821=>"100010001",
  43822=>"110000101",
  43823=>"100110101",
  43824=>"000000010",
  43825=>"101110001",
  43826=>"000110011",
  43827=>"100101110",
  43828=>"101100011",
  43829=>"010001100",
  43830=>"100110011",
  43831=>"110000010",
  43832=>"010000111",
  43833=>"001101100",
  43834=>"000101001",
  43835=>"100000011",
  43836=>"101001010",
  43837=>"110010010",
  43838=>"111000000",
  43839=>"000110000",
  43840=>"110110011",
  43841=>"101110001",
  43842=>"110010010",
  43843=>"011111010",
  43844=>"010100000",
  43845=>"111001100",
  43846=>"100000101",
  43847=>"101001100",
  43848=>"000011000",
  43849=>"110011010",
  43850=>"010000110",
  43851=>"001101111",
  43852=>"111111110",
  43853=>"010010010",
  43854=>"110000110",
  43855=>"100011000",
  43856=>"001100110",
  43857=>"100011001",
  43858=>"100011011",
  43859=>"111001010",
  43860=>"111010000",
  43861=>"100101101",
  43862=>"000100100",
  43863=>"111101100",
  43864=>"111010111",
  43865=>"010101001",
  43866=>"010000000",
  43867=>"111010011",
  43868=>"011011011",
  43869=>"111111001",
  43870=>"000000011",
  43871=>"011010100",
  43872=>"000101111",
  43873=>"101100111",
  43874=>"001011011",
  43875=>"101100000",
  43876=>"110101101",
  43877=>"111100111",
  43878=>"010001110",
  43879=>"011110001",
  43880=>"110100000",
  43881=>"100011110",
  43882=>"011110001",
  43883=>"111001110",
  43884=>"110010000",
  43885=>"011100000",
  43886=>"101100111",
  43887=>"011100110",
  43888=>"000000000",
  43889=>"111110100",
  43890=>"000011100",
  43891=>"101001010",
  43892=>"110000010",
  43893=>"110010010",
  43894=>"010111011",
  43895=>"001110111",
  43896=>"100001101",
  43897=>"011010101",
  43898=>"010010100",
  43899=>"101010100",
  43900=>"000100110",
  43901=>"110001101",
  43902=>"000000011",
  43903=>"011101001",
  43904=>"110101111",
  43905=>"100100111",
  43906=>"110101010",
  43907=>"100011101",
  43908=>"000000011",
  43909=>"100000100",
  43910=>"101110111",
  43911=>"100010110",
  43912=>"000011100",
  43913=>"100000000",
  43914=>"011000011",
  43915=>"111101011",
  43916=>"001001111",
  43917=>"110101101",
  43918=>"000101100",
  43919=>"001110100",
  43920=>"111111101",
  43921=>"001101000",
  43922=>"110100001",
  43923=>"001100111",
  43924=>"100000000",
  43925=>"001101001",
  43926=>"011101111",
  43927=>"011101010",
  43928=>"001000110",
  43929=>"011110010",
  43930=>"000111110",
  43931=>"010100101",
  43932=>"000000110",
  43933=>"010001000",
  43934=>"000100110",
  43935=>"011111001",
  43936=>"101100110",
  43937=>"101010000",
  43938=>"000111111",
  43939=>"011011100",
  43940=>"001110011",
  43941=>"111100101",
  43942=>"100000011",
  43943=>"001111111",
  43944=>"010100100",
  43945=>"000011000",
  43946=>"001100111",
  43947=>"111001000",
  43948=>"110101010",
  43949=>"010000101",
  43950=>"111001001",
  43951=>"011000111",
  43952=>"011010101",
  43953=>"001011101",
  43954=>"010000010",
  43955=>"100100010",
  43956=>"110010010",
  43957=>"111111101",
  43958=>"001001110",
  43959=>"110111111",
  43960=>"011000000",
  43961=>"100000111",
  43962=>"100010111",
  43963=>"111011110",
  43964=>"100010001",
  43965=>"001111001",
  43966=>"110101010",
  43967=>"000000100",
  43968=>"010100010",
  43969=>"110100110",
  43970=>"001100111",
  43971=>"001011111",
  43972=>"111010101",
  43973=>"101001000",
  43974=>"001100111",
  43975=>"100100000",
  43976=>"110110111",
  43977=>"011101100",
  43978=>"100111011",
  43979=>"000110011",
  43980=>"110110110",
  43981=>"101100110",
  43982=>"010000000",
  43983=>"001000010",
  43984=>"111100010",
  43985=>"111001011",
  43986=>"010000001",
  43987=>"110101001",
  43988=>"101101000",
  43989=>"001101001",
  43990=>"000101010",
  43991=>"011001011",
  43992=>"101000101",
  43993=>"111111110",
  43994=>"100101001",
  43995=>"111011010",
  43996=>"111101111",
  43997=>"000011111",
  43998=>"010010101",
  43999=>"111011111",
  44000=>"111111111",
  44001=>"000001110",
  44002=>"111101101",
  44003=>"000001001",
  44004=>"000010101",
  44005=>"011110110",
  44006=>"111010110",
  44007=>"011010001",
  44008=>"000110010",
  44009=>"111101110",
  44010=>"100011100",
  44011=>"100101101",
  44012=>"111101110",
  44013=>"011010111",
  44014=>"001000110",
  44015=>"111010110",
  44016=>"111111100",
  44017=>"101100010",
  44018=>"110110111",
  44019=>"111100100",
  44020=>"000010001",
  44021=>"101111011",
  44022=>"000010100",
  44023=>"101111001",
  44024=>"010100100",
  44025=>"011011110",
  44026=>"101000001",
  44027=>"010001000",
  44028=>"000001110",
  44029=>"011100100",
  44030=>"100011010",
  44031=>"001000101",
  44032=>"001110101",
  44033=>"110111001",
  44034=>"111000011",
  44035=>"000111000",
  44036=>"010010100",
  44037=>"000000111",
  44038=>"010101000",
  44039=>"111101001",
  44040=>"110101010",
  44041=>"110010100",
  44042=>"010101000",
  44043=>"100110011",
  44044=>"010001110",
  44045=>"111100011",
  44046=>"001001010",
  44047=>"110011000",
  44048=>"011100001",
  44049=>"100001111",
  44050=>"111000000",
  44051=>"110110111",
  44052=>"011100011",
  44053=>"111000110",
  44054=>"000100000",
  44055=>"010000001",
  44056=>"011011010",
  44057=>"011001111",
  44058=>"111101101",
  44059=>"000010101",
  44060=>"001001011",
  44061=>"000111111",
  44062=>"110010110",
  44063=>"010000101",
  44064=>"000010010",
  44065=>"010001011",
  44066=>"110101000",
  44067=>"111100101",
  44068=>"011110101",
  44069=>"100000100",
  44070=>"100101010",
  44071=>"110001111",
  44072=>"010101111",
  44073=>"001000001",
  44074=>"000110100",
  44075=>"101100111",
  44076=>"011010011",
  44077=>"001110010",
  44078=>"010000001",
  44079=>"110110001",
  44080=>"101100001",
  44081=>"011000111",
  44082=>"011010100",
  44083=>"110100011",
  44084=>"110001110",
  44085=>"011111000",
  44086=>"110011100",
  44087=>"111101010",
  44088=>"000011101",
  44089=>"111111010",
  44090=>"000000010",
  44091=>"000001000",
  44092=>"000011010",
  44093=>"011011111",
  44094=>"101101101",
  44095=>"010011101",
  44096=>"010101111",
  44097=>"000001111",
  44098=>"100101111",
  44099=>"100001101",
  44100=>"100011011",
  44101=>"110101110",
  44102=>"110111110",
  44103=>"110101011",
  44104=>"111110001",
  44105=>"010000101",
  44106=>"011011111",
  44107=>"011011110",
  44108=>"000101000",
  44109=>"100100010",
  44110=>"101111010",
  44111=>"110110110",
  44112=>"101011101",
  44113=>"010001010",
  44114=>"000111111",
  44115=>"110000010",
  44116=>"000111101",
  44117=>"001101101",
  44118=>"011110011",
  44119=>"011110111",
  44120=>"100111100",
  44121=>"010001100",
  44122=>"000010110",
  44123=>"000001010",
  44124=>"101111111",
  44125=>"010111001",
  44126=>"010011111",
  44127=>"100011110",
  44128=>"000001011",
  44129=>"001101101",
  44130=>"001111001",
  44131=>"100001011",
  44132=>"001001101",
  44133=>"110101011",
  44134=>"001111000",
  44135=>"000101000",
  44136=>"000000110",
  44137=>"011100010",
  44138=>"000000011",
  44139=>"010011011",
  44140=>"001011011",
  44141=>"001001010",
  44142=>"110111010",
  44143=>"100111100",
  44144=>"011101000",
  44145=>"000001000",
  44146=>"101000000",
  44147=>"110111110",
  44148=>"101001011",
  44149=>"111110110",
  44150=>"011010010",
  44151=>"110100001",
  44152=>"000110110",
  44153=>"001101010",
  44154=>"101000000",
  44155=>"100001000",
  44156=>"100001110",
  44157=>"001011100",
  44158=>"001011101",
  44159=>"010110011",
  44160=>"111101101",
  44161=>"101000100",
  44162=>"100101101",
  44163=>"100001101",
  44164=>"101011101",
  44165=>"101010001",
  44166=>"001100011",
  44167=>"101111011",
  44168=>"010110110",
  44169=>"001101101",
  44170=>"001100100",
  44171=>"000011111",
  44172=>"110110001",
  44173=>"101000011",
  44174=>"011111101",
  44175=>"010100001",
  44176=>"000010001",
  44177=>"111010110",
  44178=>"110111110",
  44179=>"010101011",
  44180=>"111000110",
  44181=>"001000111",
  44182=>"001111000",
  44183=>"111001110",
  44184=>"111110100",
  44185=>"111100001",
  44186=>"000010011",
  44187=>"110000100",
  44188=>"110011100",
  44189=>"010111001",
  44190=>"000110010",
  44191=>"011011110",
  44192=>"111111011",
  44193=>"111101101",
  44194=>"101000011",
  44195=>"101000100",
  44196=>"111011101",
  44197=>"001100011",
  44198=>"000000001",
  44199=>"110101101",
  44200=>"111001001",
  44201=>"000000000",
  44202=>"111010110",
  44203=>"000110101",
  44204=>"111110110",
  44205=>"111001000",
  44206=>"111100100",
  44207=>"010100011",
  44208=>"000101001",
  44209=>"100111110",
  44210=>"100111001",
  44211=>"110001001",
  44212=>"010111111",
  44213=>"100101000",
  44214=>"111100010",
  44215=>"111110110",
  44216=>"011110011",
  44217=>"011111001",
  44218=>"011110000",
  44219=>"000011010",
  44220=>"011001111",
  44221=>"010001111",
  44222=>"101100011",
  44223=>"110000000",
  44224=>"101111101",
  44225=>"101011000",
  44226=>"000000001",
  44227=>"001100111",
  44228=>"001000101",
  44229=>"110101001",
  44230=>"100111111",
  44231=>"100001001",
  44232=>"000011001",
  44233=>"111010100",
  44234=>"011001110",
  44235=>"010100100",
  44236=>"111101110",
  44237=>"111001001",
  44238=>"010000111",
  44239=>"010010101",
  44240=>"011100010",
  44241=>"111111011",
  44242=>"110010111",
  44243=>"011111111",
  44244=>"101100000",
  44245=>"100011100",
  44246=>"010101101",
  44247=>"011001101",
  44248=>"011100110",
  44249=>"001111101",
  44250=>"101001111",
  44251=>"101100011",
  44252=>"100010101",
  44253=>"000110100",
  44254=>"001010101",
  44255=>"011010110",
  44256=>"100011010",
  44257=>"101011010",
  44258=>"111001001",
  44259=>"010001110",
  44260=>"001110001",
  44261=>"100010010",
  44262=>"110001101",
  44263=>"000111001",
  44264=>"101111110",
  44265=>"100001001",
  44266=>"000101011",
  44267=>"100011100",
  44268=>"100100000",
  44269=>"111101010",
  44270=>"100110100",
  44271=>"001110111",
  44272=>"010111110",
  44273=>"111111101",
  44274=>"000010000",
  44275=>"000101101",
  44276=>"111101110",
  44277=>"111111100",
  44278=>"001110110",
  44279=>"100100000",
  44280=>"101111110",
  44281=>"011111111",
  44282=>"010011100",
  44283=>"100100100",
  44284=>"011010000",
  44285=>"000111000",
  44286=>"101010110",
  44287=>"010011011",
  44288=>"110100011",
  44289=>"100001101",
  44290=>"110011001",
  44291=>"000100110",
  44292=>"000110000",
  44293=>"010010010",
  44294=>"000101001",
  44295=>"001101111",
  44296=>"111001101",
  44297=>"010111011",
  44298=>"111101110",
  44299=>"101001000",
  44300=>"001111000",
  44301=>"100000010",
  44302=>"000010001",
  44303=>"010110100",
  44304=>"000001111",
  44305=>"110001011",
  44306=>"100011100",
  44307=>"111110000",
  44308=>"111111010",
  44309=>"001111000",
  44310=>"100000101",
  44311=>"110010001",
  44312=>"101101000",
  44313=>"111100001",
  44314=>"111011110",
  44315=>"100111111",
  44316=>"000010111",
  44317=>"111000010",
  44318=>"110010100",
  44319=>"011101001",
  44320=>"000110001",
  44321=>"101000011",
  44322=>"000000001",
  44323=>"101111111",
  44324=>"001100111",
  44325=>"010001011",
  44326=>"001100101",
  44327=>"101101101",
  44328=>"110010110",
  44329=>"000101110",
  44330=>"101101001",
  44331=>"111101011",
  44332=>"010011110",
  44333=>"111010101",
  44334=>"101000001",
  44335=>"101010100",
  44336=>"010000011",
  44337=>"110001011",
  44338=>"110011100",
  44339=>"010000111",
  44340=>"110000010",
  44341=>"111101100",
  44342=>"001000100",
  44343=>"100111000",
  44344=>"101101111",
  44345=>"100011101",
  44346=>"010110110",
  44347=>"110101101",
  44348=>"001111001",
  44349=>"100010000",
  44350=>"101011011",
  44351=>"100100000",
  44352=>"000110111",
  44353=>"000000100",
  44354=>"010010000",
  44355=>"111111100",
  44356=>"000001011",
  44357=>"010100101",
  44358=>"100110001",
  44359=>"100011000",
  44360=>"110111001",
  44361=>"011100000",
  44362=>"011010111",
  44363=>"001101111",
  44364=>"101000001",
  44365=>"110111111",
  44366=>"110011011",
  44367=>"100011111",
  44368=>"001010011",
  44369=>"001111000",
  44370=>"111001011",
  44371=>"110101101",
  44372=>"110111110",
  44373=>"011000001",
  44374=>"111010100",
  44375=>"110011110",
  44376=>"001101111",
  44377=>"110111101",
  44378=>"001011101",
  44379=>"010100000",
  44380=>"011111000",
  44381=>"001001111",
  44382=>"001111000",
  44383=>"000110010",
  44384=>"010111000",
  44385=>"111000001",
  44386=>"001001110",
  44387=>"001001110",
  44388=>"011111100",
  44389=>"100101011",
  44390=>"110011001",
  44391=>"101011100",
  44392=>"100101010",
  44393=>"100101001",
  44394=>"101101001",
  44395=>"110000101",
  44396=>"100111001",
  44397=>"110101111",
  44398=>"001100001",
  44399=>"011001101",
  44400=>"000101110",
  44401=>"100010100",
  44402=>"111100101",
  44403=>"011011000",
  44404=>"001010011",
  44405=>"100111001",
  44406=>"011100000",
  44407=>"010011001",
  44408=>"011110001",
  44409=>"101111100",
  44410=>"010000100",
  44411=>"100010111",
  44412=>"010110111",
  44413=>"100110010",
  44414=>"010101000",
  44415=>"001011000",
  44416=>"001010001",
  44417=>"001000110",
  44418=>"011110111",
  44419=>"000000110",
  44420=>"110101111",
  44421=>"001110100",
  44422=>"110101011",
  44423=>"000010110",
  44424=>"100000000",
  44425=>"111010010",
  44426=>"111100111",
  44427=>"011110111",
  44428=>"011011010",
  44429=>"000101110",
  44430=>"010101111",
  44431=>"110110101",
  44432=>"001110111",
  44433=>"100010010",
  44434=>"010101100",
  44435=>"011101111",
  44436=>"110111111",
  44437=>"010101110",
  44438=>"010111011",
  44439=>"001001010",
  44440=>"010001010",
  44441=>"101111011",
  44442=>"100111011",
  44443=>"001000000",
  44444=>"010011011",
  44445=>"110011000",
  44446=>"010110101",
  44447=>"000110010",
  44448=>"101011100",
  44449=>"011011111",
  44450=>"111110010",
  44451=>"111101111",
  44452=>"111001101",
  44453=>"010011101",
  44454=>"110011000",
  44455=>"110001001",
  44456=>"100110000",
  44457=>"011111000",
  44458=>"000011000",
  44459=>"100100010",
  44460=>"010000011",
  44461=>"110101001",
  44462=>"111010000",
  44463=>"010110100",
  44464=>"110100000",
  44465=>"101000100",
  44466=>"001010110",
  44467=>"011110001",
  44468=>"001101001",
  44469=>"101000110",
  44470=>"011100011",
  44471=>"011000110",
  44472=>"001001001",
  44473=>"101100110",
  44474=>"100110000",
  44475=>"100101011",
  44476=>"001111100",
  44477=>"101001110",
  44478=>"111100001",
  44479=>"111001001",
  44480=>"010000110",
  44481=>"001101110",
  44482=>"101111001",
  44483=>"011100111",
  44484=>"001010010",
  44485=>"100000110",
  44486=>"000000100",
  44487=>"110110001",
  44488=>"100101100",
  44489=>"001010111",
  44490=>"011010000",
  44491=>"111101000",
  44492=>"111101101",
  44493=>"010101000",
  44494=>"101000111",
  44495=>"111111111",
  44496=>"100010100",
  44497=>"011011111",
  44498=>"100101110",
  44499=>"011000001",
  44500=>"010011100",
  44501=>"110010000",
  44502=>"100000000",
  44503=>"001010010",
  44504=>"011111101",
  44505=>"110100010",
  44506=>"111110001",
  44507=>"111011110",
  44508=>"010100100",
  44509=>"110011110",
  44510=>"101100000",
  44511=>"101001101",
  44512=>"111110110",
  44513=>"100000110",
  44514=>"001011100",
  44515=>"110011101",
  44516=>"010001011",
  44517=>"111011111",
  44518=>"111101111",
  44519=>"111010101",
  44520=>"011000100",
  44521=>"100010000",
  44522=>"010001010",
  44523=>"100001100",
  44524=>"001011000",
  44525=>"000101100",
  44526=>"000110011",
  44527=>"110011100",
  44528=>"011000011",
  44529=>"011101101",
  44530=>"101100100",
  44531=>"010111001",
  44532=>"101001110",
  44533=>"100110000",
  44534=>"010000100",
  44535=>"100000001",
  44536=>"000000010",
  44537=>"011101111",
  44538=>"001010100",
  44539=>"111110110",
  44540=>"011001111",
  44541=>"000110111",
  44542=>"100001110",
  44543=>"001000011",
  44544=>"110011010",
  44545=>"100101101",
  44546=>"000001010",
  44547=>"110001010",
  44548=>"100001110",
  44549=>"000111100",
  44550=>"001100110",
  44551=>"010010001",
  44552=>"010010100",
  44553=>"000111001",
  44554=>"001011111",
  44555=>"101000010",
  44556=>"001100110",
  44557=>"100111000",
  44558=>"000000011",
  44559=>"101001111",
  44560=>"011010101",
  44561=>"010111000",
  44562=>"111010110",
  44563=>"111111010",
  44564=>"110100111",
  44565=>"000011000",
  44566=>"010111011",
  44567=>"111110000",
  44568=>"010100011",
  44569=>"011111111",
  44570=>"010001110",
  44571=>"111111111",
  44572=>"101100100",
  44573=>"100011011",
  44574=>"001011111",
  44575=>"101001101",
  44576=>"010110100",
  44577=>"110100100",
  44578=>"001110000",
  44579=>"101111100",
  44580=>"110111110",
  44581=>"010001010",
  44582=>"010111000",
  44583=>"100111001",
  44584=>"100000110",
  44585=>"111101011",
  44586=>"100110011",
  44587=>"110100111",
  44588=>"000011001",
  44589=>"011101001",
  44590=>"010011000",
  44591=>"111000001",
  44592=>"110111010",
  44593=>"011100111",
  44594=>"111111111",
  44595=>"101011011",
  44596=>"101011101",
  44597=>"100010101",
  44598=>"001111111",
  44599=>"000101001",
  44600=>"110100111",
  44601=>"100110001",
  44602=>"111000000",
  44603=>"100100101",
  44604=>"111111101",
  44605=>"001001000",
  44606=>"010011110",
  44607=>"100101011",
  44608=>"010111001",
  44609=>"000000001",
  44610=>"010011010",
  44611=>"110111111",
  44612=>"111000100",
  44613=>"111111110",
  44614=>"110111101",
  44615=>"100010010",
  44616=>"000111000",
  44617=>"110000001",
  44618=>"000110101",
  44619=>"101011001",
  44620=>"001101010",
  44621=>"010111010",
  44622=>"101001001",
  44623=>"011101001",
  44624=>"000001001",
  44625=>"110001111",
  44626=>"110000010",
  44627=>"101001111",
  44628=>"011101011",
  44629=>"001011101",
  44630=>"101001000",
  44631=>"010001101",
  44632=>"000111001",
  44633=>"011110000",
  44634=>"001001001",
  44635=>"000101000",
  44636=>"111010001",
  44637=>"001110100",
  44638=>"001011110",
  44639=>"010111000",
  44640=>"001000001",
  44641=>"010000000",
  44642=>"011001010",
  44643=>"110011101",
  44644=>"011010000",
  44645=>"101101100",
  44646=>"011010111",
  44647=>"001110001",
  44648=>"100001101",
  44649=>"110100011",
  44650=>"100001111",
  44651=>"101110111",
  44652=>"110110100",
  44653=>"110110110",
  44654=>"110111100",
  44655=>"101111000",
  44656=>"000100111",
  44657=>"100001110",
  44658=>"111001110",
  44659=>"111101011",
  44660=>"011110000",
  44661=>"011010011",
  44662=>"110000100",
  44663=>"100000001",
  44664=>"010011000",
  44665=>"100001100",
  44666=>"100010001",
  44667=>"100111111",
  44668=>"101010010",
  44669=>"101101000",
  44670=>"010111100",
  44671=>"100011010",
  44672=>"010110011",
  44673=>"110000011",
  44674=>"010111111",
  44675=>"010000110",
  44676=>"001011011",
  44677=>"001001100",
  44678=>"011100011",
  44679=>"001001000",
  44680=>"010101110",
  44681=>"000010110",
  44682=>"011011001",
  44683=>"110011011",
  44684=>"000000110",
  44685=>"111000000",
  44686=>"111110010",
  44687=>"110000100",
  44688=>"011011000",
  44689=>"001100100",
  44690=>"001011100",
  44691=>"010010000",
  44692=>"000011101",
  44693=>"001001011",
  44694=>"101001010",
  44695=>"101101010",
  44696=>"111011100",
  44697=>"111000101",
  44698=>"111001000",
  44699=>"010101001",
  44700=>"001010001",
  44701=>"010111010",
  44702=>"001000000",
  44703=>"011101111",
  44704=>"011101110",
  44705=>"101010111",
  44706=>"001101001",
  44707=>"010110110",
  44708=>"000101100",
  44709=>"100100111",
  44710=>"111100000",
  44711=>"011100100",
  44712=>"010110101",
  44713=>"011110001",
  44714=>"111001011",
  44715=>"010000001",
  44716=>"111010010",
  44717=>"101001100",
  44718=>"010011001",
  44719=>"111001111",
  44720=>"000111010",
  44721=>"111000110",
  44722=>"011000011",
  44723=>"110100010",
  44724=>"011111011",
  44725=>"100100011",
  44726=>"111011101",
  44727=>"110010100",
  44728=>"110001011",
  44729=>"100010011",
  44730=>"100001101",
  44731=>"000111111",
  44732=>"001011001",
  44733=>"001010001",
  44734=>"000110000",
  44735=>"100100010",
  44736=>"000111101",
  44737=>"100110110",
  44738=>"011111100",
  44739=>"001011100",
  44740=>"010010001",
  44741=>"101101010",
  44742=>"010011110",
  44743=>"100110000",
  44744=>"000000001",
  44745=>"111011000",
  44746=>"000011111",
  44747=>"001011101",
  44748=>"000101101",
  44749=>"110000011",
  44750=>"011011100",
  44751=>"110000011",
  44752=>"011011011",
  44753=>"001100011",
  44754=>"111001110",
  44755=>"000100111",
  44756=>"010101010",
  44757=>"101101000",
  44758=>"011111110",
  44759=>"000000101",
  44760=>"001111010",
  44761=>"010000001",
  44762=>"101100000",
  44763=>"100110001",
  44764=>"101100111",
  44765=>"101110010",
  44766=>"100010011",
  44767=>"000011100",
  44768=>"110010000",
  44769=>"011101111",
  44770=>"010011000",
  44771=>"011011100",
  44772=>"001011101",
  44773=>"100011111",
  44774=>"001001100",
  44775=>"000001000",
  44776=>"101000111",
  44777=>"100000010",
  44778=>"111000011",
  44779=>"110001111",
  44780=>"000011100",
  44781=>"001001001",
  44782=>"110111110",
  44783=>"011010100",
  44784=>"000001010",
  44785=>"100101101",
  44786=>"100111101",
  44787=>"110001101",
  44788=>"011011100",
  44789=>"110001000",
  44790=>"011011010",
  44791=>"101010001",
  44792=>"110101000",
  44793=>"110010111",
  44794=>"001110101",
  44795=>"000011010",
  44796=>"110000010",
  44797=>"111010011",
  44798=>"111010011",
  44799=>"000101000",
  44800=>"011001010",
  44801=>"000011000",
  44802=>"010011111",
  44803=>"001110101",
  44804=>"000110011",
  44805=>"111000100",
  44806=>"011100100",
  44807=>"100011000",
  44808=>"100000010",
  44809=>"010100001",
  44810=>"110100111",
  44811=>"010111111",
  44812=>"111100011",
  44813=>"101110101",
  44814=>"000110101",
  44815=>"010011111",
  44816=>"001101111",
  44817=>"010110010",
  44818=>"010100100",
  44819=>"111100010",
  44820=>"010111001",
  44821=>"001110001",
  44822=>"101111001",
  44823=>"011000100",
  44824=>"000001000",
  44825=>"101001001",
  44826=>"000110100",
  44827=>"010000111",
  44828=>"000010100",
  44829=>"110111010",
  44830=>"000000110",
  44831=>"010000000",
  44832=>"100101110",
  44833=>"110101010",
  44834=>"100111011",
  44835=>"001011111",
  44836=>"001011011",
  44837=>"100110011",
  44838=>"111011001",
  44839=>"011100101",
  44840=>"001101100",
  44841=>"001010100",
  44842=>"000100000",
  44843=>"111100010",
  44844=>"111011011",
  44845=>"101010111",
  44846=>"101011001",
  44847=>"001000010",
  44848=>"100111011",
  44849=>"110000110",
  44850=>"010100001",
  44851=>"110000100",
  44852=>"000101000",
  44853=>"100110110",
  44854=>"011010101",
  44855=>"011010110",
  44856=>"111011001",
  44857=>"000010111",
  44858=>"000111101",
  44859=>"111011110",
  44860=>"110000001",
  44861=>"001011001",
  44862=>"010010110",
  44863=>"011001101",
  44864=>"100111010",
  44865=>"001110110",
  44866=>"001010011",
  44867=>"001100000",
  44868=>"011000101",
  44869=>"011001010",
  44870=>"110011010",
  44871=>"000000010",
  44872=>"011001101",
  44873=>"111000100",
  44874=>"010111111",
  44875=>"011101011",
  44876=>"011100010",
  44877=>"101110101",
  44878=>"010000000",
  44879=>"110011010",
  44880=>"111101110",
  44881=>"110100111",
  44882=>"111000011",
  44883=>"000010010",
  44884=>"100000110",
  44885=>"010111010",
  44886=>"101011110",
  44887=>"010110100",
  44888=>"010011000",
  44889=>"010100000",
  44890=>"111001011",
  44891=>"111011000",
  44892=>"111000010",
  44893=>"101100100",
  44894=>"000000000",
  44895=>"000100110",
  44896=>"110001111",
  44897=>"011100001",
  44898=>"001010111",
  44899=>"001000101",
  44900=>"000100110",
  44901=>"010101111",
  44902=>"110011100",
  44903=>"010111010",
  44904=>"001011000",
  44905=>"001110000",
  44906=>"010011101",
  44907=>"010011010",
  44908=>"011010010",
  44909=>"000100110",
  44910=>"001110001",
  44911=>"111010101",
  44912=>"001010001",
  44913=>"110100000",
  44914=>"010001101",
  44915=>"000011110",
  44916=>"101010001",
  44917=>"100110011",
  44918=>"010111110",
  44919=>"010110011",
  44920=>"111110111",
  44921=>"011110010",
  44922=>"111011010",
  44923=>"111011000",
  44924=>"011110010",
  44925=>"101100100",
  44926=>"010001011",
  44927=>"111011011",
  44928=>"101111111",
  44929=>"000110111",
  44930=>"000010000",
  44931=>"101111011",
  44932=>"001010000",
  44933=>"110000100",
  44934=>"100001101",
  44935=>"100001010",
  44936=>"010111010",
  44937=>"101100000",
  44938=>"001111000",
  44939=>"101001010",
  44940=>"000111011",
  44941=>"000100001",
  44942=>"001110010",
  44943=>"000111110",
  44944=>"001001000",
  44945=>"000011001",
  44946=>"010010110",
  44947=>"000010011",
  44948=>"011100101",
  44949=>"001111011",
  44950=>"110001010",
  44951=>"000010100",
  44952=>"101111000",
  44953=>"100000101",
  44954=>"100111011",
  44955=>"011110001",
  44956=>"011110110",
  44957=>"110001101",
  44958=>"101010011",
  44959=>"011000101",
  44960=>"101110001",
  44961=>"100111000",
  44962=>"000010000",
  44963=>"111011010",
  44964=>"110010110",
  44965=>"010101111",
  44966=>"111111010",
  44967=>"111110000",
  44968=>"101110000",
  44969=>"110110101",
  44970=>"100010111",
  44971=>"011100000",
  44972=>"110010001",
  44973=>"111011010",
  44974=>"101110101",
  44975=>"010001110",
  44976=>"101010011",
  44977=>"001100011",
  44978=>"100110011",
  44979=>"010100001",
  44980=>"011011101",
  44981=>"111110111",
  44982=>"111110100",
  44983=>"001110110",
  44984=>"000110000",
  44985=>"101000010",
  44986=>"110111000",
  44987=>"111111011",
  44988=>"000111001",
  44989=>"101100001",
  44990=>"100101001",
  44991=>"010001010",
  44992=>"001001101",
  44993=>"001100110",
  44994=>"101111011",
  44995=>"101110010",
  44996=>"110001011",
  44997=>"011011000",
  44998=>"111110001",
  44999=>"011001111",
  45000=>"101001110",
  45001=>"000000000",
  45002=>"010010001",
  45003=>"110100111",
  45004=>"100001111",
  45005=>"110011100",
  45006=>"100000111",
  45007=>"101100100",
  45008=>"001110100",
  45009=>"010000110",
  45010=>"100001011",
  45011=>"000100000",
  45012=>"000010101",
  45013=>"000101010",
  45014=>"110100111",
  45015=>"000011100",
  45016=>"010010101",
  45017=>"010101010",
  45018=>"111110001",
  45019=>"111100000",
  45020=>"111010000",
  45021=>"010010011",
  45022=>"101011111",
  45023=>"011110000",
  45024=>"101011001",
  45025=>"111001000",
  45026=>"100110001",
  45027=>"100010000",
  45028=>"100100001",
  45029=>"100000001",
  45030=>"100101100",
  45031=>"001100010",
  45032=>"100100111",
  45033=>"001010010",
  45034=>"101001100",
  45035=>"101100010",
  45036=>"001100110",
  45037=>"111001100",
  45038=>"101110110",
  45039=>"101010011",
  45040=>"000000101",
  45041=>"110011000",
  45042=>"010000010",
  45043=>"011100000",
  45044=>"000100001",
  45045=>"110011010",
  45046=>"000100000",
  45047=>"001111001",
  45048=>"110111101",
  45049=>"111011101",
  45050=>"111000100",
  45051=>"101011110",
  45052=>"101000010",
  45053=>"101100001",
  45054=>"001110100",
  45055=>"001111000",
  45056=>"100001111",
  45057=>"000110110",
  45058=>"101111011",
  45059=>"001000101",
  45060=>"011001111",
  45061=>"000001110",
  45062=>"000111110",
  45063=>"001111001",
  45064=>"111010000",
  45065=>"111000100",
  45066=>"111010000",
  45067=>"100000101",
  45068=>"100001000",
  45069=>"010111010",
  45070=>"111010110",
  45071=>"111111100",
  45072=>"001100111",
  45073=>"001100100",
  45074=>"110010101",
  45075=>"111110101",
  45076=>"110101001",
  45077=>"110011100",
  45078=>"111111100",
  45079=>"000101010",
  45080=>"100011101",
  45081=>"001101110",
  45082=>"000011011",
  45083=>"011111101",
  45084=>"111011011",
  45085=>"101100010",
  45086=>"101110010",
  45087=>"000101100",
  45088=>"110100011",
  45089=>"110110001",
  45090=>"101100001",
  45091=>"101000000",
  45092=>"110000011",
  45093=>"100100101",
  45094=>"000010011",
  45095=>"001010111",
  45096=>"101101111",
  45097=>"111000111",
  45098=>"100100111",
  45099=>"001110000",
  45100=>"000101010",
  45101=>"000100110",
  45102=>"000010011",
  45103=>"001101110",
  45104=>"100110001",
  45105=>"100101110",
  45106=>"011110100",
  45107=>"111000000",
  45108=>"100000001",
  45109=>"000100001",
  45110=>"110100110",
  45111=>"111001110",
  45112=>"000010110",
  45113=>"101100111",
  45114=>"100010110",
  45115=>"011000101",
  45116=>"110011100",
  45117=>"001010111",
  45118=>"101110110",
  45119=>"100100001",
  45120=>"000100000",
  45121=>"111010011",
  45122=>"001000100",
  45123=>"001011111",
  45124=>"000011111",
  45125=>"011110010",
  45126=>"101110011",
  45127=>"000010010",
  45128=>"101000000",
  45129=>"010101000",
  45130=>"110110000",
  45131=>"111100110",
  45132=>"010110101",
  45133=>"010011101",
  45134=>"001010001",
  45135=>"101000000",
  45136=>"110000111",
  45137=>"000000010",
  45138=>"111000001",
  45139=>"001001101",
  45140=>"010001001",
  45141=>"000100111",
  45142=>"110001111",
  45143=>"110011111",
  45144=>"000111001",
  45145=>"100101011",
  45146=>"111100000",
  45147=>"000110110",
  45148=>"000111011",
  45149=>"101100011",
  45150=>"001100101",
  45151=>"000100110",
  45152=>"000100111",
  45153=>"001011000",
  45154=>"000010101",
  45155=>"000101000",
  45156=>"101101011",
  45157=>"001000111",
  45158=>"000011111",
  45159=>"001111111",
  45160=>"011110111",
  45161=>"100110011",
  45162=>"100000000",
  45163=>"010101001",
  45164=>"111110000",
  45165=>"010110010",
  45166=>"001100000",
  45167=>"110000100",
  45168=>"100000000",
  45169=>"010111011",
  45170=>"110011110",
  45171=>"110100000",
  45172=>"010000100",
  45173=>"001001000",
  45174=>"111001000",
  45175=>"111000111",
  45176=>"101110010",
  45177=>"101100100",
  45178=>"011000101",
  45179=>"110111000",
  45180=>"110100101",
  45181=>"000000000",
  45182=>"001001110",
  45183=>"000110101",
  45184=>"000000001",
  45185=>"111100111",
  45186=>"001001100",
  45187=>"010110000",
  45188=>"000000100",
  45189=>"010100100",
  45190=>"000100100",
  45191=>"001010111",
  45192=>"111011111",
  45193=>"101000001",
  45194=>"100001000",
  45195=>"111001111",
  45196=>"000100111",
  45197=>"001011000",
  45198=>"111001100",
  45199=>"000110110",
  45200=>"010010101",
  45201=>"000111010",
  45202=>"010001010",
  45203=>"010101111",
  45204=>"101010001",
  45205=>"100010010",
  45206=>"000100111",
  45207=>"000100010",
  45208=>"001100001",
  45209=>"011111001",
  45210=>"101100001",
  45211=>"111001111",
  45212=>"111001110",
  45213=>"010111000",
  45214=>"111001001",
  45215=>"110111010",
  45216=>"111111000",
  45217=>"011000100",
  45218=>"100000110",
  45219=>"100110111",
  45220=>"101100010",
  45221=>"111011100",
  45222=>"011001111",
  45223=>"100110000",
  45224=>"010011111",
  45225=>"001111000",
  45226=>"010011100",
  45227=>"000110011",
  45228=>"000001110",
  45229=>"100110111",
  45230=>"010110101",
  45231=>"101000100",
  45232=>"101000011",
  45233=>"011000010",
  45234=>"111110110",
  45235=>"101100000",
  45236=>"110110111",
  45237=>"000001111",
  45238=>"110110101",
  45239=>"010110111",
  45240=>"100001000",
  45241=>"010000101",
  45242=>"001001010",
  45243=>"001001000",
  45244=>"101001000",
  45245=>"110000001",
  45246=>"011101101",
  45247=>"110111110",
  45248=>"011000110",
  45249=>"010111000",
  45250=>"110101000",
  45251=>"111111111",
  45252=>"001110100",
  45253=>"111100001",
  45254=>"001010010",
  45255=>"101110001",
  45256=>"000001101",
  45257=>"000000010",
  45258=>"010100000",
  45259=>"111111101",
  45260=>"100110111",
  45261=>"010000010",
  45262=>"100111000",
  45263=>"001000001",
  45264=>"110000101",
  45265=>"111011111",
  45266=>"100011011",
  45267=>"000011010",
  45268=>"110100101",
  45269=>"000010001",
  45270=>"111101100",
  45271=>"110111001",
  45272=>"010000100",
  45273=>"001100011",
  45274=>"100001101",
  45275=>"000001110",
  45276=>"010101011",
  45277=>"000100111",
  45278=>"100111101",
  45279=>"101101011",
  45280=>"100111000",
  45281=>"001101011",
  45282=>"111001000",
  45283=>"100111000",
  45284=>"110011100",
  45285=>"111010111",
  45286=>"010000100",
  45287=>"001000000",
  45288=>"010011000",
  45289=>"000000111",
  45290=>"101001001",
  45291=>"010000111",
  45292=>"111100011",
  45293=>"100001110",
  45294=>"011000111",
  45295=>"111000001",
  45296=>"111001100",
  45297=>"010001110",
  45298=>"000000110",
  45299=>"101100000",
  45300=>"010000011",
  45301=>"011110011",
  45302=>"011111001",
  45303=>"001101111",
  45304=>"000011100",
  45305=>"010100101",
  45306=>"110001111",
  45307=>"010010010",
  45308=>"000100000",
  45309=>"000010010",
  45310=>"000010000",
  45311=>"101111010",
  45312=>"111001100",
  45313=>"100001110",
  45314=>"000011001",
  45315=>"111011100",
  45316=>"000111000",
  45317=>"100100001",
  45318=>"100000101",
  45319=>"001111001",
  45320=>"000010010",
  45321=>"010011000",
  45322=>"000000001",
  45323=>"001000000",
  45324=>"001001011",
  45325=>"101100010",
  45326=>"010001001",
  45327=>"100100100",
  45328=>"001011010",
  45329=>"000110010",
  45330=>"110111000",
  45331=>"110101110",
  45332=>"110110000",
  45333=>"001101110",
  45334=>"100110011",
  45335=>"100110011",
  45336=>"010111101",
  45337=>"001111111",
  45338=>"010000101",
  45339=>"001010110",
  45340=>"001000110",
  45341=>"111000001",
  45342=>"011000111",
  45343=>"000110011",
  45344=>"011111101",
  45345=>"101110110",
  45346=>"111110111",
  45347=>"010100111",
  45348=>"100001000",
  45349=>"110010100",
  45350=>"000100001",
  45351=>"011010001",
  45352=>"111000100",
  45353=>"100101000",
  45354=>"000110111",
  45355=>"010111001",
  45356=>"110010110",
  45357=>"001101100",
  45358=>"000101111",
  45359=>"100011011",
  45360=>"100010101",
  45361=>"101101100",
  45362=>"101111101",
  45363=>"111111110",
  45364=>"001110010",
  45365=>"011111111",
  45366=>"001001001",
  45367=>"000100110",
  45368=>"100001010",
  45369=>"001000100",
  45370=>"001011111",
  45371=>"101001010",
  45372=>"001111111",
  45373=>"101011101",
  45374=>"010010010",
  45375=>"100001100",
  45376=>"101101101",
  45377=>"101010001",
  45378=>"000101011",
  45379=>"101101011",
  45380=>"001000111",
  45381=>"111011001",
  45382=>"110001001",
  45383=>"100011010",
  45384=>"011101100",
  45385=>"001000000",
  45386=>"011000010",
  45387=>"011000001",
  45388=>"110000100",
  45389=>"111000001",
  45390=>"000010000",
  45391=>"000010010",
  45392=>"110001110",
  45393=>"010101011",
  45394=>"011001111",
  45395=>"111101110",
  45396=>"111011111",
  45397=>"110001110",
  45398=>"100100100",
  45399=>"010101101",
  45400=>"100101101",
  45401=>"100100001",
  45402=>"110010001",
  45403=>"001010100",
  45404=>"001111110",
  45405=>"000001100",
  45406=>"100001010",
  45407=>"011011011",
  45408=>"011110000",
  45409=>"010111010",
  45410=>"110000110",
  45411=>"011010000",
  45412=>"000010111",
  45413=>"111000001",
  45414=>"000100010",
  45415=>"011000110",
  45416=>"101001001",
  45417=>"101101111",
  45418=>"011110000",
  45419=>"111110000",
  45420=>"101110000",
  45421=>"111111011",
  45422=>"101010000",
  45423=>"111111100",
  45424=>"000000011",
  45425=>"101001001",
  45426=>"100011000",
  45427=>"000001001",
  45428=>"001000100",
  45429=>"100100110",
  45430=>"100101011",
  45431=>"010101001",
  45432=>"101111100",
  45433=>"011001101",
  45434=>"010010010",
  45435=>"000110001",
  45436=>"000111000",
  45437=>"011010101",
  45438=>"011111111",
  45439=>"110100000",
  45440=>"010010101",
  45441=>"111111010",
  45442=>"010111110",
  45443=>"011011101",
  45444=>"101110010",
  45445=>"000001100",
  45446=>"111110100",
  45447=>"010111101",
  45448=>"000111001",
  45449=>"011011001",
  45450=>"011101000",
  45451=>"111010111",
  45452=>"100101010",
  45453=>"011111101",
  45454=>"101010110",
  45455=>"100010110",
  45456=>"110011101",
  45457=>"000001001",
  45458=>"111010101",
  45459=>"101010010",
  45460=>"001110000",
  45461=>"010010100",
  45462=>"110100010",
  45463=>"011100010",
  45464=>"111000000",
  45465=>"111111010",
  45466=>"111101001",
  45467=>"000100100",
  45468=>"000100100",
  45469=>"001011001",
  45470=>"111000110",
  45471=>"010000101",
  45472=>"001011001",
  45473=>"111000111",
  45474=>"110010100",
  45475=>"001100111",
  45476=>"011001100",
  45477=>"110010010",
  45478=>"110001001",
  45479=>"010000100",
  45480=>"010110011",
  45481=>"011111001",
  45482=>"101000111",
  45483=>"111001100",
  45484=>"111010011",
  45485=>"010100110",
  45486=>"011110101",
  45487=>"010110001",
  45488=>"000111000",
  45489=>"110110111",
  45490=>"000100000",
  45491=>"011001000",
  45492=>"000100101",
  45493=>"110101101",
  45494=>"010111110",
  45495=>"001100001",
  45496=>"011011101",
  45497=>"010011011",
  45498=>"111100001",
  45499=>"100001101",
  45500=>"110010111",
  45501=>"000001010",
  45502=>"110110100",
  45503=>"001000100",
  45504=>"101001001",
  45505=>"011000100",
  45506=>"101010001",
  45507=>"011111000",
  45508=>"111101010",
  45509=>"001001011",
  45510=>"111000000",
  45511=>"000101001",
  45512=>"111111010",
  45513=>"111110011",
  45514=>"001100111",
  45515=>"100111001",
  45516=>"110011110",
  45517=>"000110110",
  45518=>"000011011",
  45519=>"101000111",
  45520=>"011111110",
  45521=>"000011111",
  45522=>"111011100",
  45523=>"011000100",
  45524=>"011100111",
  45525=>"010000111",
  45526=>"001110011",
  45527=>"001101010",
  45528=>"001010001",
  45529=>"111000001",
  45530=>"011000000",
  45531=>"111001111",
  45532=>"001011100",
  45533=>"111111100",
  45534=>"001100000",
  45535=>"100110111",
  45536=>"010010110",
  45537=>"100100111",
  45538=>"110011000",
  45539=>"110101100",
  45540=>"001011110",
  45541=>"100000111",
  45542=>"100010000",
  45543=>"011100110",
  45544=>"101110000",
  45545=>"110111111",
  45546=>"100000101",
  45547=>"010100100",
  45548=>"100010000",
  45549=>"100110000",
  45550=>"001001000",
  45551=>"000101001",
  45552=>"110100100",
  45553=>"011100000",
  45554=>"100101010",
  45555=>"001010111",
  45556=>"110011111",
  45557=>"000110100",
  45558=>"010111010",
  45559=>"100101101",
  45560=>"000000011",
  45561=>"110011100",
  45562=>"000110101",
  45563=>"010011011",
  45564=>"101111010",
  45565=>"110011010",
  45566=>"001010010",
  45567=>"101111000",
  45568=>"001000000",
  45569=>"011100010",
  45570=>"010000001",
  45571=>"001100011",
  45572=>"100101010",
  45573=>"000010101",
  45574=>"100101001",
  45575=>"100010100",
  45576=>"110000011",
  45577=>"001100010",
  45578=>"001100111",
  45579=>"010101001",
  45580=>"100111101",
  45581=>"011111110",
  45582=>"000010111",
  45583=>"100101010",
  45584=>"011011101",
  45585=>"110111100",
  45586=>"000001000",
  45587=>"110000101",
  45588=>"111101000",
  45589=>"110001111",
  45590=>"010110110",
  45591=>"110100101",
  45592=>"100010000",
  45593=>"011111001",
  45594=>"000000011",
  45595=>"111111101",
  45596=>"101011010",
  45597=>"110011101",
  45598=>"001110100",
  45599=>"010011010",
  45600=>"100011111",
  45601=>"001000101",
  45602=>"000000100",
  45603=>"101100000",
  45604=>"111011010",
  45605=>"010001011",
  45606=>"111100100",
  45607=>"000110001",
  45608=>"101001110",
  45609=>"001010100",
  45610=>"000101010",
  45611=>"101000001",
  45612=>"010010110",
  45613=>"010001111",
  45614=>"101101010",
  45615=>"110011001",
  45616=>"011111000",
  45617=>"000110111",
  45618=>"000110100",
  45619=>"101010111",
  45620=>"111111110",
  45621=>"011100010",
  45622=>"110111001",
  45623=>"100110011",
  45624=>"101000000",
  45625=>"010000101",
  45626=>"000111110",
  45627=>"101111100",
  45628=>"100011000",
  45629=>"000010000",
  45630=>"100010010",
  45631=>"100111000",
  45632=>"001010001",
  45633=>"110000001",
  45634=>"000011100",
  45635=>"010111001",
  45636=>"111000000",
  45637=>"011010110",
  45638=>"001110011",
  45639=>"001010101",
  45640=>"001111100",
  45641=>"011100001",
  45642=>"001111011",
  45643=>"011100111",
  45644=>"001011010",
  45645=>"101000010",
  45646=>"110101001",
  45647=>"101001011",
  45648=>"001011011",
  45649=>"110110101",
  45650=>"010100011",
  45651=>"010000100",
  45652=>"011001110",
  45653=>"010100000",
  45654=>"000001011",
  45655=>"000110101",
  45656=>"110011111",
  45657=>"101100000",
  45658=>"100100001",
  45659=>"011111100",
  45660=>"110100001",
  45661=>"001101001",
  45662=>"011001011",
  45663=>"011011100",
  45664=>"001000101",
  45665=>"001010100",
  45666=>"111011000",
  45667=>"101000100",
  45668=>"111100000",
  45669=>"000100001",
  45670=>"110010111",
  45671=>"110010001",
  45672=>"011001101",
  45673=>"000100011",
  45674=>"010010001",
  45675=>"001000000",
  45676=>"011010001",
  45677=>"111000100",
  45678=>"110010111",
  45679=>"110111010",
  45680=>"100110000",
  45681=>"111100110",
  45682=>"101001010",
  45683=>"000011110",
  45684=>"001110111",
  45685=>"000000111",
  45686=>"001001101",
  45687=>"001101111",
  45688=>"100011001",
  45689=>"011111100",
  45690=>"100111001",
  45691=>"111010011",
  45692=>"000101101",
  45693=>"110110010",
  45694=>"001110100",
  45695=>"011010010",
  45696=>"100010010",
  45697=>"101101001",
  45698=>"111000000",
  45699=>"001010100",
  45700=>"111100010",
  45701=>"100000000",
  45702=>"100110110",
  45703=>"111010000",
  45704=>"000011100",
  45705=>"000110011",
  45706=>"111100000",
  45707=>"010010110",
  45708=>"000000110",
  45709=>"001100100",
  45710=>"100101010",
  45711=>"000010100",
  45712=>"000000011",
  45713=>"011110111",
  45714=>"110111101",
  45715=>"001101110",
  45716=>"000111110",
  45717=>"111000101",
  45718=>"000100111",
  45719=>"010110100",
  45720=>"111100011",
  45721=>"101111000",
  45722=>"010101111",
  45723=>"010101010",
  45724=>"000011110",
  45725=>"110001010",
  45726=>"011110011",
  45727=>"000111110",
  45728=>"011111111",
  45729=>"111011111",
  45730=>"011101010",
  45731=>"110001110",
  45732=>"110110011",
  45733=>"111111011",
  45734=>"111010010",
  45735=>"010110000",
  45736=>"111100111",
  45737=>"000000110",
  45738=>"011111010",
  45739=>"000001001",
  45740=>"110000100",
  45741=>"001000000",
  45742=>"001110011",
  45743=>"100010000",
  45744=>"101001101",
  45745=>"001010011",
  45746=>"010100011",
  45747=>"000100100",
  45748=>"001001011",
  45749=>"010100101",
  45750=>"010001001",
  45751=>"011100000",
  45752=>"100111101",
  45753=>"101001100",
  45754=>"000010100",
  45755=>"000100111",
  45756=>"100100111",
  45757=>"001011001",
  45758=>"111010010",
  45759=>"100110101",
  45760=>"110010111",
  45761=>"001001000",
  45762=>"000100000",
  45763=>"011010010",
  45764=>"111111111",
  45765=>"011111111",
  45766=>"101011011",
  45767=>"001000110",
  45768=>"000010010",
  45769=>"111000010",
  45770=>"010110001",
  45771=>"010001010",
  45772=>"100010101",
  45773=>"000010001",
  45774=>"111001110",
  45775=>"110000110",
  45776=>"100101000",
  45777=>"010000010",
  45778=>"110111000",
  45779=>"011000100",
  45780=>"101111000",
  45781=>"001000110",
  45782=>"101001110",
  45783=>"011100110",
  45784=>"010101011",
  45785=>"001001000",
  45786=>"100001100",
  45787=>"111011101",
  45788=>"010111011",
  45789=>"000011010",
  45790=>"011011111",
  45791=>"110110111",
  45792=>"101001101",
  45793=>"011100100",
  45794=>"100111111",
  45795=>"110101111",
  45796=>"011001011",
  45797=>"111111101",
  45798=>"000101010",
  45799=>"101110001",
  45800=>"100000001",
  45801=>"001111011",
  45802=>"011000000",
  45803=>"000000000",
  45804=>"000011010",
  45805=>"001000111",
  45806=>"111000100",
  45807=>"111010111",
  45808=>"001001101",
  45809=>"011010011",
  45810=>"101101000",
  45811=>"110010101",
  45812=>"111000010",
  45813=>"111100101",
  45814=>"100010101",
  45815=>"110110010",
  45816=>"110001100",
  45817=>"111111111",
  45818=>"000101001",
  45819=>"001000001",
  45820=>"001011110",
  45821=>"000110001",
  45822=>"110001001",
  45823=>"110110011",
  45824=>"111001010",
  45825=>"100010110",
  45826=>"011000010",
  45827=>"100100000",
  45828=>"111000001",
  45829=>"010010011",
  45830=>"101011101",
  45831=>"100101101",
  45832=>"001010110",
  45833=>"100111000",
  45834=>"111111111",
  45835=>"010011110",
  45836=>"000010100",
  45837=>"011000110",
  45838=>"111100101",
  45839=>"011101111",
  45840=>"001100000",
  45841=>"100111001",
  45842=>"111001011",
  45843=>"110000100",
  45844=>"101011001",
  45845=>"111101011",
  45846=>"011011011",
  45847=>"111010111",
  45848=>"110111000",
  45849=>"000000101",
  45850=>"110011010",
  45851=>"001001111",
  45852=>"000000111",
  45853=>"111000101",
  45854=>"000110101",
  45855=>"111101011",
  45856=>"101101111",
  45857=>"011001101",
  45858=>"011010110",
  45859=>"101001011",
  45860=>"101010000",
  45861=>"110100110",
  45862=>"101010000",
  45863=>"100100100",
  45864=>"111011001",
  45865=>"101001001",
  45866=>"011010000",
  45867=>"111110011",
  45868=>"101110011",
  45869=>"011100100",
  45870=>"011011010",
  45871=>"001000011",
  45872=>"001001101",
  45873=>"000000110",
  45874=>"000101000",
  45875=>"100110011",
  45876=>"010011001",
  45877=>"101010100",
  45878=>"001011000",
  45879=>"110111101",
  45880=>"101111000",
  45881=>"000101111",
  45882=>"001101011",
  45883=>"010101010",
  45884=>"101000100",
  45885=>"111110001",
  45886=>"000000001",
  45887=>"000101101",
  45888=>"100000000",
  45889=>"011100000",
  45890=>"101001111",
  45891=>"000000001",
  45892=>"100111111",
  45893=>"110100011",
  45894=>"100111111",
  45895=>"111000001",
  45896=>"000110001",
  45897=>"010000011",
  45898=>"111110011",
  45899=>"011001011",
  45900=>"110000001",
  45901=>"110110101",
  45902=>"100010010",
  45903=>"100100100",
  45904=>"110000110",
  45905=>"100101100",
  45906=>"010011101",
  45907=>"000111111",
  45908=>"100001111",
  45909=>"111111001",
  45910=>"111100011",
  45911=>"010110011",
  45912=>"010011110",
  45913=>"000111100",
  45914=>"010011011",
  45915=>"111000100",
  45916=>"010100011",
  45917=>"100011000",
  45918=>"001011110",
  45919=>"100000010",
  45920=>"011000010",
  45921=>"000001011",
  45922=>"111000111",
  45923=>"100111111",
  45924=>"110011110",
  45925=>"110111010",
  45926=>"001100111",
  45927=>"010000011",
  45928=>"011000101",
  45929=>"101100000",
  45930=>"001010111",
  45931=>"100101011",
  45932=>"001110000",
  45933=>"100011100",
  45934=>"001110001",
  45935=>"010000101",
  45936=>"110011101",
  45937=>"011010010",
  45938=>"010100000",
  45939=>"101001100",
  45940=>"100100110",
  45941=>"011001001",
  45942=>"101110000",
  45943=>"010000001",
  45944=>"010110110",
  45945=>"101001111",
  45946=>"011011110",
  45947=>"110100111",
  45948=>"000010100",
  45949=>"110011001",
  45950=>"110111000",
  45951=>"000001111",
  45952=>"011010010",
  45953=>"000111110",
  45954=>"101100000",
  45955=>"110010111",
  45956=>"001001111",
  45957=>"010100101",
  45958=>"100101100",
  45959=>"100000011",
  45960=>"000001100",
  45961=>"010111001",
  45962=>"000000011",
  45963=>"111101010",
  45964=>"110000100",
  45965=>"001011010",
  45966=>"000001000",
  45967=>"000001100",
  45968=>"110101010",
  45969=>"010001010",
  45970=>"000000111",
  45971=>"000000111",
  45972=>"100100110",
  45973=>"001001010",
  45974=>"000111001",
  45975=>"011001110",
  45976=>"101001110",
  45977=>"110001101",
  45978=>"000010110",
  45979=>"110110111",
  45980=>"110110001",
  45981=>"110110110",
  45982=>"111001000",
  45983=>"111001000",
  45984=>"110110001",
  45985=>"011000001",
  45986=>"010101110",
  45987=>"011000100",
  45988=>"110111100",
  45989=>"101111111",
  45990=>"001101110",
  45991=>"010010010",
  45992=>"000101111",
  45993=>"000010010",
  45994=>"010001111",
  45995=>"100111011",
  45996=>"000001000",
  45997=>"100000111",
  45998=>"011101000",
  45999=>"001110000",
  46000=>"011100011",
  46001=>"010101001",
  46002=>"000100001",
  46003=>"100001000",
  46004=>"111011000",
  46005=>"110111110",
  46006=>"001011000",
  46007=>"000110100",
  46008=>"101000100",
  46009=>"001111011",
  46010=>"101100010",
  46011=>"100011110",
  46012=>"100111001",
  46013=>"000101111",
  46014=>"001111000",
  46015=>"100001000",
  46016=>"110101001",
  46017=>"011001100",
  46018=>"100001001",
  46019=>"000001111",
  46020=>"101001110",
  46021=>"100111010",
  46022=>"101101110",
  46023=>"110100001",
  46024=>"000010011",
  46025=>"001110010",
  46026=>"101100111",
  46027=>"001100100",
  46028=>"000010100",
  46029=>"001000001",
  46030=>"000000100",
  46031=>"001001010",
  46032=>"110111111",
  46033=>"110100001",
  46034=>"010000011",
  46035=>"000101000",
  46036=>"110100011",
  46037=>"010000010",
  46038=>"001011100",
  46039=>"111100111",
  46040=>"111111100",
  46041=>"001011011",
  46042=>"101000010",
  46043=>"010111101",
  46044=>"001000111",
  46045=>"000011101",
  46046=>"001001000",
  46047=>"000000001",
  46048=>"001111011",
  46049=>"011011010",
  46050=>"101111001",
  46051=>"000000101",
  46052=>"000010010",
  46053=>"010101101",
  46054=>"111001000",
  46055=>"110101000",
  46056=>"100001000",
  46057=>"010100000",
  46058=>"010100001",
  46059=>"110100110",
  46060=>"100110000",
  46061=>"100010111",
  46062=>"000011100",
  46063=>"000101100",
  46064=>"101001100",
  46065=>"000011010",
  46066=>"011000011",
  46067=>"101100110",
  46068=>"101111010",
  46069=>"000101010",
  46070=>"111011111",
  46071=>"101010111",
  46072=>"011100100",
  46073=>"111101000",
  46074=>"100110000",
  46075=>"110101001",
  46076=>"101100101",
  46077=>"011001101",
  46078=>"111011010",
  46079=>"110100001",
  46080=>"111110111",
  46081=>"100110111",
  46082=>"011011100",
  46083=>"000111011",
  46084=>"110100011",
  46085=>"101010100",
  46086=>"101100101",
  46087=>"111110010",
  46088=>"000000100",
  46089=>"100100011",
  46090=>"111110010",
  46091=>"110100001",
  46092=>"101110000",
  46093=>"110110001",
  46094=>"100010010",
  46095=>"011111001",
  46096=>"111011100",
  46097=>"111101111",
  46098=>"100111000",
  46099=>"110111100",
  46100=>"111010101",
  46101=>"000110111",
  46102=>"011011110",
  46103=>"110000000",
  46104=>"111100110",
  46105=>"100101111",
  46106=>"110100000",
  46107=>"001101011",
  46108=>"101101100",
  46109=>"011110000",
  46110=>"001111001",
  46111=>"010000100",
  46112=>"100000101",
  46113=>"110011100",
  46114=>"111001000",
  46115=>"111001111",
  46116=>"010011010",
  46117=>"101010010",
  46118=>"101011110",
  46119=>"001010011",
  46120=>"001001001",
  46121=>"000100000",
  46122=>"010011010",
  46123=>"100000110",
  46124=>"101110000",
  46125=>"110000011",
  46126=>"001110011",
  46127=>"100000111",
  46128=>"011010101",
  46129=>"110101111",
  46130=>"011100001",
  46131=>"100000000",
  46132=>"001101101",
  46133=>"111100100",
  46134=>"001101011",
  46135=>"010111110",
  46136=>"100100001",
  46137=>"001100111",
  46138=>"001111011",
  46139=>"111011100",
  46140=>"011001001",
  46141=>"001100100",
  46142=>"111101011",
  46143=>"001001101",
  46144=>"101010011",
  46145=>"011001011",
  46146=>"000101111",
  46147=>"010100000",
  46148=>"110001010",
  46149=>"000000111",
  46150=>"110111001",
  46151=>"010010101",
  46152=>"000000001",
  46153=>"110000001",
  46154=>"110111001",
  46155=>"010011001",
  46156=>"111011010",
  46157=>"000100011",
  46158=>"011101000",
  46159=>"011100101",
  46160=>"111110010",
  46161=>"010000010",
  46162=>"101100001",
  46163=>"110100101",
  46164=>"111111001",
  46165=>"010000001",
  46166=>"110111110",
  46167=>"100101001",
  46168=>"110011100",
  46169=>"010011010",
  46170=>"011001110",
  46171=>"101001001",
  46172=>"000011111",
  46173=>"001000001",
  46174=>"001111101",
  46175=>"100000010",
  46176=>"111101110",
  46177=>"011100001",
  46178=>"000110010",
  46179=>"100101000",
  46180=>"110100110",
  46181=>"101001100",
  46182=>"100001011",
  46183=>"011011110",
  46184=>"101010101",
  46185=>"011110110",
  46186=>"000101101",
  46187=>"110100100",
  46188=>"110101010",
  46189=>"010011010",
  46190=>"010110000",
  46191=>"101000111",
  46192=>"011010010",
  46193=>"100001110",
  46194=>"101010100",
  46195=>"000000100",
  46196=>"001011101",
  46197=>"011111111",
  46198=>"100111001",
  46199=>"111101111",
  46200=>"001011100",
  46201=>"101000110",
  46202=>"110100000",
  46203=>"001011000",
  46204=>"111110100",
  46205=>"100000001",
  46206=>"111001111",
  46207=>"101001100",
  46208=>"111011010",
  46209=>"101001000",
  46210=>"001110000",
  46211=>"100010001",
  46212=>"001100010",
  46213=>"001001111",
  46214=>"101001111",
  46215=>"110100100",
  46216=>"010111101",
  46217=>"011011011",
  46218=>"110111101",
  46219=>"000111011",
  46220=>"100010111",
  46221=>"111010011",
  46222=>"010001011",
  46223=>"100011100",
  46224=>"001001101",
  46225=>"001000100",
  46226=>"100101100",
  46227=>"011010001",
  46228=>"010001011",
  46229=>"110001111",
  46230=>"011111001",
  46231=>"011001100",
  46232=>"111000001",
  46233=>"000000010",
  46234=>"101100111",
  46235=>"100111110",
  46236=>"100110011",
  46237=>"011110000",
  46238=>"111000111",
  46239=>"111001010",
  46240=>"101111000",
  46241=>"100101100",
  46242=>"011000111",
  46243=>"111101110",
  46244=>"000011011",
  46245=>"000111110",
  46246=>"100011000",
  46247=>"000101000",
  46248=>"111101111",
  46249=>"100101010",
  46250=>"101000000",
  46251=>"001100101",
  46252=>"100010111",
  46253=>"010111101",
  46254=>"001110110",
  46255=>"001111001",
  46256=>"111011001",
  46257=>"011000000",
  46258=>"001101011",
  46259=>"001010100",
  46260=>"011101001",
  46261=>"110010111",
  46262=>"010101111",
  46263=>"011010110",
  46264=>"011010110",
  46265=>"100010011",
  46266=>"001100010",
  46267=>"101011100",
  46268=>"111110111",
  46269=>"000011110",
  46270=>"100111010",
  46271=>"111001100",
  46272=>"011100001",
  46273=>"001001101",
  46274=>"111111110",
  46275=>"111111001",
  46276=>"110011001",
  46277=>"010001000",
  46278=>"110111100",
  46279=>"011001101",
  46280=>"001010011",
  46281=>"001100100",
  46282=>"011100011",
  46283=>"100011010",
  46284=>"000101111",
  46285=>"100010100",
  46286=>"000100011",
  46287=>"101110100",
  46288=>"011110110",
  46289=>"111011010",
  46290=>"010000010",
  46291=>"001011001",
  46292=>"110111000",
  46293=>"010001000",
  46294=>"000111100",
  46295=>"111011010",
  46296=>"001000011",
  46297=>"010011011",
  46298=>"000010011",
  46299=>"101111111",
  46300=>"000101111",
  46301=>"000001011",
  46302=>"101111111",
  46303=>"000110001",
  46304=>"011111100",
  46305=>"000000110",
  46306=>"111000011",
  46307=>"001001000",
  46308=>"011100101",
  46309=>"111101101",
  46310=>"101101111",
  46311=>"100001110",
  46312=>"110001000",
  46313=>"110001100",
  46314=>"100110101",
  46315=>"101100010",
  46316=>"010001101",
  46317=>"111000011",
  46318=>"110110011",
  46319=>"000001110",
  46320=>"111000000",
  46321=>"010010000",
  46322=>"001101110",
  46323=>"111100111",
  46324=>"101111000",
  46325=>"101111000",
  46326=>"000001111",
  46327=>"100011011",
  46328=>"101011100",
  46329=>"111010010",
  46330=>"010011010",
  46331=>"000101111",
  46332=>"101000000",
  46333=>"010001100",
  46334=>"000010111",
  46335=>"000111010",
  46336=>"011000011",
  46337=>"010001110",
  46338=>"001010111",
  46339=>"001101010",
  46340=>"101001110",
  46341=>"111010000",
  46342=>"011000001",
  46343=>"100101111",
  46344=>"100011001",
  46345=>"000101010",
  46346=>"010111010",
  46347=>"110001100",
  46348=>"111111100",
  46349=>"110001111",
  46350=>"100111000",
  46351=>"100001011",
  46352=>"110000010",
  46353=>"000100110",
  46354=>"000000011",
  46355=>"110110011",
  46356=>"001100101",
  46357=>"111101110",
  46358=>"111111010",
  46359=>"000000111",
  46360=>"011101001",
  46361=>"111101100",
  46362=>"000101111",
  46363=>"001010101",
  46364=>"101101000",
  46365=>"010111011",
  46366=>"110111111",
  46367=>"011100110",
  46368=>"011111111",
  46369=>"010101011",
  46370=>"111100101",
  46371=>"001010110",
  46372=>"111110011",
  46373=>"011010111",
  46374=>"110010101",
  46375=>"111001101",
  46376=>"010000001",
  46377=>"001010111",
  46378=>"001001010",
  46379=>"101010010",
  46380=>"010001110",
  46381=>"001010101",
  46382=>"101000101",
  46383=>"110010101",
  46384=>"000001000",
  46385=>"111001101",
  46386=>"110011110",
  46387=>"001111110",
  46388=>"101111111",
  46389=>"000010111",
  46390=>"111100011",
  46391=>"001101000",
  46392=>"011100011",
  46393=>"001101111",
  46394=>"110101011",
  46395=>"100011110",
  46396=>"001010100",
  46397=>"011011001",
  46398=>"010011010",
  46399=>"111000001",
  46400=>"010000111",
  46401=>"110001000",
  46402=>"100101001",
  46403=>"001111010",
  46404=>"011001111",
  46405=>"111001001",
  46406=>"000001000",
  46407=>"101011111",
  46408=>"010100101",
  46409=>"110010110",
  46410=>"011110101",
  46411=>"010001001",
  46412=>"110001000",
  46413=>"110000010",
  46414=>"010110010",
  46415=>"000010101",
  46416=>"001101010",
  46417=>"011100100",
  46418=>"110010000",
  46419=>"110111000",
  46420=>"011001010",
  46421=>"000101101",
  46422=>"010001101",
  46423=>"000110110",
  46424=>"100111001",
  46425=>"000100001",
  46426=>"111100100",
  46427=>"010000101",
  46428=>"000001100",
  46429=>"101110111",
  46430=>"101011001",
  46431=>"111011110",
  46432=>"000100000",
  46433=>"111010101",
  46434=>"110001110",
  46435=>"111001111",
  46436=>"100010111",
  46437=>"010000001",
  46438=>"111000100",
  46439=>"011011001",
  46440=>"111000000",
  46441=>"100110101",
  46442=>"111001001",
  46443=>"111101011",
  46444=>"111111011",
  46445=>"101101011",
  46446=>"011010100",
  46447=>"000011011",
  46448=>"100110001",
  46449=>"011100100",
  46450=>"011100100",
  46451=>"111010100",
  46452=>"010110000",
  46453=>"001111001",
  46454=>"010011010",
  46455=>"001001100",
  46456=>"111011000",
  46457=>"100110111",
  46458=>"101101011",
  46459=>"000101111",
  46460=>"101100011",
  46461=>"111000111",
  46462=>"011001000",
  46463=>"001011011",
  46464=>"000000100",
  46465=>"110000110",
  46466=>"111111000",
  46467=>"010100000",
  46468=>"100011100",
  46469=>"001010110",
  46470=>"001101101",
  46471=>"010001000",
  46472=>"101001101",
  46473=>"111111010",
  46474=>"100100011",
  46475=>"110000100",
  46476=>"011000110",
  46477=>"001100011",
  46478=>"100011101",
  46479=>"110001010",
  46480=>"110100111",
  46481=>"111000010",
  46482=>"111000011",
  46483=>"011000110",
  46484=>"001101111",
  46485=>"000110010",
  46486=>"100000011",
  46487=>"011110001",
  46488=>"100110110",
  46489=>"111110101",
  46490=>"101110101",
  46491=>"111001000",
  46492=>"110101101",
  46493=>"001100000",
  46494=>"000010110",
  46495=>"101001011",
  46496=>"010110111",
  46497=>"011001100",
  46498=>"100010100",
  46499=>"111010111",
  46500=>"000110000",
  46501=>"110110010",
  46502=>"110001111",
  46503=>"100101001",
  46504=>"101111000",
  46505=>"110110001",
  46506=>"010110011",
  46507=>"010100011",
  46508=>"100011011",
  46509=>"111111001",
  46510=>"011010010",
  46511=>"100100100",
  46512=>"111101000",
  46513=>"000111001",
  46514=>"100100011",
  46515=>"011001010",
  46516=>"000101101",
  46517=>"111010111",
  46518=>"011100111",
  46519=>"011110010",
  46520=>"111001010",
  46521=>"101010000",
  46522=>"001010110",
  46523=>"111011101",
  46524=>"111100111",
  46525=>"010100000",
  46526=>"110101111",
  46527=>"001011111",
  46528=>"100110110",
  46529=>"001111010",
  46530=>"000111101",
  46531=>"111110101",
  46532=>"100010010",
  46533=>"110111000",
  46534=>"010010110",
  46535=>"100000100",
  46536=>"001100110",
  46537=>"001111010",
  46538=>"101111001",
  46539=>"101100010",
  46540=>"000110010",
  46541=>"111001101",
  46542=>"100010011",
  46543=>"010101011",
  46544=>"000111000",
  46545=>"110001000",
  46546=>"010100001",
  46547=>"100111101",
  46548=>"011100011",
  46549=>"010101100",
  46550=>"100101110",
  46551=>"100010111",
  46552=>"000000101",
  46553=>"111001100",
  46554=>"101111011",
  46555=>"000101001",
  46556=>"001111000",
  46557=>"010000101",
  46558=>"100011110",
  46559=>"010000010",
  46560=>"000101110",
  46561=>"110101110",
  46562=>"100111111",
  46563=>"001011010",
  46564=>"001000001",
  46565=>"010001010",
  46566=>"011011101",
  46567=>"011110100",
  46568=>"111110000",
  46569=>"100010101",
  46570=>"110011101",
  46571=>"001001100",
  46572=>"001110100",
  46573=>"100110010",
  46574=>"111111111",
  46575=>"001101011",
  46576=>"110010110",
  46577=>"010010010",
  46578=>"100100111",
  46579=>"000100001",
  46580=>"111110110",
  46581=>"000011010",
  46582=>"101010110",
  46583=>"010100110",
  46584=>"011100000",
  46585=>"010011000",
  46586=>"010101000",
  46587=>"010010000",
  46588=>"100000001",
  46589=>"100010010",
  46590=>"000011000",
  46591=>"011000101",
  46592=>"110101101",
  46593=>"110101001",
  46594=>"111000111",
  46595=>"001100111",
  46596=>"011110110",
  46597=>"110000110",
  46598=>"010111110",
  46599=>"011111110",
  46600=>"011101110",
  46601=>"110011011",
  46602=>"111101001",
  46603=>"111111010",
  46604=>"111111000",
  46605=>"010010101",
  46606=>"100110000",
  46607=>"001000011",
  46608=>"101011100",
  46609=>"001100110",
  46610=>"001001001",
  46611=>"011000110",
  46612=>"000101011",
  46613=>"111111011",
  46614=>"000001011",
  46615=>"010011101",
  46616=>"010001100",
  46617=>"000100101",
  46618=>"010100111",
  46619=>"110110001",
  46620=>"111011001",
  46621=>"110111011",
  46622=>"010001011",
  46623=>"011011010",
  46624=>"110000101",
  46625=>"000100010",
  46626=>"000110110",
  46627=>"000011111",
  46628=>"111110001",
  46629=>"111011111",
  46630=>"100001001",
  46631=>"101100111",
  46632=>"100011100",
  46633=>"111010110",
  46634=>"000101011",
  46635=>"000001011",
  46636=>"111001000",
  46637=>"110101101",
  46638=>"110001000",
  46639=>"010111011",
  46640=>"111001111",
  46641=>"100101111",
  46642=>"000101110",
  46643=>"100100100",
  46644=>"110110100",
  46645=>"110000010",
  46646=>"110010010",
  46647=>"111101111",
  46648=>"110000000",
  46649=>"011111111",
  46650=>"111000011",
  46651=>"100100100",
  46652=>"000001010",
  46653=>"101001100",
  46654=>"001100000",
  46655=>"101101010",
  46656=>"010110100",
  46657=>"101111000",
  46658=>"010000101",
  46659=>"110110111",
  46660=>"000110011",
  46661=>"101000011",
  46662=>"111100100",
  46663=>"101101110",
  46664=>"010110101",
  46665=>"111111000",
  46666=>"101101011",
  46667=>"000010000",
  46668=>"011010101",
  46669=>"010100010",
  46670=>"100110111",
  46671=>"010001001",
  46672=>"001010000",
  46673=>"111001110",
  46674=>"000001011",
  46675=>"000110111",
  46676=>"110111111",
  46677=>"101100010",
  46678=>"010000011",
  46679=>"100100111",
  46680=>"001001101",
  46681=>"100010110",
  46682=>"101110100",
  46683=>"011000100",
  46684=>"101010001",
  46685=>"001001011",
  46686=>"010100000",
  46687=>"100011110",
  46688=>"111100001",
  46689=>"001000011",
  46690=>"101101001",
  46691=>"100000110",
  46692=>"001111000",
  46693=>"010000100",
  46694=>"101000010",
  46695=>"111000000",
  46696=>"110101001",
  46697=>"100110111",
  46698=>"001110101",
  46699=>"110001000",
  46700=>"111101110",
  46701=>"010001110",
  46702=>"001110000",
  46703=>"011010000",
  46704=>"100110110",
  46705=>"010111010",
  46706=>"101001010",
  46707=>"111010101",
  46708=>"101111111",
  46709=>"001101111",
  46710=>"000010011",
  46711=>"001011001",
  46712=>"100010000",
  46713=>"110110100",
  46714=>"101110111",
  46715=>"010111100",
  46716=>"000110101",
  46717=>"011000111",
  46718=>"001011010",
  46719=>"011111011",
  46720=>"100001001",
  46721=>"001000001",
  46722=>"111000111",
  46723=>"110100100",
  46724=>"111011000",
  46725=>"010000010",
  46726=>"101001111",
  46727=>"100010100",
  46728=>"100111110",
  46729=>"001010000",
  46730=>"111101110",
  46731=>"111000001",
  46732=>"011011111",
  46733=>"101000011",
  46734=>"110001111",
  46735=>"000100101",
  46736=>"101111001",
  46737=>"111001100",
  46738=>"101000101",
  46739=>"110110010",
  46740=>"101010101",
  46741=>"011010000",
  46742=>"100000011",
  46743=>"011000101",
  46744=>"000111101",
  46745=>"101011111",
  46746=>"000011110",
  46747=>"001110111",
  46748=>"101000000",
  46749=>"100000101",
  46750=>"100101000",
  46751=>"100001111",
  46752=>"110100111",
  46753=>"111100100",
  46754=>"000001101",
  46755=>"010011100",
  46756=>"000100110",
  46757=>"111110010",
  46758=>"111111110",
  46759=>"101101000",
  46760=>"011111100",
  46761=>"011010101",
  46762=>"010001101",
  46763=>"101100111",
  46764=>"011010001",
  46765=>"111010101",
  46766=>"001110111",
  46767=>"000010100",
  46768=>"000111101",
  46769=>"010110110",
  46770=>"111000001",
  46771=>"110101101",
  46772=>"111010010",
  46773=>"101100000",
  46774=>"111101111",
  46775=>"011001010",
  46776=>"000001011",
  46777=>"100011101",
  46778=>"001001111",
  46779=>"011000000",
  46780=>"110110010",
  46781=>"011111101",
  46782=>"000100110",
  46783=>"111001000",
  46784=>"000101101",
  46785=>"111011111",
  46786=>"110001100",
  46787=>"110000011",
  46788=>"001111100",
  46789=>"110000000",
  46790=>"011101001",
  46791=>"011110010",
  46792=>"000000111",
  46793=>"100010001",
  46794=>"100000000",
  46795=>"111001100",
  46796=>"110110010",
  46797=>"010101100",
  46798=>"010000011",
  46799=>"100000011",
  46800=>"100100010",
  46801=>"000010010",
  46802=>"101000000",
  46803=>"110000100",
  46804=>"010011110",
  46805=>"110110111",
  46806=>"001000111",
  46807=>"010111100",
  46808=>"000010101",
  46809=>"010101100",
  46810=>"001111111",
  46811=>"010100101",
  46812=>"101001110",
  46813=>"000001000",
  46814=>"000010000",
  46815=>"101011011",
  46816=>"001010110",
  46817=>"101110001",
  46818=>"110100111",
  46819=>"001001010",
  46820=>"010100110",
  46821=>"100111100",
  46822=>"110101111",
  46823=>"001010000",
  46824=>"100000101",
  46825=>"100001001",
  46826=>"110011001",
  46827=>"010010110",
  46828=>"101000001",
  46829=>"111000100",
  46830=>"100010001",
  46831=>"100000111",
  46832=>"011101110",
  46833=>"000001100",
  46834=>"110000100",
  46835=>"100011000",
  46836=>"001100010",
  46837=>"000111000",
  46838=>"001101111",
  46839=>"101000100",
  46840=>"101100000",
  46841=>"000101111",
  46842=>"110010011",
  46843=>"001100110",
  46844=>"100101100",
  46845=>"010011011",
  46846=>"101101100",
  46847=>"110000111",
  46848=>"010001000",
  46849=>"010000101",
  46850=>"111100101",
  46851=>"011110111",
  46852=>"100111110",
  46853=>"111100011",
  46854=>"111001110",
  46855=>"010100110",
  46856=>"111010101",
  46857=>"000100110",
  46858=>"011010011",
  46859=>"101100100",
  46860=>"000101110",
  46861=>"001010100",
  46862=>"011100000",
  46863=>"101101000",
  46864=>"100100101",
  46865=>"001010101",
  46866=>"011010001",
  46867=>"011001000",
  46868=>"000001000",
  46869=>"001101100",
  46870=>"110011010",
  46871=>"000000011",
  46872=>"101001100",
  46873=>"001000100",
  46874=>"110010111",
  46875=>"001101100",
  46876=>"110101101",
  46877=>"101111110",
  46878=>"000010000",
  46879=>"101100000",
  46880=>"111011001",
  46881=>"100011000",
  46882=>"100010111",
  46883=>"101001110",
  46884=>"011111001",
  46885=>"011001001",
  46886=>"011110010",
  46887=>"110101001",
  46888=>"000011100",
  46889=>"111111000",
  46890=>"111010010",
  46891=>"001110111",
  46892=>"111101000",
  46893=>"000110111",
  46894=>"001101000",
  46895=>"000010100",
  46896=>"010001100",
  46897=>"110110100",
  46898=>"101011011",
  46899=>"110110100",
  46900=>"101011111",
  46901=>"110000001",
  46902=>"010110010",
  46903=>"011101111",
  46904=>"101111101",
  46905=>"000001101",
  46906=>"000111001",
  46907=>"110010110",
  46908=>"110111100",
  46909=>"010001110",
  46910=>"010010100",
  46911=>"011000100",
  46912=>"111101001",
  46913=>"011110100",
  46914=>"010000001",
  46915=>"101000111",
  46916=>"000110000",
  46917=>"110100110",
  46918=>"011010010",
  46919=>"000010011",
  46920=>"110011000",
  46921=>"100100010",
  46922=>"100111111",
  46923=>"001001001",
  46924=>"000000111",
  46925=>"111101010",
  46926=>"110101001",
  46927=>"110000001",
  46928=>"111111010",
  46929=>"110011110",
  46930=>"000000000",
  46931=>"001110010",
  46932=>"011011011",
  46933=>"010001100",
  46934=>"001100010",
  46935=>"110101100",
  46936=>"010001000",
  46937=>"001111001",
  46938=>"111001001",
  46939=>"010101111",
  46940=>"100111000",
  46941=>"000101000",
  46942=>"110010000",
  46943=>"011001000",
  46944=>"011000110",
  46945=>"101110100",
  46946=>"100010101",
  46947=>"100001100",
  46948=>"011110111",
  46949=>"110110000",
  46950=>"111011011",
  46951=>"000010010",
  46952=>"011011001",
  46953=>"110101111",
  46954=>"000001010",
  46955=>"010101110",
  46956=>"111101100",
  46957=>"111100100",
  46958=>"010011010",
  46959=>"010100101",
  46960=>"000000010",
  46961=>"001100110",
  46962=>"110101010",
  46963=>"000011000",
  46964=>"011101000",
  46965=>"001111011",
  46966=>"101100011",
  46967=>"000011111",
  46968=>"111111101",
  46969=>"011001100",
  46970=>"000001011",
  46971=>"000100101",
  46972=>"110001000",
  46973=>"000110111",
  46974=>"000001000",
  46975=>"110111100",
  46976=>"100100011",
  46977=>"111011100",
  46978=>"110111111",
  46979=>"100101011",
  46980=>"111100010",
  46981=>"011001011",
  46982=>"001000110",
  46983=>"100110001",
  46984=>"110011011",
  46985=>"110011100",
  46986=>"101010000",
  46987=>"011110101",
  46988=>"100110001",
  46989=>"010010010",
  46990=>"000100001",
  46991=>"001000001",
  46992=>"101001000",
  46993=>"111111001",
  46994=>"110001011",
  46995=>"111000011",
  46996=>"100101010",
  46997=>"100110100",
  46998=>"001011010",
  46999=>"001100110",
  47000=>"010000110",
  47001=>"010011010",
  47002=>"010010010",
  47003=>"010001111",
  47004=>"111110001",
  47005=>"110010000",
  47006=>"110011011",
  47007=>"100101111",
  47008=>"110111011",
  47009=>"001010011",
  47010=>"001100000",
  47011=>"000100101",
  47012=>"101111001",
  47013=>"111011010",
  47014=>"100001100",
  47015=>"100110101",
  47016=>"001001111",
  47017=>"100111101",
  47018=>"110110100",
  47019=>"010010010",
  47020=>"101001001",
  47021=>"011101000",
  47022=>"101101010",
  47023=>"111110110",
  47024=>"101001001",
  47025=>"000010011",
  47026=>"000010011",
  47027=>"000111000",
  47028=>"000000110",
  47029=>"000000110",
  47030=>"111000101",
  47031=>"101100110",
  47032=>"110111111",
  47033=>"001101011",
  47034=>"000000011",
  47035=>"010101001",
  47036=>"100100011",
  47037=>"100100110",
  47038=>"101110111",
  47039=>"011101000",
  47040=>"001000001",
  47041=>"111000111",
  47042=>"010100101",
  47043=>"000011000",
  47044=>"100010000",
  47045=>"010111010",
  47046=>"000011111",
  47047=>"001011101",
  47048=>"101100100",
  47049=>"110100001",
  47050=>"011111001",
  47051=>"010101000",
  47052=>"001010011",
  47053=>"001111011",
  47054=>"000001011",
  47055=>"111001111",
  47056=>"011111110",
  47057=>"110001111",
  47058=>"001100100",
  47059=>"110101111",
  47060=>"011001110",
  47061=>"001101000",
  47062=>"100111100",
  47063=>"010101110",
  47064=>"001010010",
  47065=>"001011011",
  47066=>"010000010",
  47067=>"000001010",
  47068=>"111110111",
  47069=>"100000100",
  47070=>"110010010",
  47071=>"100100101",
  47072=>"101111110",
  47073=>"100001000",
  47074=>"000101000",
  47075=>"011001011",
  47076=>"100101001",
  47077=>"000001001",
  47078=>"000100100",
  47079=>"110100100",
  47080=>"110110111",
  47081=>"000000101",
  47082=>"011010101",
  47083=>"110011111",
  47084=>"010010000",
  47085=>"011110100",
  47086=>"110010001",
  47087=>"001111011",
  47088=>"011001101",
  47089=>"001001011",
  47090=>"111110000",
  47091=>"000000101",
  47092=>"101010011",
  47093=>"000000000",
  47094=>"100000100",
  47095=>"101000000",
  47096=>"010011101",
  47097=>"001010101",
  47098=>"010011111",
  47099=>"100111111",
  47100=>"001111101",
  47101=>"101101000",
  47102=>"100110110",
  47103=>"111000010",
  47104=>"000110100",
  47105=>"111101001",
  47106=>"110111111",
  47107=>"110101111",
  47108=>"011101000",
  47109=>"000110010",
  47110=>"101011111",
  47111=>"111011001",
  47112=>"110000100",
  47113=>"000001011",
  47114=>"100100000",
  47115=>"111101111",
  47116=>"001010110",
  47117=>"111010000",
  47118=>"011010000",
  47119=>"101001110",
  47120=>"100011111",
  47121=>"011001010",
  47122=>"011010000",
  47123=>"001001101",
  47124=>"000001010",
  47125=>"110011000",
  47126=>"011110100",
  47127=>"010001101",
  47128=>"000110100",
  47129=>"101000101",
  47130=>"111010111",
  47131=>"101111011",
  47132=>"111010111",
  47133=>"111000100",
  47134=>"001111001",
  47135=>"100101000",
  47136=>"000010011",
  47137=>"010110100",
  47138=>"001000000",
  47139=>"001001000",
  47140=>"011000000",
  47141=>"111000101",
  47142=>"111000101",
  47143=>"000011110",
  47144=>"000000001",
  47145=>"000110000",
  47146=>"111010110",
  47147=>"110100000",
  47148=>"001011100",
  47149=>"111000111",
  47150=>"101110101",
  47151=>"000111001",
  47152=>"010101000",
  47153=>"011011011",
  47154=>"111110110",
  47155=>"010011010",
  47156=>"010010100",
  47157=>"101001011",
  47158=>"100000110",
  47159=>"010010101",
  47160=>"011010101",
  47161=>"010101101",
  47162=>"110101011",
  47163=>"101101100",
  47164=>"011010000",
  47165=>"001111101",
  47166=>"110001000",
  47167=>"000110000",
  47168=>"011001010",
  47169=>"111011000",
  47170=>"011000111",
  47171=>"011010101",
  47172=>"011111100",
  47173=>"011110100",
  47174=>"100101011",
  47175=>"111111010",
  47176=>"000100101",
  47177=>"110010000",
  47178=>"111110000",
  47179=>"000001111",
  47180=>"101101000",
  47181=>"111111100",
  47182=>"011000000",
  47183=>"001001011",
  47184=>"110011010",
  47185=>"101010110",
  47186=>"010110101",
  47187=>"100000110",
  47188=>"111000011",
  47189=>"111010110",
  47190=>"100001111",
  47191=>"101101110",
  47192=>"010011001",
  47193=>"110101011",
  47194=>"110011011",
  47195=>"101001010",
  47196=>"110101111",
  47197=>"110100101",
  47198=>"111110000",
  47199=>"011110111",
  47200=>"110000111",
  47201=>"110010011",
  47202=>"010100010",
  47203=>"111111010",
  47204=>"010001111",
  47205=>"110011100",
  47206=>"110011001",
  47207=>"101110110",
  47208=>"100000001",
  47209=>"010011010",
  47210=>"111010100",
  47211=>"100110001",
  47212=>"011100110",
  47213=>"101001010",
  47214=>"001001011",
  47215=>"100000000",
  47216=>"111111110",
  47217=>"000100011",
  47218=>"011011101",
  47219=>"111101101",
  47220=>"101011111",
  47221=>"110000110",
  47222=>"001100111",
  47223=>"100000001",
  47224=>"010100000",
  47225=>"111001010",
  47226=>"111000000",
  47227=>"111101001",
  47228=>"000011010",
  47229=>"000001011",
  47230=>"110010000",
  47231=>"111111010",
  47232=>"000000111",
  47233=>"001010101",
  47234=>"001001111",
  47235=>"111101010",
  47236=>"111010100",
  47237=>"000101111",
  47238=>"100110110",
  47239=>"000111011",
  47240=>"010010011",
  47241=>"000101100",
  47242=>"100001000",
  47243=>"110110110",
  47244=>"111010001",
  47245=>"100100100",
  47246=>"101101010",
  47247=>"010011011",
  47248=>"000111011",
  47249=>"011100000",
  47250=>"001001110",
  47251=>"011010001",
  47252=>"100011101",
  47253=>"101010111",
  47254=>"100011001",
  47255=>"000000100",
  47256=>"100101100",
  47257=>"100011011",
  47258=>"011100110",
  47259=>"001011101",
  47260=>"111110101",
  47261=>"000100101",
  47262=>"101111010",
  47263=>"111000000",
  47264=>"000000101",
  47265=>"110001100",
  47266=>"100001111",
  47267=>"001010001",
  47268=>"110111110",
  47269=>"110101110",
  47270=>"010010000",
  47271=>"001010101",
  47272=>"111111011",
  47273=>"001001111",
  47274=>"010100011",
  47275=>"000011011",
  47276=>"001001011",
  47277=>"010101111",
  47278=>"101111001",
  47279=>"100100011",
  47280=>"101101011",
  47281=>"000000010",
  47282=>"110110111",
  47283=>"001001111",
  47284=>"011010111",
  47285=>"010010100",
  47286=>"001010111",
  47287=>"111011000",
  47288=>"010111001",
  47289=>"100010111",
  47290=>"000110000",
  47291=>"100101101",
  47292=>"110100111",
  47293=>"011011100",
  47294=>"111101000",
  47295=>"011100001",
  47296=>"111100001",
  47297=>"111011110",
  47298=>"111011110",
  47299=>"100000110",
  47300=>"100010001",
  47301=>"111111011",
  47302=>"000001101",
  47303=>"101111001",
  47304=>"001001001",
  47305=>"111010110",
  47306=>"111101101",
  47307=>"001110100",
  47308=>"001111010",
  47309=>"100111001",
  47310=>"100011110",
  47311=>"110000101",
  47312=>"000001000",
  47313=>"001011010",
  47314=>"101101100",
  47315=>"010110000",
  47316=>"000010000",
  47317=>"000100101",
  47318=>"001000110",
  47319=>"001000111",
  47320=>"101010011",
  47321=>"101011010",
  47322=>"101001101",
  47323=>"100110011",
  47324=>"101111101",
  47325=>"101100001",
  47326=>"000110111",
  47327=>"011011000",
  47328=>"001111100",
  47329=>"110010110",
  47330=>"101110010",
  47331=>"101001100",
  47332=>"111111001",
  47333=>"001001010",
  47334=>"100111100",
  47335=>"100000011",
  47336=>"010100011",
  47337=>"010100000",
  47338=>"110101011",
  47339=>"001001011",
  47340=>"100000100",
  47341=>"101010111",
  47342=>"011011100",
  47343=>"001000001",
  47344=>"000110000",
  47345=>"110100101",
  47346=>"001000000",
  47347=>"101111111",
  47348=>"101011011",
  47349=>"000010111",
  47350=>"010110000",
  47351=>"011111111",
  47352=>"110010001",
  47353=>"100000111",
  47354=>"011010110",
  47355=>"110011000",
  47356=>"111001001",
  47357=>"100100101",
  47358=>"011110110",
  47359=>"011110110",
  47360=>"001111001",
  47361=>"010011100",
  47362=>"001111000",
  47363=>"011001100",
  47364=>"001010010",
  47365=>"010011011",
  47366=>"100101110",
  47367=>"110100111",
  47368=>"011001111",
  47369=>"101001000",
  47370=>"010001000",
  47371=>"111011000",
  47372=>"111011001",
  47373=>"111101001",
  47374=>"011011001",
  47375=>"111100000",
  47376=>"010101001",
  47377=>"110110001",
  47378=>"000101100",
  47379=>"111100111",
  47380=>"100011110",
  47381=>"110111101",
  47382=>"001111011",
  47383=>"111111101",
  47384=>"110000101",
  47385=>"101011001",
  47386=>"001010101",
  47387=>"111001011",
  47388=>"000001111",
  47389=>"100000000",
  47390=>"001010001",
  47391=>"000100001",
  47392=>"100001010",
  47393=>"111100000",
  47394=>"000111111",
  47395=>"000111010",
  47396=>"001011101",
  47397=>"101100001",
  47398=>"001010101",
  47399=>"011110111",
  47400=>"010110111",
  47401=>"000000001",
  47402=>"011100111",
  47403=>"101111010",
  47404=>"110010000",
  47405=>"100100001",
  47406=>"010110111",
  47407=>"010100011",
  47408=>"010110000",
  47409=>"100000110",
  47410=>"010101000",
  47411=>"001001000",
  47412=>"011101010",
  47413=>"001100101",
  47414=>"111000101",
  47415=>"010101000",
  47416=>"000000010",
  47417=>"111011011",
  47418=>"110001100",
  47419=>"000001101",
  47420=>"111101110",
  47421=>"000110100",
  47422=>"111110001",
  47423=>"111110001",
  47424=>"000001101",
  47425=>"101011111",
  47426=>"001101111",
  47427=>"000100011",
  47428=>"011111101",
  47429=>"111100110",
  47430=>"010110011",
  47431=>"001100100",
  47432=>"110110010",
  47433=>"000001000",
  47434=>"000110011",
  47435=>"101111100",
  47436=>"011001001",
  47437=>"010111110",
  47438=>"001010110",
  47439=>"101101010",
  47440=>"110100000",
  47441=>"101011001",
  47442=>"100111111",
  47443=>"011111101",
  47444=>"111100111",
  47445=>"110000011",
  47446=>"100110001",
  47447=>"010111110",
  47448=>"100111110",
  47449=>"101000110",
  47450=>"100110101",
  47451=>"101011000",
  47452=>"111011001",
  47453=>"101110111",
  47454=>"000000100",
  47455=>"101000110",
  47456=>"110101111",
  47457=>"100111110",
  47458=>"011001100",
  47459=>"000110110",
  47460=>"111011101",
  47461=>"000101100",
  47462=>"001110010",
  47463=>"001111001",
  47464=>"110100001",
  47465=>"000110110",
  47466=>"010010100",
  47467=>"000000001",
  47468=>"100010101",
  47469=>"011011001",
  47470=>"000000001",
  47471=>"001100111",
  47472=>"000001011",
  47473=>"011001000",
  47474=>"101110100",
  47475=>"001011011",
  47476=>"110010101",
  47477=>"110001000",
  47478=>"011111001",
  47479=>"100101101",
  47480=>"101100101",
  47481=>"001011001",
  47482=>"011110000",
  47483=>"101111101",
  47484=>"110101001",
  47485=>"010011111",
  47486=>"101011111",
  47487=>"000000110",
  47488=>"000000000",
  47489=>"000100100",
  47490=>"111101111",
  47491=>"001011100",
  47492=>"001111111",
  47493=>"110000010",
  47494=>"111110100",
  47495=>"010011110",
  47496=>"001000000",
  47497=>"000101101",
  47498=>"110100011",
  47499=>"101111010",
  47500=>"000111101",
  47501=>"010010110",
  47502=>"011101001",
  47503=>"011001110",
  47504=>"000010101",
  47505=>"000110000",
  47506=>"101100001",
  47507=>"011010101",
  47508=>"110101101",
  47509=>"100100111",
  47510=>"011011110",
  47511=>"110100111",
  47512=>"011100011",
  47513=>"001010011",
  47514=>"110011001",
  47515=>"100001001",
  47516=>"001011000",
  47517=>"100001101",
  47518=>"010000110",
  47519=>"111100000",
  47520=>"110010010",
  47521=>"000001110",
  47522=>"111000011",
  47523=>"001111110",
  47524=>"111111000",
  47525=>"010011111",
  47526=>"001000000",
  47527=>"001000110",
  47528=>"110110111",
  47529=>"101001100",
  47530=>"010101010",
  47531=>"100110101",
  47532=>"111100011",
  47533=>"100110000",
  47534=>"011000100",
  47535=>"001100011",
  47536=>"000011110",
  47537=>"111001110",
  47538=>"010010110",
  47539=>"010110000",
  47540=>"011101101",
  47541=>"100100100",
  47542=>"001111010",
  47543=>"010001010",
  47544=>"111110010",
  47545=>"010011110",
  47546=>"001101001",
  47547=>"011111110",
  47548=>"111110110",
  47549=>"111000101",
  47550=>"010011101",
  47551=>"010101110",
  47552=>"000001100",
  47553=>"101111111",
  47554=>"100011000",
  47555=>"000011011",
  47556=>"010000111",
  47557=>"010000101",
  47558=>"100001010",
  47559=>"100001000",
  47560=>"001001111",
  47561=>"111010101",
  47562=>"000000011",
  47563=>"010010001",
  47564=>"001011000",
  47565=>"100001000",
  47566=>"110011001",
  47567=>"100001000",
  47568=>"111001100",
  47569=>"011001001",
  47570=>"001110100",
  47571=>"111001100",
  47572=>"010110000",
  47573=>"000010100",
  47574=>"011101000",
  47575=>"010000010",
  47576=>"100111011",
  47577=>"000011101",
  47578=>"101100000",
  47579=>"000010101",
  47580=>"100011000",
  47581=>"101111110",
  47582=>"010100110",
  47583=>"001011010",
  47584=>"001101111",
  47585=>"100100000",
  47586=>"111101000",
  47587=>"110111011",
  47588=>"111101100",
  47589=>"110100010",
  47590=>"001010001",
  47591=>"110110101",
  47592=>"110111011",
  47593=>"101110110",
  47594=>"000110100",
  47595=>"000000001",
  47596=>"100111010",
  47597=>"101011011",
  47598=>"110111101",
  47599=>"001111011",
  47600=>"100111101",
  47601=>"100011101",
  47602=>"111111010",
  47603=>"110010010",
  47604=>"000111100",
  47605=>"010100000",
  47606=>"011011011",
  47607=>"100111000",
  47608=>"101101101",
  47609=>"010011001",
  47610=>"111000101",
  47611=>"101011000",
  47612=>"001000100",
  47613=>"001000110",
  47614=>"111101111",
  47615=>"010100001",
  47616=>"000111110",
  47617=>"010010001",
  47618=>"010111010",
  47619=>"101111000",
  47620=>"110000011",
  47621=>"111110010",
  47622=>"010010101",
  47623=>"000101001",
  47624=>"010101100",
  47625=>"001111110",
  47626=>"111110111",
  47627=>"100100001",
  47628=>"100001010",
  47629=>"010011001",
  47630=>"100001110",
  47631=>"010111001",
  47632=>"101010011",
  47633=>"100110100",
  47634=>"100100001",
  47635=>"101100001",
  47636=>"001000110",
  47637=>"110000101",
  47638=>"111100100",
  47639=>"110101110",
  47640=>"000001010",
  47641=>"101001000",
  47642=>"001001110",
  47643=>"110011001",
  47644=>"001100110",
  47645=>"111010100",
  47646=>"000111001",
  47647=>"111110000",
  47648=>"101100111",
  47649=>"100110111",
  47650=>"110001000",
  47651=>"001101010",
  47652=>"111011010",
  47653=>"001000001",
  47654=>"111010100",
  47655=>"100111010",
  47656=>"100001100",
  47657=>"110011011",
  47658=>"011000100",
  47659=>"111010010",
  47660=>"111001110",
  47661=>"001011000",
  47662=>"001001100",
  47663=>"110011101",
  47664=>"010101011",
  47665=>"010100011",
  47666=>"100011010",
  47667=>"011000101",
  47668=>"011010000",
  47669=>"110010010",
  47670=>"000100100",
  47671=>"110000001",
  47672=>"000101010",
  47673=>"010100110",
  47674=>"101110001",
  47675=>"100111111",
  47676=>"010000001",
  47677=>"110001100",
  47678=>"111000000",
  47679=>"111101010",
  47680=>"110000111",
  47681=>"111100100",
  47682=>"111111101",
  47683=>"000001111",
  47684=>"110011001",
  47685=>"010001101",
  47686=>"001010001",
  47687=>"110010000",
  47688=>"001111101",
  47689=>"101010110",
  47690=>"010110010",
  47691=>"010101000",
  47692=>"101011100",
  47693=>"010010011",
  47694=>"111110011",
  47695=>"000110011",
  47696=>"100100001",
  47697=>"101100110",
  47698=>"101000001",
  47699=>"100000011",
  47700=>"000001111",
  47701=>"000001000",
  47702=>"000001101",
  47703=>"011110001",
  47704=>"110011110",
  47705=>"101110000",
  47706=>"001000100",
  47707=>"000101010",
  47708=>"000010110",
  47709=>"110001101",
  47710=>"011000101",
  47711=>"100101001",
  47712=>"000100000",
  47713=>"000100001",
  47714=>"111111100",
  47715=>"011011011",
  47716=>"110010111",
  47717=>"101111100",
  47718=>"101110010",
  47719=>"010110000",
  47720=>"001110101",
  47721=>"100100000",
  47722=>"000011111",
  47723=>"010101100",
  47724=>"011110100",
  47725=>"010011110",
  47726=>"010001111",
  47727=>"011101000",
  47728=>"010101110",
  47729=>"110110011",
  47730=>"101100101",
  47731=>"011101010",
  47732=>"011110000",
  47733=>"001101010",
  47734=>"111010110",
  47735=>"110101110",
  47736=>"010000000",
  47737=>"010010100",
  47738=>"001011011",
  47739=>"011011001",
  47740=>"001001010",
  47741=>"110110000",
  47742=>"110110000",
  47743=>"111010001",
  47744=>"111101000",
  47745=>"000100010",
  47746=>"110100111",
  47747=>"001000011",
  47748=>"001010100",
  47749=>"100101000",
  47750=>"110001010",
  47751=>"111001100",
  47752=>"011010011",
  47753=>"000010110",
  47754=>"101001111",
  47755=>"010111001",
  47756=>"111110101",
  47757=>"111001010",
  47758=>"100110110",
  47759=>"101010100",
  47760=>"010101100",
  47761=>"100000010",
  47762=>"100111101",
  47763=>"111010011",
  47764=>"011001101",
  47765=>"011011111",
  47766=>"010110010",
  47767=>"100101000",
  47768=>"001000110",
  47769=>"000010100",
  47770=>"110110011",
  47771=>"001000010",
  47772=>"101110001",
  47773=>"000110011",
  47774=>"010011001",
  47775=>"100010000",
  47776=>"001001100",
  47777=>"100110000",
  47778=>"100011111",
  47779=>"101010101",
  47780=>"000001010",
  47781=>"011111000",
  47782=>"100000110",
  47783=>"010000101",
  47784=>"110000110",
  47785=>"010111111",
  47786=>"000010010",
  47787=>"111000100",
  47788=>"000010101",
  47789=>"101000101",
  47790=>"111000111",
  47791=>"010011001",
  47792=>"101110000",
  47793=>"010110000",
  47794=>"010110000",
  47795=>"011111100",
  47796=>"111011010",
  47797=>"111010110",
  47798=>"111000110",
  47799=>"001001101",
  47800=>"010101011",
  47801=>"000101110",
  47802=>"001000000",
  47803=>"101010101",
  47804=>"100010111",
  47805=>"101101010",
  47806=>"000101110",
  47807=>"110101111",
  47808=>"111001010",
  47809=>"100010110",
  47810=>"001000011",
  47811=>"011000100",
  47812=>"100001010",
  47813=>"000110010",
  47814=>"000010100",
  47815=>"011010101",
  47816=>"101110101",
  47817=>"011111111",
  47818=>"111001001",
  47819=>"000001100",
  47820=>"100110000",
  47821=>"111010101",
  47822=>"111011111",
  47823=>"111010111",
  47824=>"001111111",
  47825=>"111110010",
  47826=>"011100100",
  47827=>"101101110",
  47828=>"101001010",
  47829=>"100101101",
  47830=>"010010100",
  47831=>"100100111",
  47832=>"100100101",
  47833=>"110001111",
  47834=>"100001011",
  47835=>"000011101",
  47836=>"001001001",
  47837=>"110011111",
  47838=>"011001111",
  47839=>"001100110",
  47840=>"011011100",
  47841=>"000011110",
  47842=>"001111100",
  47843=>"101011110",
  47844=>"010101100",
  47845=>"101110001",
  47846=>"001010001",
  47847=>"110001100",
  47848=>"100010010",
  47849=>"000101111",
  47850=>"111011111",
  47851=>"010000100",
  47852=>"000110111",
  47853=>"100100011",
  47854=>"111110101",
  47855=>"000011011",
  47856=>"110111011",
  47857=>"110010100",
  47858=>"010010001",
  47859=>"001011110",
  47860=>"010000111",
  47861=>"111111101",
  47862=>"111010101",
  47863=>"101111110",
  47864=>"001110101",
  47865=>"011000100",
  47866=>"100101111",
  47867=>"010110011",
  47868=>"001011010",
  47869=>"111001001",
  47870=>"011101111",
  47871=>"100111010",
  47872=>"110110011",
  47873=>"011001010",
  47874=>"111010101",
  47875=>"000000100",
  47876=>"100011111",
  47877=>"000000110",
  47878=>"001110011",
  47879=>"111100111",
  47880=>"001000101",
  47881=>"000001111",
  47882=>"011110111",
  47883=>"011100101",
  47884=>"011011000",
  47885=>"110000101",
  47886=>"000100010",
  47887=>"101010011",
  47888=>"000010111",
  47889=>"110110100",
  47890=>"011100111",
  47891=>"011000010",
  47892=>"101101100",
  47893=>"101001111",
  47894=>"010100101",
  47895=>"101100101",
  47896=>"001100101",
  47897=>"000100000",
  47898=>"111111111",
  47899=>"000010000",
  47900=>"001100000",
  47901=>"011001000",
  47902=>"101010011",
  47903=>"010100111",
  47904=>"110000101",
  47905=>"011010001",
  47906=>"011100001",
  47907=>"111000100",
  47908=>"101010011",
  47909=>"010011010",
  47910=>"010111100",
  47911=>"011110001",
  47912=>"110110100",
  47913=>"111101101",
  47914=>"100010100",
  47915=>"110011101",
  47916=>"101100110",
  47917=>"111001000",
  47918=>"111110000",
  47919=>"110111001",
  47920=>"101110000",
  47921=>"101000101",
  47922=>"001101010",
  47923=>"101111011",
  47924=>"110111111",
  47925=>"111100111",
  47926=>"000000010",
  47927=>"101101101",
  47928=>"111010010",
  47929=>"101001110",
  47930=>"011010000",
  47931=>"110101000",
  47932=>"110100111",
  47933=>"101110101",
  47934=>"111110111",
  47935=>"111011000",
  47936=>"111000111",
  47937=>"101110110",
  47938=>"101011010",
  47939=>"010000001",
  47940=>"110111001",
  47941=>"010010111",
  47942=>"000000110",
  47943=>"101001110",
  47944=>"001000001",
  47945=>"001000010",
  47946=>"101001001",
  47947=>"110101001",
  47948=>"110101110",
  47949=>"100101101",
  47950=>"001000000",
  47951=>"101100001",
  47952=>"000010000",
  47953=>"101110000",
  47954=>"100010010",
  47955=>"001001001",
  47956=>"110110001",
  47957=>"111011111",
  47958=>"100011011",
  47959=>"100100110",
  47960=>"001000101",
  47961=>"001101010",
  47962=>"110011100",
  47963=>"001000100",
  47964=>"000001100",
  47965=>"000000000",
  47966=>"011000011",
  47967=>"000111001",
  47968=>"100111111",
  47969=>"100100011",
  47970=>"110100011",
  47971=>"110110111",
  47972=>"001101100",
  47973=>"001001110",
  47974=>"111001100",
  47975=>"110100100",
  47976=>"000100110",
  47977=>"001011000",
  47978=>"110011000",
  47979=>"010100111",
  47980=>"000001010",
  47981=>"001000001",
  47982=>"010000110",
  47983=>"111111100",
  47984=>"010010010",
  47985=>"000000010",
  47986=>"001101011",
  47987=>"011010010",
  47988=>"010000101",
  47989=>"101001101",
  47990=>"011111111",
  47991=>"101001011",
  47992=>"000000000",
  47993=>"100010111",
  47994=>"001101000",
  47995=>"001010001",
  47996=>"110100010",
  47997=>"001010010",
  47998=>"001100000",
  47999=>"110101111",
  48000=>"101010100",
  48001=>"000110110",
  48002=>"001001100",
  48003=>"010010011",
  48004=>"111110100",
  48005=>"111000001",
  48006=>"010111111",
  48007=>"110110100",
  48008=>"011011110",
  48009=>"110110100",
  48010=>"010010101",
  48011=>"111011101",
  48012=>"010011111",
  48013=>"100001111",
  48014=>"101011010",
  48015=>"111100010",
  48016=>"101100100",
  48017=>"000010000",
  48018=>"000001111",
  48019=>"011111101",
  48020=>"111100110",
  48021=>"110010011",
  48022=>"100110001",
  48023=>"010010111",
  48024=>"001001100",
  48025=>"001100010",
  48026=>"011000000",
  48027=>"011011101",
  48028=>"010010100",
  48029=>"000101001",
  48030=>"010101001",
  48031=>"001001111",
  48032=>"101000111",
  48033=>"101110111",
  48034=>"001001011",
  48035=>"000100000",
  48036=>"101011101",
  48037=>"001111111",
  48038=>"011001101",
  48039=>"110001111",
  48040=>"100000101",
  48041=>"011011101",
  48042=>"111000100",
  48043=>"010010001",
  48044=>"001000100",
  48045=>"001011000",
  48046=>"100010010",
  48047=>"111001001",
  48048=>"000100010",
  48049=>"101010001",
  48050=>"110100110",
  48051=>"010100111",
  48052=>"101101101",
  48053=>"111000101",
  48054=>"010000110",
  48055=>"010001011",
  48056=>"110000010",
  48057=>"011010101",
  48058=>"100000010",
  48059=>"010101010",
  48060=>"010010110",
  48061=>"100010111",
  48062=>"001100001",
  48063=>"011011000",
  48064=>"001111101",
  48065=>"010000111",
  48066=>"101100000",
  48067=>"011000110",
  48068=>"110000110",
  48069=>"110110000",
  48070=>"111111011",
  48071=>"111100011",
  48072=>"000001111",
  48073=>"100011100",
  48074=>"110001000",
  48075=>"100010101",
  48076=>"011011001",
  48077=>"100001010",
  48078=>"011001010",
  48079=>"100110000",
  48080=>"010100111",
  48081=>"110011100",
  48082=>"111011111",
  48083=>"010011010",
  48084=>"000100100",
  48085=>"101000000",
  48086=>"001101001",
  48087=>"100011100",
  48088=>"001001100",
  48089=>"000010101",
  48090=>"001000000",
  48091=>"101100101",
  48092=>"001001110",
  48093=>"011100001",
  48094=>"001000110",
  48095=>"011110100",
  48096=>"011110011",
  48097=>"011101100",
  48098=>"001100011",
  48099=>"001111000",
  48100=>"111101000",
  48101=>"000000001",
  48102=>"000010001",
  48103=>"000101110",
  48104=>"000000110",
  48105=>"111100110",
  48106=>"001110011",
  48107=>"000010001",
  48108=>"010110111",
  48109=>"100000011",
  48110=>"001100000",
  48111=>"100001110",
  48112=>"111011101",
  48113=>"111111011",
  48114=>"000000111",
  48115=>"100000010",
  48116=>"000011011",
  48117=>"011001000",
  48118=>"001110001",
  48119=>"111101101",
  48120=>"000001010",
  48121=>"111101111",
  48122=>"001011101",
  48123=>"000101111",
  48124=>"100010110",
  48125=>"000010000",
  48126=>"111100000",
  48127=>"110000110",
  48128=>"011000110",
  48129=>"111011111",
  48130=>"011111110",
  48131=>"101011010",
  48132=>"101101100",
  48133=>"100111010",
  48134=>"101101100",
  48135=>"111101110",
  48136=>"001001010",
  48137=>"000001000",
  48138=>"101000100",
  48139=>"110011101",
  48140=>"011111100",
  48141=>"110110011",
  48142=>"010011001",
  48143=>"101101000",
  48144=>"011000011",
  48145=>"100001111",
  48146=>"001101110",
  48147=>"000100011",
  48148=>"010000000",
  48149=>"000000000",
  48150=>"111001111",
  48151=>"110000010",
  48152=>"110000001",
  48153=>"001101001",
  48154=>"101101010",
  48155=>"011100100",
  48156=>"011111111",
  48157=>"110111011",
  48158=>"100101010",
  48159=>"111010110",
  48160=>"110000111",
  48161=>"101010101",
  48162=>"111101111",
  48163=>"000000111",
  48164=>"111101100",
  48165=>"001100000",
  48166=>"000101011",
  48167=>"110011001",
  48168=>"110010010",
  48169=>"101111110",
  48170=>"000001000",
  48171=>"110100000",
  48172=>"110111001",
  48173=>"000001001",
  48174=>"010000000",
  48175=>"100011000",
  48176=>"101010110",
  48177=>"000000101",
  48178=>"101010011",
  48179=>"000111000",
  48180=>"010001000",
  48181=>"010010110",
  48182=>"110110100",
  48183=>"101100111",
  48184=>"001000100",
  48185=>"101010010",
  48186=>"000101011",
  48187=>"010100110",
  48188=>"000001100",
  48189=>"010001000",
  48190=>"000101000",
  48191=>"010110011",
  48192=>"111011000",
  48193=>"000010010",
  48194=>"000010111",
  48195=>"000110111",
  48196=>"000000111",
  48197=>"000001100",
  48198=>"110000011",
  48199=>"001000001",
  48200=>"111001100",
  48201=>"000111111",
  48202=>"100101100",
  48203=>"110000110",
  48204=>"101010100",
  48205=>"001110111",
  48206=>"100111000",
  48207=>"000010000",
  48208=>"011101001",
  48209=>"111101100",
  48210=>"101111111",
  48211=>"000110110",
  48212=>"100100011",
  48213=>"101110011",
  48214=>"011101100",
  48215=>"000000111",
  48216=>"110111101",
  48217=>"111010011",
  48218=>"110010100",
  48219=>"010010000",
  48220=>"001001000",
  48221=>"100111101",
  48222=>"001001110",
  48223=>"101000100",
  48224=>"000110101",
  48225=>"101001000",
  48226=>"010110100",
  48227=>"111101111",
  48228=>"010000001",
  48229=>"011111011",
  48230=>"001101000",
  48231=>"010111010",
  48232=>"011000010",
  48233=>"011010101",
  48234=>"100111110",
  48235=>"111001110",
  48236=>"001001000",
  48237=>"101110010",
  48238=>"011111010",
  48239=>"011010010",
  48240=>"001001001",
  48241=>"001111111",
  48242=>"001110101",
  48243=>"111000110",
  48244=>"111010011",
  48245=>"110111011",
  48246=>"101011011",
  48247=>"110100111",
  48248=>"111000110",
  48249=>"101010000",
  48250=>"110101000",
  48251=>"101111000",
  48252=>"110100110",
  48253=>"011010000",
  48254=>"011101111",
  48255=>"001101010",
  48256=>"111011000",
  48257=>"111010100",
  48258=>"010100100",
  48259=>"011011111",
  48260=>"000000100",
  48261=>"011000110",
  48262=>"100100100",
  48263=>"101110100",
  48264=>"000101000",
  48265=>"111100001",
  48266=>"000011010",
  48267=>"010011101",
  48268=>"101110101",
  48269=>"011101011",
  48270=>"101000110",
  48271=>"010101011",
  48272=>"110111100",
  48273=>"111111010",
  48274=>"110010111",
  48275=>"001001001",
  48276=>"011000000",
  48277=>"001001010",
  48278=>"100000111",
  48279=>"101010011",
  48280=>"101101111",
  48281=>"000100001",
  48282=>"111001010",
  48283=>"000011110",
  48284=>"101100000",
  48285=>"001010001",
  48286=>"100010000",
  48287=>"001000110",
  48288=>"100111100",
  48289=>"111001011",
  48290=>"101101000",
  48291=>"100000101",
  48292=>"010100011",
  48293=>"010110001",
  48294=>"011000100",
  48295=>"110001100",
  48296=>"001111000",
  48297=>"110011010",
  48298=>"100100111",
  48299=>"101100001",
  48300=>"010101111",
  48301=>"111100010",
  48302=>"111001000",
  48303=>"010010101",
  48304=>"010000000",
  48305=>"010000011",
  48306=>"001000110",
  48307=>"000011100",
  48308=>"001100011",
  48309=>"110000001",
  48310=>"001011110",
  48311=>"101111010",
  48312=>"101111001",
  48313=>"100111010",
  48314=>"001010111",
  48315=>"001001011",
  48316=>"100111100",
  48317=>"010000001",
  48318=>"111101010",
  48319=>"011111101",
  48320=>"001000010",
  48321=>"001011101",
  48322=>"100100001",
  48323=>"000010011",
  48324=>"011101000",
  48325=>"101110000",
  48326=>"111101100",
  48327=>"001011111",
  48328=>"111011111",
  48329=>"101011101",
  48330=>"000001010",
  48331=>"100011001",
  48332=>"111011010",
  48333=>"101110011",
  48334=>"100011000",
  48335=>"101001100",
  48336=>"000000101",
  48337=>"101111100",
  48338=>"000001101",
  48339=>"110101100",
  48340=>"000001011",
  48341=>"111001001",
  48342=>"101110100",
  48343=>"101000110",
  48344=>"010111100",
  48345=>"000000110",
  48346=>"100101010",
  48347=>"011001110",
  48348=>"001000110",
  48349=>"111011101",
  48350=>"001111110",
  48351=>"101010001",
  48352=>"000000011",
  48353=>"101001100",
  48354=>"111011100",
  48355=>"101001100",
  48356=>"100110100",
  48357=>"101101001",
  48358=>"001111000",
  48359=>"001101111",
  48360=>"011111010",
  48361=>"100101001",
  48362=>"011111000",
  48363=>"001001111",
  48364=>"011010011",
  48365=>"111000010",
  48366=>"011001000",
  48367=>"110000101",
  48368=>"110010000",
  48369=>"101101001",
  48370=>"100000000",
  48371=>"001000010",
  48372=>"100111001",
  48373=>"000000010",
  48374=>"101100010",
  48375=>"100110101",
  48376=>"000000001",
  48377=>"011101100",
  48378=>"011100100",
  48379=>"101101100",
  48380=>"001001110",
  48381=>"000110110",
  48382=>"111100111",
  48383=>"101111011",
  48384=>"011000110",
  48385=>"111110001",
  48386=>"111010111",
  48387=>"111111101",
  48388=>"111110101",
  48389=>"001111010",
  48390=>"010000011",
  48391=>"100011110",
  48392=>"011010001",
  48393=>"001001001",
  48394=>"001011001",
  48395=>"000100001",
  48396=>"000000000",
  48397=>"110101011",
  48398=>"011101011",
  48399=>"000011101",
  48400=>"110111100",
  48401=>"111001101",
  48402=>"111010100",
  48403=>"010110001",
  48404=>"000010110",
  48405=>"000011001",
  48406=>"010110111",
  48407=>"111110101",
  48408=>"111100010",
  48409=>"000100010",
  48410=>"011111101",
  48411=>"001111100",
  48412=>"010010110",
  48413=>"111100100",
  48414=>"011011110",
  48415=>"000110001",
  48416=>"000100001",
  48417=>"101011110",
  48418=>"110001000",
  48419=>"100010001",
  48420=>"111011010",
  48421=>"111001011",
  48422=>"000111100",
  48423=>"001110001",
  48424=>"101010010",
  48425=>"100100010",
  48426=>"110110110",
  48427=>"100101001",
  48428=>"111001000",
  48429=>"101111000",
  48430=>"001000101",
  48431=>"000101001",
  48432=>"001010011",
  48433=>"111110111",
  48434=>"001010110",
  48435=>"000001011",
  48436=>"010001110",
  48437=>"010101011",
  48438=>"100100101",
  48439=>"011010011",
  48440=>"000010101",
  48441=>"111001010",
  48442=>"010001000",
  48443=>"111010000",
  48444=>"111000010",
  48445=>"110011010",
  48446=>"001110001",
  48447=>"001111000",
  48448=>"001000110",
  48449=>"100000100",
  48450=>"101000010",
  48451=>"111110110",
  48452=>"010100111",
  48453=>"001110000",
  48454=>"101001111",
  48455=>"110001010",
  48456=>"110010010",
  48457=>"001001000",
  48458=>"110011000",
  48459=>"001101000",
  48460=>"010010111",
  48461=>"111101111",
  48462=>"111100110",
  48463=>"111111100",
  48464=>"101010110",
  48465=>"111011111",
  48466=>"111010011",
  48467=>"111010111",
  48468=>"011001000",
  48469=>"100101010",
  48470=>"110111010",
  48471=>"110111100",
  48472=>"010001001",
  48473=>"100000111",
  48474=>"001110000",
  48475=>"101000000",
  48476=>"011010100",
  48477=>"110011011",
  48478=>"110110011",
  48479=>"000110001",
  48480=>"110001010",
  48481=>"010100010",
  48482=>"000011101",
  48483=>"000000110",
  48484=>"100010100",
  48485=>"101011010",
  48486=>"100010101",
  48487=>"001010111",
  48488=>"100000100",
  48489=>"000000000",
  48490=>"001001011",
  48491=>"000111110",
  48492=>"010001000",
  48493=>"101110111",
  48494=>"000100000",
  48495=>"101111001",
  48496=>"011001000",
  48497=>"000100001",
  48498=>"001000111",
  48499=>"001101110",
  48500=>"101010000",
  48501=>"011000000",
  48502=>"010000111",
  48503=>"111000100",
  48504=>"011101111",
  48505=>"110110010",
  48506=>"010101001",
  48507=>"000001011",
  48508=>"100111110",
  48509=>"111101111",
  48510=>"100111010",
  48511=>"011100100",
  48512=>"001100101",
  48513=>"011000011",
  48514=>"001001011",
  48515=>"010001000",
  48516=>"011010111",
  48517=>"001111111",
  48518=>"111101011",
  48519=>"101010110",
  48520=>"010111110",
  48521=>"001101101",
  48522=>"101100000",
  48523=>"111010010",
  48524=>"101001100",
  48525=>"100000010",
  48526=>"100100100",
  48527=>"010001010",
  48528=>"001001011",
  48529=>"101101000",
  48530=>"110111000",
  48531=>"101010010",
  48532=>"010010101",
  48533=>"110000010",
  48534=>"001100011",
  48535=>"110110001",
  48536=>"000101000",
  48537=>"000010000",
  48538=>"010101001",
  48539=>"000000000",
  48540=>"000011101",
  48541=>"010111000",
  48542=>"000110010",
  48543=>"010011111",
  48544=>"100011010",
  48545=>"111110011",
  48546=>"111001000",
  48547=>"000011100",
  48548=>"010100001",
  48549=>"101000001",
  48550=>"000100110",
  48551=>"100101000",
  48552=>"011000101",
  48553=>"110010011",
  48554=>"010100011",
  48555=>"100101100",
  48556=>"000001110",
  48557=>"100011110",
  48558=>"010110110",
  48559=>"100010000",
  48560=>"001101101",
  48561=>"100000000",
  48562=>"001011111",
  48563=>"011010000",
  48564=>"010000100",
  48565=>"100110100",
  48566=>"100011101",
  48567=>"110010001",
  48568=>"110100000",
  48569=>"100110011",
  48570=>"111011000",
  48571=>"110000101",
  48572=>"000001001",
  48573=>"111101010",
  48574=>"101010111",
  48575=>"101100001",
  48576=>"011000101",
  48577=>"010100011",
  48578=>"001110010",
  48579=>"110001001",
  48580=>"100010101",
  48581=>"010111100",
  48582=>"110100010",
  48583=>"101111001",
  48584=>"000001100",
  48585=>"011100101",
  48586=>"111011000",
  48587=>"111000001",
  48588=>"111010101",
  48589=>"010011110",
  48590=>"001110100",
  48591=>"001100000",
  48592=>"100110010",
  48593=>"111010010",
  48594=>"110111011",
  48595=>"110111101",
  48596=>"100001111",
  48597=>"001001010",
  48598=>"000110011",
  48599=>"001100001",
  48600=>"000100110",
  48601=>"001000000",
  48602=>"111010001",
  48603=>"001100101",
  48604=>"110000101",
  48605=>"011010000",
  48606=>"100001100",
  48607=>"010010101",
  48608=>"001000000",
  48609=>"010000101",
  48610=>"100100111",
  48611=>"010100100",
  48612=>"101010101",
  48613=>"001010100",
  48614=>"100101011",
  48615=>"000100110",
  48616=>"100111110",
  48617=>"000110011",
  48618=>"111011100",
  48619=>"001000111",
  48620=>"001111110",
  48621=>"011010000",
  48622=>"001100000",
  48623=>"101101111",
  48624=>"011011111",
  48625=>"010000011",
  48626=>"001001000",
  48627=>"001000110",
  48628=>"110111101",
  48629=>"111000011",
  48630=>"011010010",
  48631=>"110110000",
  48632=>"110110000",
  48633=>"100010111",
  48634=>"110100100",
  48635=>"100100011",
  48636=>"001000101",
  48637=>"100100010",
  48638=>"101101000",
  48639=>"000011011",
  48640=>"111011100",
  48641=>"101000110",
  48642=>"110111101",
  48643=>"001100011",
  48644=>"100110111",
  48645=>"000100011",
  48646=>"001100001",
  48647=>"110010101",
  48648=>"101000110",
  48649=>"101100101",
  48650=>"100101110",
  48651=>"010010100",
  48652=>"000000011",
  48653=>"111110000",
  48654=>"001101011",
  48655=>"010110101",
  48656=>"011100111",
  48657=>"001111000",
  48658=>"010001001",
  48659=>"001101001",
  48660=>"001100101",
  48661=>"110010001",
  48662=>"001111100",
  48663=>"011010011",
  48664=>"010100001",
  48665=>"001100101",
  48666=>"010001101",
  48667=>"111110011",
  48668=>"011001001",
  48669=>"010000100",
  48670=>"000001111",
  48671=>"110010110",
  48672=>"010100010",
  48673=>"001110110",
  48674=>"001111001",
  48675=>"011110000",
  48676=>"010101011",
  48677=>"000111110",
  48678=>"101011001",
  48679=>"110011101",
  48680=>"111000000",
  48681=>"000110001",
  48682=>"010101100",
  48683=>"111011010",
  48684=>"001001000",
  48685=>"001001100",
  48686=>"010100101",
  48687=>"100000101",
  48688=>"111100011",
  48689=>"101011100",
  48690=>"000110001",
  48691=>"010001000",
  48692=>"111000011",
  48693=>"001100000",
  48694=>"100000000",
  48695=>"010001110",
  48696=>"101100101",
  48697=>"111100000",
  48698=>"001000101",
  48699=>"100101001",
  48700=>"000101001",
  48701=>"100010110",
  48702=>"001100111",
  48703=>"101000101",
  48704=>"000100101",
  48705=>"100001001",
  48706=>"100110101",
  48707=>"100101111",
  48708=>"100000101",
  48709=>"011000001",
  48710=>"100110001",
  48711=>"101010010",
  48712=>"101010011",
  48713=>"011010010",
  48714=>"110000000",
  48715=>"011011110",
  48716=>"111001001",
  48717=>"100001001",
  48718=>"100000000",
  48719=>"010110100",
  48720=>"010000000",
  48721=>"000110000",
  48722=>"000100010",
  48723=>"000000001",
  48724=>"010010010",
  48725=>"010101100",
  48726=>"000001111",
  48727=>"111101100",
  48728=>"011001101",
  48729=>"011011100",
  48730=>"010111110",
  48731=>"001000101",
  48732=>"001000110",
  48733=>"000000001",
  48734=>"000101011",
  48735=>"010100000",
  48736=>"111001111",
  48737=>"100101010",
  48738=>"110111111",
  48739=>"110000110",
  48740=>"110001101",
  48741=>"111100110",
  48742=>"111101111",
  48743=>"101000111",
  48744=>"000101000",
  48745=>"100111000",
  48746=>"001100101",
  48747=>"011100000",
  48748=>"101011010",
  48749=>"101000000",
  48750=>"111011010",
  48751=>"110111111",
  48752=>"010110101",
  48753=>"100000000",
  48754=>"001011111",
  48755=>"010000111",
  48756=>"001100011",
  48757=>"111001000",
  48758=>"110010000",
  48759=>"000010011",
  48760=>"000000100",
  48761=>"101101000",
  48762=>"010100100",
  48763=>"010000101",
  48764=>"001110111",
  48765=>"010100100",
  48766=>"001000110",
  48767=>"011111101",
  48768=>"110011101",
  48769=>"101101100",
  48770=>"010101110",
  48771=>"100000000",
  48772=>"010001010",
  48773=>"100011110",
  48774=>"001101010",
  48775=>"101100011",
  48776=>"100101010",
  48777=>"001011001",
  48778=>"110110101",
  48779=>"001000101",
  48780=>"000001000",
  48781=>"100000000",
  48782=>"110101001",
  48783=>"001110000",
  48784=>"101000101",
  48785=>"010101011",
  48786=>"001011111",
  48787=>"000100110",
  48788=>"101100101",
  48789=>"101001100",
  48790=>"101100110",
  48791=>"101111010",
  48792=>"100010100",
  48793=>"101111110",
  48794=>"111110100",
  48795=>"111011011",
  48796=>"000001001",
  48797=>"010010001",
  48798=>"001011110",
  48799=>"111000011",
  48800=>"010101000",
  48801=>"011110001",
  48802=>"001000010",
  48803=>"110000100",
  48804=>"001100110",
  48805=>"100010010",
  48806=>"111011000",
  48807=>"000100000",
  48808=>"000011000",
  48809=>"111000000",
  48810=>"000011000",
  48811=>"100010100",
  48812=>"111010001",
  48813=>"000011110",
  48814=>"010101011",
  48815=>"010111101",
  48816=>"001100111",
  48817=>"011100011",
  48818=>"000101110",
  48819=>"100100001",
  48820=>"101111101",
  48821=>"010111001",
  48822=>"011001111",
  48823=>"001101111",
  48824=>"101011000",
  48825=>"011111000",
  48826=>"010110110",
  48827=>"100000010",
  48828=>"000100001",
  48829=>"011001010",
  48830=>"010101110",
  48831=>"010010101",
  48832=>"001100100",
  48833=>"010100010",
  48834=>"010101100",
  48835=>"000011001",
  48836=>"100000100",
  48837=>"100011000",
  48838=>"001110011",
  48839=>"110010110",
  48840=>"101011000",
  48841=>"001111000",
  48842=>"000100011",
  48843=>"010111010",
  48844=>"000111001",
  48845=>"001000111",
  48846=>"100001100",
  48847=>"000110000",
  48848=>"010110101",
  48849=>"011110111",
  48850=>"111110011",
  48851=>"000100101",
  48852=>"010110110",
  48853=>"101011011",
  48854=>"101111111",
  48855=>"101000110",
  48856=>"000001110",
  48857=>"101010101",
  48858=>"010010000",
  48859=>"110001001",
  48860=>"001001000",
  48861=>"001011010",
  48862=>"100011000",
  48863=>"001000010",
  48864=>"110001100",
  48865=>"000110100",
  48866=>"111101110",
  48867=>"011001111",
  48868=>"101010010",
  48869=>"110100000",
  48870=>"011010101",
  48871=>"000100111",
  48872=>"011100101",
  48873=>"011011111",
  48874=>"111010001",
  48875=>"001001110",
  48876=>"010111100",
  48877=>"110011000",
  48878=>"111110001",
  48879=>"001001001",
  48880=>"011101110",
  48881=>"001110101",
  48882=>"111110111",
  48883=>"111010101",
  48884=>"010000010",
  48885=>"001100100",
  48886=>"110001110",
  48887=>"101010100",
  48888=>"100011101",
  48889=>"000000101",
  48890=>"010110100",
  48891=>"010001110",
  48892=>"111101111",
  48893=>"000001011",
  48894=>"111100011",
  48895=>"111101000",
  48896=>"101110111",
  48897=>"011000101",
  48898=>"001010111",
  48899=>"001001100",
  48900=>"001111001",
  48901=>"011001101",
  48902=>"110011011",
  48903=>"011011011",
  48904=>"111101011",
  48905=>"111001010",
  48906=>"010111101",
  48907=>"010111100",
  48908=>"000100111",
  48909=>"101010000",
  48910=>"110110001",
  48911=>"010000001",
  48912=>"110101000",
  48913=>"001000101",
  48914=>"100100110",
  48915=>"010011110",
  48916=>"001110001",
  48917=>"100100110",
  48918=>"110000000",
  48919=>"011111111",
  48920=>"111010100",
  48921=>"000000100",
  48922=>"100111101",
  48923=>"110010001",
  48924=>"000101101",
  48925=>"000011010",
  48926=>"001001000",
  48927=>"111001000",
  48928=>"000000100",
  48929=>"011110111",
  48930=>"101011100",
  48931=>"000000110",
  48932=>"100100111",
  48933=>"001100010",
  48934=>"000011011",
  48935=>"011001100",
  48936=>"010010001",
  48937=>"010010111",
  48938=>"001001001",
  48939=>"100110010",
  48940=>"111010010",
  48941=>"110100001",
  48942=>"010010000",
  48943=>"011011000",
  48944=>"000101110",
  48945=>"011110111",
  48946=>"100001110",
  48947=>"101110101",
  48948=>"000101000",
  48949=>"100100101",
  48950=>"001011100",
  48951=>"011001100",
  48952=>"111010100",
  48953=>"000101100",
  48954=>"000100011",
  48955=>"010010111",
  48956=>"010010111",
  48957=>"001000100",
  48958=>"110011110",
  48959=>"110110101",
  48960=>"110001001",
  48961=>"010011100",
  48962=>"100010010",
  48963=>"000000100",
  48964=>"001011000",
  48965=>"111000000",
  48966=>"101110010",
  48967=>"000000111",
  48968=>"111111110",
  48969=>"001011111",
  48970=>"111011111",
  48971=>"100010001",
  48972=>"011011011",
  48973=>"010111011",
  48974=>"000100011",
  48975=>"000000111",
  48976=>"100100101",
  48977=>"001010010",
  48978=>"110110000",
  48979=>"111001010",
  48980=>"111100001",
  48981=>"100010110",
  48982=>"100000011",
  48983=>"000100110",
  48984=>"001101011",
  48985=>"101111011",
  48986=>"010111001",
  48987=>"101100101",
  48988=>"110100000",
  48989=>"001001101",
  48990=>"010010100",
  48991=>"001000000",
  48992=>"111110111",
  48993=>"100010101",
  48994=>"010111000",
  48995=>"110010011",
  48996=>"111011100",
  48997=>"100100010",
  48998=>"101111000",
  48999=>"000010001",
  49000=>"110010100",
  49001=>"010000100",
  49002=>"000111101",
  49003=>"111111110",
  49004=>"111011001",
  49005=>"000011101",
  49006=>"000001010",
  49007=>"110001001",
  49008=>"100110111",
  49009=>"001001000",
  49010=>"001000000",
  49011=>"001000001",
  49012=>"001010000",
  49013=>"000001110",
  49014=>"000011000",
  49015=>"011000101",
  49016=>"010110011",
  49017=>"010011100",
  49018=>"111111111",
  49019=>"110111111",
  49020=>"010100001",
  49021=>"011100001",
  49022=>"100010010",
  49023=>"001101011",
  49024=>"001000111",
  49025=>"000110010",
  49026=>"001001111",
  49027=>"001000000",
  49028=>"000001100",
  49029=>"000010011",
  49030=>"011011010",
  49031=>"000101010",
  49032=>"110001111",
  49033=>"010001111",
  49034=>"101100010",
  49035=>"001000110",
  49036=>"110011110",
  49037=>"010000010",
  49038=>"100100111",
  49039=>"100101100",
  49040=>"000110110",
  49041=>"100100000",
  49042=>"011010000",
  49043=>"010100001",
  49044=>"001011000",
  49045=>"010100111",
  49046=>"011111111",
  49047=>"010100011",
  49048=>"001010101",
  49049=>"101000000",
  49050=>"101001010",
  49051=>"101111101",
  49052=>"110100111",
  49053=>"100000110",
  49054=>"100001000",
  49055=>"011011111",
  49056=>"001101001",
  49057=>"001011100",
  49058=>"000110111",
  49059=>"001001110",
  49060=>"100111000",
  49061=>"111000100",
  49062=>"110101000",
  49063=>"001000111",
  49064=>"001010111",
  49065=>"001000101",
  49066=>"101011110",
  49067=>"111000001",
  49068=>"101110011",
  49069=>"101001100",
  49070=>"110110100",
  49071=>"010011100",
  49072=>"010110010",
  49073=>"111011110",
  49074=>"101110010",
  49075=>"011011000",
  49076=>"100000101",
  49077=>"001110000",
  49078=>"111011000",
  49079=>"111011010",
  49080=>"111101011",
  49081=>"001010000",
  49082=>"110011111",
  49083=>"100110011",
  49084=>"100010000",
  49085=>"010011110",
  49086=>"110000000",
  49087=>"111000010",
  49088=>"010100111",
  49089=>"111001001",
  49090=>"010101010",
  49091=>"111101010",
  49092=>"010011110",
  49093=>"010010011",
  49094=>"010001001",
  49095=>"100010011",
  49096=>"000001111",
  49097=>"000100100",
  49098=>"111111010",
  49099=>"001110011",
  49100=>"110100111",
  49101=>"011000001",
  49102=>"101011100",
  49103=>"100000110",
  49104=>"010111100",
  49105=>"000000110",
  49106=>"110011000",
  49107=>"101101101",
  49108=>"101010001",
  49109=>"001010011",
  49110=>"000110001",
  49111=>"110011110",
  49112=>"000000100",
  49113=>"011011000",
  49114=>"000100000",
  49115=>"001101010",
  49116=>"110110010",
  49117=>"010101001",
  49118=>"100110000",
  49119=>"111100000",
  49120=>"001011101",
  49121=>"011001010",
  49122=>"101111110",
  49123=>"010010100",
  49124=>"010101000",
  49125=>"010111110",
  49126=>"010111011",
  49127=>"010110110",
  49128=>"001011001",
  49129=>"011010010",
  49130=>"001101101",
  49131=>"110001001",
  49132=>"010100100",
  49133=>"100100101",
  49134=>"000110000",
  49135=>"101111101",
  49136=>"110010011",
  49137=>"001011111",
  49138=>"110011110",
  49139=>"100010000",
  49140=>"101010001",
  49141=>"010111111",
  49142=>"010000100",
  49143=>"010011101",
  49144=>"111101000",
  49145=>"111000100",
  49146=>"001101010",
  49147=>"111100010",
  49148=>"101111101",
  49149=>"100001011",
  49150=>"100001111",
  49151=>"111011110",
  49152=>"000000011",
  49153=>"111111000",
  49154=>"111011011",
  49155=>"111111010",
  49156=>"100101001",
  49157=>"001011101",
  49158=>"100011111",
  49159=>"100000010",
  49160=>"010100100",
  49161=>"100011000",
  49162=>"000111111",
  49163=>"010110010",
  49164=>"000101001",
  49165=>"110010111",
  49166=>"000010000",
  49167=>"110001111",
  49168=>"100011011",
  49169=>"000010001",
  49170=>"100000000",
  49171=>"110100100",
  49172=>"110101100",
  49173=>"011010111",
  49174=>"101100000",
  49175=>"001010100",
  49176=>"001110011",
  49177=>"010101000",
  49178=>"010000110",
  49179=>"011110111",
  49180=>"011101011",
  49181=>"100101101",
  49182=>"001000100",
  49183=>"111110011",
  49184=>"111110111",
  49185=>"100100011",
  49186=>"001001010",
  49187=>"101010001",
  49188=>"000110101",
  49189=>"100001010",
  49190=>"111100111",
  49191=>"000000101",
  49192=>"011110000",
  49193=>"000001010",
  49194=>"010000001",
  49195=>"011000100",
  49196=>"000011101",
  49197=>"111111001",
  49198=>"110000100",
  49199=>"100011101",
  49200=>"010101101",
  49201=>"000111111",
  49202=>"100100001",
  49203=>"111111011",
  49204=>"001011001",
  49205=>"100101110",
  49206=>"011010011",
  49207=>"110011100",
  49208=>"101101001",
  49209=>"101001110",
  49210=>"011001101",
  49211=>"000101110",
  49212=>"000010001",
  49213=>"110010001",
  49214=>"101010100",
  49215=>"110100100",
  49216=>"101000010",
  49217=>"111001000",
  49218=>"001011001",
  49219=>"111010101",
  49220=>"101001111",
  49221=>"000011110",
  49222=>"001000100",
  49223=>"010111110",
  49224=>"011100000",
  49225=>"101010110",
  49226=>"110010001",
  49227=>"110011111",
  49228=>"000001100",
  49229=>"010011111",
  49230=>"100001001",
  49231=>"000101000",
  49232=>"101101010",
  49233=>"000110010",
  49234=>"100100101",
  49235=>"001010110",
  49236=>"000000101",
  49237=>"101001011",
  49238=>"111100100",
  49239=>"001010001",
  49240=>"111001100",
  49241=>"111111101",
  49242=>"111100101",
  49243=>"110000111",
  49244=>"111101111",
  49245=>"000110111",
  49246=>"000000101",
  49247=>"100011011",
  49248=>"010111100",
  49249=>"001000100",
  49250=>"101010100",
  49251=>"001000100",
  49252=>"011101111",
  49253=>"111010001",
  49254=>"001010011",
  49255=>"100001111",
  49256=>"100010000",
  49257=>"001010011",
  49258=>"011011111",
  49259=>"010010110",
  49260=>"000001000",
  49261=>"111111001",
  49262=>"010000011",
  49263=>"111111100",
  49264=>"011100010",
  49265=>"010110100",
  49266=>"000101110",
  49267=>"010101010",
  49268=>"101110001",
  49269=>"100000001",
  49270=>"101111011",
  49271=>"011000101",
  49272=>"010011011",
  49273=>"010010010",
  49274=>"000010011",
  49275=>"110110111",
  49276=>"111001010",
  49277=>"011000011",
  49278=>"100010101",
  49279=>"101100011",
  49280=>"001000001",
  49281=>"110010100",
  49282=>"010010101",
  49283=>"001100101",
  49284=>"110110001",
  49285=>"000101011",
  49286=>"000000000",
  49287=>"011011110",
  49288=>"110100110",
  49289=>"110000111",
  49290=>"001111011",
  49291=>"000001110",
  49292=>"110110111",
  49293=>"111011001",
  49294=>"011111001",
  49295=>"011011000",
  49296=>"011010000",
  49297=>"101100100",
  49298=>"000000101",
  49299=>"010000001",
  49300=>"011110010",
  49301=>"101111010",
  49302=>"011100101",
  49303=>"000101111",
  49304=>"010101111",
  49305=>"000100000",
  49306=>"100100110",
  49307=>"001010110",
  49308=>"001111001",
  49309=>"001001101",
  49310=>"111100101",
  49311=>"110001010",
  49312=>"100001011",
  49313=>"000110110",
  49314=>"101101011",
  49315=>"111001111",
  49316=>"111111011",
  49317=>"010101111",
  49318=>"001010001",
  49319=>"101110000",
  49320=>"001100011",
  49321=>"011001001",
  49322=>"101100111",
  49323=>"000010010",
  49324=>"111101011",
  49325=>"001110110",
  49326=>"111010101",
  49327=>"100001111",
  49328=>"110010011",
  49329=>"001001010",
  49330=>"011001000",
  49331=>"011101000",
  49332=>"001000010",
  49333=>"011100001",
  49334=>"001010000",
  49335=>"101100100",
  49336=>"010000010",
  49337=>"101101010",
  49338=>"011100100",
  49339=>"101001111",
  49340=>"111111100",
  49341=>"001111010",
  49342=>"000001101",
  49343=>"000010001",
  49344=>"001100110",
  49345=>"010000101",
  49346=>"000010001",
  49347=>"110100011",
  49348=>"100010000",
  49349=>"111000100",
  49350=>"111101011",
  49351=>"001010001",
  49352=>"111001001",
  49353=>"011010100",
  49354=>"110100010",
  49355=>"010111110",
  49356=>"010000111",
  49357=>"010101110",
  49358=>"011011010",
  49359=>"000011110",
  49360=>"011111111",
  49361=>"000010011",
  49362=>"100001010",
  49363=>"101000100",
  49364=>"010010011",
  49365=>"010011111",
  49366=>"110111111",
  49367=>"111000101",
  49368=>"011000100",
  49369=>"001011110",
  49370=>"110000000",
  49371=>"011000010",
  49372=>"101110101",
  49373=>"101000001",
  49374=>"110111000",
  49375=>"101111111",
  49376=>"111100000",
  49377=>"100110110",
  49378=>"000011011",
  49379=>"101101110",
  49380=>"100111101",
  49381=>"000101111",
  49382=>"111010000",
  49383=>"001001111",
  49384=>"110100011",
  49385=>"010000110",
  49386=>"111101111",
  49387=>"001001101",
  49388=>"100110011",
  49389=>"010100100",
  49390=>"110001010",
  49391=>"100001111",
  49392=>"101010101",
  49393=>"011101010",
  49394=>"110000010",
  49395=>"010011100",
  49396=>"010000100",
  49397=>"101101000",
  49398=>"101011110",
  49399=>"110011000",
  49400=>"010111001",
  49401=>"000011010",
  49402=>"100101001",
  49403=>"011001001",
  49404=>"111110011",
  49405=>"101110011",
  49406=>"110101110",
  49407=>"010110111",
  49408=>"101101011",
  49409=>"111011011",
  49410=>"000011110",
  49411=>"111100010",
  49412=>"001101001",
  49413=>"010111000",
  49414=>"111111010",
  49415=>"001100101",
  49416=>"111011110",
  49417=>"111101000",
  49418=>"010111001",
  49419=>"001000000",
  49420=>"101011010",
  49421=>"111001010",
  49422=>"110010100",
  49423=>"000101110",
  49424=>"110100111",
  49425=>"111110010",
  49426=>"011100110",
  49427=>"001100001",
  49428=>"010100001",
  49429=>"111010110",
  49430=>"001010110",
  49431=>"001001100",
  49432=>"110111111",
  49433=>"010111101",
  49434=>"001001110",
  49435=>"100111111",
  49436=>"101000000",
  49437=>"000010111",
  49438=>"110110100",
  49439=>"100011100",
  49440=>"001101001",
  49441=>"001011010",
  49442=>"100101011",
  49443=>"011100001",
  49444=>"001111111",
  49445=>"000011110",
  49446=>"001110100",
  49447=>"111111001",
  49448=>"011101001",
  49449=>"101001100",
  49450=>"111000101",
  49451=>"000000110",
  49452=>"101101000",
  49453=>"010000001",
  49454=>"001110010",
  49455=>"110000010",
  49456=>"100000101",
  49457=>"010011110",
  49458=>"100011001",
  49459=>"101101010",
  49460=>"000000100",
  49461=>"000100100",
  49462=>"000010100",
  49463=>"110100001",
  49464=>"111111101",
  49465=>"110111001",
  49466=>"111001000",
  49467=>"101111101",
  49468=>"011101101",
  49469=>"001101100",
  49470=>"010001101",
  49471=>"101101101",
  49472=>"011000000",
  49473=>"101100000",
  49474=>"010110111",
  49475=>"010100111",
  49476=>"010110001",
  49477=>"010111111",
  49478=>"001001100",
  49479=>"011011001",
  49480=>"111011110",
  49481=>"111110111",
  49482=>"001110110",
  49483=>"101111100",
  49484=>"000000011",
  49485=>"100011110",
  49486=>"100011101",
  49487=>"100111011",
  49488=>"001010100",
  49489=>"001110001",
  49490=>"011101000",
  49491=>"101001101",
  49492=>"101000101",
  49493=>"100100000",
  49494=>"100110101",
  49495=>"100100101",
  49496=>"111010111",
  49497=>"010011111",
  49498=>"101100010",
  49499=>"000000011",
  49500=>"000000110",
  49501=>"001100010",
  49502=>"100101011",
  49503=>"010001110",
  49504=>"101011101",
  49505=>"001101000",
  49506=>"100100011",
  49507=>"100100000",
  49508=>"001000010",
  49509=>"110010100",
  49510=>"111011000",
  49511=>"111110011",
  49512=>"000000101",
  49513=>"000011010",
  49514=>"011010000",
  49515=>"110010110",
  49516=>"001001110",
  49517=>"010100001",
  49518=>"101100100",
  49519=>"111100110",
  49520=>"001111110",
  49521=>"000111010",
  49522=>"111100101",
  49523=>"110100111",
  49524=>"111111001",
  49525=>"111110011",
  49526=>"101001001",
  49527=>"011011011",
  49528=>"010101101",
  49529=>"111111010",
  49530=>"111100111",
  49531=>"010111110",
  49532=>"110110011",
  49533=>"010010010",
  49534=>"000010110",
  49535=>"000101010",
  49536=>"100000101",
  49537=>"001110011",
  49538=>"000101110",
  49539=>"100010000",
  49540=>"000001110",
  49541=>"110101101",
  49542=>"011011101",
  49543=>"100110010",
  49544=>"100000001",
  49545=>"001000110",
  49546=>"100111110",
  49547=>"011010101",
  49548=>"100010101",
  49549=>"111010100",
  49550=>"000101010",
  49551=>"011110000",
  49552=>"000100001",
  49553=>"000000000",
  49554=>"011100001",
  49555=>"001101100",
  49556=>"010000010",
  49557=>"111111001",
  49558=>"000001110",
  49559=>"110101000",
  49560=>"101100011",
  49561=>"000111011",
  49562=>"011111101",
  49563=>"101100100",
  49564=>"100111000",
  49565=>"100101010",
  49566=>"000101011",
  49567=>"001011100",
  49568=>"001101101",
  49569=>"111111000",
  49570=>"011010111",
  49571=>"010010001",
  49572=>"111110111",
  49573=>"010000001",
  49574=>"101001010",
  49575=>"100000011",
  49576=>"100110001",
  49577=>"101011100",
  49578=>"010000110",
  49579=>"111101110",
  49580=>"000110010",
  49581=>"010011001",
  49582=>"111110100",
  49583=>"000000000",
  49584=>"111011001",
  49585=>"101110100",
  49586=>"100010011",
  49587=>"001010010",
  49588=>"100101010",
  49589=>"111110011",
  49590=>"001101110",
  49591=>"110111000",
  49592=>"111000001",
  49593=>"111010001",
  49594=>"101010110",
  49595=>"001110011",
  49596=>"000001010",
  49597=>"011011101",
  49598=>"111101010",
  49599=>"111101110",
  49600=>"001101100",
  49601=>"101110001",
  49602=>"010100110",
  49603=>"001111111",
  49604=>"000000100",
  49605=>"000101110",
  49606=>"001000010",
  49607=>"001111111",
  49608=>"111110100",
  49609=>"000001011",
  49610=>"101101000",
  49611=>"010011000",
  49612=>"000010101",
  49613=>"011101010",
  49614=>"010100010",
  49615=>"111101111",
  49616=>"001110111",
  49617=>"010100000",
  49618=>"001001011",
  49619=>"100101100",
  49620=>"110000011",
  49621=>"010101110",
  49622=>"010010101",
  49623=>"010011000",
  49624=>"011001100",
  49625=>"101100111",
  49626=>"110010010",
  49627=>"111000011",
  49628=>"001001101",
  49629=>"000011111",
  49630=>"100101011",
  49631=>"010111110",
  49632=>"110001100",
  49633=>"010000001",
  49634=>"100010101",
  49635=>"001101011",
  49636=>"100100000",
  49637=>"000101010",
  49638=>"111011010",
  49639=>"010000100",
  49640=>"100010110",
  49641=>"010100010",
  49642=>"001010111",
  49643=>"101111101",
  49644=>"110110101",
  49645=>"010101000",
  49646=>"100011001",
  49647=>"111100000",
  49648=>"101001101",
  49649=>"011100110",
  49650=>"101001110",
  49651=>"010000101",
  49652=>"010101101",
  49653=>"000011010",
  49654=>"011011111",
  49655=>"010000001",
  49656=>"100001011",
  49657=>"010011000",
  49658=>"110101000",
  49659=>"010100110",
  49660=>"001101111",
  49661=>"011101101",
  49662=>"101111111",
  49663=>"101010101",
  49664=>"011000111",
  49665=>"010100110",
  49666=>"111010011",
  49667=>"011101100",
  49668=>"011111011",
  49669=>"001110001",
  49670=>"101010000",
  49671=>"011010010",
  49672=>"100111001",
  49673=>"111110100",
  49674=>"100010100",
  49675=>"000000101",
  49676=>"010010011",
  49677=>"110101001",
  49678=>"000100111",
  49679=>"010101011",
  49680=>"111101110",
  49681=>"010100011",
  49682=>"011011011",
  49683=>"011110111",
  49684=>"011000001",
  49685=>"000010110",
  49686=>"110010010",
  49687=>"010100111",
  49688=>"110000001",
  49689=>"010110101",
  49690=>"000011110",
  49691=>"100000110",
  49692=>"011001110",
  49693=>"001110000",
  49694=>"011010000",
  49695=>"010101001",
  49696=>"110001011",
  49697=>"011110100",
  49698=>"110010111",
  49699=>"000100000",
  49700=>"010111001",
  49701=>"110101011",
  49702=>"010100110",
  49703=>"001000111",
  49704=>"100000101",
  49705=>"000110000",
  49706=>"000100010",
  49707=>"010001110",
  49708=>"100001101",
  49709=>"101100101",
  49710=>"000010100",
  49711=>"010000010",
  49712=>"001101110",
  49713=>"110011100",
  49714=>"110010101",
  49715=>"000011101",
  49716=>"011101111",
  49717=>"101101000",
  49718=>"010101011",
  49719=>"101011001",
  49720=>"101011101",
  49721=>"010110001",
  49722=>"010100011",
  49723=>"111110011",
  49724=>"110001101",
  49725=>"000101010",
  49726=>"001111101",
  49727=>"000100010",
  49728=>"010111111",
  49729=>"010001101",
  49730=>"001000000",
  49731=>"000101011",
  49732=>"001011011",
  49733=>"101011011",
  49734=>"011100000",
  49735=>"000111001",
  49736=>"000100001",
  49737=>"000010011",
  49738=>"001100111",
  49739=>"110010011",
  49740=>"111100110",
  49741=>"000010000",
  49742=>"000011010",
  49743=>"101011100",
  49744=>"011010000",
  49745=>"101010111",
  49746=>"001101101",
  49747=>"000001011",
  49748=>"100100110",
  49749=>"100010100",
  49750=>"111101010",
  49751=>"001010011",
  49752=>"100111100",
  49753=>"001000011",
  49754=>"101110111",
  49755=>"011101001",
  49756=>"001011001",
  49757=>"101100001",
  49758=>"011010111",
  49759=>"000110100",
  49760=>"010011001",
  49761=>"111001111",
  49762=>"101111110",
  49763=>"001011111",
  49764=>"001100001",
  49765=>"000101100",
  49766=>"001100001",
  49767=>"001111011",
  49768=>"100000100",
  49769=>"011000110",
  49770=>"001110001",
  49771=>"010101000",
  49772=>"101010010",
  49773=>"010111101",
  49774=>"101111010",
  49775=>"110110111",
  49776=>"111000111",
  49777=>"110001110",
  49778=>"111111110",
  49779=>"101011100",
  49780=>"000011010",
  49781=>"011001010",
  49782=>"101100101",
  49783=>"000110100",
  49784=>"110110101",
  49785=>"100111101",
  49786=>"101110001",
  49787=>"001010110",
  49788=>"101011111",
  49789=>"000010000",
  49790=>"000111001",
  49791=>"100111001",
  49792=>"010101000",
  49793=>"111111000",
  49794=>"110101000",
  49795=>"011110010",
  49796=>"110111010",
  49797=>"101010111",
  49798=>"011101000",
  49799=>"000001001",
  49800=>"000110010",
  49801=>"010110100",
  49802=>"010001000",
  49803=>"010100000",
  49804=>"000111100",
  49805=>"101001011",
  49806=>"100111011",
  49807=>"110111010",
  49808=>"001001000",
  49809=>"000100100",
  49810=>"101110110",
  49811=>"110111101",
  49812=>"010111111",
  49813=>"010111100",
  49814=>"111000000",
  49815=>"111000010",
  49816=>"011010001",
  49817=>"101101101",
  49818=>"000001101",
  49819=>"010001101",
  49820=>"011110101",
  49821=>"111000000",
  49822=>"001101010",
  49823=>"000011110",
  49824=>"101111111",
  49825=>"011010011",
  49826=>"001011000",
  49827=>"001100000",
  49828=>"100100011",
  49829=>"111100100",
  49830=>"010100101",
  49831=>"111000000",
  49832=>"000010010",
  49833=>"011010101",
  49834=>"001010010",
  49835=>"100110011",
  49836=>"010001011",
  49837=>"010110000",
  49838=>"111110110",
  49839=>"000100011",
  49840=>"101100100",
  49841=>"010001010",
  49842=>"011111011",
  49843=>"111000101",
  49844=>"001000010",
  49845=>"110010110",
  49846=>"011101111",
  49847=>"110110010",
  49848=>"001110000",
  49849=>"010001010",
  49850=>"011111110",
  49851=>"110100101",
  49852=>"000011111",
  49853=>"101100111",
  49854=>"000010011",
  49855=>"111010001",
  49856=>"001010110",
  49857=>"001110110",
  49858=>"100111100",
  49859=>"110110110",
  49860=>"111110100",
  49861=>"010010010",
  49862=>"101001111",
  49863=>"100111111",
  49864=>"110110100",
  49865=>"001100101",
  49866=>"111011111",
  49867=>"111000011",
  49868=>"001110001",
  49869=>"100000111",
  49870=>"100010110",
  49871=>"100111111",
  49872=>"100101101",
  49873=>"101111011",
  49874=>"000101111",
  49875=>"110000000",
  49876=>"111110010",
  49877=>"110011001",
  49878=>"001010011",
  49879=>"101001110",
  49880=>"010000011",
  49881=>"100010110",
  49882=>"110110010",
  49883=>"010111011",
  49884=>"000001011",
  49885=>"000110101",
  49886=>"010001111",
  49887=>"010000100",
  49888=>"010111100",
  49889=>"101111101",
  49890=>"111000100",
  49891=>"011001000",
  49892=>"101000011",
  49893=>"101100010",
  49894=>"111010111",
  49895=>"100110000",
  49896=>"001000111",
  49897=>"001111010",
  49898=>"100100110",
  49899=>"001011010",
  49900=>"010000011",
  49901=>"100111011",
  49902=>"101001111",
  49903=>"111100111",
  49904=>"110100100",
  49905=>"101100001",
  49906=>"111010101",
  49907=>"100001110",
  49908=>"111011101",
  49909=>"110101100",
  49910=>"100000000",
  49911=>"100101000",
  49912=>"000000000",
  49913=>"101001011",
  49914=>"110001011",
  49915=>"101010110",
  49916=>"111110011",
  49917=>"000000000",
  49918=>"110110110",
  49919=>"100100100",
  49920=>"010110001",
  49921=>"001101100",
  49922=>"011000001",
  49923=>"111000010",
  49924=>"101011000",
  49925=>"101110100",
  49926=>"111001001",
  49927=>"100001000",
  49928=>"111000110",
  49929=>"110011110",
  49930=>"000101001",
  49931=>"110001011",
  49932=>"110100000",
  49933=>"000000101",
  49934=>"110111100",
  49935=>"000011110",
  49936=>"111001110",
  49937=>"000110001",
  49938=>"101010010",
  49939=>"101001100",
  49940=>"100101100",
  49941=>"101011011",
  49942=>"100101101",
  49943=>"100110011",
  49944=>"001011101",
  49945=>"011100000",
  49946=>"110101100",
  49947=>"001101001",
  49948=>"001011010",
  49949=>"010110111",
  49950=>"001111001",
  49951=>"011100111",
  49952=>"101111000",
  49953=>"001111100",
  49954=>"011010101",
  49955=>"000010111",
  49956=>"010000101",
  49957=>"111100101",
  49958=>"100001101",
  49959=>"001001011",
  49960=>"000110010",
  49961=>"100101000",
  49962=>"011001101",
  49963=>"010111011",
  49964=>"100011111",
  49965=>"010000000",
  49966=>"010101011",
  49967=>"110110111",
  49968=>"000010100",
  49969=>"100010111",
  49970=>"110000011",
  49971=>"010101110",
  49972=>"011111001",
  49973=>"111000010",
  49974=>"000001000",
  49975=>"000001000",
  49976=>"000000101",
  49977=>"110000001",
  49978=>"011101110",
  49979=>"010101101",
  49980=>"011110010",
  49981=>"101011001",
  49982=>"001111000",
  49983=>"101101000",
  49984=>"100011111",
  49985=>"011000111",
  49986=>"011111000",
  49987=>"010101111",
  49988=>"001101110",
  49989=>"101011010",
  49990=>"001100110",
  49991=>"100010011",
  49992=>"100101111",
  49993=>"101011110",
  49994=>"001110110",
  49995=>"001110011",
  49996=>"110101000",
  49997=>"110101101",
  49998=>"001101001",
  49999=>"000000010",
  50000=>"110000101",
  50001=>"101000110",
  50002=>"101011011",
  50003=>"100000101",
  50004=>"000101110",
  50005=>"111110001",
  50006=>"111100010",
  50007=>"001000000",
  50008=>"110111100",
  50009=>"001000101",
  50010=>"101001111",
  50011=>"111011010",
  50012=>"111110111",
  50013=>"010001110",
  50014=>"001011100",
  50015=>"110001100",
  50016=>"110100011",
  50017=>"000111010",
  50018=>"010011110",
  50019=>"000100011",
  50020=>"010101000",
  50021=>"011110101",
  50022=>"110101001",
  50023=>"101110111",
  50024=>"111010110",
  50025=>"101111111",
  50026=>"001000111",
  50027=>"110001001",
  50028=>"000111011",
  50029=>"111011001",
  50030=>"011011100",
  50031=>"000011101",
  50032=>"000001111",
  50033=>"111001100",
  50034=>"010010001",
  50035=>"100001010",
  50036=>"011100000",
  50037=>"111010010",
  50038=>"110110111",
  50039=>"000100010",
  50040=>"100000111",
  50041=>"111101000",
  50042=>"001011010",
  50043=>"100000001",
  50044=>"101001111",
  50045=>"000011000",
  50046=>"011101011",
  50047=>"111000010",
  50048=>"100110101",
  50049=>"111010000",
  50050=>"111000001",
  50051=>"000001101",
  50052=>"110000000",
  50053=>"010000010",
  50054=>"001010101",
  50055=>"111101010",
  50056=>"111000011",
  50057=>"111001011",
  50058=>"111111111",
  50059=>"110101100",
  50060=>"100101100",
  50061=>"101011101",
  50062=>"111001011",
  50063=>"001010010",
  50064=>"100111001",
  50065=>"010011101",
  50066=>"001111101",
  50067=>"011101011",
  50068=>"101101101",
  50069=>"011001011",
  50070=>"001110100",
  50071=>"100110000",
  50072=>"011101011",
  50073=>"011111011",
  50074=>"000110000",
  50075=>"010000011",
  50076=>"100001011",
  50077=>"110101101",
  50078=>"101111001",
  50079=>"101001101",
  50080=>"000010001",
  50081=>"000111110",
  50082=>"100110001",
  50083=>"011101111",
  50084=>"100110010",
  50085=>"110000111",
  50086=>"101000111",
  50087=>"100001100",
  50088=>"001001001",
  50089=>"110001101",
  50090=>"001010100",
  50091=>"001101101",
  50092=>"001011101",
  50093=>"000110001",
  50094=>"010101101",
  50095=>"010000000",
  50096=>"111011100",
  50097=>"101100001",
  50098=>"111001110",
  50099=>"000100011",
  50100=>"001111110",
  50101=>"110000001",
  50102=>"000000100",
  50103=>"110111010",
  50104=>"001111000",
  50105=>"010000001",
  50106=>"111000010",
  50107=>"110110100",
  50108=>"001011111",
  50109=>"101001011",
  50110=>"111111101",
  50111=>"110101100",
  50112=>"011000100",
  50113=>"111010111",
  50114=>"000010010",
  50115=>"111110111",
  50116=>"110011010",
  50117=>"011110110",
  50118=>"111100000",
  50119=>"010010001",
  50120=>"000001010",
  50121=>"111111111",
  50122=>"110001011",
  50123=>"111011101",
  50124=>"011101010",
  50125=>"001000010",
  50126=>"111010011",
  50127=>"100111100",
  50128=>"010110111",
  50129=>"000000001",
  50130=>"001010111",
  50131=>"000001010",
  50132=>"010000001",
  50133=>"001000010",
  50134=>"111000110",
  50135=>"000001100",
  50136=>"010110100",
  50137=>"010001101",
  50138=>"001011100",
  50139=>"111111010",
  50140=>"111110110",
  50141=>"011011001",
  50142=>"101100100",
  50143=>"010111011",
  50144=>"010000000",
  50145=>"011101000",
  50146=>"110001010",
  50147=>"110001111",
  50148=>"111110000",
  50149=>"010010001",
  50150=>"100000010",
  50151=>"110101001",
  50152=>"100110101",
  50153=>"000101001",
  50154=>"011110100",
  50155=>"111010110",
  50156=>"100101111",
  50157=>"011100010",
  50158=>"111011100",
  50159=>"010101111",
  50160=>"100110010",
  50161=>"010110011",
  50162=>"001010101",
  50163=>"000111000",
  50164=>"101111010",
  50165=>"001101101",
  50166=>"110000100",
  50167=>"111101111",
  50168=>"001101001",
  50169=>"110001110",
  50170=>"000011111",
  50171=>"010010101",
  50172=>"011001000",
  50173=>"011000000",
  50174=>"010100110",
  50175=>"001011010",
  50176=>"100100010",
  50177=>"000110010",
  50178=>"001100111",
  50179=>"111101100",
  50180=>"001110101",
  50181=>"010100011",
  50182=>"110001110",
  50183=>"110111100",
  50184=>"001100010",
  50185=>"110100111",
  50186=>"100100001",
  50187=>"100000101",
  50188=>"001010110",
  50189=>"101000000",
  50190=>"110101111",
  50191=>"010010101",
  50192=>"110010100",
  50193=>"111000101",
  50194=>"000010011",
  50195=>"001101001",
  50196=>"011110011",
  50197=>"101110101",
  50198=>"100110111",
  50199=>"100000101",
  50200=>"010110101",
  50201=>"110010010",
  50202=>"111001111",
  50203=>"111011110",
  50204=>"000100101",
  50205=>"000110000",
  50206=>"001100111",
  50207=>"000001100",
  50208=>"111001111",
  50209=>"000000011",
  50210=>"010010101",
  50211=>"111001101",
  50212=>"101101001",
  50213=>"111010100",
  50214=>"100100011",
  50215=>"001111001",
  50216=>"110001101",
  50217=>"000010011",
  50218=>"000001101",
  50219=>"111101110",
  50220=>"111101101",
  50221=>"110111101",
  50222=>"110011100",
  50223=>"100000110",
  50224=>"010101011",
  50225=>"010001001",
  50226=>"101010000",
  50227=>"110111101",
  50228=>"101110100",
  50229=>"000000000",
  50230=>"110101110",
  50231=>"111101001",
  50232=>"010100111",
  50233=>"010010100",
  50234=>"011100011",
  50235=>"000101101",
  50236=>"100100101",
  50237=>"111100111",
  50238=>"000011000",
  50239=>"010110101",
  50240=>"011000011",
  50241=>"000010101",
  50242=>"100110001",
  50243=>"000000001",
  50244=>"100011001",
  50245=>"111000000",
  50246=>"111101100",
  50247=>"100100000",
  50248=>"000110101",
  50249=>"010000101",
  50250=>"011010101",
  50251=>"010110101",
  50252=>"000001000",
  50253=>"101000011",
  50254=>"010010001",
  50255=>"100110111",
  50256=>"111010110",
  50257=>"111100111",
  50258=>"111111001",
  50259=>"000110111",
  50260=>"110000110",
  50261=>"001001111",
  50262=>"101111011",
  50263=>"001000010",
  50264=>"100110000",
  50265=>"010111001",
  50266=>"100011010",
  50267=>"001100110",
  50268=>"100001101",
  50269=>"011000111",
  50270=>"001010100",
  50271=>"010010000",
  50272=>"111100110",
  50273=>"001110111",
  50274=>"111010000",
  50275=>"010011011",
  50276=>"011011010",
  50277=>"010101001",
  50278=>"111110100",
  50279=>"010001011",
  50280=>"010010000",
  50281=>"011100011",
  50282=>"100100110",
  50283=>"111010100",
  50284=>"111010010",
  50285=>"000011111",
  50286=>"010100011",
  50287=>"100001011",
  50288=>"101000010",
  50289=>"111110100",
  50290=>"111101100",
  50291=>"110000000",
  50292=>"111110100",
  50293=>"100111111",
  50294=>"011100101",
  50295=>"010111010",
  50296=>"100101111",
  50297=>"100111100",
  50298=>"001100100",
  50299=>"111000100",
  50300=>"010010001",
  50301=>"010011101",
  50302=>"000001000",
  50303=>"000110111",
  50304=>"100111101",
  50305=>"000000110",
  50306=>"011000110",
  50307=>"000000000",
  50308=>"001011110",
  50309=>"011001000",
  50310=>"101110101",
  50311=>"011101000",
  50312=>"111100010",
  50313=>"000011000",
  50314=>"101010000",
  50315=>"001100001",
  50316=>"111111000",
  50317=>"100001110",
  50318=>"101010111",
  50319=>"011110101",
  50320=>"001100000",
  50321=>"101011101",
  50322=>"101001111",
  50323=>"010100111",
  50324=>"111101111",
  50325=>"101001010",
  50326=>"111010011",
  50327=>"100000010",
  50328=>"110100001",
  50329=>"111110110",
  50330=>"000101001",
  50331=>"111110101",
  50332=>"010010000",
  50333=>"011011010",
  50334=>"100011000",
  50335=>"001010001",
  50336=>"101011101",
  50337=>"111001010",
  50338=>"111001101",
  50339=>"111100100",
  50340=>"000011111",
  50341=>"000000100",
  50342=>"010011000",
  50343=>"000001000",
  50344=>"000000110",
  50345=>"101110010",
  50346=>"001001110",
  50347=>"111011011",
  50348=>"000110011",
  50349=>"101001100",
  50350=>"100111010",
  50351=>"101110000",
  50352=>"001101111",
  50353=>"010000100",
  50354=>"001000001",
  50355=>"001000011",
  50356=>"001000011",
  50357=>"111111100",
  50358=>"110101111",
  50359=>"111000101",
  50360=>"111111000",
  50361=>"001010110",
  50362=>"001001000",
  50363=>"001001111",
  50364=>"011110101",
  50365=>"010000100",
  50366=>"111001101",
  50367=>"001110110",
  50368=>"100110110",
  50369=>"111011101",
  50370=>"110010110",
  50371=>"000100010",
  50372=>"010110111",
  50373=>"000001111",
  50374=>"110111001",
  50375=>"100010101",
  50376=>"100011000",
  50377=>"000100000",
  50378=>"101100011",
  50379=>"101001010",
  50380=>"010000110",
  50381=>"110111110",
  50382=>"001010100",
  50383=>"110010110",
  50384=>"111001111",
  50385=>"000010010",
  50386=>"011011110",
  50387=>"100001001",
  50388=>"011110001",
  50389=>"101000011",
  50390=>"110011011",
  50391=>"011011010",
  50392=>"010001110",
  50393=>"111100001",
  50394=>"000010101",
  50395=>"111100101",
  50396=>"110111100",
  50397=>"000000001",
  50398=>"100111001",
  50399=>"111011000",
  50400=>"000001101",
  50401=>"110110111",
  50402=>"111111010",
  50403=>"111110110",
  50404=>"011011001",
  50405=>"100110101",
  50406=>"110101001",
  50407=>"111010000",
  50408=>"001100001",
  50409=>"111011001",
  50410=>"010111011",
  50411=>"000100101",
  50412=>"101110010",
  50413=>"110100111",
  50414=>"101011011",
  50415=>"101001000",
  50416=>"110100000",
  50417=>"100010110",
  50418=>"000010111",
  50419=>"101000010",
  50420=>"100110000",
  50421=>"001011011",
  50422=>"011111011",
  50423=>"001110001",
  50424=>"110111001",
  50425=>"110010101",
  50426=>"111101010",
  50427=>"010000101",
  50428=>"010101101",
  50429=>"100111001",
  50430=>"110100001",
  50431=>"110101101",
  50432=>"110010110",
  50433=>"011000100",
  50434=>"111101110",
  50435=>"110100010",
  50436=>"111110011",
  50437=>"110111110",
  50438=>"000001110",
  50439=>"010001101",
  50440=>"000100001",
  50441=>"010001001",
  50442=>"001101000",
  50443=>"100100101",
  50444=>"101001111",
  50445=>"100010010",
  50446=>"110011001",
  50447=>"111010000",
  50448=>"100111111",
  50449=>"100001101",
  50450=>"010111111",
  50451=>"101111110",
  50452=>"110001011",
  50453=>"000100000",
  50454=>"110010010",
  50455=>"111000000",
  50456=>"111000100",
  50457=>"000000011",
  50458=>"111110011",
  50459=>"001101101",
  50460=>"110010101",
  50461=>"001110000",
  50462=>"110000011",
  50463=>"100101001",
  50464=>"000100101",
  50465=>"000000000",
  50466=>"011100001",
  50467=>"101111001",
  50468=>"001000010",
  50469=>"001100101",
  50470=>"101100010",
  50471=>"001101001",
  50472=>"010101100",
  50473=>"110001001",
  50474=>"101111110",
  50475=>"011101001",
  50476=>"001010101",
  50477=>"011010000",
  50478=>"101100001",
  50479=>"110110100",
  50480=>"011101100",
  50481=>"011101010",
  50482=>"000001100",
  50483=>"001000000",
  50484=>"001101000",
  50485=>"010100100",
  50486=>"001101111",
  50487=>"001110101",
  50488=>"111000011",
  50489=>"101011010",
  50490=>"100100101",
  50491=>"100001001",
  50492=>"111111001",
  50493=>"100111000",
  50494=>"001110100",
  50495=>"100000111",
  50496=>"111001111",
  50497=>"110000000",
  50498=>"001110000",
  50499=>"010001010",
  50500=>"110110010",
  50501=>"110101110",
  50502=>"101000100",
  50503=>"100101100",
  50504=>"001111010",
  50505=>"100100101",
  50506=>"111000001",
  50507=>"011110011",
  50508=>"011001101",
  50509=>"110010011",
  50510=>"101001000",
  50511=>"011110111",
  50512=>"101000111",
  50513=>"110101111",
  50514=>"010111110",
  50515=>"000011001",
  50516=>"110010001",
  50517=>"000011011",
  50518=>"001110110",
  50519=>"010010100",
  50520=>"111000101",
  50521=>"011000011",
  50522=>"110101101",
  50523=>"011010001",
  50524=>"010001111",
  50525=>"011100000",
  50526=>"101100000",
  50527=>"000010010",
  50528=>"001001110",
  50529=>"111111111",
  50530=>"110000001",
  50531=>"001100000",
  50532=>"110010110",
  50533=>"001000101",
  50534=>"111101111",
  50535=>"110111111",
  50536=>"010001101",
  50537=>"001101101",
  50538=>"000010010",
  50539=>"101100010",
  50540=>"011110101",
  50541=>"001110001",
  50542=>"100111001",
  50543=>"110011111",
  50544=>"000100001",
  50545=>"101111000",
  50546=>"111010010",
  50547=>"111110110",
  50548=>"101001110",
  50549=>"101110011",
  50550=>"001001011",
  50551=>"110100100",
  50552=>"000100001",
  50553=>"001001010",
  50554=>"000101000",
  50555=>"111001100",
  50556=>"110101111",
  50557=>"011001101",
  50558=>"001111001",
  50559=>"111100100",
  50560=>"011011001",
  50561=>"011011000",
  50562=>"101100100",
  50563=>"000010111",
  50564=>"000010111",
  50565=>"000101001",
  50566=>"011111000",
  50567=>"000010001",
  50568=>"101010000",
  50569=>"011100110",
  50570=>"100101111",
  50571=>"001000010",
  50572=>"001111011",
  50573=>"111101000",
  50574=>"110101001",
  50575=>"101110111",
  50576=>"011111111",
  50577=>"001001101",
  50578=>"110000100",
  50579=>"011111110",
  50580=>"001110011",
  50581=>"011000010",
  50582=>"010010010",
  50583=>"100111010",
  50584=>"000111100",
  50585=>"101011111",
  50586=>"110000010",
  50587=>"101101101",
  50588=>"111100111",
  50589=>"000100100",
  50590=>"000110011",
  50591=>"100101001",
  50592=>"100011001",
  50593=>"000111001",
  50594=>"001000111",
  50595=>"001111000",
  50596=>"001010101",
  50597=>"100100011",
  50598=>"011101001",
  50599=>"000111010",
  50600=>"111000100",
  50601=>"011111010",
  50602=>"000000010",
  50603=>"101110000",
  50604=>"010111001",
  50605=>"011010000",
  50606=>"111001001",
  50607=>"110110010",
  50608=>"100101011",
  50609=>"001000100",
  50610=>"000101010",
  50611=>"101001011",
  50612=>"100011011",
  50613=>"101110110",
  50614=>"010100010",
  50615=>"110100011",
  50616=>"101010111",
  50617=>"000000001",
  50618=>"010110101",
  50619=>"011100010",
  50620=>"110110011",
  50621=>"100010011",
  50622=>"111110111",
  50623=>"100001010",
  50624=>"100101011",
  50625=>"001000010",
  50626=>"101010000",
  50627=>"010010111",
  50628=>"010011001",
  50629=>"000000000",
  50630=>"010000000",
  50631=>"010000110",
  50632=>"010101010",
  50633=>"110110001",
  50634=>"110010011",
  50635=>"101111011",
  50636=>"011010110",
  50637=>"000010110",
  50638=>"001100110",
  50639=>"011001110",
  50640=>"010100011",
  50641=>"001001000",
  50642=>"011011010",
  50643=>"111010100",
  50644=>"000110111",
  50645=>"111101111",
  50646=>"110110011",
  50647=>"110010011",
  50648=>"110011011",
  50649=>"111000011",
  50650=>"101010101",
  50651=>"111101001",
  50652=>"111110011",
  50653=>"000100010",
  50654=>"101000111",
  50655=>"111110011",
  50656=>"110000011",
  50657=>"101011101",
  50658=>"001101010",
  50659=>"110001001",
  50660=>"101010000",
  50661=>"001111110",
  50662=>"010101101",
  50663=>"111101011",
  50664=>"111010110",
  50665=>"101111000",
  50666=>"100100011",
  50667=>"100010111",
  50668=>"000000000",
  50669=>"001010000",
  50670=>"010010100",
  50671=>"100101000",
  50672=>"110001010",
  50673=>"010110101",
  50674=>"100100111",
  50675=>"001111000",
  50676=>"100110110",
  50677=>"111111101",
  50678=>"101111111",
  50679=>"000110010",
  50680=>"000000011",
  50681=>"100100010",
  50682=>"111001011",
  50683=>"100111011",
  50684=>"011110111",
  50685=>"010001000",
  50686=>"111101000",
  50687=>"111010110",
  50688=>"111011101",
  50689=>"110101100",
  50690=>"001111000",
  50691=>"100101011",
  50692=>"111110010",
  50693=>"001011111",
  50694=>"001110100",
  50695=>"011000100",
  50696=>"011110001",
  50697=>"101111000",
  50698=>"011000001",
  50699=>"000001001",
  50700=>"001001111",
  50701=>"001110101",
  50702=>"101100111",
  50703=>"101100100",
  50704=>"100000101",
  50705=>"111010101",
  50706=>"101001011",
  50707=>"010000101",
  50708=>"111111000",
  50709=>"110000111",
  50710=>"110011100",
  50711=>"100000011",
  50712=>"101010101",
  50713=>"000110100",
  50714=>"111101011",
  50715=>"011111101",
  50716=>"010010100",
  50717=>"100101100",
  50718=>"111001001",
  50719=>"000111111",
  50720=>"011010111",
  50721=>"111100101",
  50722=>"010000001",
  50723=>"001100111",
  50724=>"100011000",
  50725=>"000110100",
  50726=>"011011110",
  50727=>"101000110",
  50728=>"111101000",
  50729=>"001100100",
  50730=>"111110100",
  50731=>"000010110",
  50732=>"010100001",
  50733=>"111001111",
  50734=>"111011011",
  50735=>"000000111",
  50736=>"001000011",
  50737=>"101000000",
  50738=>"000101011",
  50739=>"111000111",
  50740=>"000000110",
  50741=>"111101000",
  50742=>"011110101",
  50743=>"111100101",
  50744=>"010101001",
  50745=>"111010111",
  50746=>"000100010",
  50747=>"111010111",
  50748=>"010111011",
  50749=>"111010111",
  50750=>"110111111",
  50751=>"000110110",
  50752=>"111100010",
  50753=>"000101011",
  50754=>"100111000",
  50755=>"000001010",
  50756=>"000101101",
  50757=>"111000111",
  50758=>"100000010",
  50759=>"010011101",
  50760=>"100000111",
  50761=>"001111101",
  50762=>"000000100",
  50763=>"111101110",
  50764=>"001100000",
  50765=>"000101011",
  50766=>"101001110",
  50767=>"101010011",
  50768=>"010010111",
  50769=>"101100101",
  50770=>"101000101",
  50771=>"000010100",
  50772=>"110001101",
  50773=>"110111111",
  50774=>"111001111",
  50775=>"001010111",
  50776=>"010001000",
  50777=>"110010101",
  50778=>"100000000",
  50779=>"000000010",
  50780=>"110011101",
  50781=>"000100100",
  50782=>"011110101",
  50783=>"100001010",
  50784=>"011010000",
  50785=>"001100110",
  50786=>"100001101",
  50787=>"010111111",
  50788=>"101101100",
  50789=>"011000111",
  50790=>"101010000",
  50791=>"101111110",
  50792=>"001000011",
  50793=>"111000001",
  50794=>"110000000",
  50795=>"010011100",
  50796=>"110000001",
  50797=>"011101001",
  50798=>"111111110",
  50799=>"001110111",
  50800=>"000101101",
  50801=>"000000000",
  50802=>"111001110",
  50803=>"011111111",
  50804=>"011011100",
  50805=>"111000111",
  50806=>"110011111",
  50807=>"100000011",
  50808=>"010001010",
  50809=>"101011001",
  50810=>"101000001",
  50811=>"001000111",
  50812=>"000000001",
  50813=>"000000111",
  50814=>"101010100",
  50815=>"010001111",
  50816=>"001100010",
  50817=>"001111000",
  50818=>"101001111",
  50819=>"010110111",
  50820=>"100011100",
  50821=>"101010100",
  50822=>"110010110",
  50823=>"101111100",
  50824=>"111011111",
  50825=>"000001000",
  50826=>"110100110",
  50827=>"100100101",
  50828=>"000000100",
  50829=>"100100000",
  50830=>"011000100",
  50831=>"111101100",
  50832=>"001111010",
  50833=>"110001010",
  50834=>"001010100",
  50835=>"101100011",
  50836=>"101100100",
  50837=>"100100010",
  50838=>"001001010",
  50839=>"001011100",
  50840=>"110000011",
  50841=>"110111111",
  50842=>"010011010",
  50843=>"001000001",
  50844=>"111011010",
  50845=>"101010000",
  50846=>"111010010",
  50847=>"101000110",
  50848=>"001000010",
  50849=>"010001010",
  50850=>"101011110",
  50851=>"110100111",
  50852=>"010000111",
  50853=>"000010110",
  50854=>"010001000",
  50855=>"000100010",
  50856=>"000100011",
  50857=>"101110110",
  50858=>"101000001",
  50859=>"000111101",
  50860=>"100001010",
  50861=>"011101000",
  50862=>"111001011",
  50863=>"000000011",
  50864=>"100010101",
  50865=>"111100000",
  50866=>"010001001",
  50867=>"100000011",
  50868=>"010101111",
  50869=>"100110110",
  50870=>"010011110",
  50871=>"110101111",
  50872=>"101111001",
  50873=>"011000001",
  50874=>"011111111",
  50875=>"101101001",
  50876=>"000100000",
  50877=>"001110010",
  50878=>"000101011",
  50879=>"011000110",
  50880=>"110111010",
  50881=>"110101011",
  50882=>"000010111",
  50883=>"110011111",
  50884=>"111010000",
  50885=>"100010110",
  50886=>"011010110",
  50887=>"001001100",
  50888=>"011000000",
  50889=>"111111100",
  50890=>"010000000",
  50891=>"100100111",
  50892=>"000001001",
  50893=>"000101100",
  50894=>"110001000",
  50895=>"010010001",
  50896=>"000010110",
  50897=>"110110010",
  50898=>"000110110",
  50899=>"010001011",
  50900=>"011010111",
  50901=>"111001010",
  50902=>"100100000",
  50903=>"111111011",
  50904=>"010010010",
  50905=>"100001001",
  50906=>"111111110",
  50907=>"111100100",
  50908=>"100110110",
  50909=>"010101010",
  50910=>"100000000",
  50911=>"111101110",
  50912=>"100000100",
  50913=>"000000010",
  50914=>"000001000",
  50915=>"111010010",
  50916=>"101000010",
  50917=>"001111001",
  50918=>"010011010",
  50919=>"010101000",
  50920=>"010111100",
  50921=>"111111100",
  50922=>"000111010",
  50923=>"001110110",
  50924=>"001110100",
  50925=>"100010010",
  50926=>"001001010",
  50927=>"011011011",
  50928=>"001000100",
  50929=>"011000011",
  50930=>"111000110",
  50931=>"111100011",
  50932=>"001011011",
  50933=>"010010110",
  50934=>"010001010",
  50935=>"011100111",
  50936=>"011011110",
  50937=>"011110101",
  50938=>"100100000",
  50939=>"100100011",
  50940=>"111010101",
  50941=>"011101001",
  50942=>"111011110",
  50943=>"000001100",
  50944=>"111110111",
  50945=>"010100100",
  50946=>"100000000",
  50947=>"001100111",
  50948=>"100011111",
  50949=>"101001010",
  50950=>"100001001",
  50951=>"011001011",
  50952=>"110000001",
  50953=>"111111011",
  50954=>"101101010",
  50955=>"010110111",
  50956=>"000010101",
  50957=>"111011010",
  50958=>"001100101",
  50959=>"001111000",
  50960=>"001001111",
  50961=>"010110001",
  50962=>"100010010",
  50963=>"110000001",
  50964=>"101111101",
  50965=>"010011010",
  50966=>"111111111",
  50967=>"010110000",
  50968=>"101011011",
  50969=>"001011011",
  50970=>"100110100",
  50971=>"010011101",
  50972=>"010011101",
  50973=>"101000010",
  50974=>"110011101",
  50975=>"111001101",
  50976=>"010011101",
  50977=>"111011011",
  50978=>"000111110",
  50979=>"110110011",
  50980=>"111101100",
  50981=>"111100101",
  50982=>"111110110",
  50983=>"000101111",
  50984=>"011010000",
  50985=>"001010101",
  50986=>"011111110",
  50987=>"001111100",
  50988=>"001011011",
  50989=>"000010101",
  50990=>"111101111",
  50991=>"010101010",
  50992=>"011010111",
  50993=>"110101001",
  50994=>"101011101",
  50995=>"010001100",
  50996=>"011011010",
  50997=>"011111100",
  50998=>"111101101",
  50999=>"101111100",
  51000=>"011000000",
  51001=>"101100110",
  51002=>"000111100",
  51003=>"011110011",
  51004=>"100001001",
  51005=>"000111101",
  51006=>"110111000",
  51007=>"010011111",
  51008=>"010100001",
  51009=>"000001011",
  51010=>"000110110",
  51011=>"101001001",
  51012=>"100111111",
  51013=>"101101010",
  51014=>"111101111",
  51015=>"001100011",
  51016=>"110111011",
  51017=>"011100101",
  51018=>"010111111",
  51019=>"111010100",
  51020=>"011011000",
  51021=>"100001000",
  51022=>"110011011",
  51023=>"110101111",
  51024=>"111111111",
  51025=>"010011010",
  51026=>"011100100",
  51027=>"011000110",
  51028=>"111010111",
  51029=>"010110001",
  51030=>"101111010",
  51031=>"010111000",
  51032=>"001101001",
  51033=>"110010001",
  51034=>"111010010",
  51035=>"110010101",
  51036=>"110001011",
  51037=>"011010100",
  51038=>"111100000",
  51039=>"001000000",
  51040=>"101010011",
  51041=>"110101101",
  51042=>"101010111",
  51043=>"001110110",
  51044=>"010100001",
  51045=>"010111000",
  51046=>"110110011",
  51047=>"111011010",
  51048=>"110010001",
  51049=>"010010000",
  51050=>"001000110",
  51051=>"111111111",
  51052=>"011010100",
  51053=>"001010001",
  51054=>"101111110",
  51055=>"100011000",
  51056=>"101001101",
  51057=>"000000110",
  51058=>"101100111",
  51059=>"010010010",
  51060=>"011000000",
  51061=>"001110110",
  51062=>"111100100",
  51063=>"001001111",
  51064=>"000110100",
  51065=>"100101110",
  51066=>"111111100",
  51067=>"110100111",
  51068=>"010001111",
  51069=>"001001011",
  51070=>"010111100",
  51071=>"111110000",
  51072=>"110100010",
  51073=>"110100011",
  51074=>"010011010",
  51075=>"010111001",
  51076=>"110010101",
  51077=>"011001000",
  51078=>"101111111",
  51079=>"110000101",
  51080=>"000110010",
  51081=>"111011011",
  51082=>"101010011",
  51083=>"111111111",
  51084=>"000001101",
  51085=>"000000100",
  51086=>"100001101",
  51087=>"100100100",
  51088=>"111110110",
  51089=>"101101111",
  51090=>"111001111",
  51091=>"000100111",
  51092=>"110100111",
  51093=>"011100011",
  51094=>"000100000",
  51095=>"000110010",
  51096=>"110111011",
  51097=>"000010000",
  51098=>"010100000",
  51099=>"101000011",
  51100=>"110111110",
  51101=>"000100100",
  51102=>"111001001",
  51103=>"010011001",
  51104=>"001111100",
  51105=>"101010111",
  51106=>"000000101",
  51107=>"010001010",
  51108=>"000000010",
  51109=>"110000101",
  51110=>"010011000",
  51111=>"001000010",
  51112=>"010001110",
  51113=>"010010011",
  51114=>"100100001",
  51115=>"001110111",
  51116=>"110010001",
  51117=>"101111110",
  51118=>"000111101",
  51119=>"100100001",
  51120=>"010000000",
  51121=>"001100001",
  51122=>"011001001",
  51123=>"110111111",
  51124=>"000110100",
  51125=>"101101010",
  51126=>"001011011",
  51127=>"110110011",
  51128=>"111111110",
  51129=>"001111011",
  51130=>"100001000",
  51131=>"100111101",
  51132=>"111100111",
  51133=>"111010001",
  51134=>"111001010",
  51135=>"111111001",
  51136=>"101000101",
  51137=>"011000101",
  51138=>"100000011",
  51139=>"100110011",
  51140=>"110111101",
  51141=>"010101001",
  51142=>"001001010",
  51143=>"000011001",
  51144=>"100100110",
  51145=>"001011110",
  51146=>"101110010",
  51147=>"001111111",
  51148=>"001011100",
  51149=>"100110111",
  51150=>"011000110",
  51151=>"001010111",
  51152=>"110110110",
  51153=>"000000110",
  51154=>"011000001",
  51155=>"001011000",
  51156=>"101001111",
  51157=>"101111011",
  51158=>"110100111",
  51159=>"000010001",
  51160=>"101010101",
  51161=>"110000101",
  51162=>"000010100",
  51163=>"010010011",
  51164=>"010101010",
  51165=>"100010011",
  51166=>"100110001",
  51167=>"111110111",
  51168=>"010110110",
  51169=>"111101010",
  51170=>"000011100",
  51171=>"000110101",
  51172=>"101111011",
  51173=>"010100100",
  51174=>"100001010",
  51175=>"110100000",
  51176=>"000011011",
  51177=>"110100111",
  51178=>"000010100",
  51179=>"000100111",
  51180=>"111111101",
  51181=>"101001010",
  51182=>"111010110",
  51183=>"111101010",
  51184=>"111101011",
  51185=>"000111111",
  51186=>"111010101",
  51187=>"010111011",
  51188=>"100001100",
  51189=>"100111111",
  51190=>"110011101",
  51191=>"000010100",
  51192=>"001100111",
  51193=>"101001011",
  51194=>"101010010",
  51195=>"101011000",
  51196=>"100110001",
  51197=>"110111100",
  51198=>"101010101",
  51199=>"101100011",
  51200=>"110010111",
  51201=>"000101001",
  51202=>"001001110",
  51203=>"010100110",
  51204=>"001010000",
  51205=>"011011011",
  51206=>"011111110",
  51207=>"010101100",
  51208=>"010100011",
  51209=>"011101101",
  51210=>"001110101",
  51211=>"010011110",
  51212=>"100100100",
  51213=>"111000111",
  51214=>"001110100",
  51215=>"111011110",
  51216=>"010100010",
  51217=>"110011110",
  51218=>"010010110",
  51219=>"100111000",
  51220=>"010101100",
  51221=>"101100001",
  51222=>"001110111",
  51223=>"100101100",
  51224=>"110001101",
  51225=>"000110111",
  51226=>"100010011",
  51227=>"010000111",
  51228=>"010011111",
  51229=>"100100000",
  51230=>"010100011",
  51231=>"100110100",
  51232=>"111000011",
  51233=>"101011100",
  51234=>"001000100",
  51235=>"000111000",
  51236=>"110001110",
  51237=>"101110001",
  51238=>"111100110",
  51239=>"000001100",
  51240=>"101111000",
  51241=>"010100001",
  51242=>"010001111",
  51243=>"101110010",
  51244=>"001111101",
  51245=>"011111101",
  51246=>"000011010",
  51247=>"001001111",
  51248=>"011011000",
  51249=>"101011111",
  51250=>"000100001",
  51251=>"101110111",
  51252=>"010000000",
  51253=>"111111101",
  51254=>"000011111",
  51255=>"000010101",
  51256=>"001101011",
  51257=>"100010111",
  51258=>"000010101",
  51259=>"010111101",
  51260=>"101001011",
  51261=>"100100000",
  51262=>"010011011",
  51263=>"110101001",
  51264=>"100010110",
  51265=>"010000000",
  51266=>"010011000",
  51267=>"000000011",
  51268=>"101100111",
  51269=>"101011010",
  51270=>"000001101",
  51271=>"110101000",
  51272=>"111000011",
  51273=>"010111000",
  51274=>"110010100",
  51275=>"001000011",
  51276=>"000100000",
  51277=>"000011100",
  51278=>"101001110",
  51279=>"111100101",
  51280=>"010011000",
  51281=>"011111010",
  51282=>"000000010",
  51283=>"010110011",
  51284=>"100101011",
  51285=>"010011101",
  51286=>"101110010",
  51287=>"101000000",
  51288=>"011101111",
  51289=>"001110010",
  51290=>"101010000",
  51291=>"011000010",
  51292=>"111010011",
  51293=>"000001000",
  51294=>"101100010",
  51295=>"100001000",
  51296=>"000011001",
  51297=>"000010101",
  51298=>"010011111",
  51299=>"100111011",
  51300=>"101101110",
  51301=>"010111010",
  51302=>"101111111",
  51303=>"011011000",
  51304=>"001100100",
  51305=>"111000111",
  51306=>"000010001",
  51307=>"001011110",
  51308=>"000001001",
  51309=>"011111001",
  51310=>"001100001",
  51311=>"000101011",
  51312=>"000101101",
  51313=>"101001000",
  51314=>"011011110",
  51315=>"010110010",
  51316=>"111111011",
  51317=>"001011010",
  51318=>"101011010",
  51319=>"000101010",
  51320=>"000101110",
  51321=>"010011010",
  51322=>"101001000",
  51323=>"000010111",
  51324=>"101101011",
  51325=>"110010010",
  51326=>"110101101",
  51327=>"010110010",
  51328=>"000101000",
  51329=>"010101001",
  51330=>"000001001",
  51331=>"011101111",
  51332=>"110001000",
  51333=>"010100001",
  51334=>"011001111",
  51335=>"111100101",
  51336=>"111100101",
  51337=>"011100000",
  51338=>"100101010",
  51339=>"011000101",
  51340=>"001101000",
  51341=>"000101101",
  51342=>"100110111",
  51343=>"111101110",
  51344=>"100111000",
  51345=>"111101000",
  51346=>"010111110",
  51347=>"110111111",
  51348=>"010101111",
  51349=>"101000000",
  51350=>"100011010",
  51351=>"101010101",
  51352=>"001001000",
  51353=>"111001011",
  51354=>"111001010",
  51355=>"110001111",
  51356=>"111110111",
  51357=>"010010101",
  51358=>"001111001",
  51359=>"100110010",
  51360=>"001101010",
  51361=>"101110110",
  51362=>"010010001",
  51363=>"100010111",
  51364=>"001110001",
  51365=>"101101100",
  51366=>"010111010",
  51367=>"110100000",
  51368=>"011001110",
  51369=>"101111111",
  51370=>"010010011",
  51371=>"111100100",
  51372=>"100011100",
  51373=>"011111011",
  51374=>"000111111",
  51375=>"110001100",
  51376=>"001111100",
  51377=>"001010001",
  51378=>"011000111",
  51379=>"010101000",
  51380=>"010101111",
  51381=>"111011000",
  51382=>"010111011",
  51383=>"001111000",
  51384=>"011100111",
  51385=>"001000000",
  51386=>"100110110",
  51387=>"110100111",
  51388=>"000101001",
  51389=>"100001001",
  51390=>"110000010",
  51391=>"101011100",
  51392=>"000001000",
  51393=>"110111110",
  51394=>"000100111",
  51395=>"101110110",
  51396=>"101101010",
  51397=>"101001000",
  51398=>"110111000",
  51399=>"010110000",
  51400=>"010011111",
  51401=>"101011000",
  51402=>"100110111",
  51403=>"000100111",
  51404=>"111000000",
  51405=>"000101100",
  51406=>"011100111",
  51407=>"010001110",
  51408=>"111110101",
  51409=>"001101101",
  51410=>"110000111",
  51411=>"101010101",
  51412=>"001100100",
  51413=>"110011101",
  51414=>"000111101",
  51415=>"101010000",
  51416=>"001000011",
  51417=>"000010100",
  51418=>"010000001",
  51419=>"110110111",
  51420=>"100111110",
  51421=>"111101001",
  51422=>"110111111",
  51423=>"001111011",
  51424=>"100011011",
  51425=>"000010100",
  51426=>"111111011",
  51427=>"010110000",
  51428=>"000110001",
  51429=>"000100011",
  51430=>"001001011",
  51431=>"101101000",
  51432=>"000010111",
  51433=>"101111011",
  51434=>"111011111",
  51435=>"110000000",
  51436=>"111101110",
  51437=>"010110001",
  51438=>"010010000",
  51439=>"001000011",
  51440=>"011101100",
  51441=>"000110011",
  51442=>"101011100",
  51443=>"010111101",
  51444=>"100001000",
  51445=>"110010011",
  51446=>"100100100",
  51447=>"111111111",
  51448=>"000111101",
  51449=>"001010011",
  51450=>"111101111",
  51451=>"111011001",
  51452=>"001000000",
  51453=>"001100111",
  51454=>"011001110",
  51455=>"101111100",
  51456=>"101100001",
  51457=>"110000000",
  51458=>"100001101",
  51459=>"110001111",
  51460=>"000111000",
  51461=>"111100100",
  51462=>"000000101",
  51463=>"000001001",
  51464=>"000011100",
  51465=>"001101000",
  51466=>"010100011",
  51467=>"100000000",
  51468=>"001100001",
  51469=>"001000001",
  51470=>"110111100",
  51471=>"010100111",
  51472=>"001010011",
  51473=>"000001011",
  51474=>"100110011",
  51475=>"100101011",
  51476=>"010001011",
  51477=>"011010000",
  51478=>"000101010",
  51479=>"010100100",
  51480=>"010100001",
  51481=>"101110111",
  51482=>"110110001",
  51483=>"000111001",
  51484=>"010111111",
  51485=>"000110000",
  51486=>"000111011",
  51487=>"000011101",
  51488=>"000100100",
  51489=>"000011110",
  51490=>"000101100",
  51491=>"110000110",
  51492=>"001011110",
  51493=>"011110111",
  51494=>"010000000",
  51495=>"001000110",
  51496=>"111111110",
  51497=>"010000011",
  51498=>"010111011",
  51499=>"101110000",
  51500=>"001101011",
  51501=>"100000110",
  51502=>"001010101",
  51503=>"110101110",
  51504=>"000011101",
  51505=>"110000000",
  51506=>"010010111",
  51507=>"000011110",
  51508=>"100000100",
  51509=>"100010110",
  51510=>"001110000",
  51511=>"010011111",
  51512=>"110011110",
  51513=>"000001000",
  51514=>"110110100",
  51515=>"001010001",
  51516=>"110001111",
  51517=>"010011101",
  51518=>"011011011",
  51519=>"000000000",
  51520=>"111111101",
  51521=>"110101001",
  51522=>"001001111",
  51523=>"010010001",
  51524=>"110100110",
  51525=>"000011110",
  51526=>"101001110",
  51527=>"101110100",
  51528=>"000011110",
  51529=>"000010001",
  51530=>"101001001",
  51531=>"010110001",
  51532=>"010111101",
  51533=>"000110110",
  51534=>"011100000",
  51535=>"011010001",
  51536=>"010011011",
  51537=>"001101001",
  51538=>"100011110",
  51539=>"101111111",
  51540=>"010001110",
  51541=>"000011111",
  51542=>"000101100",
  51543=>"011001111",
  51544=>"001011100",
  51545=>"010111010",
  51546=>"000110110",
  51547=>"100110010",
  51548=>"000110111",
  51549=>"110101101",
  51550=>"101010001",
  51551=>"110010100",
  51552=>"101110011",
  51553=>"011101001",
  51554=>"000001010",
  51555=>"101000110",
  51556=>"011100100",
  51557=>"110000011",
  51558=>"001101001",
  51559=>"001111011",
  51560=>"101100111",
  51561=>"000000111",
  51562=>"101101010",
  51563=>"100011111",
  51564=>"000110010",
  51565=>"110000101",
  51566=>"000011001",
  51567=>"110010110",
  51568=>"010111111",
  51569=>"100101001",
  51570=>"001101011",
  51571=>"110010001",
  51572=>"010111000",
  51573=>"011001111",
  51574=>"101101001",
  51575=>"011001110",
  51576=>"111111111",
  51577=>"010001101",
  51578=>"111010000",
  51579=>"011100001",
  51580=>"011100001",
  51581=>"000101100",
  51582=>"101010101",
  51583=>"111111010",
  51584=>"101110100",
  51585=>"000110001",
  51586=>"110011001",
  51587=>"010111111",
  51588=>"000011101",
  51589=>"011101100",
  51590=>"100011110",
  51591=>"111011110",
  51592=>"101000100",
  51593=>"101100001",
  51594=>"001100010",
  51595=>"010001010",
  51596=>"111000000",
  51597=>"000111000",
  51598=>"101101100",
  51599=>"101110100",
  51600=>"100011110",
  51601=>"000100000",
  51602=>"000011011",
  51603=>"001100001",
  51604=>"100111000",
  51605=>"100000010",
  51606=>"111001111",
  51607=>"011011000",
  51608=>"011011010",
  51609=>"110111000",
  51610=>"011111010",
  51611=>"101001101",
  51612=>"111101111",
  51613=>"101100111",
  51614=>"011111110",
  51615=>"000110100",
  51616=>"000111010",
  51617=>"100110001",
  51618=>"001000101",
  51619=>"110110010",
  51620=>"101010011",
  51621=>"101101011",
  51622=>"000001011",
  51623=>"110011111",
  51624=>"100100011",
  51625=>"000001001",
  51626=>"011111111",
  51627=>"010001101",
  51628=>"011101100",
  51629=>"001001100",
  51630=>"110001011",
  51631=>"000101100",
  51632=>"010101000",
  51633=>"001010111",
  51634=>"100001000",
  51635=>"001001101",
  51636=>"011110000",
  51637=>"101000100",
  51638=>"110000111",
  51639=>"001110101",
  51640=>"110101111",
  51641=>"000100100",
  51642=>"001000100",
  51643=>"010101011",
  51644=>"100001111",
  51645=>"111001010",
  51646=>"110111111",
  51647=>"111111100",
  51648=>"100011000",
  51649=>"001010111",
  51650=>"001111100",
  51651=>"111111111",
  51652=>"000010000",
  51653=>"111111011",
  51654=>"111001100",
  51655=>"011001010",
  51656=>"000111001",
  51657=>"111100010",
  51658=>"000000001",
  51659=>"111000101",
  51660=>"000000011",
  51661=>"100101010",
  51662=>"101111100",
  51663=>"110100101",
  51664=>"001111000",
  51665=>"010000000",
  51666=>"110010000",
  51667=>"011100100",
  51668=>"101111011",
  51669=>"001111100",
  51670=>"011111011",
  51671=>"101000100",
  51672=>"111011111",
  51673=>"111111100",
  51674=>"001001001",
  51675=>"101110110",
  51676=>"111000100",
  51677=>"010001001",
  51678=>"100000010",
  51679=>"111001001",
  51680=>"111101001",
  51681=>"100001110",
  51682=>"100111111",
  51683=>"000000010",
  51684=>"011001110",
  51685=>"011001101",
  51686=>"010100011",
  51687=>"000101000",
  51688=>"010011001",
  51689=>"010010111",
  51690=>"110000001",
  51691=>"101011010",
  51692=>"100011111",
  51693=>"100000000",
  51694=>"101111110",
  51695=>"010011100",
  51696=>"110001111",
  51697=>"100100011",
  51698=>"101000111",
  51699=>"101101000",
  51700=>"101101111",
  51701=>"011011110",
  51702=>"111100100",
  51703=>"001101010",
  51704=>"001000110",
  51705=>"101000011",
  51706=>"010110100",
  51707=>"110110111",
  51708=>"110010111",
  51709=>"110101101",
  51710=>"010101110",
  51711=>"010111000",
  51712=>"100010100",
  51713=>"100001010",
  51714=>"111010001",
  51715=>"000100001",
  51716=>"011100110",
  51717=>"100111101",
  51718=>"001010011",
  51719=>"111001010",
  51720=>"010010100",
  51721=>"010000000",
  51722=>"001101110",
  51723=>"111101010",
  51724=>"000101111",
  51725=>"011110111",
  51726=>"000010111",
  51727=>"011000010",
  51728=>"000111101",
  51729=>"010101010",
  51730=>"111100101",
  51731=>"110001010",
  51732=>"111010111",
  51733=>"100010010",
  51734=>"111101011",
  51735=>"101000010",
  51736=>"100010100",
  51737=>"101010101",
  51738=>"001001111",
  51739=>"010011001",
  51740=>"111110110",
  51741=>"000001101",
  51742=>"100100011",
  51743=>"000011010",
  51744=>"110111010",
  51745=>"110110011",
  51746=>"001000010",
  51747=>"000010100",
  51748=>"110111101",
  51749=>"100010101",
  51750=>"111011000",
  51751=>"111001000",
  51752=>"101110110",
  51753=>"100001000",
  51754=>"000100101",
  51755=>"000100111",
  51756=>"001001111",
  51757=>"010101001",
  51758=>"110101100",
  51759=>"011100001",
  51760=>"001000001",
  51761=>"101100101",
  51762=>"011101111",
  51763=>"110110010",
  51764=>"011000101",
  51765=>"011101011",
  51766=>"001100111",
  51767=>"010100001",
  51768=>"001001100",
  51769=>"011110010",
  51770=>"000001100",
  51771=>"000110110",
  51772=>"110111111",
  51773=>"110001000",
  51774=>"001101101",
  51775=>"001110000",
  51776=>"011001110",
  51777=>"011101000",
  51778=>"100101011",
  51779=>"100101101",
  51780=>"010000000",
  51781=>"001001011",
  51782=>"110000001",
  51783=>"000100010",
  51784=>"111100111",
  51785=>"000110001",
  51786=>"110100101",
  51787=>"111001110",
  51788=>"000111111",
  51789=>"010101100",
  51790=>"010110010",
  51791=>"111010000",
  51792=>"000100101",
  51793=>"100101101",
  51794=>"001000011",
  51795=>"111101000",
  51796=>"000000111",
  51797=>"011010000",
  51798=>"101110000",
  51799=>"110100010",
  51800=>"101011111",
  51801=>"100000010",
  51802=>"101011111",
  51803=>"101011010",
  51804=>"000001100",
  51805=>"011011011",
  51806=>"001011100",
  51807=>"001110000",
  51808=>"000001101",
  51809=>"110100000",
  51810=>"010001110",
  51811=>"011110100",
  51812=>"101011111",
  51813=>"111111001",
  51814=>"001100010",
  51815=>"010101111",
  51816=>"000100000",
  51817=>"000101111",
  51818=>"001111000",
  51819=>"101000110",
  51820=>"100101000",
  51821=>"111110101",
  51822=>"000000110",
  51823=>"100010111",
  51824=>"001010000",
  51825=>"011000000",
  51826=>"011111101",
  51827=>"011100100",
  51828=>"011001001",
  51829=>"001011001",
  51830=>"101101010",
  51831=>"110111000",
  51832=>"001100110",
  51833=>"110011001",
  51834=>"101000100",
  51835=>"110101010",
  51836=>"111101000",
  51837=>"111110010",
  51838=>"100010000",
  51839=>"010011100",
  51840=>"101100000",
  51841=>"111010111",
  51842=>"110010100",
  51843=>"000101110",
  51844=>"010011110",
  51845=>"001001001",
  51846=>"011001000",
  51847=>"011011010",
  51848=>"110011110",
  51849=>"101000001",
  51850=>"011111110",
  51851=>"101010110",
  51852=>"111110111",
  51853=>"100111101",
  51854=>"001001001",
  51855=>"100000101",
  51856=>"011110101",
  51857=>"100101101",
  51858=>"010100001",
  51859=>"100011100",
  51860=>"101111000",
  51861=>"011100101",
  51862=>"010101100",
  51863=>"101101000",
  51864=>"101101100",
  51865=>"100101101",
  51866=>"100011110",
  51867=>"000110111",
  51868=>"100000111",
  51869=>"111001101",
  51870=>"000001001",
  51871=>"110101101",
  51872=>"111101111",
  51873=>"001000101",
  51874=>"011100001",
  51875=>"110111110",
  51876=>"011001000",
  51877=>"111000001",
  51878=>"001101101",
  51879=>"110111110",
  51880=>"000011100",
  51881=>"100000011",
  51882=>"001100110",
  51883=>"101110001",
  51884=>"010011000",
  51885=>"111010110",
  51886=>"000000000",
  51887=>"010010011",
  51888=>"000010000",
  51889=>"011100101",
  51890=>"001110111",
  51891=>"101111111",
  51892=>"001111011",
  51893=>"110111110",
  51894=>"100101110",
  51895=>"000010100",
  51896=>"011100110",
  51897=>"101101011",
  51898=>"100011010",
  51899=>"100111010",
  51900=>"110100000",
  51901=>"000000000",
  51902=>"000100010",
  51903=>"001011011",
  51904=>"110100001",
  51905=>"111100111",
  51906=>"010101101",
  51907=>"010000000",
  51908=>"101011010",
  51909=>"101001101",
  51910=>"010000000",
  51911=>"101101101",
  51912=>"010001000",
  51913=>"010000100",
  51914=>"101010110",
  51915=>"100010100",
  51916=>"010010100",
  51917=>"010110010",
  51918=>"000011001",
  51919=>"001010100",
  51920=>"101100111",
  51921=>"100100110",
  51922=>"010101111",
  51923=>"101001110",
  51924=>"011001000",
  51925=>"000011101",
  51926=>"000001001",
  51927=>"101010001",
  51928=>"011010011",
  51929=>"010010100",
  51930=>"001000101",
  51931=>"001100110",
  51932=>"100101110",
  51933=>"101011111",
  51934=>"100100111",
  51935=>"010000010",
  51936=>"101000110",
  51937=>"110110000",
  51938=>"100001110",
  51939=>"110011010",
  51940=>"011110101",
  51941=>"010010010",
  51942=>"000011100",
  51943=>"000010001",
  51944=>"001001111",
  51945=>"001101101",
  51946=>"110100000",
  51947=>"111101100",
  51948=>"000000111",
  51949=>"000001001",
  51950=>"000001110",
  51951=>"100001000",
  51952=>"111001101",
  51953=>"001010010",
  51954=>"011001100",
  51955=>"110100111",
  51956=>"001010111",
  51957=>"101110011",
  51958=>"011110111",
  51959=>"111001100",
  51960=>"010000101",
  51961=>"101011000",
  51962=>"010001011",
  51963=>"011110111",
  51964=>"011000110",
  51965=>"110000001",
  51966=>"100000011",
  51967=>"011011010",
  51968=>"111101001",
  51969=>"000000101",
  51970=>"010011101",
  51971=>"000010110",
  51972=>"010000000",
  51973=>"110001011",
  51974=>"110010100",
  51975=>"100011110",
  51976=>"111111010",
  51977=>"000011010",
  51978=>"101011011",
  51979=>"110110111",
  51980=>"010101110",
  51981=>"011010001",
  51982=>"111000111",
  51983=>"001001111",
  51984=>"111110000",
  51985=>"000100010",
  51986=>"100001011",
  51987=>"101110000",
  51988=>"100011100",
  51989=>"011000110",
  51990=>"101100001",
  51991=>"100100000",
  51992=>"100000000",
  51993=>"001100011",
  51994=>"001010111",
  51995=>"110011101",
  51996=>"101110100",
  51997=>"110000000",
  51998=>"100110000",
  51999=>"100001000",
  52000=>"011111100",
  52001=>"111011000",
  52002=>"101110010",
  52003=>"110000011",
  52004=>"111110011",
  52005=>"101001101",
  52006=>"100000001",
  52007=>"000000101",
  52008=>"110010000",
  52009=>"000001000",
  52010=>"111100000",
  52011=>"001001111",
  52012=>"111100000",
  52013=>"110010000",
  52014=>"001001111",
  52015=>"001111111",
  52016=>"000001111",
  52017=>"001001000",
  52018=>"001000001",
  52019=>"101101110",
  52020=>"111111100",
  52021=>"001001010",
  52022=>"011000000",
  52023=>"010001110",
  52024=>"111000110",
  52025=>"110001011",
  52026=>"011111100",
  52027=>"101000001",
  52028=>"010100111",
  52029=>"110000010",
  52030=>"110111001",
  52031=>"101000100",
  52032=>"010111110",
  52033=>"000010111",
  52034=>"010110001",
  52035=>"110011001",
  52036=>"100001010",
  52037=>"000001010",
  52038=>"111100100",
  52039=>"111001110",
  52040=>"001101111",
  52041=>"101010000",
  52042=>"001010011",
  52043=>"010000011",
  52044=>"111101111",
  52045=>"000000100",
  52046=>"110111000",
  52047=>"001000100",
  52048=>"111011010",
  52049=>"000011101",
  52050=>"100111011",
  52051=>"111001111",
  52052=>"101100011",
  52053=>"000110111",
  52054=>"101111111",
  52055=>"001101000",
  52056=>"001000000",
  52057=>"001011000",
  52058=>"100111100",
  52059=>"010111010",
  52060=>"101001110",
  52061=>"101100111",
  52062=>"111111111",
  52063=>"010010010",
  52064=>"010110100",
  52065=>"110000010",
  52066=>"001001101",
  52067=>"011000010",
  52068=>"110100101",
  52069=>"010100011",
  52070=>"011110010",
  52071=>"000111110",
  52072=>"100010001",
  52073=>"111011111",
  52074=>"011101111",
  52075=>"100101001",
  52076=>"111101100",
  52077=>"110001110",
  52078=>"011010000",
  52079=>"011100011",
  52080=>"101001100",
  52081=>"101110111",
  52082=>"001101011",
  52083=>"101000010",
  52084=>"001010101",
  52085=>"000100111",
  52086=>"111111011",
  52087=>"010100100",
  52088=>"101101100",
  52089=>"001111000",
  52090=>"110100010",
  52091=>"010110001",
  52092=>"011000111",
  52093=>"000101111",
  52094=>"111001100",
  52095=>"110000010",
  52096=>"010011011",
  52097=>"111101000",
  52098=>"110000011",
  52099=>"101100010",
  52100=>"111110001",
  52101=>"010001000",
  52102=>"010000101",
  52103=>"001000011",
  52104=>"100011101",
  52105=>"100111010",
  52106=>"111111110",
  52107=>"110000111",
  52108=>"101010011",
  52109=>"011010110",
  52110=>"111010001",
  52111=>"010011010",
  52112=>"001001111",
  52113=>"010110011",
  52114=>"101000110",
  52115=>"100111110",
  52116=>"111101011",
  52117=>"101001010",
  52118=>"100000111",
  52119=>"011001010",
  52120=>"010100010",
  52121=>"010011001",
  52122=>"010100110",
  52123=>"011100111",
  52124=>"001100110",
  52125=>"010110001",
  52126=>"010110000",
  52127=>"100100001",
  52128=>"110100001",
  52129=>"110110110",
  52130=>"001101000",
  52131=>"100110110",
  52132=>"110111101",
  52133=>"001010000",
  52134=>"110001111",
  52135=>"100100011",
  52136=>"111110101",
  52137=>"000001100",
  52138=>"001110011",
  52139=>"000100110",
  52140=>"110000111",
  52141=>"010000000",
  52142=>"000000000",
  52143=>"111111100",
  52144=>"010011000",
  52145=>"101111010",
  52146=>"001110110",
  52147=>"010101101",
  52148=>"111100000",
  52149=>"000110000",
  52150=>"110101010",
  52151=>"000111100",
  52152=>"011000011",
  52153=>"100010010",
  52154=>"010011010",
  52155=>"011111011",
  52156=>"001011000",
  52157=>"100000001",
  52158=>"111100101",
  52159=>"001110100",
  52160=>"000101101",
  52161=>"001100111",
  52162=>"001100100",
  52163=>"110001011",
  52164=>"111110011",
  52165=>"110110011",
  52166=>"101111111",
  52167=>"011111111",
  52168=>"101110000",
  52169=>"111001010",
  52170=>"101111010",
  52171=>"110011000",
  52172=>"101110101",
  52173=>"110001001",
  52174=>"111000111",
  52175=>"011000101",
  52176=>"010101111",
  52177=>"111100011",
  52178=>"000101100",
  52179=>"100110100",
  52180=>"000001110",
  52181=>"011001101",
  52182=>"011011100",
  52183=>"101011001",
  52184=>"101011101",
  52185=>"001001100",
  52186=>"101001000",
  52187=>"100101001",
  52188=>"101110101",
  52189=>"111110100",
  52190=>"000100011",
  52191=>"110100011",
  52192=>"101011011",
  52193=>"011101010",
  52194=>"011110100",
  52195=>"011000001",
  52196=>"101011000",
  52197=>"001001001",
  52198=>"100111110",
  52199=>"010011100",
  52200=>"110100111",
  52201=>"100010001",
  52202=>"010000001",
  52203=>"000001100",
  52204=>"011000001",
  52205=>"000100000",
  52206=>"011101010",
  52207=>"000010010",
  52208=>"010011110",
  52209=>"100100000",
  52210=>"000100111",
  52211=>"110000010",
  52212=>"011010111",
  52213=>"001000111",
  52214=>"110110010",
  52215=>"100000001",
  52216=>"010110101",
  52217=>"000100011",
  52218=>"001001011",
  52219=>"000111011",
  52220=>"100001101",
  52221=>"101111010",
  52222=>"110000111",
  52223=>"011001100",
  52224=>"010111000",
  52225=>"001001111",
  52226=>"100110000",
  52227=>"011010000",
  52228=>"010001111",
  52229=>"001010110",
  52230=>"000000101",
  52231=>"111101011",
  52232=>"000000110",
  52233=>"010000100",
  52234=>"000110111",
  52235=>"100000101",
  52236=>"010000001",
  52237=>"111111010",
  52238=>"110010100",
  52239=>"010110100",
  52240=>"011101110",
  52241=>"001011000",
  52242=>"000100100",
  52243=>"000001100",
  52244=>"110110000",
  52245=>"011101110",
  52246=>"011011101",
  52247=>"100111101",
  52248=>"000001110",
  52249=>"010110001",
  52250=>"110100111",
  52251=>"110010101",
  52252=>"110101001",
  52253=>"011010100",
  52254=>"100010001",
  52255=>"011101000",
  52256=>"100001100",
  52257=>"010101100",
  52258=>"110100100",
  52259=>"000001110",
  52260=>"111111001",
  52261=>"000100111",
  52262=>"010110001",
  52263=>"100010111",
  52264=>"000000111",
  52265=>"001110110",
  52266=>"011010001",
  52267=>"111111110",
  52268=>"001001100",
  52269=>"000111111",
  52270=>"000011001",
  52271=>"111100100",
  52272=>"101001010",
  52273=>"001110001",
  52274=>"100010010",
  52275=>"010101111",
  52276=>"011111111",
  52277=>"111111111",
  52278=>"101011111",
  52279=>"000010110",
  52280=>"101101110",
  52281=>"010001100",
  52282=>"011001101",
  52283=>"010010100",
  52284=>"110111010",
  52285=>"111110000",
  52286=>"001001000",
  52287=>"100110001",
  52288=>"111011110",
  52289=>"110000000",
  52290=>"100101000",
  52291=>"101100100",
  52292=>"011111101",
  52293=>"100010111",
  52294=>"101110010",
  52295=>"100000110",
  52296=>"110111111",
  52297=>"110100100",
  52298=>"100000111",
  52299=>"100110001",
  52300=>"111011111",
  52301=>"111110111",
  52302=>"100111011",
  52303=>"000010101",
  52304=>"001000101",
  52305=>"010001101",
  52306=>"101011111",
  52307=>"001000011",
  52308=>"111001110",
  52309=>"100000001",
  52310=>"111001011",
  52311=>"011001001",
  52312=>"100001010",
  52313=>"110100011",
  52314=>"010100100",
  52315=>"111010010",
  52316=>"100110011",
  52317=>"100100000",
  52318=>"001111100",
  52319=>"100110111",
  52320=>"110000101",
  52321=>"101001101",
  52322=>"010100001",
  52323=>"110011000",
  52324=>"110010111",
  52325=>"111111111",
  52326=>"010000000",
  52327=>"011001100",
  52328=>"001100110",
  52329=>"000000110",
  52330=>"111010101",
  52331=>"011000010",
  52332=>"111011001",
  52333=>"010101011",
  52334=>"101111001",
  52335=>"001000000",
  52336=>"110110111",
  52337=>"000001011",
  52338=>"011001111",
  52339=>"000011101",
  52340=>"001011101",
  52341=>"100000001",
  52342=>"101100111",
  52343=>"111111000",
  52344=>"100111011",
  52345=>"110000010",
  52346=>"110011001",
  52347=>"100000011",
  52348=>"011110111",
  52349=>"000110101",
  52350=>"111100100",
  52351=>"010011000",
  52352=>"110010100",
  52353=>"000001101",
  52354=>"010001011",
  52355=>"000111101",
  52356=>"000010110",
  52357=>"011011110",
  52358=>"001011001",
  52359=>"110110101",
  52360=>"110000101",
  52361=>"111101000",
  52362=>"000000010",
  52363=>"110010111",
  52364=>"101000111",
  52365=>"101000011",
  52366=>"011100001",
  52367=>"000010000",
  52368=>"110000001",
  52369=>"000000110",
  52370=>"001110010",
  52371=>"010001111",
  52372=>"110001101",
  52373=>"001001000",
  52374=>"001111000",
  52375=>"011100101",
  52376=>"100001101",
  52377=>"111110101",
  52378=>"101111110",
  52379=>"000111001",
  52380=>"100010001",
  52381=>"001110111",
  52382=>"000100100",
  52383=>"001111100",
  52384=>"000111011",
  52385=>"000010000",
  52386=>"010100000",
  52387=>"100101011",
  52388=>"010101100",
  52389=>"110000011",
  52390=>"101111011",
  52391=>"101110001",
  52392=>"100001101",
  52393=>"001101001",
  52394=>"000111110",
  52395=>"110110110",
  52396=>"001011000",
  52397=>"100111000",
  52398=>"110010111",
  52399=>"011110001",
  52400=>"001000110",
  52401=>"110010001",
  52402=>"111001111",
  52403=>"001100110",
  52404=>"111111000",
  52405=>"000010000",
  52406=>"100101001",
  52407=>"000000000",
  52408=>"000011101",
  52409=>"001100010",
  52410=>"100001110",
  52411=>"101011100",
  52412=>"000001000",
  52413=>"000110001",
  52414=>"111010110",
  52415=>"100111011",
  52416=>"000010100",
  52417=>"100000000",
  52418=>"101110101",
  52419=>"011010101",
  52420=>"111101001",
  52421=>"000110101",
  52422=>"000111101",
  52423=>"101101000",
  52424=>"010000000",
  52425=>"111111111",
  52426=>"011010001",
  52427=>"100101000",
  52428=>"110110000",
  52429=>"011101110",
  52430=>"000111010",
  52431=>"010100100",
  52432=>"010001000",
  52433=>"010100000",
  52434=>"101111010",
  52435=>"101100111",
  52436=>"110000000",
  52437=>"000001010",
  52438=>"001010010",
  52439=>"001101000",
  52440=>"110011101",
  52441=>"001101101",
  52442=>"001010010",
  52443=>"101110000",
  52444=>"110101000",
  52445=>"110011100",
  52446=>"101001101",
  52447=>"001001101",
  52448=>"001101011",
  52449=>"001100000",
  52450=>"010001101",
  52451=>"101001001",
  52452=>"011101100",
  52453=>"010100000",
  52454=>"101111100",
  52455=>"000010100",
  52456=>"000000100",
  52457=>"100100010",
  52458=>"000001000",
  52459=>"001010101",
  52460=>"111000000",
  52461=>"100010000",
  52462=>"101011111",
  52463=>"111011000",
  52464=>"110111011",
  52465=>"011000000",
  52466=>"011101110",
  52467=>"000110111",
  52468=>"110100111",
  52469=>"000010001",
  52470=>"100011110",
  52471=>"111000111",
  52472=>"101111100",
  52473=>"101111111",
  52474=>"001101111",
  52475=>"011001011",
  52476=>"101101111",
  52477=>"001110100",
  52478=>"110111001",
  52479=>"001001001",
  52480=>"011110110",
  52481=>"110001010",
  52482=>"110111011",
  52483=>"010001100",
  52484=>"110101110",
  52485=>"011001110",
  52486=>"001001000",
  52487=>"010110110",
  52488=>"101100001",
  52489=>"011101100",
  52490=>"110110100",
  52491=>"001101100",
  52492=>"111111001",
  52493=>"111100011",
  52494=>"010010001",
  52495=>"011011100",
  52496=>"011111111",
  52497=>"110100110",
  52498=>"011111100",
  52499=>"010111010",
  52500=>"000010110",
  52501=>"001111001",
  52502=>"001001010",
  52503=>"000010100",
  52504=>"101000010",
  52505=>"101101010",
  52506=>"100010000",
  52507=>"110011010",
  52508=>"101110000",
  52509=>"100001000",
  52510=>"111111010",
  52511=>"000010010",
  52512=>"000110101",
  52513=>"110000100",
  52514=>"011110110",
  52515=>"010011000",
  52516=>"101100101",
  52517=>"001010001",
  52518=>"000100010",
  52519=>"101111111",
  52520=>"000011000",
  52521=>"101000001",
  52522=>"000111001",
  52523=>"000001001",
  52524=>"001011000",
  52525=>"000000100",
  52526=>"001101110",
  52527=>"010010100",
  52528=>"100101101",
  52529=>"001111000",
  52530=>"000010010",
  52531=>"110001111",
  52532=>"010100101",
  52533=>"011001110",
  52534=>"000001001",
  52535=>"001111111",
  52536=>"010110110",
  52537=>"011110000",
  52538=>"110100100",
  52539=>"101101001",
  52540=>"111100100",
  52541=>"001001011",
  52542=>"111111100",
  52543=>"010000110",
  52544=>"001101011",
  52545=>"011111100",
  52546=>"100000011",
  52547=>"110001101",
  52548=>"011010010",
  52549=>"110011010",
  52550=>"100011110",
  52551=>"010011011",
  52552=>"000001010",
  52553=>"111001001",
  52554=>"001000010",
  52555=>"110001110",
  52556=>"111111111",
  52557=>"000000001",
  52558=>"001111011",
  52559=>"111000000",
  52560=>"110100111",
  52561=>"000011100",
  52562=>"000001101",
  52563=>"001101000",
  52564=>"110100101",
  52565=>"000010001",
  52566=>"010001000",
  52567=>"100100001",
  52568=>"010001001",
  52569=>"111001000",
  52570=>"111010101",
  52571=>"101011011",
  52572=>"010100100",
  52573=>"001101000",
  52574=>"110011110",
  52575=>"001000001",
  52576=>"110001101",
  52577=>"000100001",
  52578=>"100111100",
  52579=>"011101010",
  52580=>"110111001",
  52581=>"010011010",
  52582=>"101000100",
  52583=>"111111100",
  52584=>"001010010",
  52585=>"000001000",
  52586=>"010010100",
  52587=>"000000010",
  52588=>"101110001",
  52589=>"001001110",
  52590=>"101011010",
  52591=>"011010010",
  52592=>"000101110",
  52593=>"011110010",
  52594=>"111001000",
  52595=>"010110011",
  52596=>"111010101",
  52597=>"011111111",
  52598=>"010101010",
  52599=>"100101100",
  52600=>"000011011",
  52601=>"100110100",
  52602=>"110001011",
  52603=>"111110001",
  52604=>"001111011",
  52605=>"000001100",
  52606=>"011100010",
  52607=>"110000111",
  52608=>"110011100",
  52609=>"100101110",
  52610=>"010101010",
  52611=>"111011100",
  52612=>"111101101",
  52613=>"101100110",
  52614=>"110101110",
  52615=>"000000111",
  52616=>"010010100",
  52617=>"100001000",
  52618=>"010011111",
  52619=>"000000000",
  52620=>"011000000",
  52621=>"110011000",
  52622=>"100110010",
  52623=>"100001100",
  52624=>"101011010",
  52625=>"000010010",
  52626=>"010011011",
  52627=>"011111011",
  52628=>"101001000",
  52629=>"101101010",
  52630=>"100011010",
  52631=>"100110100",
  52632=>"010100101",
  52633=>"000110100",
  52634=>"100000010",
  52635=>"000111011",
  52636=>"101101010",
  52637=>"111011011",
  52638=>"011001000",
  52639=>"010101001",
  52640=>"010110011",
  52641=>"011011101",
  52642=>"111010001",
  52643=>"111011110",
  52644=>"001000100",
  52645=>"101010010",
  52646=>"010010010",
  52647=>"111110111",
  52648=>"010000101",
  52649=>"000010010",
  52650=>"110111111",
  52651=>"101100101",
  52652=>"101100100",
  52653=>"110010111",
  52654=>"100001111",
  52655=>"001101101",
  52656=>"000000110",
  52657=>"100110000",
  52658=>"100100100",
  52659=>"000010101",
  52660=>"111011111",
  52661=>"110000001",
  52662=>"011011000",
  52663=>"101011111",
  52664=>"111000111",
  52665=>"111101001",
  52666=>"001111001",
  52667=>"110011000",
  52668=>"010100110",
  52669=>"010101011",
  52670=>"010000101",
  52671=>"100101000",
  52672=>"010000010",
  52673=>"110011101",
  52674=>"011001000",
  52675=>"000010100",
  52676=>"100011001",
  52677=>"000101111",
  52678=>"010110001",
  52679=>"010110000",
  52680=>"000111110",
  52681=>"001000010",
  52682=>"101111111",
  52683=>"011000111",
  52684=>"001110000",
  52685=>"010110100",
  52686=>"101000110",
  52687=>"000000110",
  52688=>"111011010",
  52689=>"001011010",
  52690=>"011010011",
  52691=>"110010011",
  52692=>"111000011",
  52693=>"101001110",
  52694=>"000110001",
  52695=>"010000110",
  52696=>"110110110",
  52697=>"011110010",
  52698=>"000011110",
  52699=>"110010001",
  52700=>"111111111",
  52701=>"111101010",
  52702=>"000101101",
  52703=>"111101110",
  52704=>"101111000",
  52705=>"111010010",
  52706=>"111110100",
  52707=>"110111110",
  52708=>"100001000",
  52709=>"010110010",
  52710=>"011100101",
  52711=>"101010100",
  52712=>"101101000",
  52713=>"001111001",
  52714=>"000010010",
  52715=>"000000011",
  52716=>"101000001",
  52717=>"111000111",
  52718=>"111100011",
  52719=>"000010110",
  52720=>"110011000",
  52721=>"111010011",
  52722=>"110101000",
  52723=>"110110001",
  52724=>"111101101",
  52725=>"010101001",
  52726=>"100000001",
  52727=>"100101000",
  52728=>"110110000",
  52729=>"010111011",
  52730=>"001000010",
  52731=>"001000111",
  52732=>"101101000",
  52733=>"100101101",
  52734=>"100011111",
  52735=>"101100011",
  52736=>"111011000",
  52737=>"110110001",
  52738=>"100101001",
  52739=>"111001111",
  52740=>"111111011",
  52741=>"011010001",
  52742=>"001010001",
  52743=>"001110110",
  52744=>"011101000",
  52745=>"111000010",
  52746=>"000000100",
  52747=>"101011110",
  52748=>"101100111",
  52749=>"101101110",
  52750=>"000001001",
  52751=>"101111011",
  52752=>"000010101",
  52753=>"100100110",
  52754=>"110001100",
  52755=>"001111101",
  52756=>"001001000",
  52757=>"101110001",
  52758=>"110000110",
  52759=>"111001001",
  52760=>"000010010",
  52761=>"000010000",
  52762=>"110011100",
  52763=>"101001011",
  52764=>"110100000",
  52765=>"110110011",
  52766=>"111001110",
  52767=>"111100101",
  52768=>"000010011",
  52769=>"111011011",
  52770=>"000001010",
  52771=>"110011101",
  52772=>"011110100",
  52773=>"000001001",
  52774=>"010100010",
  52775=>"110111011",
  52776=>"101011000",
  52777=>"111110011",
  52778=>"111110001",
  52779=>"110011011",
  52780=>"001000110",
  52781=>"011000001",
  52782=>"001000110",
  52783=>"000010010",
  52784=>"110110100",
  52785=>"100001001",
  52786=>"111001010",
  52787=>"110101011",
  52788=>"001100111",
  52789=>"111011000",
  52790=>"001111111",
  52791=>"101000011",
  52792=>"010100110",
  52793=>"000110000",
  52794=>"001001001",
  52795=>"011100111",
  52796=>"111111010",
  52797=>"101010110",
  52798=>"011001011",
  52799=>"110111001",
  52800=>"010101000",
  52801=>"101001111",
  52802=>"000100011",
  52803=>"100111101",
  52804=>"111111100",
  52805=>"001010100",
  52806=>"110000101",
  52807=>"001111100",
  52808=>"101010011",
  52809=>"000100111",
  52810=>"001110101",
  52811=>"000100111",
  52812=>"101111011",
  52813=>"001100001",
  52814=>"101000101",
  52815=>"010111101",
  52816=>"001000000",
  52817=>"010000100",
  52818=>"110010010",
  52819=>"001111110",
  52820=>"101001100",
  52821=>"110001011",
  52822=>"110111000",
  52823=>"000100001",
  52824=>"111111010",
  52825=>"100111000",
  52826=>"010100010",
  52827=>"101100101",
  52828=>"000100010",
  52829=>"001100101",
  52830=>"111011100",
  52831=>"010100011",
  52832=>"111111000",
  52833=>"001010001",
  52834=>"001001000",
  52835=>"111010000",
  52836=>"011101111",
  52837=>"011110101",
  52838=>"101110101",
  52839=>"000010110",
  52840=>"111001011",
  52841=>"001101101",
  52842=>"110111100",
  52843=>"100110100",
  52844=>"000001101",
  52845=>"111110000",
  52846=>"100011011",
  52847=>"101111110",
  52848=>"010110111",
  52849=>"110000100",
  52850=>"010001100",
  52851=>"010100100",
  52852=>"011110011",
  52853=>"110001100",
  52854=>"010001110",
  52855=>"010011101",
  52856=>"010110110",
  52857=>"100100110",
  52858=>"111110001",
  52859=>"010101010",
  52860=>"010001100",
  52861=>"100001101",
  52862=>"001101001",
  52863=>"111000111",
  52864=>"010011011",
  52865=>"000101110",
  52866=>"001001011",
  52867=>"101101111",
  52868=>"001101000",
  52869=>"010000000",
  52870=>"001000011",
  52871=>"111011100",
  52872=>"110110111",
  52873=>"001000110",
  52874=>"001110101",
  52875=>"101110100",
  52876=>"010011100",
  52877=>"010110011",
  52878=>"101011011",
  52879=>"110110000",
  52880=>"110000111",
  52881=>"101100111",
  52882=>"111110100",
  52883=>"000101110",
  52884=>"111010010",
  52885=>"101000111",
  52886=>"110010000",
  52887=>"001011100",
  52888=>"110101111",
  52889=>"001000001",
  52890=>"001001011",
  52891=>"110010110",
  52892=>"100001001",
  52893=>"100000001",
  52894=>"000101010",
  52895=>"000110010",
  52896=>"010111010",
  52897=>"000001000",
  52898=>"001101111",
  52899=>"100000101",
  52900=>"011000100",
  52901=>"011100000",
  52902=>"010111000",
  52903=>"111001011",
  52904=>"000110000",
  52905=>"110010111",
  52906=>"010001111",
  52907=>"000001000",
  52908=>"010111111",
  52909=>"101100111",
  52910=>"111111001",
  52911=>"101011001",
  52912=>"000001000",
  52913=>"001010100",
  52914=>"110001010",
  52915=>"001110010",
  52916=>"100110100",
  52917=>"101001011",
  52918=>"011010010",
  52919=>"011010111",
  52920=>"000001001",
  52921=>"110110101",
  52922=>"001010000",
  52923=>"011000010",
  52924=>"111110100",
  52925=>"001100101",
  52926=>"010011011",
  52927=>"001100110",
  52928=>"011111011",
  52929=>"000011110",
  52930=>"000000100",
  52931=>"010011111",
  52932=>"010011110",
  52933=>"000010011",
  52934=>"110110100",
  52935=>"111001110",
  52936=>"011000010",
  52937=>"100111010",
  52938=>"011000111",
  52939=>"110100100",
  52940=>"111111101",
  52941=>"100001000",
  52942=>"101001011",
  52943=>"000111010",
  52944=>"010100011",
  52945=>"011110010",
  52946=>"011001111",
  52947=>"100110101",
  52948=>"000110111",
  52949=>"100010111",
  52950=>"000111000",
  52951=>"000011100",
  52952=>"000000100",
  52953=>"010101100",
  52954=>"111100001",
  52955=>"100010011",
  52956=>"100101111",
  52957=>"011100101",
  52958=>"100100010",
  52959=>"110111111",
  52960=>"111101100",
  52961=>"010010111",
  52962=>"010100111",
  52963=>"001000010",
  52964=>"110110100",
  52965=>"011000011",
  52966=>"111001101",
  52967=>"101000100",
  52968=>"110100110",
  52969=>"010101011",
  52970=>"100101111",
  52971=>"001101110",
  52972=>"111110100",
  52973=>"101000101",
  52974=>"010110100",
  52975=>"000101010",
  52976=>"000111101",
  52977=>"011101101",
  52978=>"011000000",
  52979=>"100010100",
  52980=>"001001001",
  52981=>"100010000",
  52982=>"000111100",
  52983=>"010010001",
  52984=>"001101010",
  52985=>"011111001",
  52986=>"011100010",
  52987=>"110111111",
  52988=>"110011101",
  52989=>"110000010",
  52990=>"101100010",
  52991=>"101101101",
  52992=>"101000111",
  52993=>"000100000",
  52994=>"110111000",
  52995=>"001011110",
  52996=>"100010111",
  52997=>"000111011",
  52998=>"000000110",
  52999=>"001011000",
  53000=>"010010010",
  53001=>"011110101",
  53002=>"100010100",
  53003=>"010101101",
  53004=>"011010000",
  53005=>"010111011",
  53006=>"110101000",
  53007=>"100101000",
  53008=>"000001101",
  53009=>"000010110",
  53010=>"011011101",
  53011=>"000010101",
  53012=>"010111101",
  53013=>"010101011",
  53014=>"100111100",
  53015=>"011110110",
  53016=>"000010010",
  53017=>"111010001",
  53018=>"100101111",
  53019=>"010011100",
  53020=>"101111111",
  53021=>"111100100",
  53022=>"010001011",
  53023=>"000110111",
  53024=>"000100101",
  53025=>"110101001",
  53026=>"111111101",
  53027=>"010101100",
  53028=>"110010000",
  53029=>"001100001",
  53030=>"010111011",
  53031=>"001011100",
  53032=>"101001100",
  53033=>"110101111",
  53034=>"001001011",
  53035=>"101010001",
  53036=>"100110101",
  53037=>"111101011",
  53038=>"110000110",
  53039=>"000010001",
  53040=>"110100010",
  53041=>"111110111",
  53042=>"001100000",
  53043=>"011011111",
  53044=>"000100010",
  53045=>"111000010",
  53046=>"111101111",
  53047=>"100001110",
  53048=>"100001100",
  53049=>"110000001",
  53050=>"101011111",
  53051=>"011000000",
  53052=>"100111001",
  53053=>"101100001",
  53054=>"001111001",
  53055=>"111111101",
  53056=>"101010010",
  53057=>"011011011",
  53058=>"111001101",
  53059=>"001000101",
  53060=>"110111111",
  53061=>"000110101",
  53062=>"010000100",
  53063=>"001111110",
  53064=>"100010111",
  53065=>"101101100",
  53066=>"010110100",
  53067=>"001011101",
  53068=>"010010001",
  53069=>"110011000",
  53070=>"111110101",
  53071=>"100001000",
  53072=>"001001101",
  53073=>"110000000",
  53074=>"000010000",
  53075=>"001011000",
  53076=>"110001010",
  53077=>"010110100",
  53078=>"000000010",
  53079=>"011011101",
  53080=>"111101111",
  53081=>"110000111",
  53082=>"001110010",
  53083=>"110001001",
  53084=>"011000011",
  53085=>"110111101",
  53086=>"001000001",
  53087=>"011000110",
  53088=>"110001110",
  53089=>"010000101",
  53090=>"011110101",
  53091=>"010100011",
  53092=>"000100000",
  53093=>"101001101",
  53094=>"111111000",
  53095=>"001111000",
  53096=>"100011100",
  53097=>"110011010",
  53098=>"110101110",
  53099=>"000001011",
  53100=>"000000010",
  53101=>"010010010",
  53102=>"100110011",
  53103=>"110011000",
  53104=>"111011010",
  53105=>"100101111",
  53106=>"010101111",
  53107=>"111110011",
  53108=>"001110100",
  53109=>"000100000",
  53110=>"111110101",
  53111=>"011011111",
  53112=>"001010110",
  53113=>"000011100",
  53114=>"110110110",
  53115=>"111001100",
  53116=>"011101010",
  53117=>"100100000",
  53118=>"010000100",
  53119=>"111110100",
  53120=>"111110110",
  53121=>"011100111",
  53122=>"000010111",
  53123=>"111000010",
  53124=>"011101111",
  53125=>"110111001",
  53126=>"001000110",
  53127=>"000000000",
  53128=>"000101001",
  53129=>"011111110",
  53130=>"110100111",
  53131=>"101000001",
  53132=>"111111001",
  53133=>"011011011",
  53134=>"100001011",
  53135=>"010111000",
  53136=>"011110111",
  53137=>"001100111",
  53138=>"100100001",
  53139=>"100000101",
  53140=>"011010110",
  53141=>"010111010",
  53142=>"010001010",
  53143=>"100100000",
  53144=>"111110000",
  53145=>"110001100",
  53146=>"101010001",
  53147=>"111100011",
  53148=>"010110100",
  53149=>"100111110",
  53150=>"001001111",
  53151=>"101111010",
  53152=>"011101011",
  53153=>"110011001",
  53154=>"110111100",
  53155=>"011110110",
  53156=>"010100010",
  53157=>"100001011",
  53158=>"110011010",
  53159=>"001111000",
  53160=>"111001111",
  53161=>"011011011",
  53162=>"110001000",
  53163=>"100101110",
  53164=>"000001000",
  53165=>"110000111",
  53166=>"000000110",
  53167=>"101111000",
  53168=>"111100111",
  53169=>"100011101",
  53170=>"011010111",
  53171=>"110011110",
  53172=>"011010010",
  53173=>"110111111",
  53174=>"110111110",
  53175=>"010111110",
  53176=>"000011000",
  53177=>"011101100",
  53178=>"101110100",
  53179=>"100100101",
  53180=>"011000111",
  53181=>"011100001",
  53182=>"100110110",
  53183=>"011101111",
  53184=>"100110101",
  53185=>"100000000",
  53186=>"111101101",
  53187=>"011111001",
  53188=>"001110001",
  53189=>"111101101",
  53190=>"111011110",
  53191=>"011101111",
  53192=>"110001000",
  53193=>"110011001",
  53194=>"100010110",
  53195=>"100100111",
  53196=>"000110100",
  53197=>"100101100",
  53198=>"010110100",
  53199=>"011100100",
  53200=>"100111111",
  53201=>"011111110",
  53202=>"111010110",
  53203=>"101111011",
  53204=>"100001000",
  53205=>"000001100",
  53206=>"000010110",
  53207=>"010011001",
  53208=>"111110110",
  53209=>"011011001",
  53210=>"000110011",
  53211=>"100001010",
  53212=>"001100110",
  53213=>"011100001",
  53214=>"100111111",
  53215=>"010010110",
  53216=>"001100101",
  53217=>"111000110",
  53218=>"010101001",
  53219=>"000010111",
  53220=>"000000011",
  53221=>"000011110",
  53222=>"001010111",
  53223=>"011101011",
  53224=>"010100001",
  53225=>"100111110",
  53226=>"110111010",
  53227=>"110100111",
  53228=>"010010111",
  53229=>"011101010",
  53230=>"011011111",
  53231=>"001111100",
  53232=>"010000011",
  53233=>"011101110",
  53234=>"001110110",
  53235=>"001110110",
  53236=>"111001110",
  53237=>"111000001",
  53238=>"100011100",
  53239=>"001111111",
  53240=>"111110111",
  53241=>"101111101",
  53242=>"011000011",
  53243=>"001001110",
  53244=>"111001011",
  53245=>"000100110",
  53246=>"100000011",
  53247=>"111000010",
  53248=>"011111100",
  53249=>"010011000",
  53250=>"100101000",
  53251=>"011111110",
  53252=>"001100011",
  53253=>"110010100",
  53254=>"001010001",
  53255=>"110101111",
  53256=>"111110100",
  53257=>"001100101",
  53258=>"111100100",
  53259=>"010010100",
  53260=>"000010010",
  53261=>"000001111",
  53262=>"110111000",
  53263=>"011010101",
  53264=>"000000001",
  53265=>"101110110",
  53266=>"110111010",
  53267=>"011010111",
  53268=>"000110110",
  53269=>"111101100",
  53270=>"100011000",
  53271=>"000100100",
  53272=>"001011000",
  53273=>"000110100",
  53274=>"100100101",
  53275=>"100100110",
  53276=>"110111110",
  53277=>"000110010",
  53278=>"010010110",
  53279=>"111101010",
  53280=>"110111001",
  53281=>"100110011",
  53282=>"100111110",
  53283=>"011111111",
  53284=>"011110011",
  53285=>"000000000",
  53286=>"000011010",
  53287=>"011011011",
  53288=>"011111001",
  53289=>"100101101",
  53290=>"110011001",
  53291=>"011110010",
  53292=>"110101001",
  53293=>"001110101",
  53294=>"100001000",
  53295=>"011110111",
  53296=>"111101011",
  53297=>"011000011",
  53298=>"110100011",
  53299=>"111001101",
  53300=>"100101000",
  53301=>"101101011",
  53302=>"001010101",
  53303=>"001001110",
  53304=>"001111110",
  53305=>"010010000",
  53306=>"000111111",
  53307=>"001010110",
  53308=>"101011000",
  53309=>"101101000",
  53310=>"001101010",
  53311=>"010111010",
  53312=>"100010111",
  53313=>"010100011",
  53314=>"011100010",
  53315=>"101001100",
  53316=>"101111111",
  53317=>"000110111",
  53318=>"010110011",
  53319=>"111000010",
  53320=>"101101100",
  53321=>"011110000",
  53322=>"110001010",
  53323=>"011010011",
  53324=>"100011001",
  53325=>"110000001",
  53326=>"011101110",
  53327=>"010111110",
  53328=>"000001000",
  53329=>"111000111",
  53330=>"000100101",
  53331=>"101110000",
  53332=>"011111011",
  53333=>"111100111",
  53334=>"111101001",
  53335=>"000101001",
  53336=>"000010100",
  53337=>"100001110",
  53338=>"110101110",
  53339=>"100111111",
  53340=>"001110100",
  53341=>"101001011",
  53342=>"011000011",
  53343=>"000011111",
  53344=>"111100000",
  53345=>"111100001",
  53346=>"101000010",
  53347=>"001101100",
  53348=>"101100101",
  53349=>"010010110",
  53350=>"001001000",
  53351=>"000110011",
  53352=>"111010111",
  53353=>"110111010",
  53354=>"001111111",
  53355=>"110010111",
  53356=>"001111000",
  53357=>"100001101",
  53358=>"110000101",
  53359=>"110111111",
  53360=>"000110000",
  53361=>"011100011",
  53362=>"001111111",
  53363=>"111011011",
  53364=>"101000001",
  53365=>"100010010",
  53366=>"111111000",
  53367=>"000101011",
  53368=>"110111110",
  53369=>"010010000",
  53370=>"110111010",
  53371=>"101101110",
  53372=>"010110100",
  53373=>"011000100",
  53374=>"000000011",
  53375=>"011001111",
  53376=>"011010101",
  53377=>"001110100",
  53378=>"000010100",
  53379=>"010011111",
  53380=>"010101100",
  53381=>"101001111",
  53382=>"010011110",
  53383=>"110100100",
  53384=>"011011000",
  53385=>"001100010",
  53386=>"110101110",
  53387=>"010010011",
  53388=>"110100000",
  53389=>"000001001",
  53390=>"110101110",
  53391=>"111101100",
  53392=>"000010101",
  53393=>"010001111",
  53394=>"011010001",
  53395=>"000001111",
  53396=>"001011110",
  53397=>"000001110",
  53398=>"001000000",
  53399=>"010101110",
  53400=>"100010110",
  53401=>"100000001",
  53402=>"010101000",
  53403=>"111010101",
  53404=>"000011000",
  53405=>"101000001",
  53406=>"011001010",
  53407=>"101111010",
  53408=>"111111000",
  53409=>"011010100",
  53410=>"000100010",
  53411=>"010100010",
  53412=>"011000001",
  53413=>"110000100",
  53414=>"000000010",
  53415=>"101000111",
  53416=>"101111111",
  53417=>"000100111",
  53418=>"001010000",
  53419=>"110010101",
  53420=>"001010111",
  53421=>"100110100",
  53422=>"100110001",
  53423=>"100001010",
  53424=>"001100011",
  53425=>"011100000",
  53426=>"000110001",
  53427=>"101101000",
  53428=>"000011111",
  53429=>"000011110",
  53430=>"110001010",
  53431=>"001010000",
  53432=>"001100000",
  53433=>"011111011",
  53434=>"001000000",
  53435=>"110110110",
  53436=>"110100101",
  53437=>"001001110",
  53438=>"000010011",
  53439=>"111100001",
  53440=>"100111010",
  53441=>"010010110",
  53442=>"000011100",
  53443=>"000000011",
  53444=>"111101011",
  53445=>"111110111",
  53446=>"101111011",
  53447=>"010010000",
  53448=>"011100011",
  53449=>"101100111",
  53450=>"101100101",
  53451=>"110101101",
  53452=>"101100010",
  53453=>"000000111",
  53454=>"000000000",
  53455=>"011011010",
  53456=>"001110000",
  53457=>"111101101",
  53458=>"001011101",
  53459=>"100110100",
  53460=>"000100010",
  53461=>"111110100",
  53462=>"000111010",
  53463=>"110101010",
  53464=>"000010110",
  53465=>"100000000",
  53466=>"110110001",
  53467=>"000000000",
  53468=>"011111010",
  53469=>"100001110",
  53470=>"001001111",
  53471=>"000011101",
  53472=>"111001011",
  53473=>"000111000",
  53474=>"001101000",
  53475=>"011101010",
  53476=>"010011101",
  53477=>"100110100",
  53478=>"000100101",
  53479=>"011110010",
  53480=>"110101100",
  53481=>"101100001",
  53482=>"111000000",
  53483=>"100101110",
  53484=>"111111010",
  53485=>"111010111",
  53486=>"011000100",
  53487=>"010011000",
  53488=>"110001110",
  53489=>"011111110",
  53490=>"100110100",
  53491=>"100000000",
  53492=>"101000100",
  53493=>"101010110",
  53494=>"111101101",
  53495=>"100000001",
  53496=>"100110100",
  53497=>"011010001",
  53498=>"111100001",
  53499=>"110101101",
  53500=>"011011110",
  53501=>"000100101",
  53502=>"000001100",
  53503=>"100000100",
  53504=>"111111110",
  53505=>"010111100",
  53506=>"110110110",
  53507=>"101110011",
  53508=>"011110000",
  53509=>"100110111",
  53510=>"000001001",
  53511=>"001010001",
  53512=>"110110000",
  53513=>"001100010",
  53514=>"010001111",
  53515=>"110101110",
  53516=>"100011110",
  53517=>"111001001",
  53518=>"100011111",
  53519=>"101110011",
  53520=>"010010010",
  53521=>"101011001",
  53522=>"110000000",
  53523=>"011110001",
  53524=>"000110000",
  53525=>"010000011",
  53526=>"000101101",
  53527=>"001111001",
  53528=>"111100001",
  53529=>"011001000",
  53530=>"011010111",
  53531=>"110100000",
  53532=>"111001001",
  53533=>"110101000",
  53534=>"100001110",
  53535=>"010010100",
  53536=>"001110010",
  53537=>"100011101",
  53538=>"000100001",
  53539=>"000100100",
  53540=>"100001110",
  53541=>"110100110",
  53542=>"101111000",
  53543=>"111111011",
  53544=>"000100010",
  53545=>"010111100",
  53546=>"000100010",
  53547=>"010110001",
  53548=>"001110011",
  53549=>"100001011",
  53550=>"001101100",
  53551=>"001111101",
  53552=>"111101000",
  53553=>"011000100",
  53554=>"111000001",
  53555=>"010010001",
  53556=>"111110011",
  53557=>"011001100",
  53558=>"000111110",
  53559=>"001111100",
  53560=>"000000011",
  53561=>"000001000",
  53562=>"011100101",
  53563=>"010101011",
  53564=>"010011111",
  53565=>"101101111",
  53566=>"101101111",
  53567=>"110100111",
  53568=>"001011010",
  53569=>"101000000",
  53570=>"110110000",
  53571=>"000000110",
  53572=>"111101110",
  53573=>"110010111",
  53574=>"011111110",
  53575=>"010011010",
  53576=>"001001011",
  53577=>"010101101",
  53578=>"101101010",
  53579=>"111110101",
  53580=>"100010001",
  53581=>"001011010",
  53582=>"111111111",
  53583=>"011111001",
  53584=>"111111101",
  53585=>"101100010",
  53586=>"011010010",
  53587=>"110101001",
  53588=>"110101001",
  53589=>"010100010",
  53590=>"001110001",
  53591=>"000000001",
  53592=>"101010101",
  53593=>"010001111",
  53594=>"011000001",
  53595=>"100000100",
  53596=>"100000110",
  53597=>"110110000",
  53598=>"110111111",
  53599=>"010001110",
  53600=>"101110101",
  53601=>"010001000",
  53602=>"110101101",
  53603=>"010101011",
  53604=>"001000000",
  53605=>"001110111",
  53606=>"011001111",
  53607=>"011100001",
  53608=>"100010100",
  53609=>"001100111",
  53610=>"110100010",
  53611=>"100010000",
  53612=>"100111010",
  53613=>"111100111",
  53614=>"100101011",
  53615=>"011100101",
  53616=>"100100000",
  53617=>"110011101",
  53618=>"000110100",
  53619=>"111100001",
  53620=>"011110111",
  53621=>"000010010",
  53622=>"011110000",
  53623=>"011000111",
  53624=>"011010010",
  53625=>"100101101",
  53626=>"100011010",
  53627=>"101110010",
  53628=>"110100101",
  53629=>"110010101",
  53630=>"001010001",
  53631=>"111001100",
  53632=>"000110100",
  53633=>"010011101",
  53634=>"001001110",
  53635=>"000000100",
  53636=>"001110110",
  53637=>"110000001",
  53638=>"110101011",
  53639=>"111011100",
  53640=>"001011101",
  53641=>"111011110",
  53642=>"001010001",
  53643=>"010001001",
  53644=>"110001101",
  53645=>"010101011",
  53646=>"011010101",
  53647=>"001111011",
  53648=>"001111001",
  53649=>"100010110",
  53650=>"010100110",
  53651=>"001001101",
  53652=>"100101100",
  53653=>"000001001",
  53654=>"011010001",
  53655=>"001011001",
  53656=>"100000001",
  53657=>"101000010",
  53658=>"100000100",
  53659=>"001001001",
  53660=>"100001001",
  53661=>"011101010",
  53662=>"000111001",
  53663=>"111100001",
  53664=>"111110011",
  53665=>"010000000",
  53666=>"000101101",
  53667=>"000011111",
  53668=>"000101100",
  53669=>"011011011",
  53670=>"110000100",
  53671=>"010100011",
  53672=>"011111101",
  53673=>"001000011",
  53674=>"101011011",
  53675=>"001100110",
  53676=>"000111101",
  53677=>"011110000",
  53678=>"010110110",
  53679=>"101101100",
  53680=>"110010011",
  53681=>"100101101",
  53682=>"110000101",
  53683=>"000010101",
  53684=>"110000101",
  53685=>"101111100",
  53686=>"010001101",
  53687=>"001011000",
  53688=>"111111011",
  53689=>"110000011",
  53690=>"000010100",
  53691=>"001110000",
  53692=>"110000100",
  53693=>"011110001",
  53694=>"010000010",
  53695=>"011110010",
  53696=>"001111111",
  53697=>"100110101",
  53698=>"001010101",
  53699=>"110011000",
  53700=>"000100010",
  53701=>"000101011",
  53702=>"001000110",
  53703=>"110000000",
  53704=>"010001101",
  53705=>"000110000",
  53706=>"000110110",
  53707=>"000110110",
  53708=>"000001101",
  53709=>"100010001",
  53710=>"111101111",
  53711=>"100011100",
  53712=>"110000110",
  53713=>"100100100",
  53714=>"100001101",
  53715=>"011010001",
  53716=>"011111011",
  53717=>"100000110",
  53718=>"100010001",
  53719=>"000011001",
  53720=>"000101111",
  53721=>"110001000",
  53722=>"111100100",
  53723=>"111010110",
  53724=>"101000001",
  53725=>"110011001",
  53726=>"100110001",
  53727=>"001111000",
  53728=>"101110100",
  53729=>"000101111",
  53730=>"011101010",
  53731=>"111111111",
  53732=>"011000110",
  53733=>"010110110",
  53734=>"101001111",
  53735=>"000001111",
  53736=>"000010010",
  53737=>"111101110",
  53738=>"111000011",
  53739=>"011001101",
  53740=>"000000101",
  53741=>"111101110",
  53742=>"101001111",
  53743=>"001000110",
  53744=>"010100101",
  53745=>"000110001",
  53746=>"110000111",
  53747=>"110000010",
  53748=>"100010100",
  53749=>"000010010",
  53750=>"011010110",
  53751=>"100010100",
  53752=>"101101001",
  53753=>"010110011",
  53754=>"000101010",
  53755=>"101101001",
  53756=>"100000110",
  53757=>"010100001",
  53758=>"111111110",
  53759=>"100100111",
  53760=>"001011010",
  53761=>"101010101",
  53762=>"111100010",
  53763=>"100101011",
  53764=>"001111001",
  53765=>"111101010",
  53766=>"101110111",
  53767=>"101101011",
  53768=>"011100100",
  53769=>"110111010",
  53770=>"110100000",
  53771=>"111011111",
  53772=>"110001101",
  53773=>"011100101",
  53774=>"000001011",
  53775=>"000100010",
  53776=>"000000101",
  53777=>"001000011",
  53778=>"001000100",
  53779=>"111011110",
  53780=>"011000000",
  53781=>"000011101",
  53782=>"100011101",
  53783=>"100000110",
  53784=>"110000101",
  53785=>"001011001",
  53786=>"000010001",
  53787=>"101100111",
  53788=>"101001001",
  53789=>"100110101",
  53790=>"100110010",
  53791=>"101001001",
  53792=>"010000010",
  53793=>"010001000",
  53794=>"010110000",
  53795=>"101000001",
  53796=>"011000001",
  53797=>"010000011",
  53798=>"111010101",
  53799=>"010110000",
  53800=>"110111100",
  53801=>"010101111",
  53802=>"001101001",
  53803=>"001100010",
  53804=>"011010011",
  53805=>"011110111",
  53806=>"011000001",
  53807=>"101001110",
  53808=>"100101101",
  53809=>"111010011",
  53810=>"110011110",
  53811=>"000100010",
  53812=>"000000110",
  53813=>"101110001",
  53814=>"110000001",
  53815=>"001010010",
  53816=>"001000010",
  53817=>"100010001",
  53818=>"101111000",
  53819=>"001101010",
  53820=>"101010110",
  53821=>"100010100",
  53822=>"100111101",
  53823=>"111101001",
  53824=>"111101110",
  53825=>"001000111",
  53826=>"111110000",
  53827=>"111100010",
  53828=>"110000000",
  53829=>"000111001",
  53830=>"001101001",
  53831=>"001100111",
  53832=>"011110101",
  53833=>"001010011",
  53834=>"110101111",
  53835=>"100001110",
  53836=>"110001101",
  53837=>"001101111",
  53838=>"000101100",
  53839=>"111101101",
  53840=>"100101001",
  53841=>"100001001",
  53842=>"000011001",
  53843=>"110110100",
  53844=>"000110001",
  53845=>"110010001",
  53846=>"101101100",
  53847=>"010011110",
  53848=>"011001010",
  53849=>"011111100",
  53850=>"000100111",
  53851=>"111000111",
  53852=>"010101001",
  53853=>"010010101",
  53854=>"101111011",
  53855=>"110010000",
  53856=>"010010001",
  53857=>"000010011",
  53858=>"101110001",
  53859=>"000110011",
  53860=>"000010000",
  53861=>"001001000",
  53862=>"000011001",
  53863=>"111111101",
  53864=>"000010100",
  53865=>"000111010",
  53866=>"011101110",
  53867=>"100011111",
  53868=>"100111000",
  53869=>"111010110",
  53870=>"001110111",
  53871=>"000001000",
  53872=>"000000001",
  53873=>"000000011",
  53874=>"011000000",
  53875=>"011000011",
  53876=>"001111100",
  53877=>"000001110",
  53878=>"000100110",
  53879=>"110001010",
  53880=>"010011100",
  53881=>"000000101",
  53882=>"111001011",
  53883=>"110110000",
  53884=>"100000001",
  53885=>"001010011",
  53886=>"100110110",
  53887=>"000010111",
  53888=>"110100110",
  53889=>"110000110",
  53890=>"011010001",
  53891=>"101001100",
  53892=>"111001010",
  53893=>"011010010",
  53894=>"100111000",
  53895=>"010110100",
  53896=>"010001100",
  53897=>"010000110",
  53898=>"101011001",
  53899=>"010110010",
  53900=>"111101110",
  53901=>"110000100",
  53902=>"110001101",
  53903=>"100000110",
  53904=>"111100001",
  53905=>"100111000",
  53906=>"111101110",
  53907=>"001000000",
  53908=>"101111100",
  53909=>"111010100",
  53910=>"100001111",
  53911=>"011110100",
  53912=>"111101000",
  53913=>"100010011",
  53914=>"110100101",
  53915=>"110010110",
  53916=>"011011110",
  53917=>"010110000",
  53918=>"001010000",
  53919=>"111101110",
  53920=>"011111110",
  53921=>"001111011",
  53922=>"001011010",
  53923=>"000001001",
  53924=>"001100011",
  53925=>"011001011",
  53926=>"110000011",
  53927=>"001100000",
  53928=>"110111001",
  53929=>"000110011",
  53930=>"000000011",
  53931=>"111100110",
  53932=>"100100100",
  53933=>"000110100",
  53934=>"010111110",
  53935=>"110100011",
  53936=>"011101110",
  53937=>"010011111",
  53938=>"101000101",
  53939=>"100110000",
  53940=>"000101011",
  53941=>"011011111",
  53942=>"010100100",
  53943=>"001010000",
  53944=>"010011110",
  53945=>"111010100",
  53946=>"000001010",
  53947=>"001100001",
  53948=>"001100110",
  53949=>"100001010",
  53950=>"101101000",
  53951=>"100000100",
  53952=>"001110001",
  53953=>"101001100",
  53954=>"110001001",
  53955=>"000111101",
  53956=>"001000101",
  53957=>"000110010",
  53958=>"101111111",
  53959=>"111010010",
  53960=>"110100001",
  53961=>"001001100",
  53962=>"111000000",
  53963=>"011011110",
  53964=>"010011101",
  53965=>"000111110",
  53966=>"111100110",
  53967=>"000111111",
  53968=>"010010000",
  53969=>"011010001",
  53970=>"100110101",
  53971=>"011010100",
  53972=>"111011101",
  53973=>"011100001",
  53974=>"111011000",
  53975=>"011100101",
  53976=>"100100110",
  53977=>"110010001",
  53978=>"111101010",
  53979=>"110111000",
  53980=>"001101111",
  53981=>"111101101",
  53982=>"011111110",
  53983=>"000001100",
  53984=>"111000000",
  53985=>"100000110",
  53986=>"010010000",
  53987=>"001111001",
  53988=>"011001110",
  53989=>"101000000",
  53990=>"001011101",
  53991=>"101100111",
  53992=>"100100101",
  53993=>"011101000",
  53994=>"000100101",
  53995=>"000010010",
  53996=>"010010111",
  53997=>"011011110",
  53998=>"011000100",
  53999=>"001010100",
  54000=>"101001011",
  54001=>"111010000",
  54002=>"001001011",
  54003=>"100000010",
  54004=>"100101011",
  54005=>"111111001",
  54006=>"001010000",
  54007=>"001100111",
  54008=>"110001101",
  54009=>"011100100",
  54010=>"000010100",
  54011=>"000110100",
  54012=>"111000000",
  54013=>"100101000",
  54014=>"001101011",
  54015=>"011001011",
  54016=>"001101101",
  54017=>"100100010",
  54018=>"000101110",
  54019=>"010101011",
  54020=>"011101110",
  54021=>"101000000",
  54022=>"010010000",
  54023=>"111011000",
  54024=>"100000100",
  54025=>"010011110",
  54026=>"111000011",
  54027=>"010010000",
  54028=>"001100000",
  54029=>"000111100",
  54030=>"100101111",
  54031=>"001111011",
  54032=>"100000000",
  54033=>"010001000",
  54034=>"010001110",
  54035=>"110010011",
  54036=>"111001100",
  54037=>"000110010",
  54038=>"110000011",
  54039=>"001011001",
  54040=>"110010111",
  54041=>"011100100",
  54042=>"001010001",
  54043=>"100000100",
  54044=>"111111001",
  54045=>"111110100",
  54046=>"100100110",
  54047=>"001100100",
  54048=>"001111110",
  54049=>"100010010",
  54050=>"100111100",
  54051=>"110111010",
  54052=>"110101001",
  54053=>"100100010",
  54054=>"111110000",
  54055=>"110000000",
  54056=>"101010110",
  54057=>"010000101",
  54058=>"000011101",
  54059=>"100000111",
  54060=>"000001110",
  54061=>"000100010",
  54062=>"100101110",
  54063=>"011010001",
  54064=>"000101000",
  54065=>"100001010",
  54066=>"010011011",
  54067=>"101011110",
  54068=>"110101101",
  54069=>"110101101",
  54070=>"011000010",
  54071=>"100010001",
  54072=>"100110110",
  54073=>"101101001",
  54074=>"101100001",
  54075=>"010011001",
  54076=>"000111001",
  54077=>"010111001",
  54078=>"110001101",
  54079=>"011011001",
  54080=>"001001011",
  54081=>"101010001",
  54082=>"010110001",
  54083=>"011010010",
  54084=>"010110111",
  54085=>"000101000",
  54086=>"101000010",
  54087=>"001011011",
  54088=>"100101100",
  54089=>"110101000",
  54090=>"001000010",
  54091=>"001111010",
  54092=>"001011000",
  54093=>"000001000",
  54094=>"010111011",
  54095=>"110111001",
  54096=>"111011101",
  54097=>"100111001",
  54098=>"100100100",
  54099=>"011010000",
  54100=>"001111001",
  54101=>"001101001",
  54102=>"110011110",
  54103=>"001001000",
  54104=>"110000011",
  54105=>"100100000",
  54106=>"100101010",
  54107=>"001000101",
  54108=>"111001100",
  54109=>"000011011",
  54110=>"101100100",
  54111=>"001011100",
  54112=>"101100010",
  54113=>"111110110",
  54114=>"101101011",
  54115=>"011011010",
  54116=>"011011010",
  54117=>"000101110",
  54118=>"101001000",
  54119=>"011001011",
  54120=>"101010000",
  54121=>"000010000",
  54122=>"101000011",
  54123=>"110010010",
  54124=>"001110001",
  54125=>"001000001",
  54126=>"100000100",
  54127=>"101011100",
  54128=>"100010001",
  54129=>"110111000",
  54130=>"110111110",
  54131=>"011000110",
  54132=>"010000011",
  54133=>"000010111",
  54134=>"011110001",
  54135=>"011101010",
  54136=>"010001001",
  54137=>"000001001",
  54138=>"101001111",
  54139=>"100100011",
  54140=>"000000010",
  54141=>"101010010",
  54142=>"110110011",
  54143=>"110010011",
  54144=>"001001101",
  54145=>"001101111",
  54146=>"011001000",
  54147=>"100010010",
  54148=>"000101000",
  54149=>"011001101",
  54150=>"001100110",
  54151=>"111100011",
  54152=>"001011011",
  54153=>"110101101",
  54154=>"110110110",
  54155=>"100000010",
  54156=>"010011000",
  54157=>"000000111",
  54158=>"110000101",
  54159=>"010111100",
  54160=>"110010001",
  54161=>"011010101",
  54162=>"101100010",
  54163=>"111010010",
  54164=>"110010001",
  54165=>"011101101",
  54166=>"000001100",
  54167=>"011000100",
  54168=>"110101010",
  54169=>"110000100",
  54170=>"100001101",
  54171=>"001110100",
  54172=>"110010101",
  54173=>"111010110",
  54174=>"001011101",
  54175=>"000001110",
  54176=>"101111000",
  54177=>"010111011",
  54178=>"010010011",
  54179=>"111001110",
  54180=>"001010000",
  54181=>"000111110",
  54182=>"011011001",
  54183=>"110001111",
  54184=>"010100100",
  54185=>"010001001",
  54186=>"011010110",
  54187=>"111001010",
  54188=>"100101100",
  54189=>"100000010",
  54190=>"110000010",
  54191=>"011010010",
  54192=>"011011000",
  54193=>"000101101",
  54194=>"110111111",
  54195=>"101000110",
  54196=>"110001001",
  54197=>"110111111",
  54198=>"001011100",
  54199=>"000000000",
  54200=>"001100011",
  54201=>"000100100",
  54202=>"000101111",
  54203=>"111010110",
  54204=>"110001011",
  54205=>"100000101",
  54206=>"111011010",
  54207=>"000010000",
  54208=>"010011100",
  54209=>"010101100",
  54210=>"001111001",
  54211=>"110100110",
  54212=>"100110010",
  54213=>"001010011",
  54214=>"000000000",
  54215=>"001110111",
  54216=>"110011101",
  54217=>"100111010",
  54218=>"100111001",
  54219=>"010010011",
  54220=>"010111011",
  54221=>"110100000",
  54222=>"100010111",
  54223=>"101101100",
  54224=>"001101000",
  54225=>"100101110",
  54226=>"000110001",
  54227=>"000010011",
  54228=>"111010000",
  54229=>"101001001",
  54230=>"100101110",
  54231=>"011011111",
  54232=>"101001100",
  54233=>"110100011",
  54234=>"010101000",
  54235=>"001101001",
  54236=>"000001010",
  54237=>"010001000",
  54238=>"110011101",
  54239=>"001010000",
  54240=>"101011100",
  54241=>"000010101",
  54242=>"000111100",
  54243=>"110010101",
  54244=>"111000010",
  54245=>"111011010",
  54246=>"110111111",
  54247=>"000101100",
  54248=>"001000101",
  54249=>"001100111",
  54250=>"110011011",
  54251=>"110101110",
  54252=>"101110000",
  54253=>"000110000",
  54254=>"101111001",
  54255=>"010011100",
  54256=>"101001001",
  54257=>"110100110",
  54258=>"011011100",
  54259=>"010000001",
  54260=>"010000011",
  54261=>"010011101",
  54262=>"011001110",
  54263=>"011101000",
  54264=>"010011001",
  54265=>"011101101",
  54266=>"000100000",
  54267=>"001010010",
  54268=>"000100000",
  54269=>"011001111",
  54270=>"101000110",
  54271=>"011010110",
  54272=>"001000011",
  54273=>"011101110",
  54274=>"101001111",
  54275=>"111001100",
  54276=>"010011110",
  54277=>"101011111",
  54278=>"111111011",
  54279=>"010010100",
  54280=>"111000100",
  54281=>"111100011",
  54282=>"100000010",
  54283=>"110101011",
  54284=>"101100010",
  54285=>"101111011",
  54286=>"010001110",
  54287=>"111001001",
  54288=>"010010000",
  54289=>"000111101",
  54290=>"011111010",
  54291=>"011100000",
  54292=>"110011000",
  54293=>"010001110",
  54294=>"111110000",
  54295=>"111010110",
  54296=>"000000000",
  54297=>"010011001",
  54298=>"000100001",
  54299=>"010010110",
  54300=>"001101111",
  54301=>"110010110",
  54302=>"110001111",
  54303=>"100000011",
  54304=>"011101111",
  54305=>"100011001",
  54306=>"010100101",
  54307=>"101010111",
  54308=>"100001001",
  54309=>"111011010",
  54310=>"111110101",
  54311=>"000011010",
  54312=>"101000111",
  54313=>"100100011",
  54314=>"011011111",
  54315=>"000111010",
  54316=>"011000010",
  54317=>"101000010",
  54318=>"100000100",
  54319=>"110111100",
  54320=>"101110110",
  54321=>"011011000",
  54322=>"110011011",
  54323=>"000000000",
  54324=>"001001011",
  54325=>"000000100",
  54326=>"010111101",
  54327=>"110110111",
  54328=>"111000011",
  54329=>"100101001",
  54330=>"011110110",
  54331=>"001010110",
  54332=>"000000000",
  54333=>"100010000",
  54334=>"101101000",
  54335=>"100100101",
  54336=>"010101001",
  54337=>"100000000",
  54338=>"011111100",
  54339=>"000101000",
  54340=>"010101000",
  54341=>"000100001",
  54342=>"010100111",
  54343=>"001101000",
  54344=>"011011100",
  54345=>"010100010",
  54346=>"110001010",
  54347=>"001001111",
  54348=>"100010111",
  54349=>"110000110",
  54350=>"100101011",
  54351=>"100100001",
  54352=>"010011100",
  54353=>"111111100",
  54354=>"101001010",
  54355=>"001110110",
  54356=>"010010011",
  54357=>"010000110",
  54358=>"110110000",
  54359=>"100111000",
  54360=>"110011101",
  54361=>"101110010",
  54362=>"001010111",
  54363=>"010101001",
  54364=>"110100000",
  54365=>"100010100",
  54366=>"110001000",
  54367=>"100100001",
  54368=>"000110110",
  54369=>"001100101",
  54370=>"100101010",
  54371=>"100100111",
  54372=>"010011110",
  54373=>"000000000",
  54374=>"000000111",
  54375=>"100000110",
  54376=>"011001000",
  54377=>"100011101",
  54378=>"101000111",
  54379=>"001010100",
  54380=>"111110101",
  54381=>"111001110",
  54382=>"111101001",
  54383=>"011011011",
  54384=>"011110100",
  54385=>"101101011",
  54386=>"111111100",
  54387=>"111010010",
  54388=>"100101001",
  54389=>"111010010",
  54390=>"101101000",
  54391=>"110001011",
  54392=>"011010110",
  54393=>"011110110",
  54394=>"001101000",
  54395=>"111111100",
  54396=>"010000101",
  54397=>"111011000",
  54398=>"111100000",
  54399=>"001101101",
  54400=>"100100111",
  54401=>"111000001",
  54402=>"110010101",
  54403=>"100000011",
  54404=>"110101000",
  54405=>"100011101",
  54406=>"001011000",
  54407=>"110101000",
  54408=>"010001011",
  54409=>"111110001",
  54410=>"001100101",
  54411=>"110101010",
  54412=>"101000000",
  54413=>"001101110",
  54414=>"000110101",
  54415=>"101100111",
  54416=>"010011010",
  54417=>"011011111",
  54418=>"010101001",
  54419=>"010010111",
  54420=>"011000000",
  54421=>"001101010",
  54422=>"100111011",
  54423=>"001010100",
  54424=>"001001000",
  54425=>"001100111",
  54426=>"101100100",
  54427=>"000101110",
  54428=>"001101101",
  54429=>"111011000",
  54430=>"100110001",
  54431=>"000011100",
  54432=>"010110001",
  54433=>"010010101",
  54434=>"111101010",
  54435=>"000110100",
  54436=>"001100010",
  54437=>"111101100",
  54438=>"010100110",
  54439=>"111101110",
  54440=>"000101100",
  54441=>"011101111",
  54442=>"111100110",
  54443=>"011011010",
  54444=>"100100110",
  54445=>"010001001",
  54446=>"111000000",
  54447=>"101110110",
  54448=>"100000101",
  54449=>"001011011",
  54450=>"010111010",
  54451=>"110010111",
  54452=>"101010011",
  54453=>"100000000",
  54454=>"110001010",
  54455=>"000001010",
  54456=>"011110000",
  54457=>"010000001",
  54458=>"011110100",
  54459=>"001001001",
  54460=>"110111101",
  54461=>"111101011",
  54462=>"001110011",
  54463=>"011100110",
  54464=>"010010000",
  54465=>"011010100",
  54466=>"010101110",
  54467=>"110101011",
  54468=>"000001001",
  54469=>"110111101",
  54470=>"111001010",
  54471=>"010100001",
  54472=>"111100111",
  54473=>"111110010",
  54474=>"011011010",
  54475=>"110010000",
  54476=>"101010111",
  54477=>"100000011",
  54478=>"001000100",
  54479=>"111000000",
  54480=>"101111110",
  54481=>"101001010",
  54482=>"100001010",
  54483=>"111101100",
  54484=>"101110011",
  54485=>"111111100",
  54486=>"110100100",
  54487=>"010100000",
  54488=>"111001011",
  54489=>"011101101",
  54490=>"111101011",
  54491=>"100111001",
  54492=>"110111001",
  54493=>"100011101",
  54494=>"001001011",
  54495=>"001101010",
  54496=>"011111001",
  54497=>"100101011",
  54498=>"001101100",
  54499=>"101101111",
  54500=>"101000001",
  54501=>"011011011",
  54502=>"010000101",
  54503=>"111110011",
  54504=>"111001011",
  54505=>"110100100",
  54506=>"001101111",
  54507=>"001111101",
  54508=>"000100000",
  54509=>"011101001",
  54510=>"111100100",
  54511=>"001111100",
  54512=>"100010111",
  54513=>"001011011",
  54514=>"000000000",
  54515=>"001000000",
  54516=>"111101111",
  54517=>"110010011",
  54518=>"011101010",
  54519=>"110101000",
  54520=>"011000000",
  54521=>"000101101",
  54522=>"111100101",
  54523=>"101011101",
  54524=>"011011010",
  54525=>"100000111",
  54526=>"000000011",
  54527=>"001101001",
  54528=>"010101011",
  54529=>"010110000",
  54530=>"011010100",
  54531=>"101110001",
  54532=>"111100000",
  54533=>"011000000",
  54534=>"101111110",
  54535=>"111011001",
  54536=>"000001010",
  54537=>"100010000",
  54538=>"111001110",
  54539=>"001100001",
  54540=>"100111000",
  54541=>"111011010",
  54542=>"100000001",
  54543=>"000001100",
  54544=>"001100101",
  54545=>"010000011",
  54546=>"100100111",
  54547=>"001100101",
  54548=>"000111000",
  54549=>"010000001",
  54550=>"110101000",
  54551=>"101000001",
  54552=>"001110111",
  54553=>"001001011",
  54554=>"010000011",
  54555=>"001000100",
  54556=>"000001101",
  54557=>"010010111",
  54558=>"101010011",
  54559=>"100010011",
  54560=>"111011101",
  54561=>"110000001",
  54562=>"011100001",
  54563=>"011000010",
  54564=>"101010101",
  54565=>"001110001",
  54566=>"011000101",
  54567=>"010010101",
  54568=>"010011110",
  54569=>"101100110",
  54570=>"110011101",
  54571=>"111101001",
  54572=>"101101000",
  54573=>"101010100",
  54574=>"110000000",
  54575=>"101111010",
  54576=>"101101111",
  54577=>"011110001",
  54578=>"110010100",
  54579=>"001100000",
  54580=>"110101001",
  54581=>"101110111",
  54582=>"001010000",
  54583=>"101100101",
  54584=>"111111111",
  54585=>"100111100",
  54586=>"111001100",
  54587=>"001110001",
  54588=>"010111100",
  54589=>"010010010",
  54590=>"011111111",
  54591=>"010100111",
  54592=>"110100011",
  54593=>"011100010",
  54594=>"111111101",
  54595=>"001010110",
  54596=>"110100100",
  54597=>"011011101",
  54598=>"110000110",
  54599=>"001100011",
  54600=>"100100111",
  54601=>"010001100",
  54602=>"001010100",
  54603=>"010000001",
  54604=>"110001011",
  54605=>"001000001",
  54606=>"000101101",
  54607=>"011111100",
  54608=>"001100111",
  54609=>"000100110",
  54610=>"011010000",
  54611=>"111111010",
  54612=>"000010100",
  54613=>"100000011",
  54614=>"111011011",
  54615=>"001000100",
  54616=>"011010100",
  54617=>"110101001",
  54618=>"110101001",
  54619=>"000001011",
  54620=>"001100111",
  54621=>"011011001",
  54622=>"110101111",
  54623=>"111001011",
  54624=>"110001001",
  54625=>"001000000",
  54626=>"010111010",
  54627=>"100111000",
  54628=>"000011010",
  54629=>"100000011",
  54630=>"001001111",
  54631=>"010011100",
  54632=>"000111011",
  54633=>"000001111",
  54634=>"101101011",
  54635=>"100100000",
  54636=>"101100000",
  54637=>"000000101",
  54638=>"001101010",
  54639=>"010000001",
  54640=>"010101000",
  54641=>"000100000",
  54642=>"010111100",
  54643=>"001110010",
  54644=>"111101100",
  54645=>"000010000",
  54646=>"110101010",
  54647=>"000110011",
  54648=>"011010110",
  54649=>"001001101",
  54650=>"001011011",
  54651=>"010110001",
  54652=>"100111011",
  54653=>"101110101",
  54654=>"101000100",
  54655=>"111101000",
  54656=>"100100101",
  54657=>"110110001",
  54658=>"110011111",
  54659=>"010110001",
  54660=>"111001000",
  54661=>"100110110",
  54662=>"111001000",
  54663=>"101010001",
  54664=>"101101001",
  54665=>"011001011",
  54666=>"111111001",
  54667=>"001010111",
  54668=>"111101001",
  54669=>"100000000",
  54670=>"000100100",
  54671=>"011110100",
  54672=>"011010100",
  54673=>"000001001",
  54674=>"101101111",
  54675=>"110000011",
  54676=>"000110001",
  54677=>"010111110",
  54678=>"010010001",
  54679=>"000000001",
  54680=>"100111001",
  54681=>"010110001",
  54682=>"011011111",
  54683=>"101000100",
  54684=>"101111110",
  54685=>"010110110",
  54686=>"001110111",
  54687=>"001001001",
  54688=>"100010111",
  54689=>"100001100",
  54690=>"100010010",
  54691=>"000100001",
  54692=>"010100010",
  54693=>"110111110",
  54694=>"100100010",
  54695=>"111001110",
  54696=>"000111100",
  54697=>"100100111",
  54698=>"011100010",
  54699=>"111011001",
  54700=>"110100010",
  54701=>"110101010",
  54702=>"111000000",
  54703=>"110100101",
  54704=>"100000110",
  54705=>"000001010",
  54706=>"111001110",
  54707=>"110101100",
  54708=>"000100110",
  54709=>"101010001",
  54710=>"011010100",
  54711=>"110100111",
  54712=>"000110000",
  54713=>"001101110",
  54714=>"110000100",
  54715=>"000100100",
  54716=>"000111011",
  54717=>"000001110",
  54718=>"000000001",
  54719=>"111001010",
  54720=>"101101110",
  54721=>"111010101",
  54722=>"111101110",
  54723=>"010111010",
  54724=>"000000100",
  54725=>"011110111",
  54726=>"100100010",
  54727=>"001110111",
  54728=>"111111011",
  54729=>"111010011",
  54730=>"111101001",
  54731=>"000111101",
  54732=>"111101000",
  54733=>"110001010",
  54734=>"100101100",
  54735=>"011010101",
  54736=>"110001011",
  54737=>"111101000",
  54738=>"100010111",
  54739=>"010001000",
  54740=>"110111010",
  54741=>"110111011",
  54742=>"010000001",
  54743=>"011100111",
  54744=>"100100000",
  54745=>"100111011",
  54746=>"100001100",
  54747=>"110110001",
  54748=>"001100111",
  54749=>"111001100",
  54750=>"000000111",
  54751=>"111001100",
  54752=>"001111001",
  54753=>"010000010",
  54754=>"100011100",
  54755=>"101100111",
  54756=>"001011011",
  54757=>"100000000",
  54758=>"100000111",
  54759=>"110101110",
  54760=>"001001101",
  54761=>"000100111",
  54762=>"000000001",
  54763=>"110111111",
  54764=>"110111100",
  54765=>"011001100",
  54766=>"010101010",
  54767=>"101111000",
  54768=>"111110001",
  54769=>"010010000",
  54770=>"010110010",
  54771=>"011110010",
  54772=>"011000001",
  54773=>"010100100",
  54774=>"001111111",
  54775=>"101011100",
  54776=>"000010110",
  54777=>"010001111",
  54778=>"000111100",
  54779=>"010001001",
  54780=>"000000101",
  54781=>"100110010",
  54782=>"010000100",
  54783=>"001011110",
  54784=>"010000100",
  54785=>"010011100",
  54786=>"110001010",
  54787=>"001001010",
  54788=>"100011111",
  54789=>"000100110",
  54790=>"010110010",
  54791=>"001000101",
  54792=>"110001110",
  54793=>"011101111",
  54794=>"100011001",
  54795=>"000011110",
  54796=>"010101110",
  54797=>"011010000",
  54798=>"000010011",
  54799=>"001101101",
  54800=>"101111010",
  54801=>"100101110",
  54802=>"000000010",
  54803=>"111101100",
  54804=>"001011100",
  54805=>"000110011",
  54806=>"001100000",
  54807=>"111101111",
  54808=>"110011011",
  54809=>"001001011",
  54810=>"100110111",
  54811=>"110001101",
  54812=>"001001110",
  54813=>"001011111",
  54814=>"111010100",
  54815=>"110101001",
  54816=>"000011000",
  54817=>"000111101",
  54818=>"111100001",
  54819=>"010110110",
  54820=>"100101010",
  54821=>"100110010",
  54822=>"000000001",
  54823=>"011111000",
  54824=>"011110000",
  54825=>"110100001",
  54826=>"001001001",
  54827=>"001010010",
  54828=>"011111101",
  54829=>"001000001",
  54830=>"011011011",
  54831=>"110000010",
  54832=>"110100000",
  54833=>"001100110",
  54834=>"000000000",
  54835=>"100100110",
  54836=>"101011000",
  54837=>"110100111",
  54838=>"111000111",
  54839=>"111100010",
  54840=>"011001101",
  54841=>"001110101",
  54842=>"011101101",
  54843=>"100011110",
  54844=>"010000001",
  54845=>"110110011",
  54846=>"111100001",
  54847=>"101000101",
  54848=>"001110000",
  54849=>"000011011",
  54850=>"110110111",
  54851=>"011110101",
  54852=>"100010100",
  54853=>"010011010",
  54854=>"000010011",
  54855=>"100000100",
  54856=>"011101100",
  54857=>"110011001",
  54858=>"010001011",
  54859=>"111101111",
  54860=>"011110101",
  54861=>"101011011",
  54862=>"111000000",
  54863=>"111010001",
  54864=>"100010011",
  54865=>"101100101",
  54866=>"001100010",
  54867=>"011011000",
  54868=>"100011111",
  54869=>"101100100",
  54870=>"001011000",
  54871=>"110001111",
  54872=>"010001110",
  54873=>"010010000",
  54874=>"000001011",
  54875=>"100000110",
  54876=>"000111100",
  54877=>"011001011",
  54878=>"010101000",
  54879=>"010011001",
  54880=>"100000010",
  54881=>"001111110",
  54882=>"010001001",
  54883=>"001100010",
  54884=>"000100000",
  54885=>"000000010",
  54886=>"000111010",
  54887=>"110000101",
  54888=>"100001000",
  54889=>"110111100",
  54890=>"100011000",
  54891=>"110001110",
  54892=>"000011101",
  54893=>"100100100",
  54894=>"110111010",
  54895=>"010010111",
  54896=>"101010000",
  54897=>"101100000",
  54898=>"001001000",
  54899=>"111000001",
  54900=>"110101001",
  54901=>"111101100",
  54902=>"001110101",
  54903=>"110001010",
  54904=>"001001111",
  54905=>"110000110",
  54906=>"101011001",
  54907=>"011100100",
  54908=>"100010100",
  54909=>"110011100",
  54910=>"111110011",
  54911=>"101100001",
  54912=>"000011110",
  54913=>"111101111",
  54914=>"001110100",
  54915=>"101110101",
  54916=>"111100011",
  54917=>"010000111",
  54918=>"010011010",
  54919=>"001100101",
  54920=>"110010100",
  54921=>"100101111",
  54922=>"011111010",
  54923=>"000101011",
  54924=>"100110011",
  54925=>"000110011",
  54926=>"001100111",
  54927=>"000100100",
  54928=>"011110000",
  54929=>"011000111",
  54930=>"010111100",
  54931=>"001000100",
  54932=>"001010011",
  54933=>"011010011",
  54934=>"010110011",
  54935=>"010011100",
  54936=>"101101011",
  54937=>"010001011",
  54938=>"100000000",
  54939=>"100010011",
  54940=>"010000110",
  54941=>"000110000",
  54942=>"011110000",
  54943=>"111111000",
  54944=>"011100101",
  54945=>"000101100",
  54946=>"110000110",
  54947=>"010001000",
  54948=>"000001111",
  54949=>"001100000",
  54950=>"000010001",
  54951=>"011111110",
  54952=>"010000001",
  54953=>"000000010",
  54954=>"101010000",
  54955=>"101101101",
  54956=>"111001100",
  54957=>"011101010",
  54958=>"101001100",
  54959=>"101011111",
  54960=>"001010011",
  54961=>"110010011",
  54962=>"000111100",
  54963=>"010101111",
  54964=>"110110001",
  54965=>"001010011",
  54966=>"101000001",
  54967=>"110100101",
  54968=>"101110010",
  54969=>"100000001",
  54970=>"111000111",
  54971=>"111100101",
  54972=>"101111001",
  54973=>"100010001",
  54974=>"101001010",
  54975=>"000001001",
  54976=>"111111100",
  54977=>"001010000",
  54978=>"111110001",
  54979=>"101101010",
  54980=>"110001010",
  54981=>"011000100",
  54982=>"111111101",
  54983=>"000010000",
  54984=>"111010001",
  54985=>"010011100",
  54986=>"111011111",
  54987=>"101000100",
  54988=>"101110110",
  54989=>"100101111",
  54990=>"000001001",
  54991=>"110011110",
  54992=>"111111111",
  54993=>"010001101",
  54994=>"100000101",
  54995=>"011000001",
  54996=>"101010110",
  54997=>"001000010",
  54998=>"010010110",
  54999=>"001011010",
  55000=>"000101110",
  55001=>"001001110",
  55002=>"101111001",
  55003=>"000101000",
  55004=>"100010111",
  55005=>"000001001",
  55006=>"011111010",
  55007=>"101010011",
  55008=>"111000011",
  55009=>"101000100",
  55010=>"101100101",
  55011=>"111110010",
  55012=>"100000100",
  55013=>"100110000",
  55014=>"110101000",
  55015=>"110110010",
  55016=>"001000100",
  55017=>"010111001",
  55018=>"110000000",
  55019=>"000101110",
  55020=>"111010011",
  55021=>"110111100",
  55022=>"000010011",
  55023=>"001000000",
  55024=>"110001011",
  55025=>"001000010",
  55026=>"000100001",
  55027=>"100111111",
  55028=>"100111111",
  55029=>"110000011",
  55030=>"100110110",
  55031=>"111000000",
  55032=>"110010110",
  55033=>"100010100",
  55034=>"001000001",
  55035=>"011100010",
  55036=>"011101111",
  55037=>"000011111",
  55038=>"001110101",
  55039=>"000000001",
  55040=>"010111000",
  55041=>"001101101",
  55042=>"010000111",
  55043=>"011001001",
  55044=>"001101000",
  55045=>"000010011",
  55046=>"100110110",
  55047=>"000111110",
  55048=>"011001000",
  55049=>"110001100",
  55050=>"110111010",
  55051=>"101110000",
  55052=>"000101100",
  55053=>"010100101",
  55054=>"011000000",
  55055=>"110111001",
  55056=>"100001110",
  55057=>"111110001",
  55058=>"001010010",
  55059=>"111111101",
  55060=>"111010100",
  55061=>"100010100",
  55062=>"001101010",
  55063=>"101101100",
  55064=>"110100110",
  55065=>"000001011",
  55066=>"100011010",
  55067=>"111010001",
  55068=>"100101001",
  55069=>"111111001",
  55070=>"000010011",
  55071=>"110100100",
  55072=>"111111101",
  55073=>"010111000",
  55074=>"111111101",
  55075=>"001110011",
  55076=>"100001001",
  55077=>"010000111",
  55078=>"000000100",
  55079=>"101110100",
  55080=>"111110110",
  55081=>"000100000",
  55082=>"100100110",
  55083=>"110000101",
  55084=>"011111011",
  55085=>"100111001",
  55086=>"101110001",
  55087=>"011001100",
  55088=>"000000100",
  55089=>"111011111",
  55090=>"010000101",
  55091=>"001011100",
  55092=>"011000110",
  55093=>"110001101",
  55094=>"010110111",
  55095=>"011101110",
  55096=>"000100110",
  55097=>"100110100",
  55098=>"111001011",
  55099=>"000101111",
  55100=>"010000011",
  55101=>"000110100",
  55102=>"000101010",
  55103=>"110111111",
  55104=>"001111011",
  55105=>"101001101",
  55106=>"000000011",
  55107=>"111110010",
  55108=>"101010001",
  55109=>"101001000",
  55110=>"111110100",
  55111=>"010010110",
  55112=>"000010111",
  55113=>"110100101",
  55114=>"010110111",
  55115=>"110001100",
  55116=>"010110000",
  55117=>"000000110",
  55118=>"100101010",
  55119=>"110001001",
  55120=>"000110011",
  55121=>"101001010",
  55122=>"010010010",
  55123=>"000100110",
  55124=>"000101101",
  55125=>"101111000",
  55126=>"011010110",
  55127=>"110111001",
  55128=>"100101110",
  55129=>"111101101",
  55130=>"000010101",
  55131=>"110101111",
  55132=>"000000001",
  55133=>"111000000",
  55134=>"000001111",
  55135=>"101000011",
  55136=>"111101101",
  55137=>"010000011",
  55138=>"001101010",
  55139=>"110001000",
  55140=>"000000010",
  55141=>"000000011",
  55142=>"001101110",
  55143=>"100100011",
  55144=>"010000001",
  55145=>"111111101",
  55146=>"000010001",
  55147=>"110000000",
  55148=>"101000001",
  55149=>"111101011",
  55150=>"101101010",
  55151=>"101000111",
  55152=>"000111110",
  55153=>"111001101",
  55154=>"100111111",
  55155=>"111010001",
  55156=>"000000111",
  55157=>"110011110",
  55158=>"001011100",
  55159=>"101110010",
  55160=>"011000011",
  55161=>"011101000",
  55162=>"111111111",
  55163=>"110100101",
  55164=>"111101011",
  55165=>"100010111",
  55166=>"111111001",
  55167=>"000111100",
  55168=>"111110010",
  55169=>"111010111",
  55170=>"010100100",
  55171=>"110100010",
  55172=>"000011001",
  55173=>"110100111",
  55174=>"011001110",
  55175=>"001000001",
  55176=>"101001101",
  55177=>"001111111",
  55178=>"111100111",
  55179=>"110111100",
  55180=>"101000001",
  55181=>"100110101",
  55182=>"111101100",
  55183=>"111001111",
  55184=>"110010011",
  55185=>"010111001",
  55186=>"101011001",
  55187=>"010010110",
  55188=>"110111000",
  55189=>"110111001",
  55190=>"110000100",
  55191=>"011010010",
  55192=>"111101001",
  55193=>"111101000",
  55194=>"100101110",
  55195=>"011011000",
  55196=>"011111101",
  55197=>"100011001",
  55198=>"101110111",
  55199=>"010000110",
  55200=>"000000110",
  55201=>"011000100",
  55202=>"000010100",
  55203=>"000111101",
  55204=>"001111111",
  55205=>"111010011",
  55206=>"111111001",
  55207=>"011001010",
  55208=>"010101011",
  55209=>"010000111",
  55210=>"000110010",
  55211=>"000001110",
  55212=>"001100000",
  55213=>"000010101",
  55214=>"111111000",
  55215=>"011111010",
  55216=>"111100011",
  55217=>"101010010",
  55218=>"010001000",
  55219=>"010100001",
  55220=>"000111100",
  55221=>"001001110",
  55222=>"101000111",
  55223=>"110101100",
  55224=>"110101111",
  55225=>"110111001",
  55226=>"111001011",
  55227=>"101011110",
  55228=>"000101011",
  55229=>"111000000",
  55230=>"100101000",
  55231=>"000011011",
  55232=>"110010101",
  55233=>"000001111",
  55234=>"001101010",
  55235=>"110011000",
  55236=>"101000100",
  55237=>"000000101",
  55238=>"001101100",
  55239=>"100001111",
  55240=>"100011001",
  55241=>"101100111",
  55242=>"000100001",
  55243=>"100010001",
  55244=>"111101101",
  55245=>"011101010",
  55246=>"100010000",
  55247=>"111110010",
  55248=>"000000100",
  55249=>"100111111",
  55250=>"001011000",
  55251=>"111001100",
  55252=>"110010100",
  55253=>"110110100",
  55254=>"011010110",
  55255=>"111101010",
  55256=>"101110010",
  55257=>"011000100",
  55258=>"101100101",
  55259=>"000111011",
  55260=>"010001000",
  55261=>"010011011",
  55262=>"001010000",
  55263=>"001101001",
  55264=>"010001100",
  55265=>"100010000",
  55266=>"011010010",
  55267=>"110110010",
  55268=>"111001101",
  55269=>"101011110",
  55270=>"111111000",
  55271=>"001101011",
  55272=>"000001000",
  55273=>"111101110",
  55274=>"100111101",
  55275=>"010001101",
  55276=>"011100110",
  55277=>"000000101",
  55278=>"000110000",
  55279=>"011000111",
  55280=>"110010000",
  55281=>"111101011",
  55282=>"001111101",
  55283=>"011111010",
  55284=>"011101011",
  55285=>"101111111",
  55286=>"011010011",
  55287=>"111001111",
  55288=>"001111010",
  55289=>"111000110",
  55290=>"011011111",
  55291=>"001010101",
  55292=>"011100110",
  55293=>"001001000",
  55294=>"111110000",
  55295=>"110010101",
  55296=>"010001010",
  55297=>"111010100",
  55298=>"010010111",
  55299=>"001101011",
  55300=>"000000001",
  55301=>"100010011",
  55302=>"111011011",
  55303=>"110100101",
  55304=>"100111110",
  55305=>"100111011",
  55306=>"011111001",
  55307=>"110010111",
  55308=>"001100111",
  55309=>"001001110",
  55310=>"000110100",
  55311=>"111110000",
  55312=>"010000100",
  55313=>"000000100",
  55314=>"010010001",
  55315=>"010101101",
  55316=>"100001110",
  55317=>"110010011",
  55318=>"011001011",
  55319=>"000000101",
  55320=>"011010011",
  55321=>"001001001",
  55322=>"110100100",
  55323=>"011010110",
  55324=>"001101000",
  55325=>"001101011",
  55326=>"110101101",
  55327=>"010010011",
  55328=>"100000001",
  55329=>"010000000",
  55330=>"010110100",
  55331=>"001100100",
  55332=>"010110001",
  55333=>"011011001",
  55334=>"101100010",
  55335=>"111011111",
  55336=>"101010111",
  55337=>"000010000",
  55338=>"010101101",
  55339=>"010111100",
  55340=>"010010100",
  55341=>"100000101",
  55342=>"001101001",
  55343=>"111001001",
  55344=>"110011010",
  55345=>"000101110",
  55346=>"111000011",
  55347=>"100101000",
  55348=>"110100011",
  55349=>"110101000",
  55350=>"110100111",
  55351=>"110000000",
  55352=>"000101010",
  55353=>"100001000",
  55354=>"001101001",
  55355=>"000101001",
  55356=>"101000001",
  55357=>"010000011",
  55358=>"101111010",
  55359=>"111110010",
  55360=>"001010000",
  55361=>"100000100",
  55362=>"110011101",
  55363=>"101011010",
  55364=>"101110001",
  55365=>"110010010",
  55366=>"101101011",
  55367=>"110000010",
  55368=>"000010111",
  55369=>"011010001",
  55370=>"000101001",
  55371=>"001111001",
  55372=>"000000010",
  55373=>"001001110",
  55374=>"111110000",
  55375=>"000010011",
  55376=>"110100101",
  55377=>"111101110",
  55378=>"000111010",
  55379=>"000110010",
  55380=>"111011100",
  55381=>"110100111",
  55382=>"010100000",
  55383=>"000100000",
  55384=>"001110100",
  55385=>"110100100",
  55386=>"001001100",
  55387=>"110000110",
  55388=>"000101110",
  55389=>"010110100",
  55390=>"110111000",
  55391=>"111100111",
  55392=>"110110000",
  55393=>"001011110",
  55394=>"000010010",
  55395=>"101100011",
  55396=>"111110000",
  55397=>"111000011",
  55398=>"111001101",
  55399=>"111100101",
  55400=>"100100100",
  55401=>"101101010",
  55402=>"000100110",
  55403=>"101111111",
  55404=>"101100110",
  55405=>"100100100",
  55406=>"000010100",
  55407=>"101000100",
  55408=>"010100110",
  55409=>"011011001",
  55410=>"111001111",
  55411=>"001000001",
  55412=>"111011000",
  55413=>"011010011",
  55414=>"110011010",
  55415=>"100100010",
  55416=>"100000101",
  55417=>"011000100",
  55418=>"110100011",
  55419=>"100011001",
  55420=>"110110100",
  55421=>"111110110",
  55422=>"000000100",
  55423=>"011010010",
  55424=>"000111011",
  55425=>"110001100",
  55426=>"000000011",
  55427=>"010000100",
  55428=>"010010000",
  55429=>"111001011",
  55430=>"110010111",
  55431=>"001011100",
  55432=>"101001101",
  55433=>"101110100",
  55434=>"011111000",
  55435=>"001101110",
  55436=>"010001111",
  55437=>"011011111",
  55438=>"011110111",
  55439=>"101101011",
  55440=>"101100100",
  55441=>"001111111",
  55442=>"100010010",
  55443=>"011000100",
  55444=>"011011111",
  55445=>"000100100",
  55446=>"101011000",
  55447=>"001100000",
  55448=>"000100000",
  55449=>"101101111",
  55450=>"010110110",
  55451=>"111001000",
  55452=>"100100100",
  55453=>"101111110",
  55454=>"000001101",
  55455=>"011000001",
  55456=>"110000101",
  55457=>"111111011",
  55458=>"100101110",
  55459=>"001011011",
  55460=>"010000111",
  55461=>"000000010",
  55462=>"110000010",
  55463=>"100110111",
  55464=>"110101001",
  55465=>"101001011",
  55466=>"111101110",
  55467=>"010011101",
  55468=>"111010010",
  55469=>"111100011",
  55470=>"110010010",
  55471=>"100110101",
  55472=>"001010000",
  55473=>"010010100",
  55474=>"001000111",
  55475=>"110111101",
  55476=>"000110000",
  55477=>"000100110",
  55478=>"100100001",
  55479=>"010100010",
  55480=>"011001000",
  55481=>"100101001",
  55482=>"001001101",
  55483=>"001100111",
  55484=>"011111001",
  55485=>"111100111",
  55486=>"001101010",
  55487=>"101101110",
  55488=>"001001011",
  55489=>"001101011",
  55490=>"001001000",
  55491=>"111001100",
  55492=>"001011001",
  55493=>"001001110",
  55494=>"110100010",
  55495=>"000010011",
  55496=>"111110001",
  55497=>"000011110",
  55498=>"101110010",
  55499=>"100111001",
  55500=>"111001000",
  55501=>"000010010",
  55502=>"111111000",
  55503=>"110111000",
  55504=>"011111111",
  55505=>"110010101",
  55506=>"111111101",
  55507=>"101110001",
  55508=>"110000001",
  55509=>"110001000",
  55510=>"010111110",
  55511=>"010110100",
  55512=>"010000000",
  55513=>"001001000",
  55514=>"110010111",
  55515=>"100111011",
  55516=>"011110100",
  55517=>"011110110",
  55518=>"100111010",
  55519=>"111001001",
  55520=>"001110101",
  55521=>"100000100",
  55522=>"100000110",
  55523=>"110001111",
  55524=>"000101001",
  55525=>"110111111",
  55526=>"100001000",
  55527=>"001000000",
  55528=>"111101000",
  55529=>"100001001",
  55530=>"010000001",
  55531=>"000011000",
  55532=>"111101111",
  55533=>"011011000",
  55534=>"000000101",
  55535=>"010111000",
  55536=>"110000000",
  55537=>"110101010",
  55538=>"001010100",
  55539=>"110100010",
  55540=>"011010011",
  55541=>"000001001",
  55542=>"110010110",
  55543=>"010100001",
  55544=>"011101010",
  55545=>"000100001",
  55546=>"011100011",
  55547=>"001100101",
  55548=>"011000110",
  55549=>"000110000",
  55550=>"110101000",
  55551=>"111110101",
  55552=>"110101010",
  55553=>"100101000",
  55554=>"100000110",
  55555=>"010011100",
  55556=>"110100001",
  55557=>"111110110",
  55558=>"000001110",
  55559=>"111100011",
  55560=>"011010000",
  55561=>"011001111",
  55562=>"000111111",
  55563=>"101010001",
  55564=>"000101111",
  55565=>"100010010",
  55566=>"100101110",
  55567=>"110100111",
  55568=>"001001011",
  55569=>"100001000",
  55570=>"010010100",
  55571=>"000001111",
  55572=>"110111010",
  55573=>"001001111",
  55574=>"000010101",
  55575=>"000101011",
  55576=>"000100110",
  55577=>"101000010",
  55578=>"000101001",
  55579=>"011010010",
  55580=>"110010101",
  55581=>"010111110",
  55582=>"111011011",
  55583=>"010111111",
  55584=>"111010100",
  55585=>"101011011",
  55586=>"100011111",
  55587=>"000111101",
  55588=>"101111100",
  55589=>"100001000",
  55590=>"011111011",
  55591=>"001111011",
  55592=>"010100000",
  55593=>"011010110",
  55594=>"111111110",
  55595=>"000011001",
  55596=>"100001100",
  55597=>"100000110",
  55598=>"001001100",
  55599=>"010000010",
  55600=>"001100000",
  55601=>"010111101",
  55602=>"011001010",
  55603=>"001101111",
  55604=>"101011000",
  55605=>"111001001",
  55606=>"001011111",
  55607=>"101011010",
  55608=>"100001000",
  55609=>"110110010",
  55610=>"111101011",
  55611=>"011011101",
  55612=>"101110100",
  55613=>"010011110",
  55614=>"101101010",
  55615=>"111100001",
  55616=>"100100111",
  55617=>"100101010",
  55618=>"011111111",
  55619=>"000010111",
  55620=>"110101000",
  55621=>"010000010",
  55622=>"001010100",
  55623=>"001101010",
  55624=>"111011101",
  55625=>"101110111",
  55626=>"100110100",
  55627=>"001001110",
  55628=>"000011011",
  55629=>"000001001",
  55630=>"101111110",
  55631=>"011100110",
  55632=>"111000000",
  55633=>"011101010",
  55634=>"100111010",
  55635=>"010001001",
  55636=>"100100011",
  55637=>"101000001",
  55638=>"111001111",
  55639=>"010001110",
  55640=>"110100111",
  55641=>"100111100",
  55642=>"000110011",
  55643=>"101011010",
  55644=>"110110111",
  55645=>"110101001",
  55646=>"111000000",
  55647=>"100001001",
  55648=>"011001101",
  55649=>"011100010",
  55650=>"000100100",
  55651=>"001100110",
  55652=>"000010001",
  55653=>"000011001",
  55654=>"110001000",
  55655=>"101110001",
  55656=>"000000100",
  55657=>"110100111",
  55658=>"010100110",
  55659=>"110100101",
  55660=>"010001000",
  55661=>"111001111",
  55662=>"010000100",
  55663=>"100100100",
  55664=>"111110101",
  55665=>"011110001",
  55666=>"110110111",
  55667=>"111111111",
  55668=>"101100000",
  55669=>"001010010",
  55670=>"101010011",
  55671=>"101100010",
  55672=>"110001101",
  55673=>"011011111",
  55674=>"111111101",
  55675=>"100000111",
  55676=>"000000011",
  55677=>"110110011",
  55678=>"101110101",
  55679=>"010100011",
  55680=>"001010111",
  55681=>"100111001",
  55682=>"101101000",
  55683=>"100110000",
  55684=>"111110101",
  55685=>"110010100",
  55686=>"010110110",
  55687=>"110100010",
  55688=>"010000000",
  55689=>"001110111",
  55690=>"001001111",
  55691=>"001011111",
  55692=>"100001111",
  55693=>"010001010",
  55694=>"110111110",
  55695=>"001011110",
  55696=>"000000010",
  55697=>"001110100",
  55698=>"101001000",
  55699=>"101000001",
  55700=>"010100010",
  55701=>"111000000",
  55702=>"111111110",
  55703=>"101110001",
  55704=>"110110100",
  55705=>"000011000",
  55706=>"100010110",
  55707=>"011111110",
  55708=>"001001011",
  55709=>"101011001",
  55710=>"101111110",
  55711=>"011011010",
  55712=>"010100100",
  55713=>"111001000",
  55714=>"101101010",
  55715=>"011100000",
  55716=>"101110101",
  55717=>"111101100",
  55718=>"001101110",
  55719=>"001011110",
  55720=>"000101101",
  55721=>"110101101",
  55722=>"101101000",
  55723=>"010110001",
  55724=>"101110111",
  55725=>"111001010",
  55726=>"000111000",
  55727=>"100000110",
  55728=>"010011001",
  55729=>"111010001",
  55730=>"011110110",
  55731=>"010000101",
  55732=>"000000000",
  55733=>"011101110",
  55734=>"100001111",
  55735=>"000000011",
  55736=>"010010010",
  55737=>"101000000",
  55738=>"110100001",
  55739=>"111111101",
  55740=>"110001101",
  55741=>"000101101",
  55742=>"101111101",
  55743=>"110011000",
  55744=>"100101111",
  55745=>"110000100",
  55746=>"011110010",
  55747=>"001000110",
  55748=>"010000001",
  55749=>"001111000",
  55750=>"110100001",
  55751=>"100000100",
  55752=>"001010000",
  55753=>"110000001",
  55754=>"110000111",
  55755=>"110001111",
  55756=>"000001100",
  55757=>"001001100",
  55758=>"001111110",
  55759=>"111000100",
  55760=>"100110110",
  55761=>"010111000",
  55762=>"000010100",
  55763=>"111101110",
  55764=>"000110011",
  55765=>"100000100",
  55766=>"110010111",
  55767=>"100010000",
  55768=>"100110110",
  55769=>"101101010",
  55770=>"011000001",
  55771=>"000111100",
  55772=>"111110011",
  55773=>"010001100",
  55774=>"011101111",
  55775=>"100110111",
  55776=>"000100011",
  55777=>"010010100",
  55778=>"101011111",
  55779=>"001011000",
  55780=>"001011010",
  55781=>"110111000",
  55782=>"000101110",
  55783=>"011100100",
  55784=>"001011010",
  55785=>"010101101",
  55786=>"111110110",
  55787=>"100001111",
  55788=>"100100100",
  55789=>"110111101",
  55790=>"010001010",
  55791=>"111001110",
  55792=>"100110001",
  55793=>"000111010",
  55794=>"000111000",
  55795=>"011000100",
  55796=>"000001000",
  55797=>"001110100",
  55798=>"100101010",
  55799=>"010011010",
  55800=>"100011010",
  55801=>"011111010",
  55802=>"110101011",
  55803=>"111101010",
  55804=>"111100011",
  55805=>"011010111",
  55806=>"001010010",
  55807=>"101010011",
  55808=>"000100100",
  55809=>"011011011",
  55810=>"101011010",
  55811=>"100000101",
  55812=>"100110101",
  55813=>"101111000",
  55814=>"111101100",
  55815=>"010011010",
  55816=>"001101010",
  55817=>"001100110",
  55818=>"001010101",
  55819=>"000001000",
  55820=>"110000111",
  55821=>"000111010",
  55822=>"111000001",
  55823=>"100010010",
  55824=>"110011010",
  55825=>"110110010",
  55826=>"111011000",
  55827=>"100011101",
  55828=>"000100001",
  55829=>"011011010",
  55830=>"001001001",
  55831=>"110001110",
  55832=>"011111001",
  55833=>"111010100",
  55834=>"110100100",
  55835=>"011001011",
  55836=>"000101010",
  55837=>"011011100",
  55838=>"100110101",
  55839=>"100000101",
  55840=>"101010111",
  55841=>"010100010",
  55842=>"110100011",
  55843=>"111100001",
  55844=>"101110100",
  55845=>"000011010",
  55846=>"010011100",
  55847=>"010111000",
  55848=>"001101110",
  55849=>"110001010",
  55850=>"111111100",
  55851=>"011111110",
  55852=>"111001010",
  55853=>"101001000",
  55854=>"111000000",
  55855=>"101010111",
  55856=>"110010011",
  55857=>"110010101",
  55858=>"000000001",
  55859=>"101000101",
  55860=>"101110010",
  55861=>"000001001",
  55862=>"100011011",
  55863=>"011011111",
  55864=>"011100111",
  55865=>"101110101",
  55866=>"101010001",
  55867=>"010001110",
  55868=>"111111101",
  55869=>"101010000",
  55870=>"110010110",
  55871=>"000101110",
  55872=>"100010100",
  55873=>"010010000",
  55874=>"100110101",
  55875=>"000101111",
  55876=>"010011101",
  55877=>"001010001",
  55878=>"100110001",
  55879=>"101100000",
  55880=>"110011100",
  55881=>"111111000",
  55882=>"000000011",
  55883=>"010011011",
  55884=>"010011101",
  55885=>"101111100",
  55886=>"010110111",
  55887=>"101110100",
  55888=>"010101011",
  55889=>"000010001",
  55890=>"101011101",
  55891=>"011000011",
  55892=>"100110101",
  55893=>"010000100",
  55894=>"100110100",
  55895=>"000101010",
  55896=>"011110000",
  55897=>"001111001",
  55898=>"010110011",
  55899=>"101010111",
  55900=>"110000100",
  55901=>"100110110",
  55902=>"110001011",
  55903=>"000100001",
  55904=>"101111000",
  55905=>"010111100",
  55906=>"101010111",
  55907=>"110000100",
  55908=>"111001011",
  55909=>"000011101",
  55910=>"010100110",
  55911=>"111001001",
  55912=>"001000000",
  55913=>"111111010",
  55914=>"011111101",
  55915=>"110011000",
  55916=>"001010101",
  55917=>"100111101",
  55918=>"001011000",
  55919=>"001010101",
  55920=>"110000000",
  55921=>"000001110",
  55922=>"000001000",
  55923=>"000011000",
  55924=>"111000101",
  55925=>"001111000",
  55926=>"100111110",
  55927=>"011010111",
  55928=>"010001111",
  55929=>"111001100",
  55930=>"110010101",
  55931=>"001001001",
  55932=>"000000000",
  55933=>"110111100",
  55934=>"111101100",
  55935=>"001100010",
  55936=>"101011010",
  55937=>"110010011",
  55938=>"100010111",
  55939=>"100001011",
  55940=>"100000101",
  55941=>"100011010",
  55942=>"000110111",
  55943=>"111011110",
  55944=>"100100001",
  55945=>"110001000",
  55946=>"000010111",
  55947=>"101110010",
  55948=>"011100101",
  55949=>"110100001",
  55950=>"001011001",
  55951=>"110111110",
  55952=>"011101101",
  55953=>"000100110",
  55954=>"111100111",
  55955=>"100101100",
  55956=>"000100001",
  55957=>"011101011",
  55958=>"111101100",
  55959=>"111111010",
  55960=>"110110001",
  55961=>"010001100",
  55962=>"110101101",
  55963=>"000000011",
  55964=>"011110010",
  55965=>"010011111",
  55966=>"101010000",
  55967=>"000001100",
  55968=>"010110100",
  55969=>"001011000",
  55970=>"000110111",
  55971=>"110001001",
  55972=>"111100101",
  55973=>"001010110",
  55974=>"010100000",
  55975=>"100000000",
  55976=>"001010011",
  55977=>"100110000",
  55978=>"000000110",
  55979=>"110000110",
  55980=>"110011010",
  55981=>"011010001",
  55982=>"110110011",
  55983=>"100000011",
  55984=>"110110000",
  55985=>"000011000",
  55986=>"001000000",
  55987=>"001000110",
  55988=>"100011111",
  55989=>"001110110",
  55990=>"100101111",
  55991=>"001100010",
  55992=>"100110000",
  55993=>"111111000",
  55994=>"001000110",
  55995=>"011010001",
  55996=>"111101100",
  55997=>"001111011",
  55998=>"101111100",
  55999=>"111111101",
  56000=>"010001110",
  56001=>"001111111",
  56002=>"001000010",
  56003=>"000000010",
  56004=>"101101101",
  56005=>"110000010",
  56006=>"100000111",
  56007=>"111011000",
  56008=>"001111101",
  56009=>"001100101",
  56010=>"000010100",
  56011=>"101000100",
  56012=>"110111000",
  56013=>"101101011",
  56014=>"001110101",
  56015=>"110100001",
  56016=>"110000101",
  56017=>"000011001",
  56018=>"001111010",
  56019=>"001000101",
  56020=>"011000101",
  56021=>"010000010",
  56022=>"010100110",
  56023=>"000110010",
  56024=>"111000110",
  56025=>"010110101",
  56026=>"110111010",
  56027=>"000110011",
  56028=>"100101110",
  56029=>"100110110",
  56030=>"011100011",
  56031=>"010111010",
  56032=>"101001110",
  56033=>"110000010",
  56034=>"001001100",
  56035=>"000001101",
  56036=>"101010101",
  56037=>"000001000",
  56038=>"110111111",
  56039=>"110100010",
  56040=>"110010111",
  56041=>"101100110",
  56042=>"010000011",
  56043=>"100100001",
  56044=>"000001001",
  56045=>"001111010",
  56046=>"010100010",
  56047=>"001011111",
  56048=>"111011100",
  56049=>"110101001",
  56050=>"111011100",
  56051=>"110100101",
  56052=>"000011100",
  56053=>"110001001",
  56054=>"101110010",
  56055=>"001001010",
  56056=>"011000011",
  56057=>"111001101",
  56058=>"010010111",
  56059=>"010001100",
  56060=>"011111100",
  56061=>"010101001",
  56062=>"000100001",
  56063=>"001011000",
  56064=>"010010100",
  56065=>"111011001",
  56066=>"110010111",
  56067=>"000111110",
  56068=>"100111010",
  56069=>"001010010",
  56070=>"010100011",
  56071=>"000011110",
  56072=>"000011011",
  56073=>"100100111",
  56074=>"010000110",
  56075=>"000101000",
  56076=>"100101000",
  56077=>"101011011",
  56078=>"100001100",
  56079=>"000100000",
  56080=>"100011100",
  56081=>"101000000",
  56082=>"011010010",
  56083=>"101000100",
  56084=>"010000001",
  56085=>"010111111",
  56086=>"100101011",
  56087=>"001011000",
  56088=>"101000000",
  56089=>"001001101",
  56090=>"000001011",
  56091=>"000001110",
  56092=>"111101110",
  56093=>"111000111",
  56094=>"110100000",
  56095=>"111011110",
  56096=>"111000111",
  56097=>"010110111",
  56098=>"001101110",
  56099=>"000001100",
  56100=>"100011100",
  56101=>"100000001",
  56102=>"110010010",
  56103=>"001000001",
  56104=>"011010001",
  56105=>"001011110",
  56106=>"001100100",
  56107=>"110110000",
  56108=>"010011010",
  56109=>"101110010",
  56110=>"111011110",
  56111=>"110101001",
  56112=>"101000000",
  56113=>"011001010",
  56114=>"110010100",
  56115=>"111010010",
  56116=>"011010001",
  56117=>"100110001",
  56118=>"110110001",
  56119=>"011110110",
  56120=>"110111110",
  56121=>"101100100",
  56122=>"101100001",
  56123=>"110100010",
  56124=>"001001010",
  56125=>"000100101",
  56126=>"000001111",
  56127=>"001000110",
  56128=>"110101001",
  56129=>"111100111",
  56130=>"010010000",
  56131=>"001111111",
  56132=>"110010000",
  56133=>"010000110",
  56134=>"110010110",
  56135=>"101101100",
  56136=>"000010100",
  56137=>"111110010",
  56138=>"011000110",
  56139=>"001100101",
  56140=>"110011011",
  56141=>"110110100",
  56142=>"001110100",
  56143=>"000101001",
  56144=>"110101101",
  56145=>"000000001",
  56146=>"100100100",
  56147=>"101000110",
  56148=>"011011000",
  56149=>"111101111",
  56150=>"000000000",
  56151=>"010101011",
  56152=>"001110000",
  56153=>"000001001",
  56154=>"010111110",
  56155=>"100110100",
  56156=>"010011011",
  56157=>"101101101",
  56158=>"101111011",
  56159=>"001001010",
  56160=>"000001011",
  56161=>"101010111",
  56162=>"111000001",
  56163=>"100001101",
  56164=>"001000010",
  56165=>"001001000",
  56166=>"000100001",
  56167=>"010011111",
  56168=>"100101110",
  56169=>"110001011",
  56170=>"100100100",
  56171=>"011010111",
  56172=>"100110100",
  56173=>"100000011",
  56174=>"100110111",
  56175=>"110111110",
  56176=>"001010100",
  56177=>"001110111",
  56178=>"101101111",
  56179=>"001110000",
  56180=>"010000010",
  56181=>"000100101",
  56182=>"101100100",
  56183=>"100110000",
  56184=>"000101110",
  56185=>"010100001",
  56186=>"111110111",
  56187=>"011001011",
  56188=>"011000100",
  56189=>"011011100",
  56190=>"000001111",
  56191=>"101101111",
  56192=>"000010011",
  56193=>"110011011",
  56194=>"100100111",
  56195=>"001000100",
  56196=>"101100000",
  56197=>"110100001",
  56198=>"110101010",
  56199=>"110111111",
  56200=>"011111111",
  56201=>"010011100",
  56202=>"111001101",
  56203=>"000110101",
  56204=>"011011000",
  56205=>"001011000",
  56206=>"100010010",
  56207=>"100110011",
  56208=>"100000111",
  56209=>"011011100",
  56210=>"011010100",
  56211=>"101111110",
  56212=>"111001011",
  56213=>"101110101",
  56214=>"001000011",
  56215=>"101110110",
  56216=>"001110001",
  56217=>"100110101",
  56218=>"101111011",
  56219=>"101111110",
  56220=>"000000011",
  56221=>"110000010",
  56222=>"001010010",
  56223=>"101010110",
  56224=>"000011000",
  56225=>"100100100",
  56226=>"001001110",
  56227=>"000000100",
  56228=>"100100001",
  56229=>"110110111",
  56230=>"011011000",
  56231=>"110001000",
  56232=>"100110111",
  56233=>"001010110",
  56234=>"110111010",
  56235=>"010011111",
  56236=>"100111000",
  56237=>"100111100",
  56238=>"110100110",
  56239=>"101100110",
  56240=>"111001000",
  56241=>"011010111",
  56242=>"001110111",
  56243=>"110000101",
  56244=>"011101110",
  56245=>"001011000",
  56246=>"010010010",
  56247=>"111011101",
  56248=>"010101100",
  56249=>"111001110",
  56250=>"001110100",
  56251=>"010010100",
  56252=>"010110001",
  56253=>"011001000",
  56254=>"111101111",
  56255=>"100000100",
  56256=>"000101110",
  56257=>"000101010",
  56258=>"000001010",
  56259=>"101101100",
  56260=>"110101001",
  56261=>"010010011",
  56262=>"000011011",
  56263=>"100001000",
  56264=>"100000111",
  56265=>"001101000",
  56266=>"110111011",
  56267=>"001010101",
  56268=>"100101000",
  56269=>"101100100",
  56270=>"001001011",
  56271=>"001010110",
  56272=>"010000101",
  56273=>"010000001",
  56274=>"010101101",
  56275=>"110000000",
  56276=>"100000101",
  56277=>"011100000",
  56278=>"101011111",
  56279=>"101100011",
  56280=>"110000100",
  56281=>"000100010",
  56282=>"000110010",
  56283=>"110001110",
  56284=>"001010111",
  56285=>"101001011",
  56286=>"000110100",
  56287=>"010111010",
  56288=>"100101000",
  56289=>"000111010",
  56290=>"001110100",
  56291=>"001100010",
  56292=>"000001100",
  56293=>"011110011",
  56294=>"100111111",
  56295=>"101000100",
  56296=>"001100100",
  56297=>"100101110",
  56298=>"010010010",
  56299=>"011110110",
  56300=>"011010000",
  56301=>"000111110",
  56302=>"110111111",
  56303=>"001000110",
  56304=>"111101110",
  56305=>"111000100",
  56306=>"011000000",
  56307=>"101011111",
  56308=>"111110011",
  56309=>"010101100",
  56310=>"111011011",
  56311=>"101110001",
  56312=>"110010110",
  56313=>"101011100",
  56314=>"100100001",
  56315=>"101000000",
  56316=>"101001101",
  56317=>"011010000",
  56318=>"000011101",
  56319=>"010011111",
  56320=>"111001010",
  56321=>"000011111",
  56322=>"010111011",
  56323=>"100000111",
  56324=>"110111001",
  56325=>"101110100",
  56326=>"001000100",
  56327=>"101010110",
  56328=>"111001100",
  56329=>"011000110",
  56330=>"001101111",
  56331=>"100111100",
  56332=>"000000001",
  56333=>"001111100",
  56334=>"011101101",
  56335=>"010100010",
  56336=>"001001100",
  56337=>"111110000",
  56338=>"001111011",
  56339=>"010000001",
  56340=>"101011101",
  56341=>"110010111",
  56342=>"010101011",
  56343=>"100000010",
  56344=>"101100111",
  56345=>"111000001",
  56346=>"110001010",
  56347=>"111010111",
  56348=>"100000010",
  56349=>"011101110",
  56350=>"101110100",
  56351=>"111100000",
  56352=>"001101011",
  56353=>"010000110",
  56354=>"110100101",
  56355=>"100110100",
  56356=>"100111111",
  56357=>"011000111",
  56358=>"011000001",
  56359=>"111011010",
  56360=>"110011001",
  56361=>"000011011",
  56362=>"001111110",
  56363=>"010111101",
  56364=>"100000000",
  56365=>"011001010",
  56366=>"110010011",
  56367=>"011101001",
  56368=>"010101000",
  56369=>"111010000",
  56370=>"110110011",
  56371=>"010001110",
  56372=>"011000011",
  56373=>"110001011",
  56374=>"110110100",
  56375=>"011111111",
  56376=>"100101100",
  56377=>"011000010",
  56378=>"111010011",
  56379=>"001111000",
  56380=>"011000100",
  56381=>"110101111",
  56382=>"000010100",
  56383=>"011111001",
  56384=>"000111100",
  56385=>"001000010",
  56386=>"101100010",
  56387=>"101110111",
  56388=>"111000101",
  56389=>"101010110",
  56390=>"100001011",
  56391=>"010001000",
  56392=>"110111101",
  56393=>"110000011",
  56394=>"010101110",
  56395=>"110101010",
  56396=>"100000110",
  56397=>"001101110",
  56398=>"111000001",
  56399=>"001000111",
  56400=>"000001001",
  56401=>"111110111",
  56402=>"000101001",
  56403=>"000000011",
  56404=>"000101001",
  56405=>"111011110",
  56406=>"111001100",
  56407=>"010010010",
  56408=>"001111010",
  56409=>"000010100",
  56410=>"101000101",
  56411=>"011011100",
  56412=>"011000100",
  56413=>"111111001",
  56414=>"110001001",
  56415=>"110111101",
  56416=>"110000100",
  56417=>"011000011",
  56418=>"111000000",
  56419=>"010010000",
  56420=>"011100000",
  56421=>"100011110",
  56422=>"001110110",
  56423=>"100110101",
  56424=>"001100101",
  56425=>"111011111",
  56426=>"000001100",
  56427=>"100011000",
  56428=>"001111111",
  56429=>"110010101",
  56430=>"110011110",
  56431=>"111111011",
  56432=>"011000000",
  56433=>"000110011",
  56434=>"010111000",
  56435=>"010011100",
  56436=>"000000100",
  56437=>"110110000",
  56438=>"111010110",
  56439=>"011011101",
  56440=>"010111010",
  56441=>"011010000",
  56442=>"111111000",
  56443=>"000010100",
  56444=>"001001110",
  56445=>"011000100",
  56446=>"000100001",
  56447=>"101010110",
  56448=>"110110011",
  56449=>"011000110",
  56450=>"101101100",
  56451=>"100011000",
  56452=>"101011111",
  56453=>"001101001",
  56454=>"110010000",
  56455=>"010001000",
  56456=>"100001110",
  56457=>"010000110",
  56458=>"100000000",
  56459=>"001011101",
  56460=>"000000111",
  56461=>"100001001",
  56462=>"010110000",
  56463=>"011100100",
  56464=>"101010111",
  56465=>"001011010",
  56466=>"111010110",
  56467=>"100010000",
  56468=>"000011110",
  56469=>"111111011",
  56470=>"101000010",
  56471=>"010001000",
  56472=>"101011010",
  56473=>"010111111",
  56474=>"110100011",
  56475=>"100101111",
  56476=>"010011011",
  56477=>"100100000",
  56478=>"101000110",
  56479=>"000100110",
  56480=>"111010011",
  56481=>"001110000",
  56482=>"101110010",
  56483=>"101111101",
  56484=>"110100010",
  56485=>"101111110",
  56486=>"101011001",
  56487=>"111010000",
  56488=>"111110010",
  56489=>"001011101",
  56490=>"100000111",
  56491=>"100110110",
  56492=>"000001011",
  56493=>"011100100",
  56494=>"011111001",
  56495=>"100100010",
  56496=>"110111011",
  56497=>"011111010",
  56498=>"001110111",
  56499=>"000011000",
  56500=>"010101110",
  56501=>"101101111",
  56502=>"111011001",
  56503=>"011111111",
  56504=>"011101001",
  56505=>"011111011",
  56506=>"100001011",
  56507=>"101110101",
  56508=>"011011010",
  56509=>"001111101",
  56510=>"000011000",
  56511=>"111000100",
  56512=>"110110101",
  56513=>"100111101",
  56514=>"100011110",
  56515=>"010000011",
  56516=>"000010001",
  56517=>"101110101",
  56518=>"110110000",
  56519=>"010010000",
  56520=>"111010000",
  56521=>"000000101",
  56522=>"110011001",
  56523=>"110001000",
  56524=>"001011110",
  56525=>"100101000",
  56526=>"000000010",
  56527=>"000000001",
  56528=>"101000010",
  56529=>"011010001",
  56530=>"000011011",
  56531=>"011000110",
  56532=>"101001111",
  56533=>"101000100",
  56534=>"001011011",
  56535=>"011001000",
  56536=>"010010010",
  56537=>"011101010",
  56538=>"000000111",
  56539=>"110110100",
  56540=>"011101000",
  56541=>"010010010",
  56542=>"110101011",
  56543=>"110111100",
  56544=>"110111101",
  56545=>"001100100",
  56546=>"110000010",
  56547=>"000010001",
  56548=>"001010101",
  56549=>"101010101",
  56550=>"110001110",
  56551=>"100101000",
  56552=>"000100110",
  56553=>"000101100",
  56554=>"011010010",
  56555=>"100110001",
  56556=>"110001011",
  56557=>"110000111",
  56558=>"010110110",
  56559=>"001111001",
  56560=>"111000000",
  56561=>"100000000",
  56562=>"000000000",
  56563=>"110001101",
  56564=>"110001110",
  56565=>"111010001",
  56566=>"100111101",
  56567=>"110010110",
  56568=>"000011100",
  56569=>"011011001",
  56570=>"001010000",
  56571=>"010111101",
  56572=>"101001001",
  56573=>"000100110",
  56574=>"010111101",
  56575=>"000110001",
  56576=>"010110011",
  56577=>"011111100",
  56578=>"101101101",
  56579=>"011000100",
  56580=>"100011001",
  56581=>"000010111",
  56582=>"000011111",
  56583=>"000010101",
  56584=>"000011011",
  56585=>"000011111",
  56586=>"000001010",
  56587=>"101000101",
  56588=>"010101110",
  56589=>"111011010",
  56590=>"000111111",
  56591=>"110011100",
  56592=>"001110010",
  56593=>"000000101",
  56594=>"111010100",
  56595=>"001111101",
  56596=>"101000101",
  56597=>"010000111",
  56598=>"010000000",
  56599=>"010111100",
  56600=>"010111010",
  56601=>"110000111",
  56602=>"011011010",
  56603=>"011011010",
  56604=>"011100110",
  56605=>"001110010",
  56606=>"000101100",
  56607=>"000111000",
  56608=>"000000001",
  56609=>"101001000",
  56610=>"100001000",
  56611=>"001101111",
  56612=>"000000100",
  56613=>"000000101",
  56614=>"100010101",
  56615=>"010111011",
  56616=>"110100011",
  56617=>"111100111",
  56618=>"000111011",
  56619=>"010001001",
  56620=>"100000001",
  56621=>"000000011",
  56622=>"000001100",
  56623=>"011000100",
  56624=>"001011101",
  56625=>"100001111",
  56626=>"110001001",
  56627=>"001110010",
  56628=>"000001110",
  56629=>"000100001",
  56630=>"110001001",
  56631=>"100100000",
  56632=>"110101001",
  56633=>"100111100",
  56634=>"100011111",
  56635=>"110010110",
  56636=>"010111101",
  56637=>"110111111",
  56638=>"010010010",
  56639=>"001111000",
  56640=>"100000101",
  56641=>"011110010",
  56642=>"101111100",
  56643=>"010011011",
  56644=>"011011111",
  56645=>"010010010",
  56646=>"001000110",
  56647=>"011000000",
  56648=>"111011001",
  56649=>"111111010",
  56650=>"011001011",
  56651=>"111111011",
  56652=>"010011001",
  56653=>"011010011",
  56654=>"100110001",
  56655=>"011011000",
  56656=>"010100011",
  56657=>"111000111",
  56658=>"100111101",
  56659=>"010011111",
  56660=>"000111100",
  56661=>"100101111",
  56662=>"101000111",
  56663=>"010001101",
  56664=>"000101011",
  56665=>"101000001",
  56666=>"111000110",
  56667=>"001011011",
  56668=>"011110100",
  56669=>"010100101",
  56670=>"101001011",
  56671=>"010110111",
  56672=>"110111011",
  56673=>"100000100",
  56674=>"011010111",
  56675=>"100110010",
  56676=>"110111001",
  56677=>"111100100",
  56678=>"101000110",
  56679=>"010011000",
  56680=>"110110011",
  56681=>"001100110",
  56682=>"000001000",
  56683=>"010110000",
  56684=>"110101011",
  56685=>"110110101",
  56686=>"001010111",
  56687=>"110111111",
  56688=>"001110110",
  56689=>"000011000",
  56690=>"110101101",
  56691=>"110100000",
  56692=>"111001111",
  56693=>"010010001",
  56694=>"000010001",
  56695=>"010000011",
  56696=>"000100011",
  56697=>"001111011",
  56698=>"110011000",
  56699=>"100000000",
  56700=>"010010111",
  56701=>"101110100",
  56702=>"111101010",
  56703=>"111100001",
  56704=>"001101111",
  56705=>"100110010",
  56706=>"000011010",
  56707=>"011010010",
  56708=>"010101101",
  56709=>"010011010",
  56710=>"011001010",
  56711=>"111111010",
  56712=>"111010000",
  56713=>"101000111",
  56714=>"000111011",
  56715=>"010001101",
  56716=>"001110001",
  56717=>"100011011",
  56718=>"010111001",
  56719=>"000011101",
  56720=>"011101000",
  56721=>"100001001",
  56722=>"100010111",
  56723=>"110011001",
  56724=>"000000011",
  56725=>"000100100",
  56726=>"001001110",
  56727=>"000011111",
  56728=>"110100110",
  56729=>"010101111",
  56730=>"100011010",
  56731=>"101101001",
  56732=>"101101101",
  56733=>"111111000",
  56734=>"110111101",
  56735=>"010000101",
  56736=>"010001110",
  56737=>"011100100",
  56738=>"011000000",
  56739=>"011100011",
  56740=>"010000001",
  56741=>"111101000",
  56742=>"001010100",
  56743=>"000101010",
  56744=>"110100100",
  56745=>"011100001",
  56746=>"001000011",
  56747=>"010001000",
  56748=>"010100010",
  56749=>"011111110",
  56750=>"110000001",
  56751=>"000101111",
  56752=>"000010110",
  56753=>"101101010",
  56754=>"111110101",
  56755=>"100001110",
  56756=>"111100100",
  56757=>"001110100",
  56758=>"000011111",
  56759=>"101001011",
  56760=>"010110010",
  56761=>"110111010",
  56762=>"000011010",
  56763=>"111101110",
  56764=>"100011000",
  56765=>"111000110",
  56766=>"100100110",
  56767=>"010000111",
  56768=>"010100111",
  56769=>"100111111",
  56770=>"111001001",
  56771=>"011000101",
  56772=>"110010110",
  56773=>"010101111",
  56774=>"010000110",
  56775=>"101001011",
  56776=>"100100001",
  56777=>"110110100",
  56778=>"010101011",
  56779=>"101001100",
  56780=>"100000110",
  56781=>"010111110",
  56782=>"100111101",
  56783=>"111110000",
  56784=>"000000100",
  56785=>"011100110",
  56786=>"111001010",
  56787=>"111001010",
  56788=>"110110111",
  56789=>"000111000",
  56790=>"110001100",
  56791=>"110101000",
  56792=>"101010100",
  56793=>"100101100",
  56794=>"110001000",
  56795=>"000001110",
  56796=>"011000100",
  56797=>"101100001",
  56798=>"110010111",
  56799=>"111010101",
  56800=>"001010111",
  56801=>"011011110",
  56802=>"111100010",
  56803=>"001100110",
  56804=>"011100101",
  56805=>"001001010",
  56806=>"111100010",
  56807=>"110111001",
  56808=>"110100110",
  56809=>"110001111",
  56810=>"101011010",
  56811=>"000110000",
  56812=>"101001001",
  56813=>"101101111",
  56814=>"110110011",
  56815=>"010111111",
  56816=>"011110000",
  56817=>"010110101",
  56818=>"111101110",
  56819=>"101001000",
  56820=>"011110101",
  56821=>"010101011",
  56822=>"000001010",
  56823=>"100101010",
  56824=>"010010010",
  56825=>"100001101",
  56826=>"011101010",
  56827=>"100001101",
  56828=>"101001000",
  56829=>"011001101",
  56830=>"001011000",
  56831=>"111110111",
  56832=>"010010001",
  56833=>"111101111",
  56834=>"110101111",
  56835=>"111010101",
  56836=>"011011001",
  56837=>"001001001",
  56838=>"001101101",
  56839=>"011110001",
  56840=>"000110111",
  56841=>"110100011",
  56842=>"000011100",
  56843=>"011110011",
  56844=>"010110000",
  56845=>"100011010",
  56846=>"111000011",
  56847=>"010110011",
  56848=>"011110111",
  56849=>"001101101",
  56850=>"000001001",
  56851=>"101111000",
  56852=>"001011011",
  56853=>"110011000",
  56854=>"000001111",
  56855=>"100110010",
  56856=>"011011111",
  56857=>"011010100",
  56858=>"100010100",
  56859=>"111011011",
  56860=>"100001111",
  56861=>"110000110",
  56862=>"100100001",
  56863=>"001100000",
  56864=>"000011011",
  56865=>"010001100",
  56866=>"000100110",
  56867=>"100011010",
  56868=>"111101010",
  56869=>"011010110",
  56870=>"110111110",
  56871=>"011001001",
  56872=>"011101001",
  56873=>"001110111",
  56874=>"000011000",
  56875=>"111111111",
  56876=>"010000101",
  56877=>"011100011",
  56878=>"011010100",
  56879=>"001000000",
  56880=>"011011110",
  56881=>"011111111",
  56882=>"100010110",
  56883=>"010001001",
  56884=>"100101111",
  56885=>"000000011",
  56886=>"001100000",
  56887=>"101001111",
  56888=>"001010001",
  56889=>"001111010",
  56890=>"110111000",
  56891=>"111001001",
  56892=>"001000000",
  56893=>"010111101",
  56894=>"101110100",
  56895=>"001000001",
  56896=>"011101110",
  56897=>"010000000",
  56898=>"110000101",
  56899=>"000110110",
  56900=>"100111000",
  56901=>"100110000",
  56902=>"010001000",
  56903=>"111111101",
  56904=>"000101101",
  56905=>"011001101",
  56906=>"111111100",
  56907=>"000111000",
  56908=>"001100000",
  56909=>"001001110",
  56910=>"101100000",
  56911=>"110111111",
  56912=>"000000001",
  56913=>"000010101",
  56914=>"010110110",
  56915=>"011011010",
  56916=>"000001000",
  56917=>"001010101",
  56918=>"010000011",
  56919=>"011001111",
  56920=>"101111110",
  56921=>"010100011",
  56922=>"000000111",
  56923=>"010010111",
  56924=>"000100100",
  56925=>"100010111",
  56926=>"010111101",
  56927=>"000110101",
  56928=>"100001110",
  56929=>"000001001",
  56930=>"010100101",
  56931=>"010010000",
  56932=>"111100101",
  56933=>"111001101",
  56934=>"111111000",
  56935=>"000101010",
  56936=>"111101011",
  56937=>"100101000",
  56938=>"101110011",
  56939=>"010010100",
  56940=>"000000111",
  56941=>"100011110",
  56942=>"001101000",
  56943=>"000101101",
  56944=>"001011010",
  56945=>"110010100",
  56946=>"101100000",
  56947=>"011101111",
  56948=>"010101000",
  56949=>"001101111",
  56950=>"101010011",
  56951=>"101010101",
  56952=>"000101001",
  56953=>"111100010",
  56954=>"111011100",
  56955=>"010110011",
  56956=>"100111110",
  56957=>"111000010",
  56958=>"000111111",
  56959=>"011110111",
  56960=>"000010001",
  56961=>"101010101",
  56962=>"110010000",
  56963=>"011100000",
  56964=>"000101010",
  56965=>"000110010",
  56966=>"000100000",
  56967=>"101100101",
  56968=>"010110001",
  56969=>"111101010",
  56970=>"001111010",
  56971=>"111010010",
  56972=>"010000011",
  56973=>"010001111",
  56974=>"100010001",
  56975=>"000101000",
  56976=>"110010100",
  56977=>"010101001",
  56978=>"101001111",
  56979=>"010111111",
  56980=>"101111011",
  56981=>"100110100",
  56982=>"010100011",
  56983=>"101110110",
  56984=>"000000010",
  56985=>"100110000",
  56986=>"001100100",
  56987=>"110010011",
  56988=>"111101000",
  56989=>"000001000",
  56990=>"010111110",
  56991=>"001111010",
  56992=>"111001010",
  56993=>"110010110",
  56994=>"000100100",
  56995=>"101001111",
  56996=>"011011110",
  56997=>"000011110",
  56998=>"000001010",
  56999=>"000011000",
  57000=>"000011100",
  57001=>"110011110",
  57002=>"111100110",
  57003=>"100000011",
  57004=>"011101001",
  57005=>"100011010",
  57006=>"011001100",
  57007=>"010101100",
  57008=>"001001001",
  57009=>"000011101",
  57010=>"110010010",
  57011=>"000111001",
  57012=>"000101000",
  57013=>"100101101",
  57014=>"110000010",
  57015=>"001001000",
  57016=>"111101110",
  57017=>"110010100",
  57018=>"111010101",
  57019=>"001110001",
  57020=>"001001110",
  57021=>"110111101",
  57022=>"011001001",
  57023=>"001000110",
  57024=>"000011001",
  57025=>"111100001",
  57026=>"011100011",
  57027=>"100010010",
  57028=>"110010101",
  57029=>"000011010",
  57030=>"001010101",
  57031=>"101000010",
  57032=>"111011010",
  57033=>"011101101",
  57034=>"010110110",
  57035=>"001000110",
  57036=>"011000111",
  57037=>"100001101",
  57038=>"110000001",
  57039=>"101110111",
  57040=>"011001110",
  57041=>"001100000",
  57042=>"111100011",
  57043=>"101110010",
  57044=>"000011000",
  57045=>"011000101",
  57046=>"011011001",
  57047=>"111110111",
  57048=>"100010111",
  57049=>"111000000",
  57050=>"010110001",
  57051=>"110011000",
  57052=>"001010011",
  57053=>"001000110",
  57054=>"001011000",
  57055=>"000110001",
  57056=>"001101100",
  57057=>"000000100",
  57058=>"000011101",
  57059=>"101111101",
  57060=>"010010001",
  57061=>"110001100",
  57062=>"001111010",
  57063=>"101111001",
  57064=>"111111101",
  57065=>"011110011",
  57066=>"001111100",
  57067=>"011110100",
  57068=>"000011000",
  57069=>"010000110",
  57070=>"001110000",
  57071=>"100101000",
  57072=>"111000010",
  57073=>"100111000",
  57074=>"100101010",
  57075=>"111010101",
  57076=>"100000001",
  57077=>"110101101",
  57078=>"001001100",
  57079=>"100011101",
  57080=>"001000001",
  57081=>"111110001",
  57082=>"000110001",
  57083=>"101100100",
  57084=>"011100100",
  57085=>"010010100",
  57086=>"100000001",
  57087=>"100000101",
  57088=>"000001010",
  57089=>"101100111",
  57090=>"001001010",
  57091=>"000000010",
  57092=>"000111111",
  57093=>"001111001",
  57094=>"110111010",
  57095=>"001011001",
  57096=>"001100111",
  57097=>"001001111",
  57098=>"011001001",
  57099=>"110110010",
  57100=>"100111000",
  57101=>"111100011",
  57102=>"010111100",
  57103=>"010111100",
  57104=>"110110100",
  57105=>"001110110",
  57106=>"111010101",
  57107=>"100101000",
  57108=>"010100000",
  57109=>"100010111",
  57110=>"100000001",
  57111=>"001011011",
  57112=>"101101000",
  57113=>"011101010",
  57114=>"000010111",
  57115=>"101010000",
  57116=>"010010111",
  57117=>"110101111",
  57118=>"000010100",
  57119=>"111000101",
  57120=>"101111001",
  57121=>"000001100",
  57122=>"111101010",
  57123=>"010011000",
  57124=>"111111100",
  57125=>"101111100",
  57126=>"000000001",
  57127=>"100111001",
  57128=>"001100001",
  57129=>"010010000",
  57130=>"000010100",
  57131=>"110000011",
  57132=>"000000011",
  57133=>"011000110",
  57134=>"101101000",
  57135=>"000010011",
  57136=>"010110010",
  57137=>"000110010",
  57138=>"011110111",
  57139=>"111000100",
  57140=>"111010100",
  57141=>"111001010",
  57142=>"101111000",
  57143=>"110110110",
  57144=>"100001101",
  57145=>"100011101",
  57146=>"101101000",
  57147=>"100100100",
  57148=>"100000000",
  57149=>"000010011",
  57150=>"110011101",
  57151=>"110011001",
  57152=>"101110000",
  57153=>"110110110",
  57154=>"111001110",
  57155=>"010100001",
  57156=>"101010001",
  57157=>"001110000",
  57158=>"111111010",
  57159=>"110101111",
  57160=>"111110011",
  57161=>"011110010",
  57162=>"011100100",
  57163=>"101001010",
  57164=>"010100110",
  57165=>"001111000",
  57166=>"000000100",
  57167=>"100110010",
  57168=>"000110100",
  57169=>"110011111",
  57170=>"101110101",
  57171=>"010001101",
  57172=>"011101101",
  57173=>"001111111",
  57174=>"110111000",
  57175=>"110011010",
  57176=>"100111111",
  57177=>"001011010",
  57178=>"111100011",
  57179=>"101001011",
  57180=>"000010111",
  57181=>"010111010",
  57182=>"111110110",
  57183=>"101101111",
  57184=>"000000101",
  57185=>"100110101",
  57186=>"000111100",
  57187=>"110001110",
  57188=>"110001100",
  57189=>"000010010",
  57190=>"010101010",
  57191=>"000001100",
  57192=>"100100000",
  57193=>"010111110",
  57194=>"111010010",
  57195=>"011000111",
  57196=>"001000001",
  57197=>"010001010",
  57198=>"000100010",
  57199=>"100011110",
  57200=>"100100001",
  57201=>"001111010",
  57202=>"100001100",
  57203=>"000000000",
  57204=>"100111001",
  57205=>"010111111",
  57206=>"000111111",
  57207=>"100000000",
  57208=>"011100110",
  57209=>"011100011",
  57210=>"101101110",
  57211=>"000000111",
  57212=>"100010110",
  57213=>"011110111",
  57214=>"000101011",
  57215=>"101100000",
  57216=>"001001010",
  57217=>"001101010",
  57218=>"100111110",
  57219=>"110100111",
  57220=>"010101010",
  57221=>"000000111",
  57222=>"000100100",
  57223=>"011000110",
  57224=>"110100101",
  57225=>"011100010",
  57226=>"010010100",
  57227=>"001111111",
  57228=>"010011110",
  57229=>"010110001",
  57230=>"010111000",
  57231=>"000001111",
  57232=>"010010001",
  57233=>"011011111",
  57234=>"100010110",
  57235=>"111010110",
  57236=>"101100110",
  57237=>"101101111",
  57238=>"001011001",
  57239=>"010110000",
  57240=>"110001011",
  57241=>"111101111",
  57242=>"111000111",
  57243=>"001001011",
  57244=>"000101000",
  57245=>"010111011",
  57246=>"111010011",
  57247=>"000001100",
  57248=>"111011000",
  57249=>"111001010",
  57250=>"101000100",
  57251=>"000010011",
  57252=>"110001000",
  57253=>"101000101",
  57254=>"101011110",
  57255=>"000111000",
  57256=>"101010000",
  57257=>"000001001",
  57258=>"001101100",
  57259=>"100000001",
  57260=>"001001101",
  57261=>"110000101",
  57262=>"101111111",
  57263=>"101010011",
  57264=>"110101110",
  57265=>"010000010",
  57266=>"101000011",
  57267=>"000000011",
  57268=>"011111100",
  57269=>"000011000",
  57270=>"010000100",
  57271=>"110111001",
  57272=>"100001110",
  57273=>"011100111",
  57274=>"111010000",
  57275=>"011001011",
  57276=>"100110000",
  57277=>"111001111",
  57278=>"000001110",
  57279=>"011000001",
  57280=>"110010111",
  57281=>"010001010",
  57282=>"111001000",
  57283=>"010010111",
  57284=>"101111011",
  57285=>"110011010",
  57286=>"100111010",
  57287=>"011101110",
  57288=>"101101101",
  57289=>"100101010",
  57290=>"100101100",
  57291=>"010110010",
  57292=>"001101001",
  57293=>"101011010",
  57294=>"110101110",
  57295=>"010111111",
  57296=>"101001001",
  57297=>"001001000",
  57298=>"101000010",
  57299=>"101001001",
  57300=>"011110100",
  57301=>"101110001",
  57302=>"100101011",
  57303=>"010110111",
  57304=>"001111001",
  57305=>"010000111",
  57306=>"100100100",
  57307=>"110100100",
  57308=>"111000110",
  57309=>"010100011",
  57310=>"111011011",
  57311=>"101110001",
  57312=>"011110101",
  57313=>"011010010",
  57314=>"011101101",
  57315=>"101100000",
  57316=>"101000011",
  57317=>"010010011",
  57318=>"111011001",
  57319=>"111111010",
  57320=>"100100011",
  57321=>"111010001",
  57322=>"000011000",
  57323=>"110010011",
  57324=>"011001110",
  57325=>"000001000",
  57326=>"100001000",
  57327=>"001010111",
  57328=>"011100001",
  57329=>"000101101",
  57330=>"101010101",
  57331=>"011000110",
  57332=>"110111111",
  57333=>"110000010",
  57334=>"011010101",
  57335=>"100011101",
  57336=>"000010000",
  57337=>"000011101",
  57338=>"111011001",
  57339=>"010110000",
  57340=>"000111111",
  57341=>"101001011",
  57342=>"011100110",
  57343=>"000001100",
  57344=>"111111111",
  57345=>"000101101",
  57346=>"011100111",
  57347=>"001111100",
  57348=>"010110100",
  57349=>"101101111",
  57350=>"101001111",
  57351=>"101100101",
  57352=>"110110001",
  57353=>"011101100",
  57354=>"111011010",
  57355=>"011110011",
  57356=>"110101110",
  57357=>"011110011",
  57358=>"111010110",
  57359=>"011101111",
  57360=>"101100001",
  57361=>"000011001",
  57362=>"111110110",
  57363=>"011000100",
  57364=>"011101100",
  57365=>"111101111",
  57366=>"010000000",
  57367=>"001000110",
  57368=>"011100010",
  57369=>"000110001",
  57370=>"010100100",
  57371=>"110001010",
  57372=>"101010110",
  57373=>"010100101",
  57374=>"111101111",
  57375=>"010101000",
  57376=>"111111101",
  57377=>"101100111",
  57378=>"000011100",
  57379=>"111010100",
  57380=>"111110010",
  57381=>"011000101",
  57382=>"111101001",
  57383=>"110110110",
  57384=>"111101111",
  57385=>"100111000",
  57386=>"110101011",
  57387=>"100100100",
  57388=>"111011001",
  57389=>"000000100",
  57390=>"110101001",
  57391=>"011001000",
  57392=>"000111100",
  57393=>"000100010",
  57394=>"001101111",
  57395=>"111101011",
  57396=>"011011111",
  57397=>"111010111",
  57398=>"011110110",
  57399=>"110111000",
  57400=>"110000110",
  57401=>"001101000",
  57402=>"101110100",
  57403=>"100111000",
  57404=>"010001100",
  57405=>"100000101",
  57406=>"111000000",
  57407=>"010010110",
  57408=>"101000100",
  57409=>"010010011",
  57410=>"010001101",
  57411=>"101001001",
  57412=>"011101000",
  57413=>"101011110",
  57414=>"000000101",
  57415=>"101111100",
  57416=>"010010100",
  57417=>"011000110",
  57418=>"011001101",
  57419=>"110100010",
  57420=>"100110100",
  57421=>"101001101",
  57422=>"101001001",
  57423=>"101101000",
  57424=>"011111111",
  57425=>"100100100",
  57426=>"011001000",
  57427=>"000110110",
  57428=>"110111111",
  57429=>"001100011",
  57430=>"000100010",
  57431=>"001111111",
  57432=>"010010011",
  57433=>"100110101",
  57434=>"000010000",
  57435=>"001111111",
  57436=>"011100011",
  57437=>"101000010",
  57438=>"100101110",
  57439=>"111111111",
  57440=>"111101001",
  57441=>"111101001",
  57442=>"111010001",
  57443=>"111110011",
  57444=>"101111000",
  57445=>"110111111",
  57446=>"111000101",
  57447=>"000111000",
  57448=>"110110001",
  57449=>"011100011",
  57450=>"011011000",
  57451=>"001101000",
  57452=>"010100011",
  57453=>"100001111",
  57454=>"111010011",
  57455=>"101111010",
  57456=>"101001111",
  57457=>"010101110",
  57458=>"111100110",
  57459=>"100110110",
  57460=>"100011111",
  57461=>"110101101",
  57462=>"001001010",
  57463=>"111111001",
  57464=>"100100001",
  57465=>"110010000",
  57466=>"111100111",
  57467=>"101100111",
  57468=>"000010000",
  57469=>"110100010",
  57470=>"001100110",
  57471=>"110110110",
  57472=>"011001101",
  57473=>"101010110",
  57474=>"110111010",
  57475=>"111111011",
  57476=>"100011000",
  57477=>"011111101",
  57478=>"000001000",
  57479=>"100100101",
  57480=>"010111110",
  57481=>"011010101",
  57482=>"110101001",
  57483=>"000001011",
  57484=>"001010000",
  57485=>"011000001",
  57486=>"100110010",
  57487=>"010111001",
  57488=>"000111010",
  57489=>"011010011",
  57490=>"110011011",
  57491=>"110001011",
  57492=>"111101111",
  57493=>"111111111",
  57494=>"100111111",
  57495=>"111110001",
  57496=>"001101110",
  57497=>"010000011",
  57498=>"100110000",
  57499=>"001111110",
  57500=>"101000001",
  57501=>"000100001",
  57502=>"101110010",
  57503=>"110111101",
  57504=>"110111010",
  57505=>"110010010",
  57506=>"101110101",
  57507=>"010011000",
  57508=>"010011010",
  57509=>"010100001",
  57510=>"110100101",
  57511=>"110100111",
  57512=>"111001010",
  57513=>"100001111",
  57514=>"100101011",
  57515=>"110110000",
  57516=>"110011001",
  57517=>"110111011",
  57518=>"011101111",
  57519=>"100001100",
  57520=>"110000000",
  57521=>"101111001",
  57522=>"011011001",
  57523=>"101000011",
  57524=>"101110011",
  57525=>"111111011",
  57526=>"111011000",
  57527=>"011001000",
  57528=>"010011101",
  57529=>"100110001",
  57530=>"010101010",
  57531=>"010000001",
  57532=>"100010110",
  57533=>"010100111",
  57534=>"011110111",
  57535=>"111101110",
  57536=>"000011001",
  57537=>"001111010",
  57538=>"001110101",
  57539=>"001110011",
  57540=>"110100011",
  57541=>"111100000",
  57542=>"000111100",
  57543=>"111110001",
  57544=>"101111001",
  57545=>"110110011",
  57546=>"010100110",
  57547=>"100110000",
  57548=>"110110110",
  57549=>"010111100",
  57550=>"011011000",
  57551=>"110101000",
  57552=>"101001000",
  57553=>"011001001",
  57554=>"000110111",
  57555=>"100010011",
  57556=>"101000011",
  57557=>"110010100",
  57558=>"011010010",
  57559=>"111110010",
  57560=>"101010000",
  57561=>"011001010",
  57562=>"010000001",
  57563=>"111011111",
  57564=>"001111101",
  57565=>"000010101",
  57566=>"111110001",
  57567=>"101000001",
  57568=>"110111001",
  57569=>"111001100",
  57570=>"111110101",
  57571=>"001010001",
  57572=>"111110001",
  57573=>"000110011",
  57574=>"111000101",
  57575=>"010111101",
  57576=>"010100010",
  57577=>"001011111",
  57578=>"110110011",
  57579=>"101101100",
  57580=>"101110111",
  57581=>"101100001",
  57582=>"000101111",
  57583=>"011010001",
  57584=>"010001101",
  57585=>"000101010",
  57586=>"110001010",
  57587=>"001010111",
  57588=>"111100110",
  57589=>"101111100",
  57590=>"001110111",
  57591=>"011101101",
  57592=>"111001111",
  57593=>"001100011",
  57594=>"001010111",
  57595=>"000001111",
  57596=>"101011000",
  57597=>"011011110",
  57598=>"111000001",
  57599=>"010101111",
  57600=>"011011000",
  57601=>"110101010",
  57602=>"110011110",
  57603=>"101010010",
  57604=>"100010010",
  57605=>"100010001",
  57606=>"001110010",
  57607=>"010110110",
  57608=>"101101101",
  57609=>"110110111",
  57610=>"111100000",
  57611=>"110100100",
  57612=>"100110100",
  57613=>"000001100",
  57614=>"000000000",
  57615=>"111101000",
  57616=>"011001001",
  57617=>"010110000",
  57618=>"111100010",
  57619=>"111000111",
  57620=>"101100100",
  57621=>"100000110",
  57622=>"100110000",
  57623=>"111001101",
  57624=>"111010111",
  57625=>"101101011",
  57626=>"011000000",
  57627=>"010110101",
  57628=>"110111110",
  57629=>"100111010",
  57630=>"101101000",
  57631=>"000100111",
  57632=>"010111010",
  57633=>"010000001",
  57634=>"101000100",
  57635=>"010011000",
  57636=>"000011100",
  57637=>"000000111",
  57638=>"010101001",
  57639=>"001010000",
  57640=>"000001100",
  57641=>"110110110",
  57642=>"010101111",
  57643=>"101100010",
  57644=>"001110000",
  57645=>"011001111",
  57646=>"111011011",
  57647=>"001100100",
  57648=>"001000100",
  57649=>"100001011",
  57650=>"010000111",
  57651=>"000110001",
  57652=>"010100011",
  57653=>"101101000",
  57654=>"000001111",
  57655=>"001011001",
  57656=>"101111001",
  57657=>"101010111",
  57658=>"100000000",
  57659=>"010000100",
  57660=>"101101001",
  57661=>"101110110",
  57662=>"011110011",
  57663=>"011100010",
  57664=>"001111100",
  57665=>"100010111",
  57666=>"111110111",
  57667=>"001100101",
  57668=>"010111110",
  57669=>"011101000",
  57670=>"000010011",
  57671=>"101011111",
  57672=>"011111001",
  57673=>"101101111",
  57674=>"010101111",
  57675=>"101001011",
  57676=>"011110110",
  57677=>"100011100",
  57678=>"000110111",
  57679=>"000010000",
  57680=>"000111100",
  57681=>"111001000",
  57682=>"110000000",
  57683=>"100111000",
  57684=>"000110100",
  57685=>"000100101",
  57686=>"001100111",
  57687=>"110010110",
  57688=>"101001101",
  57689=>"100111001",
  57690=>"100110110",
  57691=>"001100001",
  57692=>"011111100",
  57693=>"000001010",
  57694=>"110100110",
  57695=>"001100110",
  57696=>"110111001",
  57697=>"010000110",
  57698=>"110000010",
  57699=>"000110111",
  57700=>"100100000",
  57701=>"010110000",
  57702=>"000110010",
  57703=>"110101111",
  57704=>"010110010",
  57705=>"111101001",
  57706=>"110001101",
  57707=>"001110000",
  57708=>"000010010",
  57709=>"011110011",
  57710=>"101111000",
  57711=>"010111000",
  57712=>"100100000",
  57713=>"100101000",
  57714=>"111000010",
  57715=>"000101011",
  57716=>"001110101",
  57717=>"001100000",
  57718=>"010011011",
  57719=>"110011100",
  57720=>"101010101",
  57721=>"011111010",
  57722=>"110101010",
  57723=>"101010101",
  57724=>"000001000",
  57725=>"111011111",
  57726=>"011111101",
  57727=>"111101100",
  57728=>"000101000",
  57729=>"011110000",
  57730=>"000101110",
  57731=>"001011101",
  57732=>"110100110",
  57733=>"111011000",
  57734=>"011001000",
  57735=>"000010000",
  57736=>"000101001",
  57737=>"010001000",
  57738=>"101011100",
  57739=>"011100010",
  57740=>"010101111",
  57741=>"111110010",
  57742=>"010111011",
  57743=>"011100101",
  57744=>"010010011",
  57745=>"101111100",
  57746=>"100110000",
  57747=>"100010011",
  57748=>"010011000",
  57749=>"000101110",
  57750=>"001010101",
  57751=>"110000011",
  57752=>"111000000",
  57753=>"001101111",
  57754=>"101010101",
  57755=>"111010011",
  57756=>"000111010",
  57757=>"001001011",
  57758=>"110001010",
  57759=>"010001010",
  57760=>"101100000",
  57761=>"000001010",
  57762=>"110000000",
  57763=>"100010111",
  57764=>"100001101",
  57765=>"000010111",
  57766=>"001100001",
  57767=>"011111111",
  57768=>"101011110",
  57769=>"010100101",
  57770=>"000000101",
  57771=>"010001111",
  57772=>"000010001",
  57773=>"101011010",
  57774=>"111110000",
  57775=>"010101001",
  57776=>"111101111",
  57777=>"100100000",
  57778=>"100010111",
  57779=>"111111110",
  57780=>"101110111",
  57781=>"001010101",
  57782=>"110101101",
  57783=>"000011000",
  57784=>"000111111",
  57785=>"101011001",
  57786=>"000000110",
  57787=>"001110011",
  57788=>"110000010",
  57789=>"111100100",
  57790=>"011100011",
  57791=>"000111000",
  57792=>"101111111",
  57793=>"110010100",
  57794=>"001011011",
  57795=>"001010011",
  57796=>"101110111",
  57797=>"110101100",
  57798=>"110010000",
  57799=>"001111111",
  57800=>"001111010",
  57801=>"111001100",
  57802=>"001010000",
  57803=>"000001000",
  57804=>"100000110",
  57805=>"001010100",
  57806=>"000011110",
  57807=>"011100110",
  57808=>"110111000",
  57809=>"001101100",
  57810=>"110111111",
  57811=>"101100010",
  57812=>"110100110",
  57813=>"000100111",
  57814=>"000000000",
  57815=>"100011110",
  57816=>"000111001",
  57817=>"011000100",
  57818=>"111011110",
  57819=>"110110001",
  57820=>"100100011",
  57821=>"101000000",
  57822=>"000011000",
  57823=>"000000011",
  57824=>"101011111",
  57825=>"010111000",
  57826=>"011001101",
  57827=>"110110001",
  57828=>"011000011",
  57829=>"001001101",
  57830=>"010001111",
  57831=>"111011111",
  57832=>"110111111",
  57833=>"010011001",
  57834=>"011100000",
  57835=>"100111010",
  57836=>"110100111",
  57837=>"111111001",
  57838=>"010010000",
  57839=>"011010000",
  57840=>"101001011",
  57841=>"010010010",
  57842=>"111011101",
  57843=>"100000010",
  57844=>"010000111",
  57845=>"000000000",
  57846=>"010101110",
  57847=>"000011010",
  57848=>"101001010",
  57849=>"110100110",
  57850=>"110100101",
  57851=>"100000100",
  57852=>"101101111",
  57853=>"111101101",
  57854=>"001110000",
  57855=>"111110111",
  57856=>"110001000",
  57857=>"100000010",
  57858=>"110000100",
  57859=>"100110101",
  57860=>"001100000",
  57861=>"010101000",
  57862=>"100100010",
  57863=>"000011011",
  57864=>"000010010",
  57865=>"010011111",
  57866=>"011001001",
  57867=>"010110000",
  57868=>"010110101",
  57869=>"010100000",
  57870=>"111110110",
  57871=>"011101110",
  57872=>"001110000",
  57873=>"101100100",
  57874=>"100010000",
  57875=>"101000101",
  57876=>"000110111",
  57877=>"011111110",
  57878=>"001001000",
  57879=>"010001011",
  57880=>"111010100",
  57881=>"101001101",
  57882=>"101110010",
  57883=>"000111000",
  57884=>"011111111",
  57885=>"010011111",
  57886=>"010000110",
  57887=>"110000111",
  57888=>"001001000",
  57889=>"011001000",
  57890=>"101011011",
  57891=>"001001111",
  57892=>"000100000",
  57893=>"010011011",
  57894=>"011100010",
  57895=>"011101011",
  57896=>"000000101",
  57897=>"100010100",
  57898=>"100011010",
  57899=>"011111001",
  57900=>"001000001",
  57901=>"101000000",
  57902=>"011011111",
  57903=>"111000100",
  57904=>"111001001",
  57905=>"110111110",
  57906=>"111001011",
  57907=>"000111001",
  57908=>"000111010",
  57909=>"011111111",
  57910=>"000011011",
  57911=>"111110110",
  57912=>"111000101",
  57913=>"000001001",
  57914=>"010001001",
  57915=>"010010000",
  57916=>"101101100",
  57917=>"101110111",
  57918=>"011011101",
  57919=>"101001010",
  57920=>"010000011",
  57921=>"101010011",
  57922=>"000101001",
  57923=>"011011100",
  57924=>"001010101",
  57925=>"101111000",
  57926=>"001011100",
  57927=>"010111011",
  57928=>"001010101",
  57929=>"100111000",
  57930=>"100110001",
  57931=>"101010001",
  57932=>"110011011",
  57933=>"001101010",
  57934=>"000000011",
  57935=>"010110111",
  57936=>"001111111",
  57937=>"001111001",
  57938=>"101010101",
  57939=>"110101100",
  57940=>"111001101",
  57941=>"111110001",
  57942=>"110001110",
  57943=>"110011111",
  57944=>"111100000",
  57945=>"100110101",
  57946=>"010111100",
  57947=>"111011000",
  57948=>"010000101",
  57949=>"110101001",
  57950=>"111101000",
  57951=>"000011000",
  57952=>"110010110",
  57953=>"000000110",
  57954=>"001001111",
  57955=>"111001010",
  57956=>"001110011",
  57957=>"110101111",
  57958=>"000010111",
  57959=>"101011011",
  57960=>"100010010",
  57961=>"100011001",
  57962=>"100000101",
  57963=>"111101101",
  57964=>"000011100",
  57965=>"111010000",
  57966=>"111001000",
  57967=>"100000011",
  57968=>"110001110",
  57969=>"001111011",
  57970=>"000010011",
  57971=>"011010000",
  57972=>"010000000",
  57973=>"111011110",
  57974=>"011111101",
  57975=>"110010010",
  57976=>"101010101",
  57977=>"111000010",
  57978=>"010001000",
  57979=>"010000010",
  57980=>"000000100",
  57981=>"011000100",
  57982=>"111111001",
  57983=>"100111000",
  57984=>"101001101",
  57985=>"010001001",
  57986=>"100011110",
  57987=>"101101101",
  57988=>"101101110",
  57989=>"110101111",
  57990=>"011001101",
  57991=>"010101110",
  57992=>"111101011",
  57993=>"001100000",
  57994=>"001111111",
  57995=>"001010011",
  57996=>"100100010",
  57997=>"101000101",
  57998=>"010001010",
  57999=>"010100100",
  58000=>"000111110",
  58001=>"110111000",
  58002=>"101011111",
  58003=>"101010101",
  58004=>"011010010",
  58005=>"000101000",
  58006=>"101111100",
  58007=>"011011101",
  58008=>"011011001",
  58009=>"010010110",
  58010=>"100111001",
  58011=>"001100101",
  58012=>"010011000",
  58013=>"111110111",
  58014=>"011110010",
  58015=>"101010110",
  58016=>"100100100",
  58017=>"100000001",
  58018=>"011101011",
  58019=>"001110110",
  58020=>"010001110",
  58021=>"000000100",
  58022=>"100111001",
  58023=>"000001100",
  58024=>"010000111",
  58025=>"011110111",
  58026=>"000100010",
  58027=>"000011000",
  58028=>"000101100",
  58029=>"101101101",
  58030=>"000100100",
  58031=>"101000000",
  58032=>"010110000",
  58033=>"101101000",
  58034=>"101010111",
  58035=>"001011010",
  58036=>"101000010",
  58037=>"010011010",
  58038=>"010111001",
  58039=>"010000010",
  58040=>"010100001",
  58041=>"001111011",
  58042=>"100101111",
  58043=>"010100110",
  58044=>"000001011",
  58045=>"111111100",
  58046=>"101111111",
  58047=>"010110111",
  58048=>"110110000",
  58049=>"111010110",
  58050=>"101010000",
  58051=>"110111001",
  58052=>"010111110",
  58053=>"101010011",
  58054=>"001101111",
  58055=>"010001010",
  58056=>"011000000",
  58057=>"011100111",
  58058=>"010100010",
  58059=>"110011110",
  58060=>"011001011",
  58061=>"000110011",
  58062=>"010100101",
  58063=>"001111011",
  58064=>"101100101",
  58065=>"110000100",
  58066=>"101110001",
  58067=>"011011100",
  58068=>"000000110",
  58069=>"111000000",
  58070=>"110011100",
  58071=>"101100000",
  58072=>"010100000",
  58073=>"110101001",
  58074=>"001001000",
  58075=>"010111000",
  58076=>"101101010",
  58077=>"011110111",
  58078=>"110010110",
  58079=>"010100111",
  58080=>"111000000",
  58081=>"111101111",
  58082=>"110000010",
  58083=>"000000110",
  58084=>"000110100",
  58085=>"000111011",
  58086=>"011100110",
  58087=>"010110110",
  58088=>"101011000",
  58089=>"001011100",
  58090=>"011110100",
  58091=>"011010111",
  58092=>"010111010",
  58093=>"011010101",
  58094=>"001001100",
  58095=>"001111100",
  58096=>"110101111",
  58097=>"100100000",
  58098=>"000110000",
  58099=>"000110101",
  58100=>"110010000",
  58101=>"111000001",
  58102=>"111110101",
  58103=>"011101110",
  58104=>"000100101",
  58105=>"011111101",
  58106=>"110010011",
  58107=>"101011100",
  58108=>"000101000",
  58109=>"000100111",
  58110=>"011110011",
  58111=>"101101100",
  58112=>"110111101",
  58113=>"111111110",
  58114=>"011000011",
  58115=>"111110001",
  58116=>"110010011",
  58117=>"000100111",
  58118=>"111100000",
  58119=>"000100110",
  58120=>"010100010",
  58121=>"001101011",
  58122=>"010110010",
  58123=>"100011011",
  58124=>"111110110",
  58125=>"001000001",
  58126=>"110011011",
  58127=>"110101101",
  58128=>"100011110",
  58129=>"101101100",
  58130=>"001101101",
  58131=>"111111011",
  58132=>"100101101",
  58133=>"011000001",
  58134=>"001111100",
  58135=>"000100000",
  58136=>"110100000",
  58137=>"000001000",
  58138=>"111011011",
  58139=>"100001111",
  58140=>"101011100",
  58141=>"100010101",
  58142=>"111001001",
  58143=>"010111111",
  58144=>"110101000",
  58145=>"101000010",
  58146=>"101110010",
  58147=>"101011111",
  58148=>"101011100",
  58149=>"101001111",
  58150=>"000010010",
  58151=>"110100100",
  58152=>"000111011",
  58153=>"011000011",
  58154=>"111111101",
  58155=>"010000111",
  58156=>"001010010",
  58157=>"110001001",
  58158=>"100101101",
  58159=>"111100100",
  58160=>"011111100",
  58161=>"100111111",
  58162=>"100101111",
  58163=>"000001001",
  58164=>"001111010",
  58165=>"111101011",
  58166=>"101010111",
  58167=>"010000000",
  58168=>"010010100",
  58169=>"010000100",
  58170=>"000100000",
  58171=>"000111110",
  58172=>"111011011",
  58173=>"110110111",
  58174=>"110110100",
  58175=>"101011010",
  58176=>"100011100",
  58177=>"011110000",
  58178=>"010111000",
  58179=>"000111100",
  58180=>"001100101",
  58181=>"111011101",
  58182=>"011101111",
  58183=>"000100101",
  58184=>"111110111",
  58185=>"000000110",
  58186=>"110110111",
  58187=>"011110111",
  58188=>"110100101",
  58189=>"010010000",
  58190=>"111011011",
  58191=>"101111001",
  58192=>"100101111",
  58193=>"001111101",
  58194=>"110001110",
  58195=>"111000100",
  58196=>"000000111",
  58197=>"100011001",
  58198=>"001011000",
  58199=>"010000100",
  58200=>"101110100",
  58201=>"110111000",
  58202=>"000100110",
  58203=>"101101100",
  58204=>"110010100",
  58205=>"010011011",
  58206=>"001100110",
  58207=>"111111110",
  58208=>"000011111",
  58209=>"000011111",
  58210=>"001110001",
  58211=>"011001100",
  58212=>"111010111",
  58213=>"100110110",
  58214=>"100100011",
  58215=>"001000110",
  58216=>"110111111",
  58217=>"100101001",
  58218=>"111000100",
  58219=>"001100110",
  58220=>"111101100",
  58221=>"000001001",
  58222=>"101010110",
  58223=>"011100011",
  58224=>"011010110",
  58225=>"000001001",
  58226=>"001000111",
  58227=>"000001101",
  58228=>"111000000",
  58229=>"011111010",
  58230=>"011111010",
  58231=>"001110011",
  58232=>"110111011",
  58233=>"101000001",
  58234=>"000010110",
  58235=>"111100100",
  58236=>"111101100",
  58237=>"000001010",
  58238=>"101101010",
  58239=>"110101010",
  58240=>"011101100",
  58241=>"010101110",
  58242=>"000110010",
  58243=>"101111110",
  58244=>"100100010",
  58245=>"101110101",
  58246=>"011000000",
  58247=>"001001100",
  58248=>"011000000",
  58249=>"100111010",
  58250=>"101001000",
  58251=>"001000001",
  58252=>"111000011",
  58253=>"111001111",
  58254=>"101011101",
  58255=>"000010000",
  58256=>"000100100",
  58257=>"001011101",
  58258=>"110000100",
  58259=>"010011111",
  58260=>"110000100",
  58261=>"101000001",
  58262=>"101001101",
  58263=>"011011010",
  58264=>"111110010",
  58265=>"101011000",
  58266=>"010011110",
  58267=>"000111011",
  58268=>"101011111",
  58269=>"111101000",
  58270=>"011101101",
  58271=>"110010110",
  58272=>"000001010",
  58273=>"000101110",
  58274=>"000000100",
  58275=>"101111011",
  58276=>"001001111",
  58277=>"000101100",
  58278=>"001000001",
  58279=>"101011010",
  58280=>"101001110",
  58281=>"010110100",
  58282=>"101100010",
  58283=>"011100000",
  58284=>"110001101",
  58285=>"101100010",
  58286=>"111100110",
  58287=>"111111101",
  58288=>"011010110",
  58289=>"001011011",
  58290=>"111111111",
  58291=>"011010011",
  58292=>"010000110",
  58293=>"111000010",
  58294=>"010111110",
  58295=>"110000000",
  58296=>"101001111",
  58297=>"001000000",
  58298=>"001011000",
  58299=>"010111111",
  58300=>"010001000",
  58301=>"101111101",
  58302=>"001011110",
  58303=>"101011101",
  58304=>"100101010",
  58305=>"000001110",
  58306=>"101010101",
  58307=>"111001110",
  58308=>"000011111",
  58309=>"111000111",
  58310=>"101101101",
  58311=>"111100000",
  58312=>"111101100",
  58313=>"101000010",
  58314=>"111100100",
  58315=>"101100110",
  58316=>"001101011",
  58317=>"101101000",
  58318=>"010111111",
  58319=>"101011110",
  58320=>"100010000",
  58321=>"010000101",
  58322=>"110001011",
  58323=>"110111110",
  58324=>"101011101",
  58325=>"111111100",
  58326=>"101000001",
  58327=>"101001100",
  58328=>"000000011",
  58329=>"111100100",
  58330=>"010010111",
  58331=>"110100000",
  58332=>"010001000",
  58333=>"010010101",
  58334=>"010100101",
  58335=>"110011000",
  58336=>"001001111",
  58337=>"101100001",
  58338=>"110001011",
  58339=>"011001100",
  58340=>"111111001",
  58341=>"101110111",
  58342=>"100000000",
  58343=>"010010111",
  58344=>"001010100",
  58345=>"000000010",
  58346=>"000000100",
  58347=>"100101100",
  58348=>"101010111",
  58349=>"100000011",
  58350=>"100000100",
  58351=>"011110011",
  58352=>"111011111",
  58353=>"011011010",
  58354=>"000101010",
  58355=>"001011100",
  58356=>"011100001",
  58357=>"111110000",
  58358=>"110011110",
  58359=>"101110000",
  58360=>"111100000",
  58361=>"000100001",
  58362=>"101110111",
  58363=>"001100111",
  58364=>"101010010",
  58365=>"000011100",
  58366=>"000110000",
  58367=>"100000000",
  58368=>"010110010",
  58369=>"111011101",
  58370=>"010111101",
  58371=>"010111011",
  58372=>"011110000",
  58373=>"010000010",
  58374=>"100100100",
  58375=>"101011101",
  58376=>"011001101",
  58377=>"010000001",
  58378=>"110110100",
  58379=>"010100110",
  58380=>"000010010",
  58381=>"011111100",
  58382=>"000000101",
  58383=>"000010000",
  58384=>"011111010",
  58385=>"001110001",
  58386=>"000100110",
  58387=>"010011001",
  58388=>"111001011",
  58389=>"001000000",
  58390=>"100000011",
  58391=>"010101011",
  58392=>"111101100",
  58393=>"110011011",
  58394=>"000000000",
  58395=>"000001010",
  58396=>"110000111",
  58397=>"111001100",
  58398=>"110000001",
  58399=>"001000110",
  58400=>"101101101",
  58401=>"100101011",
  58402=>"101000110",
  58403=>"011100100",
  58404=>"011010001",
  58405=>"100110101",
  58406=>"111001110",
  58407=>"001011000",
  58408=>"100101010",
  58409=>"010110110",
  58410=>"010111001",
  58411=>"011001100",
  58412=>"000001000",
  58413=>"111000000",
  58414=>"000111110",
  58415=>"100100011",
  58416=>"100010000",
  58417=>"100011010",
  58418=>"010001001",
  58419=>"101101101",
  58420=>"101000101",
  58421=>"001110010",
  58422=>"110111101",
  58423=>"011111001",
  58424=>"010001101",
  58425=>"100100001",
  58426=>"100011001",
  58427=>"011110111",
  58428=>"010001101",
  58429=>"100101110",
  58430=>"101100000",
  58431=>"001010100",
  58432=>"010011010",
  58433=>"001000010",
  58434=>"011010011",
  58435=>"101001010",
  58436=>"000000000",
  58437=>"001111100",
  58438=>"111001000",
  58439=>"110100110",
  58440=>"101110100",
  58441=>"001110001",
  58442=>"000001000",
  58443=>"011111010",
  58444=>"101001110",
  58445=>"001100110",
  58446=>"111101100",
  58447=>"011000100",
  58448=>"100001101",
  58449=>"110010111",
  58450=>"101100111",
  58451=>"111001100",
  58452=>"000010111",
  58453=>"010001000",
  58454=>"011011111",
  58455=>"110110100",
  58456=>"110100001",
  58457=>"101111110",
  58458=>"000001111",
  58459=>"110000000",
  58460=>"000101000",
  58461=>"110001111",
  58462=>"000010010",
  58463=>"000001111",
  58464=>"001001000",
  58465=>"111101001",
  58466=>"011011100",
  58467=>"100000000",
  58468=>"000000011",
  58469=>"011110110",
  58470=>"100011001",
  58471=>"011110000",
  58472=>"000101001",
  58473=>"100101000",
  58474=>"101101110",
  58475=>"100001101",
  58476=>"110000110",
  58477=>"011111100",
  58478=>"100100001",
  58479=>"101100001",
  58480=>"111000010",
  58481=>"111101001",
  58482=>"010000101",
  58483=>"001101010",
  58484=>"011111010",
  58485=>"010100001",
  58486=>"100000001",
  58487=>"010000011",
  58488=>"100001101",
  58489=>"110100101",
  58490=>"011010100",
  58491=>"100000101",
  58492=>"100101111",
  58493=>"000110111",
  58494=>"000101111",
  58495=>"000000010",
  58496=>"011000010",
  58497=>"011000111",
  58498=>"010101100",
  58499=>"010000000",
  58500=>"001101111",
  58501=>"101000110",
  58502=>"111101001",
  58503=>"010011011",
  58504=>"100110000",
  58505=>"000110110",
  58506=>"010001001",
  58507=>"010101101",
  58508=>"101001001",
  58509=>"111101011",
  58510=>"000001110",
  58511=>"010000111",
  58512=>"111101000",
  58513=>"101011101",
  58514=>"010001000",
  58515=>"101001011",
  58516=>"110010100",
  58517=>"110010100",
  58518=>"001100010",
  58519=>"111111111",
  58520=>"111100001",
  58521=>"100011101",
  58522=>"011010000",
  58523=>"001111011",
  58524=>"110010001",
  58525=>"100101000",
  58526=>"011010000",
  58527=>"110111100",
  58528=>"011111101",
  58529=>"100001010",
  58530=>"101101011",
  58531=>"110010111",
  58532=>"111001110",
  58533=>"001011010",
  58534=>"011001110",
  58535=>"111010101",
  58536=>"001011010",
  58537=>"000010001",
  58538=>"110011111",
  58539=>"011000111",
  58540=>"101101010",
  58541=>"010000111",
  58542=>"011100000",
  58543=>"110100101",
  58544=>"010001110",
  58545=>"000101011",
  58546=>"111001010",
  58547=>"000000000",
  58548=>"001100110",
  58549=>"100001000",
  58550=>"110001110",
  58551=>"110010011",
  58552=>"000111111",
  58553=>"010101111",
  58554=>"000100010",
  58555=>"111000111",
  58556=>"111000100",
  58557=>"011000111",
  58558=>"100111100",
  58559=>"100110001",
  58560=>"111111111",
  58561=>"101001011",
  58562=>"000000101",
  58563=>"100111010",
  58564=>"100111011",
  58565=>"000100011",
  58566=>"011011001",
  58567=>"100000010",
  58568=>"110110010",
  58569=>"010100101",
  58570=>"000000101",
  58571=>"110010001",
  58572=>"001101101",
  58573=>"010100100",
  58574=>"001100001",
  58575=>"001010111",
  58576=>"111101100",
  58577=>"101010001",
  58578=>"101010000",
  58579=>"100001010",
  58580=>"101001010",
  58581=>"010101100",
  58582=>"011100110",
  58583=>"011110010",
  58584=>"011100110",
  58585=>"100110101",
  58586=>"100001001",
  58587=>"010100010",
  58588=>"101000000",
  58589=>"110011100",
  58590=>"000110000",
  58591=>"010111101",
  58592=>"110110011",
  58593=>"100011110",
  58594=>"011101110",
  58595=>"010011010",
  58596=>"101100101",
  58597=>"011011001",
  58598=>"100110111",
  58599=>"101111111",
  58600=>"101101100",
  58601=>"001111111",
  58602=>"100101111",
  58603=>"110111000",
  58604=>"000101011",
  58605=>"000101000",
  58606=>"000111100",
  58607=>"011001110",
  58608=>"001100011",
  58609=>"000000000",
  58610=>"111011001",
  58611=>"010000001",
  58612=>"001001100",
  58613=>"000101111",
  58614=>"011010010",
  58615=>"011101011",
  58616=>"000001110",
  58617=>"111000110",
  58618=>"000100011",
  58619=>"100001100",
  58620=>"110101110",
  58621=>"011110100",
  58622=>"000111110",
  58623=>"000100100",
  58624=>"100101100",
  58625=>"110111001",
  58626=>"100011000",
  58627=>"011111011",
  58628=>"101111011",
  58629=>"000110110",
  58630=>"100100000",
  58631=>"110100110",
  58632=>"010010010",
  58633=>"111110101",
  58634=>"000100111",
  58635=>"000010000",
  58636=>"011010001",
  58637=>"001000100",
  58638=>"110011001",
  58639=>"001000011",
  58640=>"011101110",
  58641=>"100011101",
  58642=>"010001010",
  58643=>"110100101",
  58644=>"010110100",
  58645=>"010000010",
  58646=>"001111001",
  58647=>"011101101",
  58648=>"011001111",
  58649=>"100001100",
  58650=>"000000001",
  58651=>"010111000",
  58652=>"100100001",
  58653=>"100100111",
  58654=>"111111111",
  58655=>"110110000",
  58656=>"001011111",
  58657=>"100100101",
  58658=>"011111110",
  58659=>"011101011",
  58660=>"000101111",
  58661=>"010111011",
  58662=>"110011100",
  58663=>"111100110",
  58664=>"010011011",
  58665=>"000100001",
  58666=>"110010110",
  58667=>"110000011",
  58668=>"011100000",
  58669=>"000000001",
  58670=>"101011011",
  58671=>"000000000",
  58672=>"001001100",
  58673=>"011101101",
  58674=>"000011000",
  58675=>"100110111",
  58676=>"001101001",
  58677=>"000111010",
  58678=>"000010001",
  58679=>"110001000",
  58680=>"111110100",
  58681=>"111000111",
  58682=>"110100010",
  58683=>"111110001",
  58684=>"101100111",
  58685=>"001101010",
  58686=>"011101100",
  58687=>"100101000",
  58688=>"101001011",
  58689=>"101100101",
  58690=>"011010101",
  58691=>"101111100",
  58692=>"001010010",
  58693=>"101001010",
  58694=>"001000110",
  58695=>"100100101",
  58696=>"100010011",
  58697=>"010001000",
  58698=>"001001000",
  58699=>"010000000",
  58700=>"100110011",
  58701=>"000101001",
  58702=>"110011111",
  58703=>"001100001",
  58704=>"001001011",
  58705=>"110111111",
  58706=>"101011110",
  58707=>"010100001",
  58708=>"000110001",
  58709=>"100000101",
  58710=>"101010000",
  58711=>"111011100",
  58712=>"111101011",
  58713=>"010010110",
  58714=>"010011101",
  58715=>"110011100",
  58716=>"101011110",
  58717=>"011001111",
  58718=>"111011010",
  58719=>"111000111",
  58720=>"111110101",
  58721=>"111000100",
  58722=>"111001000",
  58723=>"010001100",
  58724=>"110110010",
  58725=>"101000000",
  58726=>"001000111",
  58727=>"011110001",
  58728=>"001101101",
  58729=>"000010101",
  58730=>"011110111",
  58731=>"011000110",
  58732=>"100101010",
  58733=>"100101111",
  58734=>"010000000",
  58735=>"010110001",
  58736=>"101100111",
  58737=>"100110001",
  58738=>"111101110",
  58739=>"000111110",
  58740=>"000100000",
  58741=>"000110110",
  58742=>"010110011",
  58743=>"100001010",
  58744=>"000000000",
  58745=>"000001000",
  58746=>"101100001",
  58747=>"100011000",
  58748=>"101101110",
  58749=>"100011111",
  58750=>"011110011",
  58751=>"101110100",
  58752=>"001110011",
  58753=>"111101010",
  58754=>"101111110",
  58755=>"101111000",
  58756=>"110111101",
  58757=>"011111000",
  58758=>"110101000",
  58759=>"100001010",
  58760=>"001011001",
  58761=>"101001110",
  58762=>"000010000",
  58763=>"010111110",
  58764=>"000001011",
  58765=>"101001001",
  58766=>"110101001",
  58767=>"111110010",
  58768=>"110010011",
  58769=>"100111110",
  58770=>"000110111",
  58771=>"111010010",
  58772=>"101000011",
  58773=>"011000101",
  58774=>"101101000",
  58775=>"110100110",
  58776=>"010101000",
  58777=>"010010011",
  58778=>"101111110",
  58779=>"011011001",
  58780=>"110100010",
  58781=>"101001001",
  58782=>"001001001",
  58783=>"000011010",
  58784=>"101110000",
  58785=>"011111000",
  58786=>"000011011",
  58787=>"011001111",
  58788=>"100101010",
  58789=>"110101100",
  58790=>"100110011",
  58791=>"100000111",
  58792=>"000010110",
  58793=>"110101000",
  58794=>"111000000",
  58795=>"100000110",
  58796=>"100001011",
  58797=>"000011010",
  58798=>"001101000",
  58799=>"001010111",
  58800=>"111011100",
  58801=>"100111010",
  58802=>"111111100",
  58803=>"000110001",
  58804=>"110001100",
  58805=>"111000011",
  58806=>"110010101",
  58807=>"011111000",
  58808=>"010101110",
  58809=>"111011010",
  58810=>"111001111",
  58811=>"011001001",
  58812=>"101111110",
  58813=>"000110110",
  58814=>"000100001",
  58815=>"110100100",
  58816=>"111111011",
  58817=>"011111000",
  58818=>"111010111",
  58819=>"100110110",
  58820=>"111000101",
  58821=>"100010100",
  58822=>"101001001",
  58823=>"101111101",
  58824=>"000000100",
  58825=>"110011011",
  58826=>"001111110",
  58827=>"011001000",
  58828=>"011000011",
  58829=>"011011011",
  58830=>"001101000",
  58831=>"001111100",
  58832=>"010111111",
  58833=>"000010100",
  58834=>"011101010",
  58835=>"000000011",
  58836=>"001011000",
  58837=>"101001101",
  58838=>"100000111",
  58839=>"101101101",
  58840=>"110000100",
  58841=>"010001000",
  58842=>"100000100",
  58843=>"111110110",
  58844=>"101010111",
  58845=>"100110001",
  58846=>"001001111",
  58847=>"101000010",
  58848=>"101110110",
  58849=>"011101101",
  58850=>"100001010",
  58851=>"000101111",
  58852=>"011000100",
  58853=>"001000101",
  58854=>"000101011",
  58855=>"111011010",
  58856=>"010101111",
  58857=>"001110100",
  58858=>"100100011",
  58859=>"011000001",
  58860=>"100000100",
  58861=>"001110000",
  58862=>"101011111",
  58863=>"000010001",
  58864=>"101001111",
  58865=>"101010111",
  58866=>"011111001",
  58867=>"101001000",
  58868=>"000110101",
  58869=>"111110000",
  58870=>"010001001",
  58871=>"110010010",
  58872=>"100101011",
  58873=>"000001011",
  58874=>"100110110",
  58875=>"101010000",
  58876=>"001110100",
  58877=>"100101110",
  58878=>"010000111",
  58879=>"110000110",
  58880=>"010101111",
  58881=>"011110111",
  58882=>"011110110",
  58883=>"000111100",
  58884=>"000011001",
  58885=>"101000100",
  58886=>"001110000",
  58887=>"101111100",
  58888=>"011000110",
  58889=>"011001101",
  58890=>"010010100",
  58891=>"010001100",
  58892=>"111011101",
  58893=>"111100101",
  58894=>"111111001",
  58895=>"011011001",
  58896=>"001001111",
  58897=>"100101001",
  58898=>"001101111",
  58899=>"111001001",
  58900=>"100101101",
  58901=>"010010011",
  58902=>"011100000",
  58903=>"010110001",
  58904=>"111100110",
  58905=>"010101011",
  58906=>"000001000",
  58907=>"101000001",
  58908=>"100000101",
  58909=>"111001100",
  58910=>"001110000",
  58911=>"111111010",
  58912=>"010001001",
  58913=>"001111001",
  58914=>"011110111",
  58915=>"011101101",
  58916=>"010100110",
  58917=>"000000000",
  58918=>"111000010",
  58919=>"011111011",
  58920=>"001011000",
  58921=>"100110111",
  58922=>"111011011",
  58923=>"110101001",
  58924=>"001010110",
  58925=>"101000110",
  58926=>"110100000",
  58927=>"011111001",
  58928=>"010110000",
  58929=>"100001010",
  58930=>"001101010",
  58931=>"100010001",
  58932=>"110000000",
  58933=>"000111001",
  58934=>"111110001",
  58935=>"010101110",
  58936=>"000001100",
  58937=>"001001000",
  58938=>"000110010",
  58939=>"010010100",
  58940=>"000100101",
  58941=>"111011110",
  58942=>"111010000",
  58943=>"011100010",
  58944=>"010101101",
  58945=>"000011101",
  58946=>"001110011",
  58947=>"010000011",
  58948=>"010110110",
  58949=>"010000110",
  58950=>"001110000",
  58951=>"000001010",
  58952=>"000011010",
  58953=>"111001010",
  58954=>"100100111",
  58955=>"000101111",
  58956=>"101100100",
  58957=>"010100001",
  58958=>"101010110",
  58959=>"111000101",
  58960=>"011101100",
  58961=>"011001111",
  58962=>"000001000",
  58963=>"000010001",
  58964=>"101000101",
  58965=>"110001111",
  58966=>"110101110",
  58967=>"011111111",
  58968=>"010101011",
  58969=>"011001011",
  58970=>"111010111",
  58971=>"101001000",
  58972=>"111111001",
  58973=>"111110010",
  58974=>"001010101",
  58975=>"001100110",
  58976=>"011010001",
  58977=>"010011010",
  58978=>"010101111",
  58979=>"001010110",
  58980=>"001100011",
  58981=>"111011110",
  58982=>"000000110",
  58983=>"001000000",
  58984=>"010001101",
  58985=>"111101110",
  58986=>"001011000",
  58987=>"010101000",
  58988=>"000010101",
  58989=>"110100110",
  58990=>"111001001",
  58991=>"101001001",
  58992=>"101111011",
  58993=>"001010110",
  58994=>"011111110",
  58995=>"101001010",
  58996=>"111101001",
  58997=>"111011010",
  58998=>"011101001",
  58999=>"111101101",
  59000=>"110010101",
  59001=>"000101011",
  59002=>"110101010",
  59003=>"000110101",
  59004=>"101100101",
  59005=>"100000111",
  59006=>"001000101",
  59007=>"010110100",
  59008=>"011101111",
  59009=>"100001010",
  59010=>"010010010",
  59011=>"001100010",
  59012=>"111101010",
  59013=>"111000000",
  59014=>"111101000",
  59015=>"011010010",
  59016=>"101101100",
  59017=>"011001011",
  59018=>"001100010",
  59019=>"010110110",
  59020=>"001000010",
  59021=>"110100011",
  59022=>"100110000",
  59023=>"001111010",
  59024=>"101100011",
  59025=>"100011111",
  59026=>"110000111",
  59027=>"111100110",
  59028=>"101100111",
  59029=>"100000100",
  59030=>"111111000",
  59031=>"100100001",
  59032=>"000000100",
  59033=>"101011000",
  59034=>"001011001",
  59035=>"010111001",
  59036=>"010011111",
  59037=>"100000101",
  59038=>"101110110",
  59039=>"110100001",
  59040=>"011011011",
  59041=>"010000100",
  59042=>"011110100",
  59043=>"100110111",
  59044=>"101101101",
  59045=>"001011101",
  59046=>"011010110",
  59047=>"101110100",
  59048=>"001000011",
  59049=>"001101110",
  59050=>"100100110",
  59051=>"101011010",
  59052=>"011001000",
  59053=>"111000000",
  59054=>"111110010",
  59055=>"011000000",
  59056=>"010000011",
  59057=>"100110111",
  59058=>"001010101",
  59059=>"000001100",
  59060=>"110101110",
  59061=>"100000010",
  59062=>"010011000",
  59063=>"011110111",
  59064=>"000100111",
  59065=>"010001011",
  59066=>"011011001",
  59067=>"110101111",
  59068=>"111011110",
  59069=>"001000110",
  59070=>"101011101",
  59071=>"000011110",
  59072=>"110110010",
  59073=>"110010111",
  59074=>"010111010",
  59075=>"110001111",
  59076=>"110110111",
  59077=>"111010001",
  59078=>"001010100",
  59079=>"010110101",
  59080=>"001010100",
  59081=>"011010100",
  59082=>"011111111",
  59083=>"100011011",
  59084=>"011110011",
  59085=>"100001101",
  59086=>"111000111",
  59087=>"010011100",
  59088=>"100101100",
  59089=>"111000110",
  59090=>"010100000",
  59091=>"001101101",
  59092=>"100011100",
  59093=>"100001100",
  59094=>"101101000",
  59095=>"110010011",
  59096=>"100000010",
  59097=>"010101001",
  59098=>"100101011",
  59099=>"010010011",
  59100=>"101100111",
  59101=>"011110110",
  59102=>"010010101",
  59103=>"101011100",
  59104=>"010101010",
  59105=>"000111111",
  59106=>"100111100",
  59107=>"110100111",
  59108=>"100010000",
  59109=>"101000110",
  59110=>"000000110",
  59111=>"010110101",
  59112=>"000100101",
  59113=>"110100010",
  59114=>"001101111",
  59115=>"010001101",
  59116=>"110011011",
  59117=>"010001010",
  59118=>"010011100",
  59119=>"011011000",
  59120=>"101111001",
  59121=>"111010000",
  59122=>"011011010",
  59123=>"101110111",
  59124=>"000011101",
  59125=>"001101010",
  59126=>"010000000",
  59127=>"010000000",
  59128=>"000010010",
  59129=>"111011001",
  59130=>"110101100",
  59131=>"110101111",
  59132=>"011001001",
  59133=>"110101111",
  59134=>"100000000",
  59135=>"101100001",
  59136=>"010100101",
  59137=>"110110010",
  59138=>"001101111",
  59139=>"111100011",
  59140=>"011111011",
  59141=>"110100011",
  59142=>"100010010",
  59143=>"110101010",
  59144=>"101001101",
  59145=>"001101001",
  59146=>"010001000",
  59147=>"001100111",
  59148=>"101010100",
  59149=>"001010001",
  59150=>"010010011",
  59151=>"000110001",
  59152=>"110101000",
  59153=>"011010000",
  59154=>"101010111",
  59155=>"000011010",
  59156=>"010011111",
  59157=>"011000010",
  59158=>"011011011",
  59159=>"001101110",
  59160=>"010011001",
  59161=>"101100001",
  59162=>"000011101",
  59163=>"111000111",
  59164=>"011110100",
  59165=>"111000101",
  59166=>"000010101",
  59167=>"010010011",
  59168=>"010001011",
  59169=>"010000011",
  59170=>"000110010",
  59171=>"010001000",
  59172=>"011111111",
  59173=>"000101010",
  59174=>"010000010",
  59175=>"101101110",
  59176=>"010011010",
  59177=>"111101001",
  59178=>"000100101",
  59179=>"010100101",
  59180=>"011001101",
  59181=>"001010101",
  59182=>"001101011",
  59183=>"100111010",
  59184=>"110110110",
  59185=>"110001001",
  59186=>"000001010",
  59187=>"000000011",
  59188=>"100100010",
  59189=>"110111010",
  59190=>"001100010",
  59191=>"000010111",
  59192=>"110010000",
  59193=>"011000000",
  59194=>"000100110",
  59195=>"001001001",
  59196=>"010000010",
  59197=>"100001000",
  59198=>"100011001",
  59199=>"110001101",
  59200=>"010100101",
  59201=>"011101010",
  59202=>"111101011",
  59203=>"101011101",
  59204=>"000111110",
  59205=>"011111110",
  59206=>"010100110",
  59207=>"001000000",
  59208=>"011011001",
  59209=>"110011010",
  59210=>"100111110",
  59211=>"000000001",
  59212=>"010011011",
  59213=>"010111110",
  59214=>"100010100",
  59215=>"011111100",
  59216=>"101011110",
  59217=>"101011000",
  59218=>"111010010",
  59219=>"110001010",
  59220=>"111000101",
  59221=>"110010010",
  59222=>"011101000",
  59223=>"101001000",
  59224=>"001001010",
  59225=>"000010011",
  59226=>"111100110",
  59227=>"111101100",
  59228=>"011100111",
  59229=>"110010010",
  59230=>"000001001",
  59231=>"000111110",
  59232=>"101011111",
  59233=>"110000010",
  59234=>"011010001",
  59235=>"010000110",
  59236=>"001001011",
  59237=>"101000011",
  59238=>"100100011",
  59239=>"010111111",
  59240=>"101001100",
  59241=>"100110111",
  59242=>"111001010",
  59243=>"111111001",
  59244=>"010110100",
  59245=>"001000000",
  59246=>"110011001",
  59247=>"011011101",
  59248=>"100011010",
  59249=>"111011010",
  59250=>"001100110",
  59251=>"001001100",
  59252=>"101000100",
  59253=>"100000100",
  59254=>"010001111",
  59255=>"110101100",
  59256=>"000111010",
  59257=>"111010011",
  59258=>"011110010",
  59259=>"101111011",
  59260=>"101010001",
  59261=>"011111110",
  59262=>"111010110",
  59263=>"110000101",
  59264=>"000101100",
  59265=>"011110010",
  59266=>"111110101",
  59267=>"000001011",
  59268=>"111011000",
  59269=>"110100000",
  59270=>"110000111",
  59271=>"010010001",
  59272=>"100000101",
  59273=>"100101001",
  59274=>"000100010",
  59275=>"010001110",
  59276=>"100111110",
  59277=>"011001111",
  59278=>"101000111",
  59279=>"111111001",
  59280=>"110000100",
  59281=>"010111110",
  59282=>"100111110",
  59283=>"011011011",
  59284=>"101000100",
  59285=>"001010111",
  59286=>"000011110",
  59287=>"000001110",
  59288=>"001001011",
  59289=>"000101010",
  59290=>"010110101",
  59291=>"110100111",
  59292=>"010011111",
  59293=>"100010010",
  59294=>"110000000",
  59295=>"101010111",
  59296=>"111101001",
  59297=>"001101110",
  59298=>"001011000",
  59299=>"000011100",
  59300=>"100011010",
  59301=>"111110100",
  59302=>"000110100",
  59303=>"101110011",
  59304=>"101010011",
  59305=>"000011100",
  59306=>"000010110",
  59307=>"110110111",
  59308=>"101101100",
  59309=>"110101001",
  59310=>"100101101",
  59311=>"111111001",
  59312=>"000110101",
  59313=>"001110010",
  59314=>"001110111",
  59315=>"010000110",
  59316=>"110001001",
  59317=>"001111101",
  59318=>"110100100",
  59319=>"011010100",
  59320=>"110101011",
  59321=>"100010010",
  59322=>"001001010",
  59323=>"001111111",
  59324=>"110001101",
  59325=>"111110001",
  59326=>"100010000",
  59327=>"001000000",
  59328=>"100011001",
  59329=>"001100011",
  59330=>"010100101",
  59331=>"010110101",
  59332=>"001000001",
  59333=>"101110101",
  59334=>"110011011",
  59335=>"010011010",
  59336=>"100011100",
  59337=>"000110110",
  59338=>"100110111",
  59339=>"111001011",
  59340=>"000010100",
  59341=>"000100001",
  59342=>"000110110",
  59343=>"101001110",
  59344=>"001010110",
  59345=>"101100000",
  59346=>"010111111",
  59347=>"011000110",
  59348=>"101000110",
  59349=>"101000001",
  59350=>"111101011",
  59351=>"001001001",
  59352=>"101100001",
  59353=>"111111101",
  59354=>"100011000",
  59355=>"111101100",
  59356=>"110010011",
  59357=>"101100010",
  59358=>"010000001",
  59359=>"011001110",
  59360=>"111010010",
  59361=>"111100001",
  59362=>"101001010",
  59363=>"101100010",
  59364=>"001011001",
  59365=>"110001100",
  59366=>"100101101",
  59367=>"011111000",
  59368=>"011110100",
  59369=>"000100100",
  59370=>"010001101",
  59371=>"110011111",
  59372=>"111100010",
  59373=>"110110110",
  59374=>"111100010",
  59375=>"100011011",
  59376=>"010101000",
  59377=>"000001100",
  59378=>"001001011",
  59379=>"100111011",
  59380=>"110110111",
  59381=>"101100010",
  59382=>"001101010",
  59383=>"111100000",
  59384=>"101010110",
  59385=>"100010110",
  59386=>"001001100",
  59387=>"010001011",
  59388=>"000101000",
  59389=>"000011010",
  59390=>"011001110",
  59391=>"011110000",
  59392=>"000011001",
  59393=>"110011111",
  59394=>"101111100",
  59395=>"111001111",
  59396=>"111000110",
  59397=>"000101010",
  59398=>"101100000",
  59399=>"001100111",
  59400=>"000011000",
  59401=>"111001101",
  59402=>"111010110",
  59403=>"011011001",
  59404=>"011010011",
  59405=>"100001001",
  59406=>"001010111",
  59407=>"000011011",
  59408=>"000001011",
  59409=>"010101010",
  59410=>"111101111",
  59411=>"100001000",
  59412=>"011001001",
  59413=>"011000100",
  59414=>"111010110",
  59415=>"001001010",
  59416=>"000001100",
  59417=>"010110000",
  59418=>"001110110",
  59419=>"000111110",
  59420=>"111000110",
  59421=>"001010001",
  59422=>"101111001",
  59423=>"101101111",
  59424=>"101101110",
  59425=>"111101111",
  59426=>"001100000",
  59427=>"010101000",
  59428=>"000110011",
  59429=>"111000000",
  59430=>"010010010",
  59431=>"011101100",
  59432=>"110000000",
  59433=>"111110010",
  59434=>"001111000",
  59435=>"010101111",
  59436=>"110001111",
  59437=>"111011100",
  59438=>"110110101",
  59439=>"100100000",
  59440=>"110111011",
  59441=>"011110110",
  59442=>"100000011",
  59443=>"101101111",
  59444=>"000100111",
  59445=>"000001110",
  59446=>"010100110",
  59447=>"011011110",
  59448=>"111110011",
  59449=>"101011001",
  59450=>"011111010",
  59451=>"000001011",
  59452=>"010011100",
  59453=>"000010100",
  59454=>"011111110",
  59455=>"100010010",
  59456=>"000010100",
  59457=>"010001110",
  59458=>"110101110",
  59459=>"001001011",
  59460=>"000100001",
  59461=>"100000001",
  59462=>"000000000",
  59463=>"101100000",
  59464=>"101001101",
  59465=>"111010101",
  59466=>"101010110",
  59467=>"100010001",
  59468=>"111001011",
  59469=>"101110010",
  59470=>"100000010",
  59471=>"000110101",
  59472=>"110000100",
  59473=>"000011000",
  59474=>"010101010",
  59475=>"111010001",
  59476=>"101101001",
  59477=>"100000101",
  59478=>"110000100",
  59479=>"000100100",
  59480=>"101100010",
  59481=>"001100000",
  59482=>"000011011",
  59483=>"000000001",
  59484=>"000110000",
  59485=>"111101000",
  59486=>"111110111",
  59487=>"011000100",
  59488=>"111001111",
  59489=>"011011001",
  59490=>"100001010",
  59491=>"101100100",
  59492=>"110010010",
  59493=>"110001001",
  59494=>"010101001",
  59495=>"001111101",
  59496=>"010001010",
  59497=>"101110111",
  59498=>"111011001",
  59499=>"111110101",
  59500=>"000001010",
  59501=>"011000010",
  59502=>"010010010",
  59503=>"000111010",
  59504=>"011011110",
  59505=>"101101011",
  59506=>"000000111",
  59507=>"011011000",
  59508=>"011001000",
  59509=>"011111001",
  59510=>"111001011",
  59511=>"111110001",
  59512=>"110111110",
  59513=>"011101011",
  59514=>"010110000",
  59515=>"010011000",
  59516=>"111001110",
  59517=>"101001100",
  59518=>"000010000",
  59519=>"010110110",
  59520=>"011010010",
  59521=>"110101001",
  59522=>"001001001",
  59523=>"001000011",
  59524=>"001001001",
  59525=>"000110111",
  59526=>"000000011",
  59527=>"111111010",
  59528=>"110000111",
  59529=>"111101110",
  59530=>"001110110",
  59531=>"101101111",
  59532=>"101101100",
  59533=>"100100101",
  59534=>"110100101",
  59535=>"101111110",
  59536=>"000000001",
  59537=>"111101001",
  59538=>"100110010",
  59539=>"000001111",
  59540=>"010101111",
  59541=>"000110100",
  59542=>"010000001",
  59543=>"000000010",
  59544=>"000010100",
  59545=>"001111111",
  59546=>"000100001",
  59547=>"001100111",
  59548=>"000101111",
  59549=>"010010100",
  59550=>"101011101",
  59551=>"000110000",
  59552=>"010011000",
  59553=>"111100111",
  59554=>"110010111",
  59555=>"001100110",
  59556=>"001110010",
  59557=>"000110000",
  59558=>"001101110",
  59559=>"001101001",
  59560=>"000110001",
  59561=>"010010010",
  59562=>"100010110",
  59563=>"110011000",
  59564=>"101110110",
  59565=>"100011000",
  59566=>"101111000",
  59567=>"001110111",
  59568=>"001111111",
  59569=>"101110111",
  59570=>"101010100",
  59571=>"111101001",
  59572=>"000001001",
  59573=>"011011110",
  59574=>"011011100",
  59575=>"111100010",
  59576=>"110100001",
  59577=>"001000001",
  59578=>"111001010",
  59579=>"001110000",
  59580=>"111111110",
  59581=>"111101101",
  59582=>"001101001",
  59583=>"000000101",
  59584=>"101011110",
  59585=>"110101010",
  59586=>"000010011",
  59587=>"111110110",
  59588=>"110101000",
  59589=>"111100001",
  59590=>"111000011",
  59591=>"010101001",
  59592=>"100110110",
  59593=>"111010011",
  59594=>"010010000",
  59595=>"011111001",
  59596=>"011111100",
  59597=>"100001100",
  59598=>"010010011",
  59599=>"110100101",
  59600=>"001110101",
  59601=>"010101011",
  59602=>"100110111",
  59603=>"001100111",
  59604=>"101111110",
  59605=>"001010100",
  59606=>"000101100",
  59607=>"101110100",
  59608=>"001001111",
  59609=>"010011111",
  59610=>"100110111",
  59611=>"000000001",
  59612=>"101110101",
  59613=>"011011001",
  59614=>"001001001",
  59615=>"110111100",
  59616=>"110100001",
  59617=>"010010000",
  59618=>"011110001",
  59619=>"011111001",
  59620=>"000011011",
  59621=>"101110100",
  59622=>"101000111",
  59623=>"000100010",
  59624=>"010100101",
  59625=>"000010111",
  59626=>"100110110",
  59627=>"000101110",
  59628=>"011011010",
  59629=>"101000100",
  59630=>"001011110",
  59631=>"100111111",
  59632=>"010001100",
  59633=>"100101111",
  59634=>"000000011",
  59635=>"000111010",
  59636=>"000100001",
  59637=>"010101101",
  59638=>"011001001",
  59639=>"001000000",
  59640=>"111111100",
  59641=>"100000100",
  59642=>"110101010",
  59643=>"111110101",
  59644=>"000111101",
  59645=>"111001001",
  59646=>"011100000",
  59647=>"011100110",
  59648=>"010100101",
  59649=>"010010100",
  59650=>"110110101",
  59651=>"110111010",
  59652=>"011011000",
  59653=>"000001100",
  59654=>"100000110",
  59655=>"111100110",
  59656=>"001001010",
  59657=>"001001110",
  59658=>"011001000",
  59659=>"001110011",
  59660=>"010111000",
  59661=>"010011001",
  59662=>"000010011",
  59663=>"000101101",
  59664=>"101111111",
  59665=>"101100101",
  59666=>"000010000",
  59667=>"000111111",
  59668=>"110100010",
  59669=>"001010001",
  59670=>"101100000",
  59671=>"101001001",
  59672=>"111000001",
  59673=>"010111110",
  59674=>"110111100",
  59675=>"010000010",
  59676=>"011000000",
  59677=>"111111011",
  59678=>"111011100",
  59679=>"101001000",
  59680=>"110010011",
  59681=>"000101111",
  59682=>"010111010",
  59683=>"001101101",
  59684=>"100111111",
  59685=>"100110101",
  59686=>"111101111",
  59687=>"100001010",
  59688=>"111011111",
  59689=>"110001100",
  59690=>"111000101",
  59691=>"011110010",
  59692=>"011101111",
  59693=>"101111000",
  59694=>"101110001",
  59695=>"101010001",
  59696=>"000011011",
  59697=>"100100011",
  59698=>"111111010",
  59699=>"111000001",
  59700=>"011111111",
  59701=>"111011000",
  59702=>"111001111",
  59703=>"100110111",
  59704=>"000000010",
  59705=>"111110111",
  59706=>"011010111",
  59707=>"000011110",
  59708=>"100101001",
  59709=>"101000000",
  59710=>"010001101",
  59711=>"110111101",
  59712=>"011111000",
  59713=>"101011001",
  59714=>"110111000",
  59715=>"000101100",
  59716=>"011011000",
  59717=>"011110010",
  59718=>"011001110",
  59719=>"111000101",
  59720=>"111110110",
  59721=>"110100111",
  59722=>"001101001",
  59723=>"110001101",
  59724=>"100100001",
  59725=>"100111101",
  59726=>"100110111",
  59727=>"001010111",
  59728=>"100000011",
  59729=>"011001001",
  59730=>"010110010",
  59731=>"110000000",
  59732=>"110010111",
  59733=>"101001010",
  59734=>"111111111",
  59735=>"001101010",
  59736=>"000000110",
  59737=>"010100001",
  59738=>"110000101",
  59739=>"011101001",
  59740=>"000110001",
  59741=>"111011100",
  59742=>"100111111",
  59743=>"111110011",
  59744=>"111100100",
  59745=>"000011110",
  59746=>"000000000",
  59747=>"011100011",
  59748=>"000010000",
  59749=>"101011110",
  59750=>"010011010",
  59751=>"101101000",
  59752=>"110011111",
  59753=>"000010100",
  59754=>"111101011",
  59755=>"101110001",
  59756=>"110101010",
  59757=>"001110111",
  59758=>"010000000",
  59759=>"111100001",
  59760=>"110001100",
  59761=>"001011100",
  59762=>"000110011",
  59763=>"110111110",
  59764=>"000011000",
  59765=>"101010111",
  59766=>"011101011",
  59767=>"110111111",
  59768=>"111100010",
  59769=>"111110011",
  59770=>"011101011",
  59771=>"100111110",
  59772=>"100111100",
  59773=>"110111010",
  59774=>"111001101",
  59775=>"010010011",
  59776=>"000111110",
  59777=>"111000111",
  59778=>"101011110",
  59779=>"101100110",
  59780=>"000101110",
  59781=>"100100110",
  59782=>"001001011",
  59783=>"011100101",
  59784=>"000000101",
  59785=>"011011001",
  59786=>"011011111",
  59787=>"111100101",
  59788=>"011111000",
  59789=>"001100101",
  59790=>"000001110",
  59791=>"000001001",
  59792=>"110111011",
  59793=>"000000000",
  59794=>"000110101",
  59795=>"100101101",
  59796=>"010000111",
  59797=>"001110110",
  59798=>"000101111",
  59799=>"101011101",
  59800=>"110010011",
  59801=>"001010010",
  59802=>"001000010",
  59803=>"010011101",
  59804=>"100111000",
  59805=>"011000001",
  59806=>"101011101",
  59807=>"010110000",
  59808=>"101010000",
  59809=>"111101010",
  59810=>"100100000",
  59811=>"000000001",
  59812=>"110011011",
  59813=>"000001001",
  59814=>"011011000",
  59815=>"001001000",
  59816=>"010110100",
  59817=>"100111000",
  59818=>"100010000",
  59819=>"111011010",
  59820=>"000011111",
  59821=>"111010100",
  59822=>"111100101",
  59823=>"011101001",
  59824=>"100010010",
  59825=>"110100001",
  59826=>"111100111",
  59827=>"000010110",
  59828=>"001011010",
  59829=>"110001110",
  59830=>"001100111",
  59831=>"111111111",
  59832=>"101111100",
  59833=>"111100111",
  59834=>"100100001",
  59835=>"001101001",
  59836=>"011111011",
  59837=>"001100010",
  59838=>"001000010",
  59839=>"100110100",
  59840=>"101110010",
  59841=>"011100011",
  59842=>"111111001",
  59843=>"101111111",
  59844=>"110101111",
  59845=>"011100111",
  59846=>"000100110",
  59847=>"111101011",
  59848=>"111110100",
  59849=>"011100111",
  59850=>"000111111",
  59851=>"011010111",
  59852=>"100011001",
  59853=>"011110010",
  59854=>"000001101",
  59855=>"011011001",
  59856=>"100111011",
  59857=>"101000010",
  59858=>"000110110",
  59859=>"111011101",
  59860=>"011011111",
  59861=>"111010111",
  59862=>"000110001",
  59863=>"010100000",
  59864=>"111111001",
  59865=>"001110000",
  59866=>"111011111",
  59867=>"111011001",
  59868=>"101101001",
  59869=>"110001101",
  59870=>"010011011",
  59871=>"110011110",
  59872=>"101000001",
  59873=>"011111000",
  59874=>"010111110",
  59875=>"110000110",
  59876=>"001100100",
  59877=>"101100111",
  59878=>"100001000",
  59879=>"101001100",
  59880=>"010000001",
  59881=>"010010111",
  59882=>"000101100",
  59883=>"111101001",
  59884=>"110011000",
  59885=>"110001101",
  59886=>"011011101",
  59887=>"010101101",
  59888=>"101010001",
  59889=>"011110010",
  59890=>"010011010",
  59891=>"110100001",
  59892=>"001000100",
  59893=>"010001101",
  59894=>"100101111",
  59895=>"110000100",
  59896=>"000000110",
  59897=>"111000001",
  59898=>"110110111",
  59899=>"010111010",
  59900=>"001110111",
  59901=>"101011111",
  59902=>"110111011",
  59903=>"111100101",
  59904=>"110011001",
  59905=>"010110001",
  59906=>"001110100",
  59907=>"111110100",
  59908=>"010111001",
  59909=>"001010100",
  59910=>"001111010",
  59911=>"110111010",
  59912=>"100001000",
  59913=>"000001001",
  59914=>"100110011",
  59915=>"111011000",
  59916=>"001110011",
  59917=>"111001001",
  59918=>"111111011",
  59919=>"000011101",
  59920=>"011111111",
  59921=>"000000011",
  59922=>"001101010",
  59923=>"100001000",
  59924=>"010001111",
  59925=>"011001101",
  59926=>"000111110",
  59927=>"111000111",
  59928=>"000010010",
  59929=>"100100011",
  59930=>"111010111",
  59931=>"000111100",
  59932=>"101111010",
  59933=>"010010101",
  59934=>"110001110",
  59935=>"001101001",
  59936=>"001111111",
  59937=>"000101001",
  59938=>"110101101",
  59939=>"001110001",
  59940=>"101000111",
  59941=>"101001100",
  59942=>"000110100",
  59943=>"110111001",
  59944=>"101011010",
  59945=>"100111010",
  59946=>"100100000",
  59947=>"100010101",
  59948=>"101100001",
  59949=>"100011100",
  59950=>"010001011",
  59951=>"101010010",
  59952=>"000010111",
  59953=>"100001011",
  59954=>"110100010",
  59955=>"000010101",
  59956=>"101110010",
  59957=>"101101110",
  59958=>"000010000",
  59959=>"111111010",
  59960=>"110110111",
  59961=>"100101011",
  59962=>"001101010",
  59963=>"111001000",
  59964=>"101010110",
  59965=>"010011110",
  59966=>"111011010",
  59967=>"101010000",
  59968=>"001001000",
  59969=>"001100001",
  59970=>"100001111",
  59971=>"010010000",
  59972=>"001010010",
  59973=>"110111111",
  59974=>"000010000",
  59975=>"111010000",
  59976=>"011011001",
  59977=>"001000110",
  59978=>"011111010",
  59979=>"111101100",
  59980=>"111001100",
  59981=>"011010000",
  59982=>"111101101",
  59983=>"011111011",
  59984=>"010101011",
  59985=>"010111011",
  59986=>"101101100",
  59987=>"001011001",
  59988=>"001011000",
  59989=>"101101000",
  59990=>"010001011",
  59991=>"101111011",
  59992=>"101110111",
  59993=>"111101000",
  59994=>"001101100",
  59995=>"000100000",
  59996=>"111001001",
  59997=>"101010111",
  59998=>"100011011",
  59999=>"010011010",
  60000=>"000000001",
  60001=>"001110101",
  60002=>"000010001",
  60003=>"001011101",
  60004=>"100100110",
  60005=>"110000010",
  60006=>"100011111",
  60007=>"111110011",
  60008=>"100110101",
  60009=>"010011110",
  60010=>"000011001",
  60011=>"010110000",
  60012=>"001011100",
  60013=>"010000110",
  60014=>"011111010",
  60015=>"111001101",
  60016=>"111111101",
  60017=>"011110100",
  60018=>"011100001",
  60019=>"001110010",
  60020=>"111101110",
  60021=>"100010100",
  60022=>"010000010",
  60023=>"101101101",
  60024=>"010001101",
  60025=>"100000010",
  60026=>"000010010",
  60027=>"000000110",
  60028=>"001001100",
  60029=>"110110101",
  60030=>"111101100",
  60031=>"111000011",
  60032=>"101001011",
  60033=>"010001101",
  60034=>"111010001",
  60035=>"101001001",
  60036=>"001011001",
  60037=>"110000101",
  60038=>"101000100",
  60039=>"000011110",
  60040=>"011010100",
  60041=>"110101111",
  60042=>"100111010",
  60043=>"000110101",
  60044=>"011111100",
  60045=>"101010011",
  60046=>"100001000",
  60047=>"101111001",
  60048=>"000110110",
  60049=>"100100111",
  60050=>"010010100",
  60051=>"110011000",
  60052=>"100111000",
  60053=>"001001110",
  60054=>"000100001",
  60055=>"110001000",
  60056=>"101011110",
  60057=>"001110000",
  60058=>"100000110",
  60059=>"001110011",
  60060=>"111100100",
  60061=>"111111000",
  60062=>"001101011",
  60063=>"110001001",
  60064=>"010110000",
  60065=>"001011001",
  60066=>"101010001",
  60067=>"010000011",
  60068=>"110011110",
  60069=>"110110111",
  60070=>"100101111",
  60071=>"110100100",
  60072=>"101001011",
  60073=>"000010000",
  60074=>"000001011",
  60075=>"110100010",
  60076=>"110100000",
  60077=>"100001001",
  60078=>"110000100",
  60079=>"001101101",
  60080=>"011001101",
  60081=>"000100111",
  60082=>"110010011",
  60083=>"011010001",
  60084=>"010001010",
  60085=>"010011001",
  60086=>"110011011",
  60087=>"101001101",
  60088=>"010000101",
  60089=>"001110001",
  60090=>"010000011",
  60091=>"100111001",
  60092=>"001010010",
  60093=>"101000100",
  60094=>"001000011",
  60095=>"101110010",
  60096=>"001111000",
  60097=>"011101111",
  60098=>"011010101",
  60099=>"111001110",
  60100=>"110000011",
  60101=>"000010011",
  60102=>"001000100",
  60103=>"000011100",
  60104=>"101011100",
  60105=>"111110111",
  60106=>"111011001",
  60107=>"011010000",
  60108=>"000000010",
  60109=>"001111001",
  60110=>"111011001",
  60111=>"011010110",
  60112=>"111101111",
  60113=>"011010000",
  60114=>"011100011",
  60115=>"001011011",
  60116=>"100000001",
  60117=>"111010101",
  60118=>"110101010",
  60119=>"010111001",
  60120=>"000001111",
  60121=>"001000010",
  60122=>"101001110",
  60123=>"000011001",
  60124=>"000011000",
  60125=>"100000011",
  60126=>"100110110",
  60127=>"110001111",
  60128=>"011110010",
  60129=>"010101011",
  60130=>"110110100",
  60131=>"111001111",
  60132=>"110001000",
  60133=>"101000100",
  60134=>"001011011",
  60135=>"000000110",
  60136=>"010010010",
  60137=>"100001110",
  60138=>"011110000",
  60139=>"010100010",
  60140=>"000011101",
  60141=>"001011111",
  60142=>"010101100",
  60143=>"000000110",
  60144=>"110010000",
  60145=>"101001010",
  60146=>"000110110",
  60147=>"111101011",
  60148=>"100010001",
  60149=>"111110011",
  60150=>"101000011",
  60151=>"001001001",
  60152=>"001000100",
  60153=>"101000000",
  60154=>"010010000",
  60155=>"111000010",
  60156=>"101101111",
  60157=>"110101100",
  60158=>"111011110",
  60159=>"111000110",
  60160=>"000010100",
  60161=>"001110100",
  60162=>"001101001",
  60163=>"000011000",
  60164=>"110000110",
  60165=>"011001111",
  60166=>"111000011",
  60167=>"000011010",
  60168=>"111011101",
  60169=>"100011010",
  60170=>"001001011",
  60171=>"101110100",
  60172=>"110010011",
  60173=>"000001001",
  60174=>"001111001",
  60175=>"110110100",
  60176=>"001011010",
  60177=>"101101101",
  60178=>"011111110",
  60179=>"000001010",
  60180=>"000110011",
  60181=>"011111010",
  60182=>"000101110",
  60183=>"111011001",
  60184=>"101000000",
  60185=>"000011100",
  60186=>"001110110",
  60187=>"000000111",
  60188=>"101100110",
  60189=>"110101100",
  60190=>"101110010",
  60191=>"001000101",
  60192=>"011011101",
  60193=>"111110110",
  60194=>"111110001",
  60195=>"110010010",
  60196=>"101001011",
  60197=>"011101110",
  60198=>"010001110",
  60199=>"110000010",
  60200=>"010000110",
  60201=>"001001000",
  60202=>"001110101",
  60203=>"100000001",
  60204=>"001111111",
  60205=>"000101000",
  60206=>"000000011",
  60207=>"000101001",
  60208=>"010100001",
  60209=>"100011010",
  60210=>"000100001",
  60211=>"000011100",
  60212=>"110111111",
  60213=>"000101100",
  60214=>"011010001",
  60215=>"101010100",
  60216=>"111010111",
  60217=>"010111001",
  60218=>"001000110",
  60219=>"000011011",
  60220=>"111011000",
  60221=>"010100100",
  60222=>"101110001",
  60223=>"011010100",
  60224=>"010110010",
  60225=>"101000101",
  60226=>"001010110",
  60227=>"010010101",
  60228=>"110000101",
  60229=>"101100001",
  60230=>"101100010",
  60231=>"001100011",
  60232=>"101100111",
  60233=>"101111000",
  60234=>"101001001",
  60235=>"111001010",
  60236=>"001000101",
  60237=>"101100101",
  60238=>"001000101",
  60239=>"111110110",
  60240=>"010010000",
  60241=>"001001011",
  60242=>"100000100",
  60243=>"110000111",
  60244=>"110000001",
  60245=>"000010111",
  60246=>"010101110",
  60247=>"001101000",
  60248=>"111010101",
  60249=>"111000011",
  60250=>"010010010",
  60251=>"111001010",
  60252=>"100110100",
  60253=>"010100110",
  60254=>"001001100",
  60255=>"101100001",
  60256=>"010111111",
  60257=>"001001001",
  60258=>"001110111",
  60259=>"000001001",
  60260=>"110101101",
  60261=>"001001101",
  60262=>"110011000",
  60263=>"000000001",
  60264=>"011000001",
  60265=>"001111100",
  60266=>"010101001",
  60267=>"111101101",
  60268=>"000001000",
  60269=>"011000001",
  60270=>"001001001",
  60271=>"011110001",
  60272=>"011111000",
  60273=>"111111101",
  60274=>"011011100",
  60275=>"011111110",
  60276=>"000101000",
  60277=>"011111110",
  60278=>"011101010",
  60279=>"110100101",
  60280=>"101010001",
  60281=>"001110110",
  60282=>"011010101",
  60283=>"100101100",
  60284=>"111101010",
  60285=>"011011110",
  60286=>"100011101",
  60287=>"101010100",
  60288=>"100111111",
  60289=>"111000101",
  60290=>"111101101",
  60291=>"010011011",
  60292=>"000010100",
  60293=>"001110010",
  60294=>"000110010",
  60295=>"010101000",
  60296=>"101100111",
  60297=>"001100001",
  60298=>"111010111",
  60299=>"101001011",
  60300=>"011001011",
  60301=>"000011100",
  60302=>"000001011",
  60303=>"111001011",
  60304=>"111101101",
  60305=>"101000011",
  60306=>"011011001",
  60307=>"111101001",
  60308=>"111000011",
  60309=>"100110010",
  60310=>"010101110",
  60311=>"000110101",
  60312=>"010000101",
  60313=>"111111110",
  60314=>"000110100",
  60315=>"101010001",
  60316=>"001100110",
  60317=>"101011000",
  60318=>"001100100",
  60319=>"100110001",
  60320=>"000001101",
  60321=>"100011011",
  60322=>"101100111",
  60323=>"000001001",
  60324=>"001010101",
  60325=>"101100010",
  60326=>"111101100",
  60327=>"011101111",
  60328=>"100110001",
  60329=>"010000010",
  60330=>"001010011",
  60331=>"100101111",
  60332=>"001100000",
  60333=>"100011100",
  60334=>"101010110",
  60335=>"001000000",
  60336=>"101000101",
  60337=>"001101001",
  60338=>"010111100",
  60339=>"110011000",
  60340=>"000100111",
  60341=>"010001100",
  60342=>"111111001",
  60343=>"001000000",
  60344=>"111001110",
  60345=>"000110011",
  60346=>"101101100",
  60347=>"110001011",
  60348=>"101111001",
  60349=>"010101101",
  60350=>"101101001",
  60351=>"101111000",
  60352=>"011110111",
  60353=>"100000010",
  60354=>"000000101",
  60355=>"110010100",
  60356=>"011010000",
  60357=>"000010111",
  60358=>"001100100",
  60359=>"111100101",
  60360=>"000101010",
  60361=>"101001111",
  60362=>"110010010",
  60363=>"111111110",
  60364=>"001110011",
  60365=>"010011100",
  60366=>"101010101",
  60367=>"111111110",
  60368=>"110011000",
  60369=>"010101110",
  60370=>"110100001",
  60371=>"110001011",
  60372=>"101110101",
  60373=>"111110111",
  60374=>"011000001",
  60375=>"111011110",
  60376=>"011100000",
  60377=>"111000101",
  60378=>"010001000",
  60379=>"100001100",
  60380=>"010100010",
  60381=>"100110001",
  60382=>"100000000",
  60383=>"000000110",
  60384=>"101100110",
  60385=>"011111101",
  60386=>"001100010",
  60387=>"000011011",
  60388=>"001100101",
  60389=>"000001010",
  60390=>"110010100",
  60391=>"000110001",
  60392=>"100010111",
  60393=>"111010010",
  60394=>"100111101",
  60395=>"010011010",
  60396=>"100001101",
  60397=>"100111010",
  60398=>"011101000",
  60399=>"111010000",
  60400=>"010001101",
  60401=>"110010010",
  60402=>"101101101",
  60403=>"100110001",
  60404=>"000100111",
  60405=>"110011011",
  60406=>"000101001",
  60407=>"011011011",
  60408=>"111001111",
  60409=>"000001111",
  60410=>"010101001",
  60411=>"110101110",
  60412=>"001001011",
  60413=>"001001001",
  60414=>"000100010",
  60415=>"111110100",
  60416=>"110111010",
  60417=>"001100000",
  60418=>"100101101",
  60419=>"111011101",
  60420=>"001101000",
  60421=>"010100110",
  60422=>"110010001",
  60423=>"011000001",
  60424=>"111011011",
  60425=>"110000111",
  60426=>"001101110",
  60427=>"100001000",
  60428=>"000000101",
  60429=>"101101101",
  60430=>"111111101",
  60431=>"101110111",
  60432=>"110010111",
  60433=>"001001011",
  60434=>"111111001",
  60435=>"101110100",
  60436=>"001110100",
  60437=>"100000010",
  60438=>"001100110",
  60439=>"100110110",
  60440=>"110110000",
  60441=>"000100101",
  60442=>"010010101",
  60443=>"001010010",
  60444=>"110000001",
  60445=>"110001110",
  60446=>"101101011",
  60447=>"100110110",
  60448=>"011000010",
  60449=>"001100011",
  60450=>"010110001",
  60451=>"000100011",
  60452=>"100001000",
  60453=>"011110110",
  60454=>"100110001",
  60455=>"110011110",
  60456=>"110111011",
  60457=>"000001000",
  60458=>"100110001",
  60459=>"101111010",
  60460=>"000100001",
  60461=>"011001001",
  60462=>"001001001",
  60463=>"100001001",
  60464=>"111011001",
  60465=>"101110100",
  60466=>"100000101",
  60467=>"010101111",
  60468=>"010000000",
  60469=>"000001111",
  60470=>"010101111",
  60471=>"111110111",
  60472=>"100100011",
  60473=>"111111111",
  60474=>"000000110",
  60475=>"100100100",
  60476=>"000001010",
  60477=>"110011001",
  60478=>"011010000",
  60479=>"000101000",
  60480=>"110001011",
  60481=>"000110001",
  60482=>"110100010",
  60483=>"010011011",
  60484=>"000110010",
  60485=>"100010010",
  60486=>"100000011",
  60487=>"111011101",
  60488=>"010001111",
  60489=>"101111110",
  60490=>"111111000",
  60491=>"011010101",
  60492=>"011001101",
  60493=>"110110111",
  60494=>"101011011",
  60495=>"101010010",
  60496=>"111000100",
  60497=>"010110101",
  60498=>"001110111",
  60499=>"101011100",
  60500=>"000100110",
  60501=>"000010111",
  60502=>"111101111",
  60503=>"010100000",
  60504=>"000001111",
  60505=>"100101000",
  60506=>"011101100",
  60507=>"100000011",
  60508=>"100011001",
  60509=>"001001000",
  60510=>"000000000",
  60511=>"110010010",
  60512=>"100000011",
  60513=>"000000001",
  60514=>"111101010",
  60515=>"000100011",
  60516=>"001111111",
  60517=>"000110111",
  60518=>"110101100",
  60519=>"000011110",
  60520=>"100010100",
  60521=>"101111010",
  60522=>"100001000",
  60523=>"001010011",
  60524=>"100101110",
  60525=>"011010111",
  60526=>"000000000",
  60527=>"000010011",
  60528=>"101001010",
  60529=>"010111101",
  60530=>"101111010",
  60531=>"100011000",
  60532=>"100010000",
  60533=>"000011110",
  60534=>"011111111",
  60535=>"110101110",
  60536=>"001100000",
  60537=>"110010011",
  60538=>"000100010",
  60539=>"111001010",
  60540=>"000101000",
  60541=>"000101100",
  60542=>"010001010",
  60543=>"010000100",
  60544=>"101000111",
  60545=>"010011011",
  60546=>"010001010",
  60547=>"100100100",
  60548=>"110000100",
  60549=>"101001010",
  60550=>"001111111",
  60551=>"001101001",
  60552=>"100101100",
  60553=>"011001001",
  60554=>"110001010",
  60555=>"100100010",
  60556=>"101111100",
  60557=>"110000110",
  60558=>"001100110",
  60559=>"001000001",
  60560=>"111000011",
  60561=>"000001011",
  60562=>"011111100",
  60563=>"110011010",
  60564=>"010111000",
  60565=>"101111001",
  60566=>"001011100",
  60567=>"011010110",
  60568=>"110011001",
  60569=>"011100111",
  60570=>"000111011",
  60571=>"010100001",
  60572=>"010101111",
  60573=>"110100011",
  60574=>"001111010",
  60575=>"110001110",
  60576=>"001001001",
  60577=>"100101101",
  60578=>"000010100",
  60579=>"000011011",
  60580=>"001110010",
  60581=>"100001111",
  60582=>"101010001",
  60583=>"110110010",
  60584=>"101010100",
  60585=>"010001100",
  60586=>"110010100",
  60587=>"110010111",
  60588=>"110101100",
  60589=>"011010110",
  60590=>"010110110",
  60591=>"111110100",
  60592=>"111110000",
  60593=>"101000000",
  60594=>"111111110",
  60595=>"010100000",
  60596=>"110110101",
  60597=>"011111011",
  60598=>"100011100",
  60599=>"110111100",
  60600=>"001001001",
  60601=>"000100100",
  60602=>"101110001",
  60603=>"100111001",
  60604=>"011010001",
  60605=>"100110111",
  60606=>"110111100",
  60607=>"011001001",
  60608=>"100001001",
  60609=>"110110101",
  60610=>"100001010",
  60611=>"110011011",
  60612=>"101000010",
  60613=>"010000111",
  60614=>"010000111",
  60615=>"011111011",
  60616=>"101110001",
  60617=>"000000111",
  60618=>"000101010",
  60619=>"000001100",
  60620=>"010101011",
  60621=>"001101101",
  60622=>"111000001",
  60623=>"001001001",
  60624=>"000000001",
  60625=>"001011011",
  60626=>"000100110",
  60627=>"011100001",
  60628=>"010000011",
  60629=>"101110100",
  60630=>"101001000",
  60631=>"010110101",
  60632=>"101110001",
  60633=>"000101110",
  60634=>"110110011",
  60635=>"000000000",
  60636=>"011010010",
  60637=>"011001110",
  60638=>"100111111",
  60639=>"111000100",
  60640=>"110001001",
  60641=>"110000000",
  60642=>"111111111",
  60643=>"000000100",
  60644=>"010100011",
  60645=>"111011110",
  60646=>"001000011",
  60647=>"000010111",
  60648=>"100001001",
  60649=>"100110111",
  60650=>"000001110",
  60651=>"101000010",
  60652=>"010110001",
  60653=>"001111000",
  60654=>"110001011",
  60655=>"011000101",
  60656=>"100110110",
  60657=>"110111110",
  60658=>"010011001",
  60659=>"110010011",
  60660=>"110111110",
  60661=>"100001011",
  60662=>"000010001",
  60663=>"001100001",
  60664=>"001011100",
  60665=>"100100100",
  60666=>"100101000",
  60667=>"010011101",
  60668=>"111001000",
  60669=>"011001110",
  60670=>"101011110",
  60671=>"111001100",
  60672=>"100011100",
  60673=>"111010011",
  60674=>"100010100",
  60675=>"001000001",
  60676=>"101111110",
  60677=>"010110011",
  60678=>"001101011",
  60679=>"011011111",
  60680=>"000101100",
  60681=>"011110111",
  60682=>"000000001",
  60683=>"000111000",
  60684=>"101000110",
  60685=>"011011010",
  60686=>"001000010",
  60687=>"001111110",
  60688=>"011100101",
  60689=>"101111110",
  60690=>"011011011",
  60691=>"110000010",
  60692=>"000011011",
  60693=>"011010001",
  60694=>"101011111",
  60695=>"101010000",
  60696=>"011011001",
  60697=>"001010000",
  60698=>"110111010",
  60699=>"001000010",
  60700=>"010100101",
  60701=>"100000011",
  60702=>"111001101",
  60703=>"011010011",
  60704=>"001000000",
  60705=>"001001101",
  60706=>"000011111",
  60707=>"110100111",
  60708=>"111000100",
  60709=>"111000101",
  60710=>"000010010",
  60711=>"010101011",
  60712=>"001101001",
  60713=>"000100010",
  60714=>"011010001",
  60715=>"110111001",
  60716=>"010010011",
  60717=>"001000011",
  60718=>"110011101",
  60719=>"100001101",
  60720=>"111101000",
  60721=>"111101011",
  60722=>"110100111",
  60723=>"000001111",
  60724=>"010101100",
  60725=>"000001110",
  60726=>"101010011",
  60727=>"011010000",
  60728=>"000111001",
  60729=>"100000001",
  60730=>"011110100",
  60731=>"111100001",
  60732=>"101000100",
  60733=>"001100100",
  60734=>"111110101",
  60735=>"111011001",
  60736=>"111010010",
  60737=>"101001110",
  60738=>"001000010",
  60739=>"110110111",
  60740=>"101011010",
  60741=>"011011001",
  60742=>"100100110",
  60743=>"101100001",
  60744=>"011110101",
  60745=>"100100111",
  60746=>"011010001",
  60747=>"010000110",
  60748=>"010111001",
  60749=>"111110001",
  60750=>"100010000",
  60751=>"111011111",
  60752=>"010100010",
  60753=>"100001101",
  60754=>"111110110",
  60755=>"001101000",
  60756=>"010100100",
  60757=>"101011110",
  60758=>"000000001",
  60759=>"100011010",
  60760=>"101001100",
  60761=>"001101110",
  60762=>"011111011",
  60763=>"010001101",
  60764=>"100110101",
  60765=>"010011010",
  60766=>"000101000",
  60767=>"100101100",
  60768=>"010100110",
  60769=>"101001001",
  60770=>"000000111",
  60771=>"001101001",
  60772=>"011011010",
  60773=>"010100000",
  60774=>"000011000",
  60775=>"101110111",
  60776=>"111110111",
  60777=>"001001010",
  60778=>"011111101",
  60779=>"110110000",
  60780=>"110100101",
  60781=>"111100111",
  60782=>"001111010",
  60783=>"011011111",
  60784=>"100110010",
  60785=>"001101001",
  60786=>"101111010",
  60787=>"000101111",
  60788=>"010000011",
  60789=>"101111000",
  60790=>"010011011",
  60791=>"111111101",
  60792=>"001101010",
  60793=>"011100100",
  60794=>"000001011",
  60795=>"101100000",
  60796=>"000010001",
  60797=>"101011011",
  60798=>"011110111",
  60799=>"001100000",
  60800=>"010101101",
  60801=>"011011110",
  60802=>"110010011",
  60803=>"010001100",
  60804=>"010011101",
  60805=>"100011001",
  60806=>"011110000",
  60807=>"110000101",
  60808=>"000010000",
  60809=>"011010111",
  60810=>"010010110",
  60811=>"100111011",
  60812=>"000101001",
  60813=>"000000011",
  60814=>"110111010",
  60815=>"111101110",
  60816=>"101011100",
  60817=>"100001111",
  60818=>"100010111",
  60819=>"001111011",
  60820=>"011000011",
  60821=>"000010100",
  60822=>"111000111",
  60823=>"011110001",
  60824=>"110001100",
  60825=>"110000000",
  60826=>"010000010",
  60827=>"000010001",
  60828=>"110011010",
  60829=>"101001000",
  60830=>"110110100",
  60831=>"000110110",
  60832=>"100000001",
  60833=>"110101011",
  60834=>"001001001",
  60835=>"001010000",
  60836=>"101011011",
  60837=>"010101010",
  60838=>"010010000",
  60839=>"010100100",
  60840=>"010011010",
  60841=>"000000011",
  60842=>"110100100",
  60843=>"101001001",
  60844=>"010111111",
  60845=>"100110010",
  60846=>"001101000",
  60847=>"111010000",
  60848=>"110101011",
  60849=>"010100011",
  60850=>"110011110",
  60851=>"001000110",
  60852=>"001100111",
  60853=>"100001000",
  60854=>"010111001",
  60855=>"011001000",
  60856=>"101000010",
  60857=>"001100010",
  60858=>"000000001",
  60859=>"001010001",
  60860=>"010110001",
  60861=>"010101010",
  60862=>"101000011",
  60863=>"110011000",
  60864=>"110101000",
  60865=>"101000000",
  60866=>"001010010",
  60867=>"101001010",
  60868=>"000000101",
  60869=>"100010011",
  60870=>"101001010",
  60871=>"110110110",
  60872=>"111010101",
  60873=>"101101000",
  60874=>"101001010",
  60875=>"010100110",
  60876=>"110111001",
  60877=>"000101001",
  60878=>"100010011",
  60879=>"110000011",
  60880=>"001001011",
  60881=>"000110010",
  60882=>"000001000",
  60883=>"011000101",
  60884=>"110110110",
  60885=>"010100001",
  60886=>"010000000",
  60887=>"011101001",
  60888=>"110100101",
  60889=>"110011110",
  60890=>"100010011",
  60891=>"101111011",
  60892=>"010100010",
  60893=>"000000110",
  60894=>"110010000",
  60895=>"100111110",
  60896=>"011000000",
  60897=>"110111111",
  60898=>"110000000",
  60899=>"011011001",
  60900=>"100011010",
  60901=>"000101100",
  60902=>"010110100",
  60903=>"010001100",
  60904=>"001110100",
  60905=>"000111001",
  60906=>"000101010",
  60907=>"101000101",
  60908=>"100010100",
  60909=>"011001010",
  60910=>"001010110",
  60911=>"111111110",
  60912=>"101010001",
  60913=>"001011111",
  60914=>"111111000",
  60915=>"010111111",
  60916=>"111110010",
  60917=>"100000101",
  60918=>"000110001",
  60919=>"011110101",
  60920=>"101000111",
  60921=>"111010011",
  60922=>"001001000",
  60923=>"100111011",
  60924=>"000001101",
  60925=>"111001010",
  60926=>"101011000",
  60927=>"011101101",
  60928=>"100110100",
  60929=>"101101101",
  60930=>"010110001",
  60931=>"001001101",
  60932=>"101011110",
  60933=>"100101100",
  60934=>"011100010",
  60935=>"001101000",
  60936=>"000000111",
  60937=>"010110101",
  60938=>"100011100",
  60939=>"110000010",
  60940=>"100111011",
  60941=>"100000111",
  60942=>"110100000",
  60943=>"110001110",
  60944=>"100011111",
  60945=>"000000010",
  60946=>"101110001",
  60947=>"111001010",
  60948=>"011010100",
  60949=>"111101101",
  60950=>"001111011",
  60951=>"111010010",
  60952=>"000001100",
  60953=>"010110010",
  60954=>"110110010",
  60955=>"110101001",
  60956=>"000001111",
  60957=>"100001011",
  60958=>"001100101",
  60959=>"100110100",
  60960=>"111011010",
  60961=>"000101111",
  60962=>"111110100",
  60963=>"000010110",
  60964=>"100110111",
  60965=>"010010100",
  60966=>"000000110",
  60967=>"011000001",
  60968=>"001111000",
  60969=>"101101010",
  60970=>"101100101",
  60971=>"110011010",
  60972=>"110000001",
  60973=>"000001110",
  60974=>"000010000",
  60975=>"001101010",
  60976=>"110011111",
  60977=>"111101111",
  60978=>"000001111",
  60979=>"000011011",
  60980=>"111100011",
  60981=>"010010111",
  60982=>"111101110",
  60983=>"010110010",
  60984=>"111000011",
  60985=>"101101011",
  60986=>"011111110",
  60987=>"011011110",
  60988=>"100100011",
  60989=>"100000101",
  60990=>"101100101",
  60991=>"010110101",
  60992=>"010101000",
  60993=>"000010010",
  60994=>"000000110",
  60995=>"010001101",
  60996=>"110101111",
  60997=>"111000100",
  60998=>"000000010",
  60999=>"010011110",
  61000=>"011010111",
  61001=>"010010110",
  61002=>"100000111",
  61003=>"100110111",
  61004=>"011111110",
  61005=>"100000001",
  61006=>"100010111",
  61007=>"101100000",
  61008=>"001011001",
  61009=>"100010000",
  61010=>"111011000",
  61011=>"001101001",
  61012=>"011001001",
  61013=>"101101000",
  61014=>"011101011",
  61015=>"000101011",
  61016=>"011000011",
  61017=>"100101001",
  61018=>"011111100",
  61019=>"001000110",
  61020=>"011101100",
  61021=>"010010111",
  61022=>"110101000",
  61023=>"101111001",
  61024=>"100000011",
  61025=>"101010010",
  61026=>"110111101",
  61027=>"000010101",
  61028=>"110101011",
  61029=>"110110111",
  61030=>"001110011",
  61031=>"001101011",
  61032=>"010100011",
  61033=>"011011111",
  61034=>"110101101",
  61035=>"000000101",
  61036=>"100100000",
  61037=>"000101100",
  61038=>"100011111",
  61039=>"011100000",
  61040=>"011100110",
  61041=>"111101010",
  61042=>"100101001",
  61043=>"000110100",
  61044=>"111010100",
  61045=>"001001000",
  61046=>"110101000",
  61047=>"011000000",
  61048=>"000101111",
  61049=>"100100100",
  61050=>"100111000",
  61051=>"001111100",
  61052=>"111100101",
  61053=>"101010000",
  61054=>"000110001",
  61055=>"010000011",
  61056=>"011010101",
  61057=>"010001011",
  61058=>"100001101",
  61059=>"101011011",
  61060=>"011010010",
  61061=>"101011000",
  61062=>"110101111",
  61063=>"001101010",
  61064=>"110010101",
  61065=>"101101000",
  61066=>"111100001",
  61067=>"110110110",
  61068=>"010101101",
  61069=>"010000000",
  61070=>"101011110",
  61071=>"010011110",
  61072=>"011011001",
  61073=>"010100000",
  61074=>"000001111",
  61075=>"010111101",
  61076=>"001011011",
  61077=>"100100111",
  61078=>"101010111",
  61079=>"101000001",
  61080=>"111101100",
  61081=>"101011101",
  61082=>"110010010",
  61083=>"001000110",
  61084=>"110100100",
  61085=>"010010011",
  61086=>"001001010",
  61087=>"011101001",
  61088=>"111101000",
  61089=>"000010111",
  61090=>"101101100",
  61091=>"000110111",
  61092=>"011100101",
  61093=>"001011110",
  61094=>"000000100",
  61095=>"000101010",
  61096=>"111011111",
  61097=>"110101100",
  61098=>"001101100",
  61099=>"110100001",
  61100=>"101010000",
  61101=>"010000011",
  61102=>"011110100",
  61103=>"001101101",
  61104=>"011001010",
  61105=>"001000001",
  61106=>"111101100",
  61107=>"110000001",
  61108=>"010011101",
  61109=>"001011111",
  61110=>"001111100",
  61111=>"001101001",
  61112=>"100101100",
  61113=>"110000010",
  61114=>"011011110",
  61115=>"101100011",
  61116=>"100010000",
  61117=>"110011101",
  61118=>"001000100",
  61119=>"001100001",
  61120=>"000111001",
  61121=>"010001101",
  61122=>"110111110",
  61123=>"111101101",
  61124=>"101101010",
  61125=>"101100101",
  61126=>"001110011",
  61127=>"001010101",
  61128=>"000000011",
  61129=>"110010110",
  61130=>"011100101",
  61131=>"100010100",
  61132=>"010001010",
  61133=>"011011011",
  61134=>"110011000",
  61135=>"111011011",
  61136=>"101111101",
  61137=>"000010100",
  61138=>"011100000",
  61139=>"010100000",
  61140=>"000000110",
  61141=>"110011111",
  61142=>"000101100",
  61143=>"000110111",
  61144=>"001111101",
  61145=>"000000000",
  61146=>"110001010",
  61147=>"110010000",
  61148=>"101001000",
  61149=>"110110110",
  61150=>"000111111",
  61151=>"010110001",
  61152=>"000011000",
  61153=>"100010010",
  61154=>"011101110",
  61155=>"000101111",
  61156=>"000111011",
  61157=>"000101001",
  61158=>"101101010",
  61159=>"101010001",
  61160=>"001010100",
  61161=>"111111001",
  61162=>"011001110",
  61163=>"101100111",
  61164=>"100011000",
  61165=>"111110011",
  61166=>"110010110",
  61167=>"000001111",
  61168=>"110010001",
  61169=>"001001000",
  61170=>"000011011",
  61171=>"011111010",
  61172=>"000000100",
  61173=>"111101111",
  61174=>"010011010",
  61175=>"110000101",
  61176=>"000110000",
  61177=>"101110110",
  61178=>"111000001",
  61179=>"101001100",
  61180=>"100010100",
  61181=>"001001100",
  61182=>"010111000",
  61183=>"011110111",
  61184=>"010111101",
  61185=>"010010111",
  61186=>"001101001",
  61187=>"000010110",
  61188=>"000000000",
  61189=>"001001010",
  61190=>"001110010",
  61191=>"001110110",
  61192=>"001000001",
  61193=>"111011000",
  61194=>"110101111",
  61195=>"110011001",
  61196=>"100001111",
  61197=>"010111111",
  61198=>"001100010",
  61199=>"101111111",
  61200=>"100000011",
  61201=>"100110001",
  61202=>"100000111",
  61203=>"111111110",
  61204=>"001100110",
  61205=>"001000100",
  61206=>"010000011",
  61207=>"010010010",
  61208=>"110101110",
  61209=>"001101000",
  61210=>"010010000",
  61211=>"101010101",
  61212=>"010100001",
  61213=>"111001001",
  61214=>"011001010",
  61215=>"110101110",
  61216=>"001001101",
  61217=>"110011100",
  61218=>"100000011",
  61219=>"011111110",
  61220=>"010101001",
  61221=>"100000011",
  61222=>"100111101",
  61223=>"001101100",
  61224=>"101100100",
  61225=>"001100001",
  61226=>"110100010",
  61227=>"011011101",
  61228=>"111011011",
  61229=>"001100101",
  61230=>"010010011",
  61231=>"111000000",
  61232=>"101110111",
  61233=>"011110000",
  61234=>"000110101",
  61235=>"011010011",
  61236=>"010111110",
  61237=>"010000010",
  61238=>"110110000",
  61239=>"001000001",
  61240=>"010111111",
  61241=>"001010110",
  61242=>"010000001",
  61243=>"011110100",
  61244=>"100010000",
  61245=>"011001011",
  61246=>"110011101",
  61247=>"010101101",
  61248=>"101011100",
  61249=>"111101100",
  61250=>"101100111",
  61251=>"001000000",
  61252=>"101000111",
  61253=>"010101100",
  61254=>"011100101",
  61255=>"001100001",
  61256=>"100011110",
  61257=>"111110000",
  61258=>"101011001",
  61259=>"100010000",
  61260=>"001110000",
  61261=>"111010111",
  61262=>"101010110",
  61263=>"001001011",
  61264=>"100010100",
  61265=>"110100110",
  61266=>"101101100",
  61267=>"000010000",
  61268=>"000000010",
  61269=>"100100100",
  61270=>"011000010",
  61271=>"110101001",
  61272=>"111111000",
  61273=>"110100111",
  61274=>"000011111",
  61275=>"100001100",
  61276=>"111100001",
  61277=>"010100110",
  61278=>"110100101",
  61279=>"000010010",
  61280=>"110010000",
  61281=>"101000011",
  61282=>"001010101",
  61283=>"011001101",
  61284=>"110011001",
  61285=>"111001011",
  61286=>"010011101",
  61287=>"010110110",
  61288=>"001010000",
  61289=>"110011111",
  61290=>"011000100",
  61291=>"010100010",
  61292=>"010101100",
  61293=>"000000110",
  61294=>"000010001",
  61295=>"101111101",
  61296=>"111111111",
  61297=>"111010100",
  61298=>"010001010",
  61299=>"111101000",
  61300=>"111000010",
  61301=>"000000100",
  61302=>"000111000",
  61303=>"100110000",
  61304=>"001111000",
  61305=>"001100101",
  61306=>"100101011",
  61307=>"001010000",
  61308=>"000010001",
  61309=>"010000000",
  61310=>"000000000",
  61311=>"101010101",
  61312=>"011001000",
  61313=>"111011000",
  61314=>"110011110",
  61315=>"000100100",
  61316=>"110100001",
  61317=>"010011111",
  61318=>"110110011",
  61319=>"111100101",
  61320=>"110100010",
  61321=>"010111101",
  61322=>"110001010",
  61323=>"111010111",
  61324=>"110011000",
  61325=>"110010000",
  61326=>"001000010",
  61327=>"101000001",
  61328=>"101101001",
  61329=>"011000011",
  61330=>"110010101",
  61331=>"110000001",
  61332=>"001111001",
  61333=>"101001000",
  61334=>"101010001",
  61335=>"011110000",
  61336=>"010101110",
  61337=>"110100000",
  61338=>"111101010",
  61339=>"101100001",
  61340=>"110111000",
  61341=>"101011001",
  61342=>"110010101",
  61343=>"011100111",
  61344=>"000010100",
  61345=>"001001000",
  61346=>"111000011",
  61347=>"101101000",
  61348=>"100001110",
  61349=>"100110100",
  61350=>"111000101",
  61351=>"011100111",
  61352=>"010101110",
  61353=>"001000000",
  61354=>"100010000",
  61355=>"000001110",
  61356=>"010010001",
  61357=>"100100011",
  61358=>"010100001",
  61359=>"011010000",
  61360=>"110101101",
  61361=>"111110010",
  61362=>"111111010",
  61363=>"101001010",
  61364=>"010001100",
  61365=>"001101010",
  61366=>"101000011",
  61367=>"110001000",
  61368=>"010001111",
  61369=>"011010000",
  61370=>"101000101",
  61371=>"011011101",
  61372=>"000000010",
  61373=>"010000011",
  61374=>"111000100",
  61375=>"001001010",
  61376=>"111111101",
  61377=>"000100101",
  61378=>"010100001",
  61379=>"001010110",
  61380=>"010101001",
  61381=>"110001010",
  61382=>"101001101",
  61383=>"000000100",
  61384=>"100100100",
  61385=>"110100111",
  61386=>"001110000",
  61387=>"101110010",
  61388=>"011100100",
  61389=>"011010010",
  61390=>"100110110",
  61391=>"111000110",
  61392=>"011110100",
  61393=>"111100001",
  61394=>"011011111",
  61395=>"011110000",
  61396=>"111110101",
  61397=>"100110110",
  61398=>"011011011",
  61399=>"111001100",
  61400=>"011010111",
  61401=>"101101101",
  61402=>"000000000",
  61403=>"101011110",
  61404=>"001010100",
  61405=>"101001110",
  61406=>"100000101",
  61407=>"001101101",
  61408=>"101111110",
  61409=>"101110101",
  61410=>"011001000",
  61411=>"110010001",
  61412=>"001000000",
  61413=>"000100110",
  61414=>"010110110",
  61415=>"101100000",
  61416=>"110100111",
  61417=>"110000011",
  61418=>"101101001",
  61419=>"110101000",
  61420=>"011111101",
  61421=>"100001000",
  61422=>"000000000",
  61423=>"000000010",
  61424=>"111011100",
  61425=>"010111111",
  61426=>"000100011",
  61427=>"100100001",
  61428=>"000011101",
  61429=>"100000000",
  61430=>"101010110",
  61431=>"011101010",
  61432=>"001011100",
  61433=>"010101011",
  61434=>"100100000",
  61435=>"010111001",
  61436=>"001111001",
  61437=>"111000101",
  61438=>"110111001",
  61439=>"111000010",
  61440=>"111110000",
  61441=>"011100100",
  61442=>"000010100",
  61443=>"000010101",
  61444=>"100011001",
  61445=>"000110011",
  61446=>"011110111",
  61447=>"011001011",
  61448=>"101110101",
  61449=>"000011101",
  61450=>"101100001",
  61451=>"011101100",
  61452=>"101111111",
  61453=>"111110011",
  61454=>"010001110",
  61455=>"111001110",
  61456=>"111110100",
  61457=>"100010010",
  61458=>"010011111",
  61459=>"001000011",
  61460=>"000100000",
  61461=>"010111111",
  61462=>"110011011",
  61463=>"111000010",
  61464=>"111100011",
  61465=>"111110101",
  61466=>"100111100",
  61467=>"101001101",
  61468=>"001000110",
  61469=>"010101011",
  61470=>"000011000",
  61471=>"101101010",
  61472=>"000111001",
  61473=>"101000110",
  61474=>"010110001",
  61475=>"010000011",
  61476=>"010110111",
  61477=>"000000011",
  61478=>"100000000",
  61479=>"110110111",
  61480=>"011111110",
  61481=>"000010000",
  61482=>"111101011",
  61483=>"110110010",
  61484=>"111110000",
  61485=>"011110110",
  61486=>"100010101",
  61487=>"100110110",
  61488=>"110001010",
  61489=>"100110011",
  61490=>"001101011",
  61491=>"011011111",
  61492=>"000110011",
  61493=>"111001010",
  61494=>"010001010",
  61495=>"110111010",
  61496=>"000001101",
  61497=>"111101000",
  61498=>"101000110",
  61499=>"111000000",
  61500=>"000000110",
  61501=>"111111111",
  61502=>"001000101",
  61503=>"010111101",
  61504=>"111010110",
  61505=>"000000100",
  61506=>"101011111",
  61507=>"100000100",
  61508=>"011001000",
  61509=>"011000001",
  61510=>"110011101",
  61511=>"010000000",
  61512=>"100010111",
  61513=>"010111011",
  61514=>"111101010",
  61515=>"111111101",
  61516=>"000000001",
  61517=>"011111111",
  61518=>"110111101",
  61519=>"101101000",
  61520=>"010000001",
  61521=>"101110110",
  61522=>"000010111",
  61523=>"110101010",
  61524=>"011011100",
  61525=>"101110100",
  61526=>"011011111",
  61527=>"101111000",
  61528=>"111010111",
  61529=>"001011110",
  61530=>"000001111",
  61531=>"010110111",
  61532=>"111100001",
  61533=>"100111111",
  61534=>"110100110",
  61535=>"100010000",
  61536=>"101101010",
  61537=>"101011001",
  61538=>"001100111",
  61539=>"100001101",
  61540=>"000010000",
  61541=>"001000111",
  61542=>"100101000",
  61543=>"011001000",
  61544=>"111011100",
  61545=>"011110100",
  61546=>"110000001",
  61547=>"100000100",
  61548=>"100011101",
  61549=>"010011011",
  61550=>"101101101",
  61551=>"111000011",
  61552=>"000110000",
  61553=>"100100110",
  61554=>"000100111",
  61555=>"100010011",
  61556=>"011011110",
  61557=>"111010110",
  61558=>"001000110",
  61559=>"101101010",
  61560=>"111000100",
  61561=>"110001100",
  61562=>"100001011",
  61563=>"111010010",
  61564=>"111000011",
  61565=>"010010101",
  61566=>"111000111",
  61567=>"011100011",
  61568=>"101000110",
  61569=>"000101000",
  61570=>"000001000",
  61571=>"000000110",
  61572=>"110010110",
  61573=>"110101000",
  61574=>"100001101",
  61575=>"111010010",
  61576=>"000010110",
  61577=>"010010110",
  61578=>"111001110",
  61579=>"010001001",
  61580=>"000110010",
  61581=>"100010000",
  61582=>"110000000",
  61583=>"011101000",
  61584=>"101000001",
  61585=>"011011011",
  61586=>"000110001",
  61587=>"010111110",
  61588=>"101100101",
  61589=>"110101010",
  61590=>"001000000",
  61591=>"111011110",
  61592=>"001100011",
  61593=>"111101010",
  61594=>"110100001",
  61595=>"000001001",
  61596=>"101011000",
  61597=>"001010101",
  61598=>"000101011",
  61599=>"011000100",
  61600=>"111111101",
  61601=>"100100100",
  61602=>"001001011",
  61603=>"001001010",
  61604=>"100111101",
  61605=>"110101110",
  61606=>"111010000",
  61607=>"000000011",
  61608=>"101111110",
  61609=>"111100100",
  61610=>"110011001",
  61611=>"000011000",
  61612=>"000011001",
  61613=>"010010110",
  61614=>"110110010",
  61615=>"101000011",
  61616=>"000011000",
  61617=>"110000100",
  61618=>"110001111",
  61619=>"110010010",
  61620=>"110111101",
  61621=>"111011101",
  61622=>"110010100",
  61623=>"011010100",
  61624=>"111000000",
  61625=>"110000101",
  61626=>"010001010",
  61627=>"111100010",
  61628=>"011100000",
  61629=>"010000110",
  61630=>"010111100",
  61631=>"111001110",
  61632=>"100000110",
  61633=>"111001100",
  61634=>"011100100",
  61635=>"000000001",
  61636=>"111011111",
  61637=>"000110000",
  61638=>"001001101",
  61639=>"110111111",
  61640=>"011100100",
  61641=>"101011011",
  61642=>"110100000",
  61643=>"111000000",
  61644=>"011010110",
  61645=>"000010011",
  61646=>"110111001",
  61647=>"011110010",
  61648=>"111100011",
  61649=>"001011100",
  61650=>"001110001",
  61651=>"111101101",
  61652=>"000100011",
  61653=>"100001000",
  61654=>"001010010",
  61655=>"101100111",
  61656=>"000001000",
  61657=>"000111001",
  61658=>"000000011",
  61659=>"011111111",
  61660=>"111100110",
  61661=>"110111111",
  61662=>"010011000",
  61663=>"111011000",
  61664=>"101010101",
  61665=>"011100011",
  61666=>"011011000",
  61667=>"110100110",
  61668=>"100110011",
  61669=>"011011101",
  61670=>"110101001",
  61671=>"110101110",
  61672=>"000101101",
  61673=>"111101111",
  61674=>"110001100",
  61675=>"100100111",
  61676=>"110101001",
  61677=>"001111010",
  61678=>"100000000",
  61679=>"000100010",
  61680=>"111111010",
  61681=>"000001100",
  61682=>"110011000",
  61683=>"110111110",
  61684=>"101001111",
  61685=>"010001111",
  61686=>"111001101",
  61687=>"010000010",
  61688=>"101111111",
  61689=>"110011001",
  61690=>"101111100",
  61691=>"010000001",
  61692=>"011100000",
  61693=>"100111110",
  61694=>"101110101",
  61695=>"001111110",
  61696=>"100000111",
  61697=>"000111010",
  61698=>"100111011",
  61699=>"011011110",
  61700=>"000011110",
  61701=>"111010111",
  61702=>"010000101",
  61703=>"000100100",
  61704=>"010101010",
  61705=>"001001011",
  61706=>"010010010",
  61707=>"011001110",
  61708=>"000001000",
  61709=>"111000100",
  61710=>"110010110",
  61711=>"111111000",
  61712=>"010010001",
  61713=>"111010110",
  61714=>"110001101",
  61715=>"001010010",
  61716=>"100011001",
  61717=>"001101101",
  61718=>"101010011",
  61719=>"101001100",
  61720=>"011001111",
  61721=>"010101100",
  61722=>"011101001",
  61723=>"010011111",
  61724=>"100110111",
  61725=>"101100001",
  61726=>"101101000",
  61727=>"100001000",
  61728=>"110000111",
  61729=>"000010110",
  61730=>"110111111",
  61731=>"010111110",
  61732=>"001001001",
  61733=>"001111000",
  61734=>"001101100",
  61735=>"100101101",
  61736=>"110100100",
  61737=>"011111001",
  61738=>"000000001",
  61739=>"010011010",
  61740=>"010101000",
  61741=>"011101101",
  61742=>"001101000",
  61743=>"010010010",
  61744=>"111001101",
  61745=>"100101101",
  61746=>"010011110",
  61747=>"111111100",
  61748=>"110100111",
  61749=>"101100111",
  61750=>"000110110",
  61751=>"010100100",
  61752=>"110000000",
  61753=>"101101011",
  61754=>"100100000",
  61755=>"010101100",
  61756=>"000000110",
  61757=>"111110110",
  61758=>"110101100",
  61759=>"000001000",
  61760=>"001111100",
  61761=>"101011100",
  61762=>"111101110",
  61763=>"111100111",
  61764=>"111110011",
  61765=>"000010100",
  61766=>"001101101",
  61767=>"001011100",
  61768=>"100101010",
  61769=>"001010011",
  61770=>"110101100",
  61771=>"001001100",
  61772=>"011100100",
  61773=>"101001110",
  61774=>"111011110",
  61775=>"001100100",
  61776=>"001000100",
  61777=>"011010100",
  61778=>"111001001",
  61779=>"010010000",
  61780=>"011000001",
  61781=>"111111111",
  61782=>"010001001",
  61783=>"000111111",
  61784=>"001001000",
  61785=>"100100101",
  61786=>"100111101",
  61787=>"111110100",
  61788=>"010100100",
  61789=>"111111100",
  61790=>"011000000",
  61791=>"101000100",
  61792=>"100100000",
  61793=>"110000101",
  61794=>"000110001",
  61795=>"001110111",
  61796=>"011111010",
  61797=>"111011011",
  61798=>"101001010",
  61799=>"010100111",
  61800=>"010000010",
  61801=>"011101100",
  61802=>"000010111",
  61803=>"000000001",
  61804=>"000101111",
  61805=>"111011110",
  61806=>"101010101",
  61807=>"101011000",
  61808=>"000001100",
  61809=>"000101100",
  61810=>"111011100",
  61811=>"111110000",
  61812=>"110011000",
  61813=>"111010010",
  61814=>"100010010",
  61815=>"000001011",
  61816=>"000000111",
  61817=>"001001110",
  61818=>"100010010",
  61819=>"000100000",
  61820=>"001001111",
  61821=>"111111011",
  61822=>"010001100",
  61823=>"111110101",
  61824=>"110100111",
  61825=>"110000100",
  61826=>"101110111",
  61827=>"111001100",
  61828=>"100110000",
  61829=>"101111111",
  61830=>"101110101",
  61831=>"000110000",
  61832=>"010000000",
  61833=>"011110001",
  61834=>"000010110",
  61835=>"101000000",
  61836=>"111111110",
  61837=>"100010100",
  61838=>"101111100",
  61839=>"101000001",
  61840=>"111111001",
  61841=>"001101100",
  61842=>"000100000",
  61843=>"011100011",
  61844=>"011101100",
  61845=>"101000110",
  61846=>"111101111",
  61847=>"100011010",
  61848=>"100010011",
  61849=>"001101001",
  61850=>"111000011",
  61851=>"000000010",
  61852=>"010100111",
  61853=>"101100000",
  61854=>"001100111",
  61855=>"110100001",
  61856=>"001110100",
  61857=>"101001010",
  61858=>"110000101",
  61859=>"100000001",
  61860=>"010110010",
  61861=>"010001100",
  61862=>"000011011",
  61863=>"101011000",
  61864=>"000100010",
  61865=>"001011011",
  61866=>"000111011",
  61867=>"101010000",
  61868=>"111110110",
  61869=>"000100011",
  61870=>"000011000",
  61871=>"010101110",
  61872=>"000011001",
  61873=>"101001001",
  61874=>"001111101",
  61875=>"101000011",
  61876=>"010000100",
  61877=>"110000010",
  61878=>"111111111",
  61879=>"101110111",
  61880=>"001011001",
  61881=>"101100001",
  61882=>"001011011",
  61883=>"110110111",
  61884=>"110000100",
  61885=>"010100000",
  61886=>"000101000",
  61887=>"010001111",
  61888=>"000000100",
  61889=>"100011011",
  61890=>"011101100",
  61891=>"001001000",
  61892=>"111111101",
  61893=>"110000010",
  61894=>"001011000",
  61895=>"000000000",
  61896=>"110010000",
  61897=>"011100111",
  61898=>"100100011",
  61899=>"100111111",
  61900=>"100010110",
  61901=>"100111101",
  61902=>"011001011",
  61903=>"011110101",
  61904=>"000100111",
  61905=>"111110010",
  61906=>"101100001",
  61907=>"011011101",
  61908=>"000010001",
  61909=>"101101110",
  61910=>"010000000",
  61911=>"000111011",
  61912=>"001011011",
  61913=>"001001001",
  61914=>"110110010",
  61915=>"001110001",
  61916=>"010001101",
  61917=>"000111001",
  61918=>"011111000",
  61919=>"001101011",
  61920=>"100110101",
  61921=>"000011111",
  61922=>"101011101",
  61923=>"110000011",
  61924=>"000011101",
  61925=>"110010011",
  61926=>"111100111",
  61927=>"010001000",
  61928=>"010101110",
  61929=>"111111010",
  61930=>"111110000",
  61931=>"100000101",
  61932=>"010010010",
  61933=>"001011111",
  61934=>"111011110",
  61935=>"111010010",
  61936=>"000100000",
  61937=>"001111010",
  61938=>"001100010",
  61939=>"010100011",
  61940=>"110110110",
  61941=>"011010011",
  61942=>"111100101",
  61943=>"111100010",
  61944=>"000010000",
  61945=>"111001001",
  61946=>"100101001",
  61947=>"001010110",
  61948=>"000011000",
  61949=>"101011100",
  61950=>"001011010",
  61951=>"110110011",
  61952=>"111001110",
  61953=>"111100011",
  61954=>"100011000",
  61955=>"001000001",
  61956=>"111011100",
  61957=>"111111111",
  61958=>"111100001",
  61959=>"101110111",
  61960=>"111111000",
  61961=>"001011000",
  61962=>"111111010",
  61963=>"010001110",
  61964=>"001000011",
  61965=>"100000100",
  61966=>"001010000",
  61967=>"000100000",
  61968=>"100111111",
  61969=>"101101100",
  61970=>"010110101",
  61971=>"101000101",
  61972=>"011110110",
  61973=>"111110000",
  61974=>"101100001",
  61975=>"101001010",
  61976=>"110101000",
  61977=>"001100101",
  61978=>"110000100",
  61979=>"100011011",
  61980=>"111100000",
  61981=>"000100111",
  61982=>"011100100",
  61983=>"001010011",
  61984=>"100101000",
  61985=>"011100110",
  61986=>"000010100",
  61987=>"000000101",
  61988=>"001101001",
  61989=>"110101001",
  61990=>"101011101",
  61991=>"101111110",
  61992=>"100110111",
  61993=>"101101101",
  61994=>"011101010",
  61995=>"011011111",
  61996=>"110011111",
  61997=>"101101010",
  61998=>"001000000",
  61999=>"000101001",
  62000=>"100000010",
  62001=>"100101111",
  62002=>"101000010",
  62003=>"011101111",
  62004=>"001010010",
  62005=>"010000101",
  62006=>"110000010",
  62007=>"111011001",
  62008=>"111000001",
  62009=>"100101101",
  62010=>"011001010",
  62011=>"001001111",
  62012=>"101011101",
  62013=>"000001001",
  62014=>"101010110",
  62015=>"010100111",
  62016=>"100010110",
  62017=>"100111010",
  62018=>"011110111",
  62019=>"100111000",
  62020=>"100000110",
  62021=>"000001001",
  62022=>"101001101",
  62023=>"000110001",
  62024=>"000101111",
  62025=>"110010111",
  62026=>"101001000",
  62027=>"110000110",
  62028=>"010001001",
  62029=>"101000101",
  62030=>"110101111",
  62031=>"001110111",
  62032=>"000000001",
  62033=>"001010001",
  62034=>"100011100",
  62035=>"000000001",
  62036=>"011011101",
  62037=>"001010101",
  62038=>"000001010",
  62039=>"111010111",
  62040=>"110100111",
  62041=>"101111111",
  62042=>"000001001",
  62043=>"001001010",
  62044=>"111010000",
  62045=>"100001001",
  62046=>"000010001",
  62047=>"111110100",
  62048=>"111001100",
  62049=>"110110101",
  62050=>"000111010",
  62051=>"101100001",
  62052=>"000111111",
  62053=>"111011111",
  62054=>"011110110",
  62055=>"000101100",
  62056=>"010011111",
  62057=>"100111111",
  62058=>"110011011",
  62059=>"101001100",
  62060=>"000010110",
  62061=>"000001000",
  62062=>"100101001",
  62063=>"001100110",
  62064=>"011100110",
  62065=>"011110100",
  62066=>"111000000",
  62067=>"001111000",
  62068=>"111101100",
  62069=>"101011010",
  62070=>"101110101",
  62071=>"101101101",
  62072=>"010100011",
  62073=>"011001010",
  62074=>"110001001",
  62075=>"111100110",
  62076=>"101000001",
  62077=>"111000110",
  62078=>"010000100",
  62079=>"010010000",
  62080=>"000100001",
  62081=>"000110111",
  62082=>"100011101",
  62083=>"001101000",
  62084=>"011101000",
  62085=>"001000000",
  62086=>"010100011",
  62087=>"010000111",
  62088=>"111011011",
  62089=>"010000000",
  62090=>"010100001",
  62091=>"001101101",
  62092=>"101110100",
  62093=>"000010010",
  62094=>"111011111",
  62095=>"101010100",
  62096=>"001101111",
  62097=>"111101111",
  62098=>"010101110",
  62099=>"100111101",
  62100=>"001011010",
  62101=>"000101001",
  62102=>"110011110",
  62103=>"000010100",
  62104=>"111110110",
  62105=>"001111000",
  62106=>"101000000",
  62107=>"010001011",
  62108=>"010000000",
  62109=>"000100111",
  62110=>"000000110",
  62111=>"101011101",
  62112=>"100111110",
  62113=>"000100111",
  62114=>"010111100",
  62115=>"011111001",
  62116=>"101000001",
  62117=>"101101101",
  62118=>"110000110",
  62119=>"010010001",
  62120=>"010111100",
  62121=>"000010110",
  62122=>"111101011",
  62123=>"001001001",
  62124=>"010001000",
  62125=>"000011010",
  62126=>"111011010",
  62127=>"100000111",
  62128=>"001101011",
  62129=>"101110110",
  62130=>"011010010",
  62131=>"111011010",
  62132=>"010010110",
  62133=>"101001000",
  62134=>"000100011",
  62135=>"011011000",
  62136=>"111110100",
  62137=>"000010000",
  62138=>"011111001",
  62139=>"101001010",
  62140=>"000110010",
  62141=>"001010000",
  62142=>"001001101",
  62143=>"000111000",
  62144=>"111011101",
  62145=>"010101100",
  62146=>"011100000",
  62147=>"001100000",
  62148=>"000000010",
  62149=>"010000101",
  62150=>"001100001",
  62151=>"001111010",
  62152=>"100001000",
  62153=>"000100111",
  62154=>"001100010",
  62155=>"010000111",
  62156=>"101100100",
  62157=>"010111111",
  62158=>"010010101",
  62159=>"001111000",
  62160=>"100000010",
  62161=>"110010100",
  62162=>"011011100",
  62163=>"101011101",
  62164=>"001001110",
  62165=>"110010100",
  62166=>"111101110",
  62167=>"011010101",
  62168=>"010110010",
  62169=>"010001100",
  62170=>"010001101",
  62171=>"100011100",
  62172=>"001111111",
  62173=>"110101100",
  62174=>"101111101",
  62175=>"110000101",
  62176=>"001111000",
  62177=>"101101111",
  62178=>"011011001",
  62179=>"010010010",
  62180=>"011010000",
  62181=>"111000100",
  62182=>"101010110",
  62183=>"000001110",
  62184=>"110010011",
  62185=>"010100000",
  62186=>"110110000",
  62187=>"110010001",
  62188=>"001010000",
  62189=>"010100101",
  62190=>"111111111",
  62191=>"101101111",
  62192=>"000000111",
  62193=>"110111110",
  62194=>"001100111",
  62195=>"100000111",
  62196=>"110000111",
  62197=>"001001100",
  62198=>"001110000",
  62199=>"110111001",
  62200=>"111011110",
  62201=>"111101100",
  62202=>"101001010",
  62203=>"000011110",
  62204=>"110110110",
  62205=>"000011010",
  62206=>"101100001",
  62207=>"101011111",
  62208=>"101110011",
  62209=>"001010010",
  62210=>"010111110",
  62211=>"010000001",
  62212=>"000001011",
  62213=>"001100000",
  62214=>"110001010",
  62215=>"100111100",
  62216=>"000010000",
  62217=>"011001111",
  62218=>"001001000",
  62219=>"010011110",
  62220=>"011110101",
  62221=>"011000100",
  62222=>"010100111",
  62223=>"001111101",
  62224=>"011110010",
  62225=>"101000101",
  62226=>"100111110",
  62227=>"011110010",
  62228=>"001101000",
  62229=>"011001011",
  62230=>"011010101",
  62231=>"001001010",
  62232=>"000001001",
  62233=>"110011000",
  62234=>"010010111",
  62235=>"100110011",
  62236=>"010000111",
  62237=>"111000100",
  62238=>"100100011",
  62239=>"001001111",
  62240=>"101011001",
  62241=>"011110000",
  62242=>"000010011",
  62243=>"110101111",
  62244=>"110001000",
  62245=>"100000100",
  62246=>"111101011",
  62247=>"100000000",
  62248=>"011111010",
  62249=>"100000010",
  62250=>"000011001",
  62251=>"010110111",
  62252=>"000001110",
  62253=>"001101111",
  62254=>"111011010",
  62255=>"101100011",
  62256=>"011000000",
  62257=>"001100110",
  62258=>"000000010",
  62259=>"110111000",
  62260=>"101101101",
  62261=>"000111101",
  62262=>"111111101",
  62263=>"011001010",
  62264=>"100000000",
  62265=>"100000110",
  62266=>"001000110",
  62267=>"100011110",
  62268=>"000101110",
  62269=>"000100111",
  62270=>"111000010",
  62271=>"001011101",
  62272=>"100001010",
  62273=>"101001001",
  62274=>"100001111",
  62275=>"111001001",
  62276=>"011000000",
  62277=>"100101011",
  62278=>"001110101",
  62279=>"101110111",
  62280=>"010011001",
  62281=>"101101101",
  62282=>"110001000",
  62283=>"111111100",
  62284=>"100101010",
  62285=>"000101110",
  62286=>"000101110",
  62287=>"011100010",
  62288=>"110101001",
  62289=>"010101101",
  62290=>"111100111",
  62291=>"111111011",
  62292=>"111011101",
  62293=>"001011011",
  62294=>"110000011",
  62295=>"010000110",
  62296=>"011001010",
  62297=>"110000110",
  62298=>"110100011",
  62299=>"111000101",
  62300=>"011100111",
  62301=>"001100101",
  62302=>"011111111",
  62303=>"100110011",
  62304=>"000010111",
  62305=>"111110111",
  62306=>"100100110",
  62307=>"011101110",
  62308=>"001110010",
  62309=>"101010000",
  62310=>"101101100",
  62311=>"001100100",
  62312=>"011101001",
  62313=>"111101111",
  62314=>"111101100",
  62315=>"000000111",
  62316=>"100010100",
  62317=>"111100001",
  62318=>"111111000",
  62319=>"110000000",
  62320=>"110000010",
  62321=>"111110010",
  62322=>"010010110",
  62323=>"101101010",
  62324=>"010100001",
  62325=>"100111010",
  62326=>"011000000",
  62327=>"100111100",
  62328=>"110100101",
  62329=>"001000011",
  62330=>"111000001",
  62331=>"111111100",
  62332=>"101101011",
  62333=>"000110111",
  62334=>"100010110",
  62335=>"000010001",
  62336=>"111011111",
  62337=>"110000111",
  62338=>"000001101",
  62339=>"110101111",
  62340=>"110011100",
  62341=>"000110011",
  62342=>"101101111",
  62343=>"011111110",
  62344=>"100010011",
  62345=>"111010101",
  62346=>"000000110",
  62347=>"000101010",
  62348=>"100011010",
  62349=>"010000000",
  62350=>"000010011",
  62351=>"010100101",
  62352=>"100000010",
  62353=>"000111011",
  62354=>"000100111",
  62355=>"001000101",
  62356=>"001011111",
  62357=>"010100011",
  62358=>"000011111",
  62359=>"010000100",
  62360=>"110000110",
  62361=>"001100010",
  62362=>"100111011",
  62363=>"110000010",
  62364=>"000110001",
  62365=>"100100101",
  62366=>"000010010",
  62367=>"100100111",
  62368=>"001011111",
  62369=>"111111111",
  62370=>"001111110",
  62371=>"000010100",
  62372=>"010011000",
  62373=>"011100000",
  62374=>"001000110",
  62375=>"001111100",
  62376=>"001101111",
  62377=>"111111100",
  62378=>"001100001",
  62379=>"110000011",
  62380=>"000101010",
  62381=>"111011010",
  62382=>"010010011",
  62383=>"100001111",
  62384=>"011111110",
  62385=>"110100011",
  62386=>"110111000",
  62387=>"111101000",
  62388=>"011111110",
  62389=>"110000001",
  62390=>"000001010",
  62391=>"111100110",
  62392=>"100100000",
  62393=>"100000111",
  62394=>"101010011",
  62395=>"110111011",
  62396=>"010010001",
  62397=>"101101000",
  62398=>"000100001",
  62399=>"100000101",
  62400=>"000100101",
  62401=>"000110100",
  62402=>"101001111",
  62403=>"111010101",
  62404=>"111010111",
  62405=>"100001111",
  62406=>"101010001",
  62407=>"010010010",
  62408=>"111101001",
  62409=>"110000010",
  62410=>"111111100",
  62411=>"010011000",
  62412=>"111111110",
  62413=>"111101010",
  62414=>"110010111",
  62415=>"000011000",
  62416=>"111100101",
  62417=>"100011010",
  62418=>"001010001",
  62419=>"001001010",
  62420=>"100001000",
  62421=>"110011110",
  62422=>"111001010",
  62423=>"101110110",
  62424=>"110010011",
  62425=>"111101001",
  62426=>"000010000",
  62427=>"101101000",
  62428=>"101000011",
  62429=>"001110000",
  62430=>"110001101",
  62431=>"111000100",
  62432=>"000001010",
  62433=>"101100100",
  62434=>"100011000",
  62435=>"000100100",
  62436=>"011001111",
  62437=>"001000001",
  62438=>"000100011",
  62439=>"000100111",
  62440=>"000000000",
  62441=>"011011001",
  62442=>"000011000",
  62443=>"110001000",
  62444=>"101011011",
  62445=>"100111010",
  62446=>"001110000",
  62447=>"011000111",
  62448=>"011010111",
  62449=>"000111111",
  62450=>"101000101",
  62451=>"100110100",
  62452=>"100000100",
  62453=>"000001010",
  62454=>"011111111",
  62455=>"100000000",
  62456=>"000100010",
  62457=>"010011100",
  62458=>"011011011",
  62459=>"000111001",
  62460=>"111110111",
  62461=>"000110011",
  62462=>"001000001",
  62463=>"001010001",
  62464=>"000111000",
  62465=>"011011110",
  62466=>"101111011",
  62467=>"011100001",
  62468=>"100001101",
  62469=>"100101011",
  62470=>"001000001",
  62471=>"011100011",
  62472=>"111100100",
  62473=>"100111111",
  62474=>"010101111",
  62475=>"101010100",
  62476=>"000101100",
  62477=>"000000010",
  62478=>"000110010",
  62479=>"111111101",
  62480=>"100010010",
  62481=>"100100100",
  62482=>"010111101",
  62483=>"101010011",
  62484=>"100111101",
  62485=>"001101110",
  62486=>"110000010",
  62487=>"001001110",
  62488=>"010101010",
  62489=>"000011000",
  62490=>"000011111",
  62491=>"101111001",
  62492=>"000000010",
  62493=>"000001100",
  62494=>"000011010",
  62495=>"101100110",
  62496=>"001001010",
  62497=>"010001110",
  62498=>"110110111",
  62499=>"100000111",
  62500=>"100101011",
  62501=>"100010011",
  62502=>"000101100",
  62503=>"001001111",
  62504=>"000111011",
  62505=>"010000011",
  62506=>"010011100",
  62507=>"110011010",
  62508=>"110010110",
  62509=>"000000110",
  62510=>"001110111",
  62511=>"000101110",
  62512=>"111011101",
  62513=>"111110000",
  62514=>"101010001",
  62515=>"000110010",
  62516=>"110001011",
  62517=>"000101101",
  62518=>"011110011",
  62519=>"001000100",
  62520=>"100110100",
  62521=>"000100011",
  62522=>"001010101",
  62523=>"111011000",
  62524=>"001101010",
  62525=>"001000101",
  62526=>"001101001",
  62527=>"101001010",
  62528=>"101000000",
  62529=>"001110000",
  62530=>"110000111",
  62531=>"101101000",
  62532=>"111000010",
  62533=>"111100000",
  62534=>"101011001",
  62535=>"111010010",
  62536=>"000000000",
  62537=>"001011011",
  62538=>"101111000",
  62539=>"001010000",
  62540=>"001100111",
  62541=>"101011001",
  62542=>"111000001",
  62543=>"011100011",
  62544=>"010000100",
  62545=>"000011100",
  62546=>"000101110",
  62547=>"000111011",
  62548=>"111110110",
  62549=>"110010110",
  62550=>"111111111",
  62551=>"000110010",
  62552=>"110110110",
  62553=>"101110100",
  62554=>"110011011",
  62555=>"100001110",
  62556=>"100000101",
  62557=>"010011000",
  62558=>"111011101",
  62559=>"110011010",
  62560=>"010011000",
  62561=>"111000000",
  62562=>"100010000",
  62563=>"000011011",
  62564=>"000011010",
  62565=>"111011101",
  62566=>"000000111",
  62567=>"111101001",
  62568=>"011100001",
  62569=>"111110101",
  62570=>"010010000",
  62571=>"110101010",
  62572=>"010100110",
  62573=>"000110111",
  62574=>"100111010",
  62575=>"011010111",
  62576=>"110011101",
  62577=>"101101101",
  62578=>"110111101",
  62579=>"111111011",
  62580=>"000100111",
  62581=>"010101100",
  62582=>"110110100",
  62583=>"011110110",
  62584=>"000011000",
  62585=>"100010000",
  62586=>"101100100",
  62587=>"010000001",
  62588=>"011111011",
  62589=>"100101111",
  62590=>"011010101",
  62591=>"100000011",
  62592=>"011001011",
  62593=>"111000010",
  62594=>"000010110",
  62595=>"111111000",
  62596=>"111111101",
  62597=>"100010110",
  62598=>"101001010",
  62599=>"110010010",
  62600=>"110110010",
  62601=>"111000100",
  62602=>"110110010",
  62603=>"111111000",
  62604=>"000001010",
  62605=>"111001110",
  62606=>"111000100",
  62607=>"001110001",
  62608=>"010000101",
  62609=>"000000101",
  62610=>"001000001",
  62611=>"011110100",
  62612=>"111110000",
  62613=>"001110101",
  62614=>"100111001",
  62615=>"100011111",
  62616=>"010100101",
  62617=>"111000111",
  62618=>"000111101",
  62619=>"110100000",
  62620=>"010011100",
  62621=>"110101110",
  62622=>"110011110",
  62623=>"110010001",
  62624=>"010101101",
  62625=>"001111001",
  62626=>"010010010",
  62627=>"000000101",
  62628=>"011000111",
  62629=>"111011100",
  62630=>"100110001",
  62631=>"011111110",
  62632=>"111100010",
  62633=>"100011010",
  62634=>"011100001",
  62635=>"011000010",
  62636=>"111111011",
  62637=>"111101001",
  62638=>"011010101",
  62639=>"011111101",
  62640=>"000000110",
  62641=>"001011000",
  62642=>"101101010",
  62643=>"100011010",
  62644=>"110010101",
  62645=>"000111110",
  62646=>"110110111",
  62647=>"101010010",
  62648=>"111101001",
  62649=>"010000010",
  62650=>"110000000",
  62651=>"110111000",
  62652=>"010011100",
  62653=>"001111011",
  62654=>"110101101",
  62655=>"110101001",
  62656=>"011000001",
  62657=>"100000000",
  62658=>"001011011",
  62659=>"010111100",
  62660=>"100111101",
  62661=>"111110110",
  62662=>"011011001",
  62663=>"011000010",
  62664=>"111110101",
  62665=>"110101111",
  62666=>"011011011",
  62667=>"001011110",
  62668=>"000100001",
  62669=>"010101001",
  62670=>"100110100",
  62671=>"011000100",
  62672=>"101000111",
  62673=>"101010010",
  62674=>"100000010",
  62675=>"100001111",
  62676=>"010001001",
  62677=>"110100000",
  62678=>"001011110",
  62679=>"111110000",
  62680=>"110001000",
  62681=>"000011000",
  62682=>"011011001",
  62683=>"111000000",
  62684=>"111110001",
  62685=>"100011101",
  62686=>"100101000",
  62687=>"010100001",
  62688=>"111011010",
  62689=>"010011001",
  62690=>"000000101",
  62691=>"101010001",
  62692=>"101011010",
  62693=>"000101010",
  62694=>"000111111",
  62695=>"011010010",
  62696=>"100000111",
  62697=>"000000000",
  62698=>"111101000",
  62699=>"000000000",
  62700=>"010000010",
  62701=>"010110100",
  62702=>"001100110",
  62703=>"000000100",
  62704=>"010100011",
  62705=>"100010100",
  62706=>"000010001",
  62707=>"010111101",
  62708=>"111100011",
  62709=>"110011010",
  62710=>"100010010",
  62711=>"001000100",
  62712=>"101110100",
  62713=>"101110101",
  62714=>"000011110",
  62715=>"010011000",
  62716=>"001000011",
  62717=>"110110010",
  62718=>"111001111",
  62719=>"100010000",
  62720=>"010001001",
  62721=>"101110100",
  62722=>"001000011",
  62723=>"110011010",
  62724=>"011011101",
  62725=>"010001010",
  62726=>"011000000",
  62727=>"100110011",
  62728=>"111101010",
  62729=>"101000111",
  62730=>"000110110",
  62731=>"100001010",
  62732=>"011011010",
  62733=>"001010001",
  62734=>"101011001",
  62735=>"000010100",
  62736=>"100111110",
  62737=>"111101001",
  62738=>"000010110",
  62739=>"111001100",
  62740=>"000101010",
  62741=>"001000101",
  62742=>"101110001",
  62743=>"111011101",
  62744=>"111101001",
  62745=>"000010010",
  62746=>"010010110",
  62747=>"100110100",
  62748=>"000100110",
  62749=>"010010111",
  62750=>"111111000",
  62751=>"101100100",
  62752=>"011110001",
  62753=>"010110011",
  62754=>"111001111",
  62755=>"110001101",
  62756=>"000001010",
  62757=>"011011110",
  62758=>"001000001",
  62759=>"101011000",
  62760=>"001011000",
  62761=>"010011010",
  62762=>"100011000",
  62763=>"011010001",
  62764=>"110001100",
  62765=>"100101111",
  62766=>"011010000",
  62767=>"001001111",
  62768=>"011110110",
  62769=>"101011111",
  62770=>"001110010",
  62771=>"000011100",
  62772=>"101110111",
  62773=>"111111101",
  62774=>"000001000",
  62775=>"001110010",
  62776=>"001011110",
  62777=>"101101100",
  62778=>"101000111",
  62779=>"010001000",
  62780=>"100001011",
  62781=>"001101100",
  62782=>"101101011",
  62783=>"000100101",
  62784=>"010001111",
  62785=>"011001000",
  62786=>"100101000",
  62787=>"110000000",
  62788=>"110001110",
  62789=>"100101010",
  62790=>"100000010",
  62791=>"101111100",
  62792=>"100010110",
  62793=>"110010010",
  62794=>"001110111",
  62795=>"111111011",
  62796=>"010111011",
  62797=>"110001001",
  62798=>"000110111",
  62799=>"111000010",
  62800=>"001111010",
  62801=>"111001110",
  62802=>"000111001",
  62803=>"101011101",
  62804=>"011101001",
  62805=>"101000010",
  62806=>"110101000",
  62807=>"001110000",
  62808=>"011001101",
  62809=>"111101000",
  62810=>"111110011",
  62811=>"001010110",
  62812=>"011100101",
  62813=>"111100100",
  62814=>"111100001",
  62815=>"010110110",
  62816=>"001001111",
  62817=>"010011001",
  62818=>"011100000",
  62819=>"101111101",
  62820=>"001010001",
  62821=>"100100000",
  62822=>"110000101",
  62823=>"101110011",
  62824=>"101111010",
  62825=>"011110101",
  62826=>"000100110",
  62827=>"000110010",
  62828=>"001100010",
  62829=>"011110010",
  62830=>"011010110",
  62831=>"001011110",
  62832=>"001010010",
  62833=>"011100100",
  62834=>"110110100",
  62835=>"100111100",
  62836=>"100011110",
  62837=>"100011011",
  62838=>"100010011",
  62839=>"000110110",
  62840=>"110100110",
  62841=>"101110101",
  62842=>"100111101",
  62843=>"010000111",
  62844=>"000000000",
  62845=>"100011010",
  62846=>"101100010",
  62847=>"011111000",
  62848=>"010100110",
  62849=>"101100011",
  62850=>"001101101",
  62851=>"100011000",
  62852=>"100110000",
  62853=>"110000001",
  62854=>"111110101",
  62855=>"001110011",
  62856=>"011111010",
  62857=>"011011000",
  62858=>"011000011",
  62859=>"010000000",
  62860=>"101110101",
  62861=>"001011011",
  62862=>"010000101",
  62863=>"011000010",
  62864=>"110111010",
  62865=>"100110010",
  62866=>"100010000",
  62867=>"000011001",
  62868=>"111110101",
  62869=>"000011100",
  62870=>"101000010",
  62871=>"100110111",
  62872=>"010011101",
  62873=>"011100111",
  62874=>"110110100",
  62875=>"010100000",
  62876=>"100100011",
  62877=>"000111100",
  62878=>"000110101",
  62879=>"010000010",
  62880=>"000111000",
  62881=>"100000100",
  62882=>"111010011",
  62883=>"001101010",
  62884=>"100000001",
  62885=>"101001110",
  62886=>"000111000",
  62887=>"001001000",
  62888=>"111010110",
  62889=>"010110001",
  62890=>"010010101",
  62891=>"100101101",
  62892=>"100011110",
  62893=>"001010000",
  62894=>"000101100",
  62895=>"111011011",
  62896=>"000111000",
  62897=>"011010111",
  62898=>"101101001",
  62899=>"010111101",
  62900=>"001111111",
  62901=>"000101111",
  62902=>"111000110",
  62903=>"100011001",
  62904=>"000111111",
  62905=>"111001100",
  62906=>"000111101",
  62907=>"110111010",
  62908=>"101111011",
  62909=>"110010100",
  62910=>"001000010",
  62911=>"111110001",
  62912=>"010010111",
  62913=>"100010110",
  62914=>"010010111",
  62915=>"000110011",
  62916=>"000001010",
  62917=>"101100100",
  62918=>"101100001",
  62919=>"110011000",
  62920=>"001001011",
  62921=>"110011011",
  62922=>"010111010",
  62923=>"111010101",
  62924=>"111000011",
  62925=>"110010111",
  62926=>"011110011",
  62927=>"100011110",
  62928=>"111110101",
  62929=>"011110011",
  62930=>"101111101",
  62931=>"011000101",
  62932=>"010001101",
  62933=>"100100010",
  62934=>"000101010",
  62935=>"111111110",
  62936=>"101100110",
  62937=>"011011110",
  62938=>"111001010",
  62939=>"100001111",
  62940=>"100011101",
  62941=>"010010000",
  62942=>"100011100",
  62943=>"011110011",
  62944=>"010110001",
  62945=>"110000010",
  62946=>"000110001",
  62947=>"011010011",
  62948=>"100010011",
  62949=>"101111000",
  62950=>"010101111",
  62951=>"101010011",
  62952=>"001110010",
  62953=>"110010011",
  62954=>"000001010",
  62955=>"001011111",
  62956=>"000011111",
  62957=>"101010100",
  62958=>"110001100",
  62959=>"001001100",
  62960=>"100100011",
  62961=>"000100000",
  62962=>"101001001",
  62963=>"111010100",
  62964=>"110101011",
  62965=>"000100001",
  62966=>"001101110",
  62967=>"101000110",
  62968=>"010000000",
  62969=>"110111000",
  62970=>"001000000",
  62971=>"000100011",
  62972=>"001000000",
  62973=>"101011000",
  62974=>"101011110",
  62975=>"110010101",
  62976=>"001010000",
  62977=>"010000110",
  62978=>"111100010",
  62979=>"110010000",
  62980=>"010110101",
  62981=>"101110110",
  62982=>"010000110",
  62983=>"111100010",
  62984=>"110111011",
  62985=>"100110001",
  62986=>"010001110",
  62987=>"011000010",
  62988=>"110001110",
  62989=>"100110110",
  62990=>"011011000",
  62991=>"111111010",
  62992=>"110110101",
  62993=>"111000100",
  62994=>"101100101",
  62995=>"101111000",
  62996=>"010101000",
  62997=>"000100000",
  62998=>"110101101",
  62999=>"000011010",
  63000=>"001101010",
  63001=>"000111010",
  63002=>"110111100",
  63003=>"110110111",
  63004=>"011000110",
  63005=>"010110000",
  63006=>"000011011",
  63007=>"100110001",
  63008=>"110100001",
  63009=>"001111111",
  63010=>"101101011",
  63011=>"001111001",
  63012=>"011111111",
  63013=>"111000100",
  63014=>"100010000",
  63015=>"111000000",
  63016=>"010000111",
  63017=>"101000011",
  63018=>"110111101",
  63019=>"000111010",
  63020=>"011000011",
  63021=>"010001111",
  63022=>"111110101",
  63023=>"111110011",
  63024=>"110010010",
  63025=>"000111101",
  63026=>"101101001",
  63027=>"100100111",
  63028=>"011000100",
  63029=>"010011010",
  63030=>"110011101",
  63031=>"000100111",
  63032=>"101101010",
  63033=>"111111000",
  63034=>"101100010",
  63035=>"000111110",
  63036=>"001011010",
  63037=>"101011000",
  63038=>"011010110",
  63039=>"101111101",
  63040=>"001101010",
  63041=>"011011011",
  63042=>"000011000",
  63043=>"100111001",
  63044=>"101011100",
  63045=>"101000101",
  63046=>"111101011",
  63047=>"110101001",
  63048=>"101001001",
  63049=>"010101001",
  63050=>"101101000",
  63051=>"110010010",
  63052=>"110110011",
  63053=>"101101010",
  63054=>"011010101",
  63055=>"111110010",
  63056=>"110110110",
  63057=>"000100101",
  63058=>"000011110",
  63059=>"001101110",
  63060=>"001111000",
  63061=>"000011000",
  63062=>"000100010",
  63063=>"000010011",
  63064=>"010000101",
  63065=>"100110000",
  63066=>"111101111",
  63067=>"101100010",
  63068=>"011001001",
  63069=>"001011001",
  63070=>"010110001",
  63071=>"100010101",
  63072=>"001000101",
  63073=>"001011000",
  63074=>"110101101",
  63075=>"001110010",
  63076=>"110001001",
  63077=>"111111001",
  63078=>"000100111",
  63079=>"011010100",
  63080=>"101000010",
  63081=>"100000001",
  63082=>"011010100",
  63083=>"100111001",
  63084=>"110101001",
  63085=>"111011010",
  63086=>"001011010",
  63087=>"001110000",
  63088=>"010110101",
  63089=>"000101011",
  63090=>"101011010",
  63091=>"101000001",
  63092=>"011001100",
  63093=>"001000001",
  63094=>"010010010",
  63095=>"101011100",
  63096=>"010111111",
  63097=>"000010000",
  63098=>"101100101",
  63099=>"110101001",
  63100=>"101001100",
  63101=>"011011000",
  63102=>"000010001",
  63103=>"101000101",
  63104=>"101001011",
  63105=>"010010001",
  63106=>"100001011",
  63107=>"010111101",
  63108=>"100101101",
  63109=>"111100011",
  63110=>"100110101",
  63111=>"100000111",
  63112=>"100000001",
  63113=>"001011110",
  63114=>"101100111",
  63115=>"000000001",
  63116=>"101101001",
  63117=>"000100110",
  63118=>"110001001",
  63119=>"110111101",
  63120=>"011000000",
  63121=>"100011010",
  63122=>"110110111",
  63123=>"011101100",
  63124=>"111000100",
  63125=>"100100111",
  63126=>"101001101",
  63127=>"101110000",
  63128=>"011011000",
  63129=>"001000111",
  63130=>"011010011",
  63131=>"000110000",
  63132=>"011110100",
  63133=>"110001111",
  63134=>"000010010",
  63135=>"001010010",
  63136=>"001111101",
  63137=>"101010110",
  63138=>"101010110",
  63139=>"011001111",
  63140=>"011101101",
  63141=>"011011111",
  63142=>"110111001",
  63143=>"000100111",
  63144=>"000010100",
  63145=>"011100000",
  63146=>"110000101",
  63147=>"010100100",
  63148=>"011000001",
  63149=>"100100000",
  63150=>"000000010",
  63151=>"110011101",
  63152=>"101110110",
  63153=>"110000010",
  63154=>"001100100",
  63155=>"111111011",
  63156=>"100010111",
  63157=>"110010000",
  63158=>"001111001",
  63159=>"111000101",
  63160=>"011100010",
  63161=>"011101110",
  63162=>"011110001",
  63163=>"000001000",
  63164=>"101000101",
  63165=>"010110000",
  63166=>"000001110",
  63167=>"001011110",
  63168=>"011100000",
  63169=>"101101001",
  63170=>"101001010",
  63171=>"000001000",
  63172=>"110101111",
  63173=>"011010111",
  63174=>"000101010",
  63175=>"011000001",
  63176=>"100000001",
  63177=>"101111100",
  63178=>"101000101",
  63179=>"001101010",
  63180=>"111111000",
  63181=>"010011111",
  63182=>"010111111",
  63183=>"001100111",
  63184=>"111111000",
  63185=>"010011001",
  63186=>"001110000",
  63187=>"001011011",
  63188=>"001000000",
  63189=>"111110001",
  63190=>"010110000",
  63191=>"011000100",
  63192=>"111100111",
  63193=>"101110101",
  63194=>"011101101",
  63195=>"100110001",
  63196=>"111001010",
  63197=>"110100010",
  63198=>"000110011",
  63199=>"100011111",
  63200=>"101110100",
  63201=>"010011001",
  63202=>"110111110",
  63203=>"011000111",
  63204=>"110011000",
  63205=>"000001110",
  63206=>"000000000",
  63207=>"010010110",
  63208=>"100111111",
  63209=>"100000110",
  63210=>"011010000",
  63211=>"111100111",
  63212=>"010111011",
  63213=>"000100100",
  63214=>"100111110",
  63215=>"001011100",
  63216=>"000101001",
  63217=>"011000110",
  63218=>"100101101",
  63219=>"010110011",
  63220=>"101010110",
  63221=>"111100101",
  63222=>"111001111",
  63223=>"100010001",
  63224=>"111110111",
  63225=>"101110101",
  63226=>"010111101",
  63227=>"100000110",
  63228=>"010010000",
  63229=>"001000001",
  63230=>"110101011",
  63231=>"111110100",
  63232=>"000100011",
  63233=>"100111110",
  63234=>"011010111",
  63235=>"000010110",
  63236=>"100000100",
  63237=>"001011010",
  63238=>"001011011",
  63239=>"010101110",
  63240=>"100010101",
  63241=>"000001111",
  63242=>"111110001",
  63243=>"110010010",
  63244=>"100111001",
  63245=>"000101010",
  63246=>"010010010",
  63247=>"100001111",
  63248=>"000100000",
  63249=>"000001101",
  63250=>"010110100",
  63251=>"110011010",
  63252=>"110010001",
  63253=>"000110000",
  63254=>"101110100",
  63255=>"011001000",
  63256=>"111100000",
  63257=>"111001001",
  63258=>"101100000",
  63259=>"011111101",
  63260=>"110001001",
  63261=>"010101100",
  63262=>"010001010",
  63263=>"100101101",
  63264=>"011000101",
  63265=>"100011000",
  63266=>"001000110",
  63267=>"001011100",
  63268=>"000100111",
  63269=>"110110000",
  63270=>"100001011",
  63271=>"001000001",
  63272=>"100010100",
  63273=>"001110001",
  63274=>"110111111",
  63275=>"000110001",
  63276=>"010110000",
  63277=>"101110011",
  63278=>"101101101",
  63279=>"000110011",
  63280=>"110010101",
  63281=>"010101101",
  63282=>"010000110",
  63283=>"001000000",
  63284=>"001110011",
  63285=>"101111101",
  63286=>"111000100",
  63287=>"000111100",
  63288=>"011101111",
  63289=>"001001010",
  63290=>"110001011",
  63291=>"110011001",
  63292=>"000111100",
  63293=>"000110010",
  63294=>"100001100",
  63295=>"001010001",
  63296=>"000011010",
  63297=>"010011101",
  63298=>"001000010",
  63299=>"010001010",
  63300=>"011110000",
  63301=>"110111000",
  63302=>"111111001",
  63303=>"100010110",
  63304=>"001010100",
  63305=>"011100000",
  63306=>"110100010",
  63307=>"001111001",
  63308=>"110011100",
  63309=>"001000100",
  63310=>"001000010",
  63311=>"100110110",
  63312=>"011110000",
  63313=>"100101000",
  63314=>"111100001",
  63315=>"011000100",
  63316=>"110010110",
  63317=>"000101100",
  63318=>"101011010",
  63319=>"000000110",
  63320=>"011100111",
  63321=>"110001111",
  63322=>"000110001",
  63323=>"000101110",
  63324=>"110101000",
  63325=>"100110001",
  63326=>"000010101",
  63327=>"001100111",
  63328=>"100101110",
  63329=>"010010010",
  63330=>"100101011",
  63331=>"110101111",
  63332=>"010010011",
  63333=>"000011000",
  63334=>"011111010",
  63335=>"101000000",
  63336=>"011011111",
  63337=>"110111111",
  63338=>"010100010",
  63339=>"011100011",
  63340=>"001110100",
  63341=>"101001010",
  63342=>"101111000",
  63343=>"111001011",
  63344=>"110100110",
  63345=>"110001101",
  63346=>"010001111",
  63347=>"101010001",
  63348=>"110111010",
  63349=>"100011000",
  63350=>"011011111",
  63351=>"001111010",
  63352=>"011000111",
  63353=>"100001001",
  63354=>"001111111",
  63355=>"110110111",
  63356=>"011001010",
  63357=>"001101010",
  63358=>"001111010",
  63359=>"010011111",
  63360=>"111101011",
  63361=>"001101101",
  63362=>"001111111",
  63363=>"010000110",
  63364=>"000010111",
  63365=>"110111100",
  63366=>"110001001",
  63367=>"011110111",
  63368=>"010101011",
  63369=>"101001001",
  63370=>"001000110",
  63371=>"110011101",
  63372=>"111001010",
  63373=>"110110010",
  63374=>"111000010",
  63375=>"111100001",
  63376=>"000000110",
  63377=>"101111100",
  63378=>"001010111",
  63379=>"011100011",
  63380=>"001001001",
  63381=>"111110110",
  63382=>"011011011",
  63383=>"010111111",
  63384=>"011001000",
  63385=>"010001001",
  63386=>"110010001",
  63387=>"000110101",
  63388=>"001011000",
  63389=>"101000101",
  63390=>"100100000",
  63391=>"110011100",
  63392=>"010100010",
  63393=>"011010101",
  63394=>"011000000",
  63395=>"111110011",
  63396=>"101110110",
  63397=>"110010110",
  63398=>"010010111",
  63399=>"000001100",
  63400=>"010011110",
  63401=>"011011100",
  63402=>"100110011",
  63403=>"111101100",
  63404=>"000100000",
  63405=>"111111111",
  63406=>"110111100",
  63407=>"101111010",
  63408=>"111100110",
  63409=>"001110001",
  63410=>"011011001",
  63411=>"110001101",
  63412=>"000010110",
  63413=>"011001000",
  63414=>"010110010",
  63415=>"110111010",
  63416=>"110010010",
  63417=>"101010101",
  63418=>"101000100",
  63419=>"100010001",
  63420=>"101000101",
  63421=>"010111100",
  63422=>"000010111",
  63423=>"100100100",
  63424=>"010110010",
  63425=>"001001010",
  63426=>"100101011",
  63427=>"011111010",
  63428=>"110010001",
  63429=>"101001011",
  63430=>"011000100",
  63431=>"101100010",
  63432=>"010011001",
  63433=>"011010001",
  63434=>"111100001",
  63435=>"110000000",
  63436=>"010000110",
  63437=>"000001000",
  63438=>"001101100",
  63439=>"011010101",
  63440=>"110101100",
  63441=>"101011010",
  63442=>"000001111",
  63443=>"001101111",
  63444=>"110011101",
  63445=>"100011011",
  63446=>"010111111",
  63447=>"101001111",
  63448=>"111110010",
  63449=>"110101001",
  63450=>"010100111",
  63451=>"100010011",
  63452=>"101101111",
  63453=>"001001001",
  63454=>"011010101",
  63455=>"011001111",
  63456=>"011101101",
  63457=>"001011100",
  63458=>"111100101",
  63459=>"010110010",
  63460=>"101101000",
  63461=>"001101001",
  63462=>"110001001",
  63463=>"001101010",
  63464=>"101110000",
  63465=>"011111000",
  63466=>"110110001",
  63467=>"000001110",
  63468=>"111000011",
  63469=>"100111100",
  63470=>"010111001",
  63471=>"000010100",
  63472=>"100100010",
  63473=>"101011000",
  63474=>"001001101",
  63475=>"010010110",
  63476=>"010011010",
  63477=>"101000110",
  63478=>"111011000",
  63479=>"010001000",
  63480=>"000100000",
  63481=>"100011001",
  63482=>"001111111",
  63483=>"100001111",
  63484=>"100001011",
  63485=>"011111011",
  63486=>"001001110",
  63487=>"110100111",
  63488=>"110011011",
  63489=>"001100111",
  63490=>"010100111",
  63491=>"010101101",
  63492=>"000010111",
  63493=>"001111101",
  63494=>"100000111",
  63495=>"111000101",
  63496=>"110111000",
  63497=>"111111001",
  63498=>"101011001",
  63499=>"110001100",
  63500=>"000000000",
  63501=>"101101111",
  63502=>"010011010",
  63503=>"000111010",
  63504=>"000101101",
  63505=>"101000001",
  63506=>"011000110",
  63507=>"010000100",
  63508=>"111101110",
  63509=>"100100010",
  63510=>"001110011",
  63511=>"000001000",
  63512=>"000000011",
  63513=>"101110100",
  63514=>"001000010",
  63515=>"101000000",
  63516=>"110001010",
  63517=>"000011110",
  63518=>"110010010",
  63519=>"000100000",
  63520=>"000101000",
  63521=>"001011100",
  63522=>"100110011",
  63523=>"011101100",
  63524=>"010100110",
  63525=>"001100110",
  63526=>"100111100",
  63527=>"101001101",
  63528=>"001111111",
  63529=>"101100110",
  63530=>"000110101",
  63531=>"101100100",
  63532=>"111111110",
  63533=>"001010111",
  63534=>"100110000",
  63535=>"101110110",
  63536=>"101111010",
  63537=>"101000000",
  63538=>"000000100",
  63539=>"011100000",
  63540=>"111000011",
  63541=>"101100011",
  63542=>"001001000",
  63543=>"111010111",
  63544=>"001010100",
  63545=>"000011110",
  63546=>"101000000",
  63547=>"100000001",
  63548=>"010111011",
  63549=>"010110100",
  63550=>"100011001",
  63551=>"000001011",
  63552=>"100000001",
  63553=>"011001011",
  63554=>"111000000",
  63555=>"000110000",
  63556=>"010011010",
  63557=>"011111111",
  63558=>"101011011",
  63559=>"100111110",
  63560=>"010110011",
  63561=>"100001001",
  63562=>"101101100",
  63563=>"010000000",
  63564=>"001100100",
  63565=>"111010100",
  63566=>"001111100",
  63567=>"000011101",
  63568=>"001110011",
  63569=>"100001011",
  63570=>"111110011",
  63571=>"111100011",
  63572=>"001000111",
  63573=>"110000011",
  63574=>"001011101",
  63575=>"101111101",
  63576=>"010100010",
  63577=>"000010001",
  63578=>"100101101",
  63579=>"010010101",
  63580=>"101011000",
  63581=>"001000001",
  63582=>"001000001",
  63583=>"101001001",
  63584=>"011110000",
  63585=>"111110100",
  63586=>"101011001",
  63587=>"110111001",
  63588=>"011001000",
  63589=>"010010100",
  63590=>"101001010",
  63591=>"101011000",
  63592=>"101011000",
  63593=>"101011000",
  63594=>"111111000",
  63595=>"001000110",
  63596=>"011111001",
  63597=>"100100101",
  63598=>"110000011",
  63599=>"010100110",
  63600=>"010011011",
  63601=>"111000111",
  63602=>"011100000",
  63603=>"010000000",
  63604=>"010001010",
  63605=>"000000001",
  63606=>"001011101",
  63607=>"010101001",
  63608=>"000010101",
  63609=>"101010001",
  63610=>"010100000",
  63611=>"101011101",
  63612=>"111010000",
  63613=>"011011000",
  63614=>"010000011",
  63615=>"011101101",
  63616=>"011010011",
  63617=>"010000010",
  63618=>"000010000",
  63619=>"001101110",
  63620=>"010100000",
  63621=>"111100101",
  63622=>"010110111",
  63623=>"000101001",
  63624=>"110101101",
  63625=>"000101001",
  63626=>"111001010",
  63627=>"110100101",
  63628=>"111010111",
  63629=>"010000100",
  63630=>"110100000",
  63631=>"011000111",
  63632=>"000011000",
  63633=>"101110111",
  63634=>"100010111",
  63635=>"010000001",
  63636=>"010100010",
  63637=>"100000110",
  63638=>"101101000",
  63639=>"010000100",
  63640=>"011000101",
  63641=>"101101111",
  63642=>"100110001",
  63643=>"011011000",
  63644=>"100101011",
  63645=>"000001100",
  63646=>"111100010",
  63647=>"000000111",
  63648=>"000001100",
  63649=>"101000100",
  63650=>"110000000",
  63651=>"010100011",
  63652=>"000111101",
  63653=>"010010110",
  63654=>"001101101",
  63655=>"010110011",
  63656=>"101010000",
  63657=>"001100010",
  63658=>"111010110",
  63659=>"001111001",
  63660=>"110000001",
  63661=>"000110010",
  63662=>"100110100",
  63663=>"110111111",
  63664=>"001100010",
  63665=>"111101000",
  63666=>"001011011",
  63667=>"001011001",
  63668=>"010111000",
  63669=>"110011100",
  63670=>"110011110",
  63671=>"111001110",
  63672=>"000000101",
  63673=>"001101111",
  63674=>"100110101",
  63675=>"111101010",
  63676=>"111110010",
  63677=>"111001101",
  63678=>"010100101",
  63679=>"010101011",
  63680=>"011111001",
  63681=>"010111001",
  63682=>"101011100",
  63683=>"111101010",
  63684=>"101110100",
  63685=>"010111010",
  63686=>"100001011",
  63687=>"001100000",
  63688=>"100111010",
  63689=>"111110011",
  63690=>"011100100",
  63691=>"111111101",
  63692=>"010110110",
  63693=>"100101101",
  63694=>"011111110",
  63695=>"000000110",
  63696=>"100000000",
  63697=>"011110110",
  63698=>"101101100",
  63699=>"001100100",
  63700=>"100010000",
  63701=>"101111100",
  63702=>"011000010",
  63703=>"010001100",
  63704=>"011011011",
  63705=>"001111011",
  63706=>"011110111",
  63707=>"000000011",
  63708=>"011110011",
  63709=>"000010101",
  63710=>"110101010",
  63711=>"000011001",
  63712=>"011100001",
  63713=>"010010101",
  63714=>"010000000",
  63715=>"111111011",
  63716=>"111101100",
  63717=>"110011100",
  63718=>"011010110",
  63719=>"001111111",
  63720=>"010001111",
  63721=>"100111011",
  63722=>"110001101",
  63723=>"111111110",
  63724=>"111011000",
  63725=>"010110010",
  63726=>"000101000",
  63727=>"110101001",
  63728=>"000100101",
  63729=>"000011000",
  63730=>"011000100",
  63731=>"100000001",
  63732=>"001100000",
  63733=>"000110011",
  63734=>"001010111",
  63735=>"101000000",
  63736=>"111011100",
  63737=>"011010001",
  63738=>"111100100",
  63739=>"111011110",
  63740=>"011111010",
  63741=>"010001110",
  63742=>"111110011",
  63743=>"101010011",
  63744=>"111000000",
  63745=>"000101010",
  63746=>"011011110",
  63747=>"111111110",
  63748=>"100010001",
  63749=>"010000101",
  63750=>"110110100",
  63751=>"100100001",
  63752=>"110011101",
  63753=>"100010111",
  63754=>"111000100",
  63755=>"011001001",
  63756=>"111011011",
  63757=>"010000111",
  63758=>"110010000",
  63759=>"001011111",
  63760=>"011011001",
  63761=>"111011110",
  63762=>"101011110",
  63763=>"000011011",
  63764=>"101110000",
  63765=>"010100011",
  63766=>"111010001",
  63767=>"001100111",
  63768=>"000011100",
  63769=>"101100000",
  63770=>"110111011",
  63771=>"000001010",
  63772=>"000001011",
  63773=>"100111001",
  63774=>"010001100",
  63775=>"111111011",
  63776=>"101000111",
  63777=>"000000100",
  63778=>"100111101",
  63779=>"000000110",
  63780=>"111101010",
  63781=>"011001100",
  63782=>"101000111",
  63783=>"010010011",
  63784=>"100001110",
  63785=>"000101000",
  63786=>"000100010",
  63787=>"010110110",
  63788=>"110001101",
  63789=>"000110110",
  63790=>"001010111",
  63791=>"100010010",
  63792=>"100001011",
  63793=>"110101111",
  63794=>"011011111",
  63795=>"111011110",
  63796=>"100011110",
  63797=>"011010011",
  63798=>"101100101",
  63799=>"101110100",
  63800=>"100101111",
  63801=>"010001101",
  63802=>"000010101",
  63803=>"001000011",
  63804=>"010111100",
  63805=>"010001000",
  63806=>"000001011",
  63807=>"001001011",
  63808=>"001011111",
  63809=>"010000100",
  63810=>"000110010",
  63811=>"011000001",
  63812=>"111111111",
  63813=>"101010100",
  63814=>"111011011",
  63815=>"010011111",
  63816=>"001001011",
  63817=>"110101000",
  63818=>"100100010",
  63819=>"011000011",
  63820=>"110001010",
  63821=>"010110110",
  63822=>"011011010",
  63823=>"001100001",
  63824=>"010010001",
  63825=>"101110110",
  63826=>"101100000",
  63827=>"100000010",
  63828=>"010011110",
  63829=>"000010111",
  63830=>"011010011",
  63831=>"000010111",
  63832=>"111110010",
  63833=>"111010101",
  63834=>"101111101",
  63835=>"000000000",
  63836=>"001011110",
  63837=>"011010011",
  63838=>"100001011",
  63839=>"101110000",
  63840=>"001101010",
  63841=>"110111001",
  63842=>"111100111",
  63843=>"001001100",
  63844=>"011101010",
  63845=>"111111011",
  63846=>"000010110",
  63847=>"000100110",
  63848=>"110010001",
  63849=>"100001010",
  63850=>"111010101",
  63851=>"100001001",
  63852=>"100001000",
  63853=>"010110111",
  63854=>"111000100",
  63855=>"111111100",
  63856=>"001100001",
  63857=>"010011001",
  63858=>"100011100",
  63859=>"101110011",
  63860=>"100111100",
  63861=>"001111100",
  63862=>"111000101",
  63863=>"000101111",
  63864=>"100000101",
  63865=>"000011010",
  63866=>"010001111",
  63867=>"010110011",
  63868=>"001001011",
  63869=>"101011011",
  63870=>"101100100",
  63871=>"001000001",
  63872=>"111111110",
  63873=>"111011010",
  63874=>"011111010",
  63875=>"111010111",
  63876=>"010010000",
  63877=>"000110000",
  63878=>"100010101",
  63879=>"001100000",
  63880=>"110001010",
  63881=>"111011011",
  63882=>"110010101",
  63883=>"010011010",
  63884=>"111011111",
  63885=>"000011010",
  63886=>"111011010",
  63887=>"001011010",
  63888=>"111011010",
  63889=>"000011001",
  63890=>"100110100",
  63891=>"000000100",
  63892=>"010110010",
  63893=>"100011100",
  63894=>"001010100",
  63895=>"111000000",
  63896=>"100000101",
  63897=>"101101101",
  63898=>"000110111",
  63899=>"011001000",
  63900=>"011001100",
  63901=>"111001010",
  63902=>"010111111",
  63903=>"110100000",
  63904=>"000000100",
  63905=>"011000101",
  63906=>"111010100",
  63907=>"100000110",
  63908=>"001111001",
  63909=>"001011011",
  63910=>"010001000",
  63911=>"101100100",
  63912=>"111001001",
  63913=>"100111100",
  63914=>"001110011",
  63915=>"000111101",
  63916=>"000100011",
  63917=>"010010001",
  63918=>"111010000",
  63919=>"110111011",
  63920=>"111001101",
  63921=>"111100101",
  63922=>"101101011",
  63923=>"100010100",
  63924=>"010000000",
  63925=>"011000000",
  63926=>"111011011",
  63927=>"011000011",
  63928=>"010001000",
  63929=>"010111010",
  63930=>"011101100",
  63931=>"101101001",
  63932=>"111011100",
  63933=>"010110000",
  63934=>"100011011",
  63935=>"100101010",
  63936=>"001011010",
  63937=>"110110011",
  63938=>"110111110",
  63939=>"101000010",
  63940=>"111100110",
  63941=>"110010101",
  63942=>"011001111",
  63943=>"111100101",
  63944=>"010100010",
  63945=>"010101110",
  63946=>"000011010",
  63947=>"111001000",
  63948=>"100111001",
  63949=>"011001010",
  63950=>"000111011",
  63951=>"000000000",
  63952=>"100100011",
  63953=>"101011101",
  63954=>"010011010",
  63955=>"100101001",
  63956=>"001001011",
  63957=>"001110000",
  63958=>"100100000",
  63959=>"100111110",
  63960=>"110010101",
  63961=>"001000001",
  63962=>"111010110",
  63963=>"000111110",
  63964=>"111111110",
  63965=>"000101101",
  63966=>"010100110",
  63967=>"001000100",
  63968=>"001110110",
  63969=>"111010000",
  63970=>"110101101",
  63971=>"000000000",
  63972=>"101110000",
  63973=>"111111111",
  63974=>"000010101",
  63975=>"001111011",
  63976=>"101111000",
  63977=>"001010101",
  63978=>"011000010",
  63979=>"111000001",
  63980=>"101101111",
  63981=>"101011011",
  63982=>"010110110",
  63983=>"101111101",
  63984=>"000100111",
  63985=>"011101101",
  63986=>"010100001",
  63987=>"101101100",
  63988=>"100100001",
  63989=>"111111010",
  63990=>"000100001",
  63991=>"110111100",
  63992=>"011101100",
  63993=>"000000101",
  63994=>"001001000",
  63995=>"111111111",
  63996=>"100111001",
  63997=>"011011011",
  63998=>"101010110",
  63999=>"111010111",
  64000=>"111100000",
  64001=>"001111101",
  64002=>"011000101",
  64003=>"111110000",
  64004=>"111111001",
  64005=>"001001111",
  64006=>"100100001",
  64007=>"110100011",
  64008=>"000010001",
  64009=>"100011110",
  64010=>"001000000",
  64011=>"000000000",
  64012=>"100000010",
  64013=>"000011111",
  64014=>"110000110",
  64015=>"110011111",
  64016=>"001100111",
  64017=>"011010001",
  64018=>"110110011",
  64019=>"101100010",
  64020=>"000011101",
  64021=>"001001100",
  64022=>"111110101",
  64023=>"111001011",
  64024=>"001110101",
  64025=>"000010001",
  64026=>"001011101",
  64027=>"110010011",
  64028=>"010111000",
  64029=>"001111101",
  64030=>"001000101",
  64031=>"101110100",
  64032=>"000101001",
  64033=>"001111101",
  64034=>"101110111",
  64035=>"111110011",
  64036=>"010100100",
  64037=>"010110011",
  64038=>"100011010",
  64039=>"000100110",
  64040=>"000001000",
  64041=>"000100000",
  64042=>"110110100",
  64043=>"101000001",
  64044=>"011110010",
  64045=>"001110101",
  64046=>"100110111",
  64047=>"101101000",
  64048=>"100110000",
  64049=>"101111110",
  64050=>"000100111",
  64051=>"000011110",
  64052=>"101101011",
  64053=>"110010011",
  64054=>"100101010",
  64055=>"100001011",
  64056=>"001110100",
  64057=>"001001100",
  64058=>"001011101",
  64059=>"000000010",
  64060=>"000111000",
  64061=>"000011011",
  64062=>"101011010",
  64063=>"000111000",
  64064=>"011011100",
  64065=>"111000101",
  64066=>"101101111",
  64067=>"111111001",
  64068=>"001000011",
  64069=>"101011110",
  64070=>"110000010",
  64071=>"100000011",
  64072=>"100011111",
  64073=>"011110110",
  64074=>"110111010",
  64075=>"011001101",
  64076=>"000100011",
  64077=>"111100101",
  64078=>"111111111",
  64079=>"110011011",
  64080=>"101011101",
  64081=>"100110110",
  64082=>"000011110",
  64083=>"100110111",
  64084=>"000001111",
  64085=>"000000010",
  64086=>"001100101",
  64087=>"110100100",
  64088=>"010111000",
  64089=>"010101111",
  64090=>"110001100",
  64091=>"110000001",
  64092=>"010011110",
  64093=>"000101111",
  64094=>"101101001",
  64095=>"010100100",
  64096=>"100000001",
  64097=>"111001100",
  64098=>"010010011",
  64099=>"110010011",
  64100=>"011011010",
  64101=>"111100101",
  64102=>"101000101",
  64103=>"101000101",
  64104=>"000000000",
  64105=>"011110100",
  64106=>"110011101",
  64107=>"100111001",
  64108=>"100001001",
  64109=>"011001110",
  64110=>"000101110",
  64111=>"100000111",
  64112=>"110001110",
  64113=>"000111111",
  64114=>"001110000",
  64115=>"001011010",
  64116=>"011101111",
  64117=>"010001111",
  64118=>"110000010",
  64119=>"100101011",
  64120=>"011010110",
  64121=>"110000100",
  64122=>"010110101",
  64123=>"010000111",
  64124=>"001010101",
  64125=>"010001001",
  64126=>"110000111",
  64127=>"110111001",
  64128=>"111000001",
  64129=>"100101010",
  64130=>"001001000",
  64131=>"111001001",
  64132=>"100001010",
  64133=>"011000100",
  64134=>"011110000",
  64135=>"101111101",
  64136=>"110110000",
  64137=>"101001110",
  64138=>"110001010",
  64139=>"111111001",
  64140=>"110000001",
  64141=>"101101000",
  64142=>"111001000",
  64143=>"111101100",
  64144=>"110001101",
  64145=>"100101110",
  64146=>"111110100",
  64147=>"011000110",
  64148=>"011001011",
  64149=>"011111010",
  64150=>"001110000",
  64151=>"010101010",
  64152=>"000011101",
  64153=>"000011000",
  64154=>"000100111",
  64155=>"101111110",
  64156=>"111010111",
  64157=>"110001101",
  64158=>"011110101",
  64159=>"001110001",
  64160=>"010000010",
  64161=>"000100101",
  64162=>"101100001",
  64163=>"010001100",
  64164=>"110010011",
  64165=>"001000000",
  64166=>"001011001",
  64167=>"010111111",
  64168=>"110001101",
  64169=>"000100000",
  64170=>"010011000",
  64171=>"111010011",
  64172=>"110110001",
  64173=>"000000010",
  64174=>"100100100",
  64175=>"111101111",
  64176=>"011111010",
  64177=>"101010010",
  64178=>"101100100",
  64179=>"010100001",
  64180=>"101101101",
  64181=>"111110011",
  64182=>"001111000",
  64183=>"101110010",
  64184=>"000001010",
  64185=>"010001000",
  64186=>"001101100",
  64187=>"110001001",
  64188=>"000110001",
  64189=>"111000000",
  64190=>"011100011",
  64191=>"100101101",
  64192=>"111110011",
  64193=>"001100000",
  64194=>"101110101",
  64195=>"111010000",
  64196=>"001011110",
  64197=>"010011000",
  64198=>"001111111",
  64199=>"111000100",
  64200=>"000000100",
  64201=>"011101011",
  64202=>"010100011",
  64203=>"101110000",
  64204=>"101011100",
  64205=>"100010001",
  64206=>"100011011",
  64207=>"010110010",
  64208=>"110000110",
  64209=>"101101101",
  64210=>"010110101",
  64211=>"011010111",
  64212=>"100101000",
  64213=>"100101001",
  64214=>"000010101",
  64215=>"011100101",
  64216=>"010000101",
  64217=>"100100000",
  64218=>"100001100",
  64219=>"010001011",
  64220=>"110000001",
  64221=>"000001000",
  64222=>"000100011",
  64223=>"100110101",
  64224=>"011010100",
  64225=>"111111000",
  64226=>"010000111",
  64227=>"110111011",
  64228=>"001110001",
  64229=>"010111100",
  64230=>"010011001",
  64231=>"000101110",
  64232=>"110101011",
  64233=>"110010011",
  64234=>"100000100",
  64235=>"001111111",
  64236=>"001011111",
  64237=>"101111100",
  64238=>"111011111",
  64239=>"000001000",
  64240=>"100111010",
  64241=>"010011111",
  64242=>"001010101",
  64243=>"001100011",
  64244=>"011110101",
  64245=>"100011100",
  64246=>"010111101",
  64247=>"111110000",
  64248=>"010000010",
  64249=>"010000111",
  64250=>"110010101",
  64251=>"010000001",
  64252=>"001100110",
  64253=>"011011001",
  64254=>"011011101",
  64255=>"110010111",
  64256=>"000010110",
  64257=>"101111011",
  64258=>"001001111",
  64259=>"010100010",
  64260=>"110010100",
  64261=>"110000001",
  64262=>"101010000",
  64263=>"101011010",
  64264=>"111100011",
  64265=>"110000101",
  64266=>"011001000",
  64267=>"011110010",
  64268=>"010001010",
  64269=>"001111110",
  64270=>"000100001",
  64271=>"010010010",
  64272=>"001100101",
  64273=>"011000100",
  64274=>"000011110",
  64275=>"100011100",
  64276=>"000101110",
  64277=>"110010000",
  64278=>"010000100",
  64279=>"101101101",
  64280=>"101100110",
  64281=>"000011000",
  64282=>"001010110",
  64283=>"101000001",
  64284=>"001000111",
  64285=>"011110101",
  64286=>"111001010",
  64287=>"110000010",
  64288=>"000110101",
  64289=>"110111101",
  64290=>"100110101",
  64291=>"100101111",
  64292=>"010110011",
  64293=>"101000111",
  64294=>"011011100",
  64295=>"001000000",
  64296=>"101100010",
  64297=>"000011001",
  64298=>"011010011",
  64299=>"001111110",
  64300=>"011100111",
  64301=>"111100100",
  64302=>"000001101",
  64303=>"011001011",
  64304=>"110010100",
  64305=>"010100001",
  64306=>"100011000",
  64307=>"110010111",
  64308=>"010101011",
  64309=>"010100010",
  64310=>"111000000",
  64311=>"010011001",
  64312=>"001110101",
  64313=>"111000111",
  64314=>"010001100",
  64315=>"111111101",
  64316=>"010011010",
  64317=>"111101010",
  64318=>"100011101",
  64319=>"111001011",
  64320=>"110011101",
  64321=>"101101000",
  64322=>"011101011",
  64323=>"111010011",
  64324=>"010011111",
  64325=>"110000111",
  64326=>"100011111",
  64327=>"100001111",
  64328=>"101011101",
  64329=>"111001010",
  64330=>"000100011",
  64331=>"100011001",
  64332=>"011011111",
  64333=>"010101111",
  64334=>"000011101",
  64335=>"011001100",
  64336=>"000000010",
  64337=>"101100101",
  64338=>"101001011",
  64339=>"011100010",
  64340=>"000101011",
  64341=>"000100101",
  64342=>"011110111",
  64343=>"011101111",
  64344=>"110100100",
  64345=>"011001101",
  64346=>"010110010",
  64347=>"001001010",
  64348=>"111100001",
  64349=>"111010110",
  64350=>"111100101",
  64351=>"100100010",
  64352=>"100000110",
  64353=>"001011001",
  64354=>"001111011",
  64355=>"010001011",
  64356=>"101101111",
  64357=>"010101010",
  64358=>"110010101",
  64359=>"010011100",
  64360=>"111011011",
  64361=>"000100111",
  64362=>"111110101",
  64363=>"101101111",
  64364=>"001010001",
  64365=>"100001111",
  64366=>"000001001",
  64367=>"000111000",
  64368=>"011100010",
  64369=>"100011100",
  64370=>"101110001",
  64371=>"110001001",
  64372=>"000111110",
  64373=>"011100101",
  64374=>"000110111",
  64375=>"101001011",
  64376=>"010000011",
  64377=>"101111101",
  64378=>"111101111",
  64379=>"011110100",
  64380=>"111111011",
  64381=>"011101001",
  64382=>"111101111",
  64383=>"100000111",
  64384=>"001100101",
  64385=>"111011000",
  64386=>"111010100",
  64387=>"110101100",
  64388=>"000100101",
  64389=>"010100110",
  64390=>"010110010",
  64391=>"101011011",
  64392=>"101110101",
  64393=>"001011011",
  64394=>"000001011",
  64395=>"100010001",
  64396=>"000111010",
  64397=>"111110101",
  64398=>"100000010",
  64399=>"101101010",
  64400=>"101001101",
  64401=>"001100010",
  64402=>"101110011",
  64403=>"110011111",
  64404=>"111111100",
  64405=>"101011001",
  64406=>"111010110",
  64407=>"111101111",
  64408=>"100111111",
  64409=>"101001111",
  64410=>"000000010",
  64411=>"100100100",
  64412=>"110000000",
  64413=>"000101001",
  64414=>"010010000",
  64415=>"001010010",
  64416=>"101011000",
  64417=>"101111000",
  64418=>"011111110",
  64419=>"100001010",
  64420=>"100001100",
  64421=>"000001101",
  64422=>"111101110",
  64423=>"111100010",
  64424=>"100011101",
  64425=>"011100101",
  64426=>"010001011",
  64427=>"110110111",
  64428=>"101001000",
  64429=>"111110001",
  64430=>"001101110",
  64431=>"110100110",
  64432=>"011000110",
  64433=>"000100011",
  64434=>"000000111",
  64435=>"100010000",
  64436=>"100110100",
  64437=>"011010100",
  64438=>"110000110",
  64439=>"110101110",
  64440=>"101000011",
  64441=>"011111100",
  64442=>"001011110",
  64443=>"110011010",
  64444=>"100101011",
  64445=>"011010001",
  64446=>"000010111",
  64447=>"001001010",
  64448=>"000111111",
  64449=>"111111001",
  64450=>"000101010",
  64451=>"001110101",
  64452=>"000001110",
  64453=>"000000111",
  64454=>"001110000",
  64455=>"111001100",
  64456=>"011000110",
  64457=>"010000111",
  64458=>"001000000",
  64459=>"001011001",
  64460=>"000101111",
  64461=>"100001011",
  64462=>"100001000",
  64463=>"001111100",
  64464=>"111011100",
  64465=>"110110001",
  64466=>"111100010",
  64467=>"100100001",
  64468=>"011011100",
  64469=>"111011111",
  64470=>"100011010",
  64471=>"100110000",
  64472=>"110011100",
  64473=>"000000100",
  64474=>"100111000",
  64475=>"100101001",
  64476=>"001011100",
  64477=>"010001110",
  64478=>"000001010",
  64479=>"101100111",
  64480=>"001011000",
  64481=>"110001001",
  64482=>"011011011",
  64483=>"001111101",
  64484=>"101011011",
  64485=>"000010000",
  64486=>"100100100",
  64487=>"000010010",
  64488=>"011101111",
  64489=>"011100100",
  64490=>"010100000",
  64491=>"111010010",
  64492=>"000110101",
  64493=>"010110110",
  64494=>"011001000",
  64495=>"010101001",
  64496=>"110011011",
  64497=>"100100111",
  64498=>"111000010",
  64499=>"010101011",
  64500=>"101110001",
  64501=>"111000000",
  64502=>"100110101",
  64503=>"100100001",
  64504=>"011000101",
  64505=>"001011010",
  64506=>"101010001",
  64507=>"010101001",
  64508=>"001101001",
  64509=>"010101000",
  64510=>"100011001",
  64511=>"000010100",
  64512=>"110001000",
  64513=>"101000110",
  64514=>"011010101",
  64515=>"010110101",
  64516=>"101000101",
  64517=>"011100010",
  64518=>"110111011",
  64519=>"101010110",
  64520=>"011101010",
  64521=>"101111100",
  64522=>"101010001",
  64523=>"011111011",
  64524=>"001011000",
  64525=>"100001101",
  64526=>"101111101",
  64527=>"010011111",
  64528=>"101011111",
  64529=>"011111111",
  64530=>"110111101",
  64531=>"101010000",
  64532=>"010111101",
  64533=>"110001011",
  64534=>"011111011",
  64535=>"000001100",
  64536=>"011101010",
  64537=>"100101001",
  64538=>"010011011",
  64539=>"100110011",
  64540=>"111000011",
  64541=>"011100001",
  64542=>"101010100",
  64543=>"111111010",
  64544=>"101001011",
  64545=>"111001001",
  64546=>"010110111",
  64547=>"111101110",
  64548=>"101111011",
  64549=>"010000100",
  64550=>"101000001",
  64551=>"111101111",
  64552=>"101011010",
  64553=>"110000101",
  64554=>"010001100",
  64555=>"111011010",
  64556=>"100000000",
  64557=>"101110111",
  64558=>"101011101",
  64559=>"000001000",
  64560=>"100001000",
  64561=>"111110110",
  64562=>"000110011",
  64563=>"000000000",
  64564=>"011010000",
  64565=>"011000010",
  64566=>"100000100",
  64567=>"110001001",
  64568=>"111111111",
  64569=>"110101110",
  64570=>"101001000",
  64571=>"111110101",
  64572=>"001100010",
  64573=>"100100010",
  64574=>"101000101",
  64575=>"001011000",
  64576=>"000111101",
  64577=>"011111010",
  64578=>"111010101",
  64579=>"101100001",
  64580=>"100100000",
  64581=>"011011000",
  64582=>"001010000",
  64583=>"011010101",
  64584=>"011010000",
  64585=>"111111001",
  64586=>"100000001",
  64587=>"000110101",
  64588=>"100101100",
  64589=>"000111010",
  64590=>"011000111",
  64591=>"100101111",
  64592=>"111010111",
  64593=>"001011111",
  64594=>"101110110",
  64595=>"010011010",
  64596=>"000010111",
  64597=>"111111011",
  64598=>"100110101",
  64599=>"001110011",
  64600=>"111011000",
  64601=>"111101001",
  64602=>"000000001",
  64603=>"111110001",
  64604=>"100000101",
  64605=>"101011010",
  64606=>"101110100",
  64607=>"110101000",
  64608=>"000111000",
  64609=>"010010000",
  64610=>"000001101",
  64611=>"001000011",
  64612=>"101000010",
  64613=>"111111011",
  64614=>"001010010",
  64615=>"100000101",
  64616=>"010000000",
  64617=>"110111110",
  64618=>"100000011",
  64619=>"110101010",
  64620=>"010011010",
  64621=>"101100011",
  64622=>"101010010",
  64623=>"011111000",
  64624=>"111100111",
  64625=>"000100000",
  64626=>"111011010",
  64627=>"111010111",
  64628=>"010111111",
  64629=>"001010000",
  64630=>"000111010",
  64631=>"011010011",
  64632=>"011111101",
  64633=>"001111111",
  64634=>"111110110",
  64635=>"011001110",
  64636=>"111011101",
  64637=>"000010011",
  64638=>"000110010",
  64639=>"010101000",
  64640=>"000111010",
  64641=>"101001110",
  64642=>"100001001",
  64643=>"101100001",
  64644=>"000101101",
  64645=>"001100111",
  64646=>"111000010",
  64647=>"001110100",
  64648=>"001010101",
  64649=>"000101111",
  64650=>"101001101",
  64651=>"111110100",
  64652=>"010100100",
  64653=>"111011010",
  64654=>"000101101",
  64655=>"011001111",
  64656=>"111111101",
  64657=>"101110010",
  64658=>"100100010",
  64659=>"001100101",
  64660=>"110110010",
  64661=>"001011100",
  64662=>"000100010",
  64663=>"101100111",
  64664=>"010001100",
  64665=>"110010001",
  64666=>"010011100",
  64667=>"100100000",
  64668=>"000010100",
  64669=>"110000101",
  64670=>"100011011",
  64671=>"010001101",
  64672=>"101010110",
  64673=>"100101001",
  64674=>"100110100",
  64675=>"011001111",
  64676=>"101000100",
  64677=>"001000011",
  64678=>"000100000",
  64679=>"011110000",
  64680=>"110001001",
  64681=>"010001001",
  64682=>"010111101",
  64683=>"101001111",
  64684=>"010001000",
  64685=>"011000001",
  64686=>"010010100",
  64687=>"111001011",
  64688=>"010110100",
  64689=>"111111111",
  64690=>"111001011",
  64691=>"111101000",
  64692=>"001110001",
  64693=>"011010011",
  64694=>"101001001",
  64695=>"000000101",
  64696=>"101101100",
  64697=>"000000000",
  64698=>"111001000",
  64699=>"100101000",
  64700=>"011010001",
  64701=>"100110010",
  64702=>"111011111",
  64703=>"001000100",
  64704=>"011110100",
  64705=>"001001000",
  64706=>"001101111",
  64707=>"110110111",
  64708=>"000101010",
  64709=>"001011010",
  64710=>"010111011",
  64711=>"010001110",
  64712=>"001101010",
  64713=>"111011010",
  64714=>"010101110",
  64715=>"001001011",
  64716=>"110011011",
  64717=>"100100110",
  64718=>"111101010",
  64719=>"010010000",
  64720=>"100010011",
  64721=>"000001010",
  64722=>"000011101",
  64723=>"110100100",
  64724=>"101001110",
  64725=>"111100100",
  64726=>"100111111",
  64727=>"001000110",
  64728=>"100110110",
  64729=>"011111101",
  64730=>"101001000",
  64731=>"011100000",
  64732=>"001100011",
  64733=>"000010000",
  64734=>"000111010",
  64735=>"100111110",
  64736=>"000111101",
  64737=>"011000101",
  64738=>"010001101",
  64739=>"111100111",
  64740=>"110000000",
  64741=>"001000111",
  64742=>"100100010",
  64743=>"010000110",
  64744=>"001011000",
  64745=>"101101111",
  64746=>"010100111",
  64747=>"000011000",
  64748=>"101011001",
  64749=>"101000110",
  64750=>"100111010",
  64751=>"010010010",
  64752=>"110101011",
  64753=>"000100011",
  64754=>"101001110",
  64755=>"011011000",
  64756=>"101111000",
  64757=>"011100000",
  64758=>"110100111",
  64759=>"011111100",
  64760=>"001000001",
  64761=>"110110000",
  64762=>"000011101",
  64763=>"111100111",
  64764=>"000101100",
  64765=>"111010011",
  64766=>"011100111",
  64767=>"101111110",
  64768=>"101000001",
  64769=>"011011110",
  64770=>"001101011",
  64771=>"001010110",
  64772=>"101100110",
  64773=>"001101010",
  64774=>"001101100",
  64775=>"100000101",
  64776=>"010001111",
  64777=>"010001010",
  64778=>"011101010",
  64779=>"100000100",
  64780=>"110011100",
  64781=>"010010001",
  64782=>"000010101",
  64783=>"111111110",
  64784=>"111000010",
  64785=>"110101101",
  64786=>"000101000",
  64787=>"001110111",
  64788=>"100110000",
  64789=>"000000100",
  64790=>"011001111",
  64791=>"101101111",
  64792=>"011010101",
  64793=>"111101001",
  64794=>"011111001",
  64795=>"101000110",
  64796=>"000101011",
  64797=>"011111111",
  64798=>"001011110",
  64799=>"010010001",
  64800=>"110110110",
  64801=>"000010110",
  64802=>"110010111",
  64803=>"010000000",
  64804=>"001010011",
  64805=>"100000001",
  64806=>"000011111",
  64807=>"100110110",
  64808=>"011110011",
  64809=>"100110011",
  64810=>"111001000",
  64811=>"100100001",
  64812=>"101111110",
  64813=>"010010000",
  64814=>"111111111",
  64815=>"101100010",
  64816=>"010111001",
  64817=>"001100010",
  64818=>"000001001",
  64819=>"101110101",
  64820=>"101011111",
  64821=>"001111110",
  64822=>"010001100",
  64823=>"100011010",
  64824=>"011001110",
  64825=>"111001010",
  64826=>"100110000",
  64827=>"110000100",
  64828=>"100011110",
  64829=>"101101011",
  64830=>"101111011",
  64831=>"010100100",
  64832=>"100100000",
  64833=>"000100100",
  64834=>"000011000",
  64835=>"001110111",
  64836=>"100001000",
  64837=>"100111010",
  64838=>"101001101",
  64839=>"011111010",
  64840=>"000001101",
  64841=>"001111010",
  64842=>"011010000",
  64843=>"001000110",
  64844=>"000010110",
  64845=>"101011101",
  64846=>"001000001",
  64847=>"000001101",
  64848=>"100010111",
  64849=>"111010101",
  64850=>"000100010",
  64851=>"001111010",
  64852=>"100000000",
  64853=>"100110101",
  64854=>"110010110",
  64855=>"111001101",
  64856=>"000000101",
  64857=>"001100111",
  64858=>"011000011",
  64859=>"100110101",
  64860=>"010101111",
  64861=>"100110010",
  64862=>"100000010",
  64863=>"111010000",
  64864=>"110111110",
  64865=>"110000000",
  64866=>"111001100",
  64867=>"000100110",
  64868=>"011110111",
  64869=>"001100101",
  64870=>"111110101",
  64871=>"010000101",
  64872=>"011000000",
  64873=>"100000110",
  64874=>"011111011",
  64875=>"010111001",
  64876=>"111110000",
  64877=>"100101000",
  64878=>"101001001",
  64879=>"011111101",
  64880=>"011001110",
  64881=>"010111001",
  64882=>"000010011",
  64883=>"010110100",
  64884=>"110100011",
  64885=>"111111000",
  64886=>"010100101",
  64887=>"110001101",
  64888=>"100100000",
  64889=>"001100101",
  64890=>"101110111",
  64891=>"101110010",
  64892=>"001101110",
  64893=>"111111000",
  64894=>"001010100",
  64895=>"011111101",
  64896=>"101110111",
  64897=>"011001011",
  64898=>"000001011",
  64899=>"111100011",
  64900=>"110011100",
  64901=>"101110000",
  64902=>"000100111",
  64903=>"100011011",
  64904=>"111110000",
  64905=>"000100000",
  64906=>"000011001",
  64907=>"010001011",
  64908=>"101110111",
  64909=>"010010111",
  64910=>"000100011",
  64911=>"010101010",
  64912=>"111101110",
  64913=>"101111010",
  64914=>"101000111",
  64915=>"011111000",
  64916=>"001001011",
  64917=>"000110001",
  64918=>"111100101",
  64919=>"011010100",
  64920=>"100010100",
  64921=>"000100101",
  64922=>"111010011",
  64923=>"000000000",
  64924=>"100011010",
  64925=>"000011100",
  64926=>"110101001",
  64927=>"100110010",
  64928=>"001011010",
  64929=>"110001001",
  64930=>"100101100",
  64931=>"000001000",
  64932=>"110111110",
  64933=>"001000111",
  64934=>"010111000",
  64935=>"000000101",
  64936=>"111011011",
  64937=>"010100001",
  64938=>"100100011",
  64939=>"111011110",
  64940=>"110101010",
  64941=>"000011010",
  64942=>"001011000",
  64943=>"100010000",
  64944=>"010100110",
  64945=>"100100101",
  64946=>"010110111",
  64947=>"101010101",
  64948=>"000011001",
  64949=>"110111100",
  64950=>"101110001",
  64951=>"100101100",
  64952=>"110000101",
  64953=>"010000000",
  64954=>"101110101",
  64955=>"011001110",
  64956=>"100000011",
  64957=>"010011110",
  64958=>"011001010",
  64959=>"001011100",
  64960=>"111001110",
  64961=>"100101100",
  64962=>"010011100",
  64963=>"111110111",
  64964=>"010000000",
  64965=>"011111111",
  64966=>"011101110",
  64967=>"000110110",
  64968=>"001000000",
  64969=>"000011111",
  64970=>"100000010",
  64971=>"011111011",
  64972=>"101011110",
  64973=>"110000000",
  64974=>"010001000",
  64975=>"000101110",
  64976=>"110000010",
  64977=>"110010111",
  64978=>"111000000",
  64979=>"011101111",
  64980=>"111000010",
  64981=>"001100000",
  64982=>"111100001",
  64983=>"010010111",
  64984=>"010011111",
  64985=>"001010110",
  64986=>"100110111",
  64987=>"001110111",
  64988=>"011000000",
  64989=>"101110001",
  64990=>"000100111",
  64991=>"011001001",
  64992=>"101110010",
  64993=>"111111011",
  64994=>"000110110",
  64995=>"001111101",
  64996=>"001010011",
  64997=>"010110001",
  64998=>"001101100",
  64999=>"000001101",
  65000=>"110010101",
  65001=>"011110111",
  65002=>"000010110",
  65003=>"111000110",
  65004=>"110110001",
  65005=>"110100001",
  65006=>"111001001",
  65007=>"111110001",
  65008=>"110110011",
  65009=>"100100000",
  65010=>"111110100",
  65011=>"111110000",
  65012=>"111001010",
  65013=>"100111101",
  65014=>"011011101",
  65015=>"100011100",
  65016=>"111100101",
  65017=>"110011010",
  65018=>"011000011",
  65019=>"011001001",
  65020=>"100101111",
  65021=>"111110001",
  65022=>"010001000",
  65023=>"110111110",
  65024=>"100010111",
  65025=>"111001111",
  65026=>"000001100",
  65027=>"110101011",
  65028=>"000100100",
  65029=>"111000011",
  65030=>"000100100",
  65031=>"101110111",
  65032=>"010110000",
  65033=>"001000100",
  65034=>"011110001",
  65035=>"100001011",
  65036=>"001110000",
  65037=>"101010100",
  65038=>"000101011",
  65039=>"111001011",
  65040=>"001111010",
  65041=>"110010011",
  65042=>"110110110",
  65043=>"110100001",
  65044=>"111001101",
  65045=>"010110110",
  65046=>"111001011",
  65047=>"010011010",
  65048=>"111111010",
  65049=>"010111011",
  65050=>"000000011",
  65051=>"101010110",
  65052=>"011101110",
  65053=>"100000101",
  65054=>"100100101",
  65055=>"100001001",
  65056=>"101011000",
  65057=>"010011100",
  65058=>"001011000",
  65059=>"000000100",
  65060=>"000010111",
  65061=>"100001111",
  65062=>"011010010",
  65063=>"101110001",
  65064=>"001000101",
  65065=>"001100110",
  65066=>"101000110",
  65067=>"101100111",
  65068=>"101110011",
  65069=>"000010010",
  65070=>"110010011",
  65071=>"000100010",
  65072=>"100011000",
  65073=>"010111111",
  65074=>"010011001",
  65075=>"101110111",
  65076=>"011000111",
  65077=>"110110101",
  65078=>"111111010",
  65079=>"000100010",
  65080=>"100101010",
  65081=>"010000101",
  65082=>"000111111",
  65083=>"101010011",
  65084=>"111011111",
  65085=>"101110000",
  65086=>"011001111",
  65087=>"011110101",
  65088=>"011110111",
  65089=>"001111000",
  65090=>"001001111",
  65091=>"101111001",
  65092=>"010111001",
  65093=>"110010100",
  65094=>"000011101",
  65095=>"001000100",
  65096=>"000100001",
  65097=>"010101110",
  65098=>"100010011",
  65099=>"111011111",
  65100=>"110110111",
  65101=>"110110000",
  65102=>"110011110",
  65103=>"001000000",
  65104=>"100111111",
  65105=>"010101101",
  65106=>"110001100",
  65107=>"011101100",
  65108=>"010001010",
  65109=>"011111001",
  65110=>"000110001",
  65111=>"001011111",
  65112=>"001100000",
  65113=>"111100000",
  65114=>"101001010",
  65115=>"110001010",
  65116=>"101100101",
  65117=>"001000011",
  65118=>"010100010",
  65119=>"110111111",
  65120=>"011110101",
  65121=>"000000001",
  65122=>"011001000",
  65123=>"110101101",
  65124=>"110111010",
  65125=>"101000011",
  65126=>"101001110",
  65127=>"100010110",
  65128=>"101010101",
  65129=>"011100110",
  65130=>"111111001",
  65131=>"001111000",
  65132=>"000000000",
  65133=>"111011011",
  65134=>"001010111",
  65135=>"010000011",
  65136=>"001101010",
  65137=>"011110100",
  65138=>"101111001",
  65139=>"001101110",
  65140=>"100110111",
  65141=>"000100000",
  65142=>"101101000",
  65143=>"000001000",
  65144=>"001000110",
  65145=>"000001111",
  65146=>"100000011",
  65147=>"000010001",
  65148=>"010011101",
  65149=>"011000111",
  65150=>"011111001",
  65151=>"101001110",
  65152=>"010000001",
  65153=>"001101101",
  65154=>"111001000",
  65155=>"111001101",
  65156=>"010110111",
  65157=>"100000100",
  65158=>"111101101",
  65159=>"110110110",
  65160=>"111101110",
  65161=>"011100110",
  65162=>"111101111",
  65163=>"000101100",
  65164=>"011100101",
  65165=>"101010100",
  65166=>"010001000",
  65167=>"011011111",
  65168=>"011001111",
  65169=>"101111111",
  65170=>"101001110",
  65171=>"111110101",
  65172=>"110011101",
  65173=>"000011010",
  65174=>"101100110",
  65175=>"011001100",
  65176=>"000101010",
  65177=>"110001101",
  65178=>"001110010",
  65179=>"011011000",
  65180=>"110011100",
  65181=>"011000001",
  65182=>"001011100",
  65183=>"100000001",
  65184=>"100000000",
  65185=>"110001000",
  65186=>"110111111",
  65187=>"111111101",
  65188=>"100011101",
  65189=>"001010110",
  65190=>"111011100",
  65191=>"000101110",
  65192=>"000000010",
  65193=>"000011000",
  65194=>"000011100",
  65195=>"001111110",
  65196=>"110110100",
  65197=>"111110111",
  65198=>"000010000",
  65199=>"000011011",
  65200=>"101011010",
  65201=>"011100110",
  65202=>"000111010",
  65203=>"011110111",
  65204=>"001000011",
  65205=>"111110011",
  65206=>"110010100",
  65207=>"100100010",
  65208=>"110111001",
  65209=>"010101011",
  65210=>"010110111",
  65211=>"101001111",
  65212=>"011111000",
  65213=>"001101011",
  65214=>"000000000",
  65215=>"011110010",
  65216=>"111100100",
  65217=>"101110100",
  65218=>"001110000",
  65219=>"101101100",
  65220=>"100010011",
  65221=>"000110100",
  65222=>"100001100",
  65223=>"110111101",
  65224=>"100101101",
  65225=>"101101101",
  65226=>"111011111",
  65227=>"001100000",
  65228=>"011111111",
  65229=>"011111111",
  65230=>"101110110",
  65231=>"110110001",
  65232=>"001001100",
  65233=>"100000000",
  65234=>"001110011",
  65235=>"100000101",
  65236=>"101110110",
  65237=>"011000111",
  65238=>"100100101",
  65239=>"101110001",
  65240=>"100110100",
  65241=>"100101010",
  65242=>"111001101",
  65243=>"010001101",
  65244=>"100100011",
  65245=>"100011000",
  65246=>"000111111",
  65247=>"110100100",
  65248=>"000100000",
  65249=>"011011010",
  65250=>"110100101",
  65251=>"011001011",
  65252=>"101100000",
  65253=>"011110101",
  65254=>"101101011",
  65255=>"010000001",
  65256=>"100101101",
  65257=>"001101001",
  65258=>"100010111",
  65259=>"111100101",
  65260=>"101001110",
  65261=>"110111101",
  65262=>"011011000",
  65263=>"010000111",
  65264=>"100110001",
  65265=>"100111110",
  65266=>"110100000",
  65267=>"001110010",
  65268=>"010001111",
  65269=>"001001111",
  65270=>"110000000",
  65271=>"000010101",
  65272=>"100111001",
  65273=>"111101110",
  65274=>"011101011",
  65275=>"111010101",
  65276=>"001001110",
  65277=>"110100000",
  65278=>"010111000",
  65279=>"111111010",
  65280=>"010111100",
  65281=>"110001101",
  65282=>"111100011",
  65283=>"001000000",
  65284=>"001001011",
  65285=>"001111111",
  65286=>"111100101",
  65287=>"010010001",
  65288=>"010000000",
  65289=>"100100101",
  65290=>"101111001",
  65291=>"111010000",
  65292=>"100100011",
  65293=>"101000011",
  65294=>"101011110",
  65295=>"001101011",
  65296=>"000101001",
  65297=>"001000001",
  65298=>"111011000",
  65299=>"010111001",
  65300=>"010011001",
  65301=>"100010110",
  65302=>"100110111",
  65303=>"001000000",
  65304=>"010100000",
  65305=>"000011010",
  65306=>"110000001",
  65307=>"110010010",
  65308=>"010110000",
  65309=>"010110111",
  65310=>"001101011",
  65311=>"000111111",
  65312=>"111011100",
  65313=>"110000010",
  65314=>"101000011",
  65315=>"010101000",
  65316=>"100000000",
  65317=>"000100100",
  65318=>"000110010",
  65319=>"100100000",
  65320=>"101110010",
  65321=>"111111010",
  65322=>"010101101",
  65323=>"101010111",
  65324=>"111000101",
  65325=>"101000001",
  65326=>"001100111",
  65327=>"010010111",
  65328=>"110110010",
  65329=>"100101100",
  65330=>"011011110",
  65331=>"010010011",
  65332=>"000111111",
  65333=>"011111011",
  65334=>"010000101",
  65335=>"100010110",
  65336=>"011111101",
  65337=>"011110001",
  65338=>"100101111",
  65339=>"001000000",
  65340=>"111100010",
  65341=>"000111001",
  65342=>"100001010",
  65343=>"010000001",
  65344=>"011011111",
  65345=>"110010110",
  65346=>"011001100",
  65347=>"000010100",
  65348=>"101111111",
  65349=>"111111101",
  65350=>"100000111",
  65351=>"111011001",
  65352=>"010110011",
  65353=>"001101100",
  65354=>"110111111",
  65355=>"011111010",
  65356=>"011010101",
  65357=>"111011110",
  65358=>"010001101",
  65359=>"100110111",
  65360=>"011111010",
  65361=>"100010010",
  65362=>"011100001",
  65363=>"011000010",
  65364=>"011110111",
  65365=>"000101000",
  65366=>"000011000",
  65367=>"100111111",
  65368=>"001011101",
  65369=>"001010000",
  65370=>"000111011",
  65371=>"111000101",
  65372=>"001000010",
  65373=>"100100100",
  65374=>"101000010",
  65375=>"000100110",
  65376=>"100011000",
  65377=>"110101010",
  65378=>"111111011",
  65379=>"111111011",
  65380=>"110000001",
  65381=>"110101001",
  65382=>"101010010",
  65383=>"001111100",
  65384=>"111000011",
  65385=>"011111001",
  65386=>"101111001",
  65387=>"001011000",
  65388=>"111011101",
  65389=>"101110010",
  65390=>"000110100",
  65391=>"000011010",
  65392=>"001101111",
  65393=>"100001000",
  65394=>"111101001",
  65395=>"110010111",
  65396=>"100010111",
  65397=>"111011100",
  65398=>"111010010",
  65399=>"111000011",
  65400=>"011110111",
  65401=>"111001010",
  65402=>"100010001",
  65403=>"011110111",
  65404=>"110011000",
  65405=>"110010010",
  65406=>"111010111",
  65407=>"011101101",
  65408=>"111001001",
  65409=>"011100000",
  65410=>"011010111",
  65411=>"011100000",
  65412=>"111100010",
  65413=>"111100101",
  65414=>"000101110",
  65415=>"001101111",
  65416=>"100000010",
  65417=>"110010011",
  65418=>"111111001",
  65419=>"101101111",
  65420=>"100100001",
  65421=>"110011001",
  65422=>"110110101",
  65423=>"000011011",
  65424=>"000110000",
  65425=>"101101111",
  65426=>"000111111",
  65427=>"100001100",
  65428=>"001101110",
  65429=>"000101001",
  65430=>"101010101",
  65431=>"011010010",
  65432=>"001000011",
  65433=>"000110001",
  65434=>"110101001",
  65435=>"010111011",
  65436=>"101001011",
  65437=>"100100000",
  65438=>"001010101",
  65439=>"000101011",
  65440=>"001000011",
  65441=>"000111011",
  65442=>"000001100",
  65443=>"101100011",
  65444=>"101110101",
  65445=>"101110110",
  65446=>"011011000",
  65447=>"110111000",
  65448=>"101011000",
  65449=>"111111001",
  65450=>"001101110",
  65451=>"001111010",
  65452=>"010100111",
  65453=>"000000101",
  65454=>"110001101",
  65455=>"010111100",
  65456=>"001110011",
  65457=>"011100001",
  65458=>"100110101",
  65459=>"100101100",
  65460=>"100011110",
  65461=>"011010101",
  65462=>"110110001",
  65463=>"101000011",
  65464=>"110000011",
  65465=>"100011001",
  65466=>"100001001",
  65467=>"110000110",
  65468=>"111001001",
  65469=>"010011111",
  65470=>"100101010",
  65471=>"000010100",
  65472=>"101011110",
  65473=>"001001011",
  65474=>"000000111",
  65475=>"001100110",
  65476=>"000001011",
  65477=>"101011110",
  65478=>"111100101",
  65479=>"111001010",
  65480=>"111000001",
  65481=>"101011101",
  65482=>"001110001",
  65483=>"100100110",
  65484=>"011110110",
  65485=>"111100010",
  65486=>"100111011",
  65487=>"011111110",
  65488=>"101010010",
  65489=>"110010000",
  65490=>"011010111",
  65491=>"110000110",
  65492=>"010001000",
  65493=>"010100101",
  65494=>"100111000",
  65495=>"111111101",
  65496=>"110110000",
  65497=>"000011011",
  65498=>"010000001",
  65499=>"100110010",
  65500=>"010010010",
  65501=>"010001011",
  65502=>"100100110",
  65503=>"101001110",
  65504=>"000101010",
  65505=>"010000010",
  65506=>"110110011",
  65507=>"101001110",
  65508=>"001111000",
  65509=>"111000111",
  65510=>"111011111",
  65511=>"110101000",
  65512=>"000011000",
  65513=>"111000000",
  65514=>"110101111",
  65515=>"000111111",
  65516=>"111100111",
  65517=>"101010011",
  65518=>"000001100",
  65519=>"001111011",
  65520=>"101011011",
  65521=>"010101000",
  65522=>"010001011",
  65523=>"100111000",
  65524=>"000110011",
  65525=>"111011101",
  65526=>"001111101",
  65527=>"111110111",
  65528=>"000100000",
  65529=>"010011110",
  65530=>"111111010",
  65531=>"110001101",
  65532=>"010001101",
  65533=>"010001101",
  65534=>"011000010",
  65535=>"010110100");

BEGIN
  weight <= ROM_content(to_integer(address));
END RTL;