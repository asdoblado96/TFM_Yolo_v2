LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L7_8_BNROM IS
  PORT (
    coefs : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    address : IN unsigned(6 DOWNTO 0));
END L7_8_BNROM;

ARCHITECTURE RTL OF L7_8_BNROM IS

  TYPE ROM_mem IS ARRAY (0 TO 127) OF STD_LOGIC_VECTOR(31 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem :=

  --Contenido bias || scale
  (0=>"1111110101101001"&"0010010011010000",
  1=>"1111011001000001"&"0010110011011101",
  2=>"1110110100100001"&"0010011011010101",
  3=>"1110110001101100"&"0010001110111110",
  4=>"1111000000101101"&"0010001101000101",
  5=>"1110010110111110"&"0010010111100011",
  6=>"1110110000110111"&"0010010101101100",
  7=>"1111001100010000"&"0010001001010010",
  8=>"1110111011111001"&"0010001110010001",
  9=>"1111010010010000"&"0010101111001010",
  10=>"1101101100011111"&"0010100110111111",
  11=>"1110011111111000"&"0010101010011111",
  12=>"1101111101011000"&"0010011100000001",
  13=>"1111001001000001"&"0010100001100100",
  14=>"1101110111100000"&"0010101100010111",
  15=>"1110111010001111"&"0010100011010110",
  16=>"1111010101110011"&"0010101110001100",
  17=>"1111011111010001"&"0010100001100111",
  18=>"1110110011111001"&"0001101010001111",
  19=>"1111000011001011"&"0010001001010011",
  20=>"1111111010010010"&"0010001011111010",
  21=>"1111011111000101"&"0010010011101100",
  22=>"0000011101011000"&"0010101111100111",
  23=>"1101111110101000"&"0010110010010010",
  24=>"1110010100101111"&"0010101001011100",
  25=>"1100101001000101"&"0010010001001111",
  26=>"1111010000001100"&"0010011101001100",
  27=>"1111101010110101"&"0010001000110100",
  28=>"1110101101111100"&"0010110100110101",
  29=>"1110101001110100"&"0010001010001101",
  30=>"1110101100011111"&"0010100000101000",
  31=>"1111100001010111"&"0010101010101001",
  32=>"1110111011111100"&"0010000011010101",
  33=>"1110111011101001"&"0010011011110001",
  34=>"1110110100001100"&"0010101000001111",
  35=>"1110011111010100"&"0010010100001001",
  36=>"1101111110100111"&"0001111110010010",
  37=>"1101011110001101"&"0011000100100000",
  38=>"1111000100100011"&"0010010101110000",
  39=>"1110111000110111"&"0010100110100001",
  40=>"1110111110101010"&"0010000101110011",
  41=>"1101001010101111"&"0010000100011100",
  42=>"1111010111110100"&"0010011000101110",
  43=>"1110101010011010"&"0010111111010100",
  44=>"1110101000010110"&"0010001110010100",
  45=>"1111000010000010"&"0010010001010011",
  46=>"1110111110110110"&"0010010000001010",
  47=>"1110010101001010"&"0010100010001011",
  48=>"1111101111110000"&"0010010100100110",
  49=>"1101110110000011"&"0010011100101110",
  50=>"1110111010100100"&"0010100011111010",
  51=>"1111011101001011"&"0010100110110011",
  52=>"1110101110000010"&"0010101110010010",
  53=>"1110110011011001"&"0010010011011100",
  54=>"1110100001110000"&"0010100101100001",
  55=>"1111011000100000"&"0010011111110010",
  56=>"1110101011001000"&"0010011010000110",
  57=>"1111111111111100"&"0010010110111111",
  58=>"1111000101011010"&"0010000011111000",
  59=>"1110111110011000"&"0010010011010110",
  60=>"1110101100110010"&"0010100110000111",
  61=>"1111100100010010"&"0010001000001101",
  62=>"1111011000110000"&"0010100001110111",
  63=>"1110110101110010"&"0010011101111110",
  64=>"1111001010101110"&"0010101001110001",
  65=>"1110111000010010"&"0010000101101100",
  66=>"1110011010001101"&"0010110010011010",
  67=>"0000001010011001"&"0010011000110111",
  68=>"1111000001001001"&"0010011101101001",
  69=>"1110010001000100"&"0010110000000110",
  70=>"1111111010010111"&"0001111111010101",
  71=>"0000000011100000"&"0010011001001001",
  72=>"1110101111101001"&"0001110111010100",
  73=>"1110110010011011"&"0010010010010111",
  74=>"1110110010001000"&"0010010110110011",
  75=>"1111101000000010"&"0010010100001010",
  76=>"1110111010100010"&"0010011001100001",
  77=>"1101000011110000"&"0010100110110101",
  78=>"1110110110100111"&"0001110100110101",
  79=>"1111010101000000"&"0010010100100000",
  80=>"1110111111101001"&"0010010001010010",
  81=>"1111000011110111"&"0010001111010110",
  82=>"1111000011100111"&"0010100101010011",
  83=>"1111011111101000"&"0010000110001011",
  84=>"1101111110000111"&"0010100011000101",
  85=>"1110101101010101"&"0010011101101110",
  86=>"1111000101111101"&"0010010010111000",
  87=>"1101101101011011"&"0010100011011001",
  88=>"1111000101011001"&"0010010100011100",
  89=>"1111000110001110"&"0010001001001011",
  90=>"1111000110010100"&"0010010100111011",
  91=>"1110001101010011"&"0010010011100100",
  92=>"1111010111100001"&"0010010101001011",
  93=>"1111010100110111"&"0010101011110100",
  94=>"1110110000000011"&"0010101000111010",
  95=>"1110110001011010"&"0010100101111100",
  96=>"1110110000001011"&"0010100010110000",
  97=>"1110111101110011"&"0010001111001000",
  98=>"1111011100110101"&"0001110011100101",
  99=>"1111010011101101"&"0010000001110000",
  100=>"1110101110010011"&"0001010011100001",
  101=>"1110111110111110"&"0010101010010001",
  102=>"1111001001101010"&"0010011000001111",
  103=>"1111010000111010"&"0010010100001000",
  104=>"1110001001011101"&"0010001101011011",
  105=>"1111011000010001"&"0010001010101100",
  106=>"1111000100101110"&"0010010010011011",
  107=>"1111100100110010"&"0010001010111110",
  108=>"1111010011010111"&"0010000011111101",
  109=>"1111001100000100"&"0010011110010101",
  110=>"1110011000110010"&"0010000110101110",
  111=>"1110100110100111"&"0010100000101000",
  112=>"1111111000000100"&"0010000000010111",
  113=>"1110111110110000"&"0010011001111000",
  114=>"1111010011010110"&"0010010110010000",
  115=>"1110011010011110"&"0010011000101101",
  116=>"0000011101010100"&"0010011000011010",
  117=>"1101110100111001"&"0010000011100101",
  118=>"1111010111101100"&"0010010111011110",
  119=>"1111000100100100"&"0010100111110010",
  120=>"1110100101010100"&"0010011111101000",
  121=>"1111000010010101"&"0010000000011111",
  122=>"1111101100001010"&"0010011010111010",
  123=>"1110101111100100"&"0010101110111010",
  124=>"1111100011110001"&"0010011000000100",
  125=>"1111011000110111"&"0010011100011000",
  126=>"1110101011100011"&"0010101110100011",
  127=>"0000000000001111"&"0010011101110101");

BEGIN
  coefs <= ROM_content(to_integer(address));
END RTL;