LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L5_2_WROM IS
    PORT (
        weight : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
        address : IN unsigned(weightsbitsAddress(5)-1 DOWNTO 0));
END L5_2_WROM;

ARCHITECTURE RTL OF L5_2_WROM IS

    TYPE ROM_mem IS ARRAY (0 TO 16383) OF STD_LOGIC_VECTOR(8 DOWNTO 0);

    CONSTANT ROM_content : ROM_mem := (
        0=>"101101110",
        1=>"111111000",
        2=>"111100000",
        3=>"010010000",
        4=>"001000000",
        5=>"000010111",
        6=>"111111111",
        7=>"000111000",
        8=>"000011111",
        9=>"010110111",
        10=>"111110000",
        11=>"011111101",
        12=>"110000111",
        13=>"110010010",
        14=>"010000011",
        15=>"001100000",
        16=>"000000011",
        17=>"100111011",
        18=>"000000001",
        19=>"111110100",
        20=>"100100000",
        21=>"000000001",
        22=>"111011000",
        23=>"111111101",
        24=>"010001000",
        25=>"000110100",
        26=>"000000001",
        27=>"000000110",
        28=>"000000111",
        29=>"000000000",
        30=>"000000011",
        31=>"100001111",
        32=>"000000011",
        33=>"000010101",
        34=>"000001001",
        35=>"100000000",
        36=>"010111101",
        37=>"000110110",
        38=>"110101101",
        39=>"111111000",
        40=>"111111000",
        41=>"101110100",
        42=>"010000001",
        43=>"000100101",
        44=>"010001001",
        45=>"000100000",
        46=>"000100101",
        47=>"110111000",
        48=>"100100000",
        49=>"111111000",
        50=>"000001001",
        51=>"011001111",
        52=>"000000100",
        53=>"000111111",
        54=>"000011111",
        55=>"101000011",
        56=>"100111000",
        57=>"000000111",
        58=>"000100100",
        59=>"100011000",
        60=>"011111000",
        61=>"011111001",
        62=>"000000111",
        63=>"100011111",
        64=>"111111000",
        65=>"011101110",
        66=>"111111110",
        67=>"101000000",
        68=>"100000010",
        69=>"011011000",
        70=>"000010000",
        71=>"111111111",
        72=>"000010110",
        73=>"111000101",
        74=>"111111000",
        75=>"000101101",
        76=>"110000101",
        77=>"001100000",
        78=>"000000110",
        79=>"111101000",
        80=>"111111000",
        81=>"111111000",
        82=>"000100111",
        83=>"000000010",
        84=>"110110101",
        85=>"111000000",
        86=>"001000011",
        87=>"000010111",
        88=>"000001000",
        89=>"001111111",
        90=>"100000110",
        91=>"111111000",
        92=>"000000111",
        93=>"110011001",
        94=>"011000000",
        95=>"111000010",
        96=>"000100110",
        97=>"111110000",
        98=>"111101000",
        99=>"111111000",
        100=>"000100100",
        101=>"000011101",
        102=>"110001000",
        103=>"110011110",
        104=>"101011001",
        105=>"001100100",
        106=>"110100110",
        107=>"101111111",
        108=>"100000001",
        109=>"011101000",
        110=>"000000011",
        111=>"000000111",
        112=>"111111101",
        113=>"111101001",
        114=>"010000000",
        115=>"000010011",
        116=>"111100000",
        117=>"111101000",
        118=>"000100010",
        119=>"000000110",
        120=>"111001000",
        121=>"001000000",
        122=>"100000100",
        123=>"000010011",
        124=>"000000111",
        125=>"000111110",
        126=>"000000100",
        127=>"011100110",
        128=>"111111101",
        129=>"110110000",
        130=>"111011111",
        131=>"110111100",
        132=>"110000110",
        133=>"100010000",
        134=>"000011001",
        135=>"001001111",
        136=>"000000000",
        137=>"000000010",
        138=>"111111000",
        139=>"111110011",
        140=>"000101111",
        141=>"110010100",
        142=>"111111001",
        143=>"000001111",
        144=>"111011111",
        145=>"000000101",
        146=>"100000011",
        147=>"111111101",
        148=>"001000111",
        149=>"000000000",
        150=>"000000000",
        151=>"111111111",
        152=>"111110111",
        153=>"111111111",
        154=>"110111000",
        155=>"011111111",
        156=>"001101110",
        157=>"001000000",
        158=>"111111011",
        159=>"010010111",
        160=>"100101111",
        161=>"100100110",
        162=>"110110110",
        163=>"000001111",
        164=>"000001111",
        165=>"001001000",
        166=>"000000000",
        167=>"001111111",
        168=>"010001111",
        169=>"111000001",
        170=>"111101101",
        171=>"010001000",
        172=>"000010011",
        173=>"000000011",
        174=>"111111101",
        175=>"000000101",
        176=>"000000100",
        177=>"110011001",
        178=>"101111111",
        179=>"000100000",
        180=>"001001111",
        181=>"000110000",
        182=>"000000111",
        183=>"111110111",
        184=>"111000000",
        185=>"111110001",
        186=>"010100101",
        187=>"110010011",
        188=>"111011000",
        189=>"111111011",
        190=>"111111101",
        191=>"111111111",
        192=>"110111001",
        193=>"101110000",
        194=>"000000000",
        195=>"111111110",
        196=>"111000000",
        197=>"000000100",
        198=>"000000111",
        199=>"111111111",
        200=>"101100111",
        201=>"000000001",
        202=>"011100101",
        203=>"111111000",
        204=>"010000111",
        205=>"010000100",
        206=>"010111111",
        207=>"000110111",
        208=>"001001100",
        209=>"000101011",
        210=>"000001111",
        211=>"000010111",
        212=>"000001011",
        213=>"110110000",
        214=>"111111000",
        215=>"000111111",
        216=>"011000100",
        217=>"111001001",
        218=>"100001101",
        219=>"110000100",
        220=>"000000001",
        221=>"111011000",
        222=>"110110100",
        223=>"111110000",
        224=>"010000000",
        225=>"000000000",
        226=>"111110000",
        227=>"111110000",
        228=>"000000001",
        229=>"100001110",
        230=>"001001100",
        231=>"000000000",
        232=>"001101101",
        233=>"110111111",
        234=>"000100001",
        235=>"111111000",
        236=>"000000011",
        237=>"000000010",
        238=>"111111011",
        239=>"110110101",
        240=>"111100000",
        241=>"010000100",
        242=>"000001111",
        243=>"000000111",
        244=>"110010000",
        245=>"000001111",
        246=>"111011101",
        247=>"111100101",
        248=>"000010000",
        249=>"001000000",
        250=>"101001001",
        251=>"000010111",
        252=>"001001101",
        253=>"000000000",
        254=>"101100100",
        255=>"111001110",
        256=>"111110000",
        257=>"111000111",
        258=>"111000000",
        259=>"100100110",
        260=>"011011100",
        261=>"000101111",
        262=>"111111000",
        263=>"001101111",
        264=>"011010100",
        265=>"011011000",
        266=>"011000000",
        267=>"111001000",
        268=>"000111111",
        269=>"110110000",
        270=>"100101111",
        271=>"110000001",
        272=>"001011110",
        273=>"110010000",
        274=>"101011111",
        275=>"110101001",
        276=>"010110110",
        277=>"000011000",
        278=>"000100101",
        279=>"101100000",
        280=>"001010111",
        281=>"100000000",
        282=>"000001110",
        283=>"000000100",
        284=>"110111111",
        285=>"000100100",
        286=>"100000110",
        287=>"000011111",
        288=>"000001111",
        289=>"101110011",
        290=>"000001101",
        291=>"101000000",
        292=>"101100101",
        293=>"111111111",
        294=>"001111111",
        295=>"000101111",
        296=>"111001001",
        297=>"011001001",
        298=>"000110110",
        299=>"100000110",
        300=>"011000000",
        301=>"111111100",
        302=>"000111101",
        303=>"111010101",
        304=>"111111101",
        305=>"000011011",
        306=>"011011110",
        307=>"111111001",
        308=>"000000110",
        309=>"111111110",
        310=>"111100000",
        311=>"010000000",
        312=>"111000000",
        313=>"111000101",
        314=>"110110100",
        315=>"000100111",
        316=>"000001000",
        317=>"001001011",
        318=>"000000000",
        319=>"110011111",
        320=>"111111110",
        321=>"000011110",
        322=>"111000010",
        323=>"000000001",
        324=>"000000010",
        325=>"100000001",
        326=>"000111000",
        327=>"010000000",
        328=>"100110111",
        329=>"000110111",
        330=>"111000010",
        331=>"111000011",
        332=>"100111111",
        333=>"000000001",
        334=>"000001111",
        335=>"000111111",
        336=>"000000111",
        337=>"001001000",
        338=>"000001011",
        339=>"111111000",
        340=>"000001000",
        341=>"110110001",
        342=>"000000111",
        343=>"010011111",
        344=>"011000000",
        345=>"101001000",
        346=>"000001110",
        347=>"011110000",
        348=>"010100011",
        349=>"011011010",
        350=>"000010111",
        351=>"011100000",
        352=>"000001011",
        353=>"110111101",
        354=>"110000100",
        355=>"110000000",
        356=>"000001111",
        357=>"000111110",
        358=>"000010000",
        359=>"110000000",
        360=>"000101111",
        361=>"000000100",
        362=>"000001110",
        363=>"000000001",
        364=>"111010000",
        365=>"010110110",
        366=>"011111111",
        367=>"111111111",
        368=>"111111000",
        369=>"000000010",
        370=>"001111110",
        371=>"000100000",
        372=>"001001001",
        373=>"000100110",
        374=>"000000111",
        375=>"100001000",
        376=>"111000101",
        377=>"111100100",
        378=>"000100111",
        379=>"111110000",
        380=>"000111111",
        381=>"000000000",
        382=>"111011111",
        383=>"000100100",
        384=>"000111111",
        385=>"010111101",
        386=>"000111111",
        387=>"111110011",
        388=>"101100110",
        389=>"111000000",
        390=>"101101111",
        391=>"000100111",
        392=>"001111110",
        393=>"100011001",
        394=>"111101110",
        395=>"000100000",
        396=>"000101110",
        397=>"111000000",
        398=>"011001000",
        399=>"000000111",
        400=>"001001011",
        401=>"001001111",
        402=>"111010111",
        403=>"000011111",
        404=>"011000000",
        405=>"000000011",
        406=>"000111111",
        407=>"110000000",
        408=>"100011110",
        409=>"100101100",
        410=>"100111100",
        411=>"100110000",
        412=>"110000000",
        413=>"111000000",
        414=>"001000000",
        415=>"010001000",
        416=>"000000111",
        417=>"111001000",
        418=>"001111001",
        419=>"100000000",
        420=>"111111000",
        421=>"010100010",
        422=>"100110011",
        423=>"000111111",
        424=>"000100101",
        425=>"000000000",
        426=>"000010100",
        427=>"011100001",
        428=>"110000100",
        429=>"100101101",
        430=>"111000010",
        431=>"000111111",
        432=>"010000000",
        433=>"000111110",
        434=>"111011100",
        435=>"000010000",
        436=>"111000000",
        437=>"101000000",
        438=>"011000100",
        439=>"000101101",
        440=>"000101110",
        441=>"111111000",
        442=>"100011010",
        443=>"001111111",
        444=>"000010110",
        445=>"000100000",
        446=>"001100000",
        447=>"111000000",
        448=>"011000010",
        449=>"000101110",
        450=>"110010001",
        451=>"000000000",
        452=>"000000001",
        453=>"100110011",
        454=>"111100110",
        455=>"111011000",
        456=>"100110011",
        457=>"111000000",
        458=>"010011000",
        459=>"000101000",
        460=>"000000000",
        461=>"011001101",
        462=>"111010000",
        463=>"000111010",
        464=>"000011100",
        465=>"000111111",
        466=>"111000000",
        467=>"111011001",
        468=>"101011011",
        469=>"000101111",
        470=>"101000110",
        471=>"111000000",
        472=>"000100100",
        473=>"111101111",
        474=>"110110011",
        475=>"101100000",
        476=>"100101100",
        477=>"000000111",
        478=>"000111111",
        479=>"111000001",
        480=>"000011010",
        481=>"100110110",
        482=>"000111111",
        483=>"000010010",
        484=>"000000000",
        485=>"000111111",
        486=>"000111111",
        487=>"010000000",
        488=>"000111111",
        489=>"100111000",
        490=>"101101111",
        491=>"000000000",
        492=>"111001000",
        493=>"001001001",
        494=>"111000000",
        495=>"111100001",
        496=>"100100100",
        497=>"010010000",
        498=>"000111010",
        499=>"111000000",
        500=>"101001110",
        501=>"000000011",
        502=>"000000001",
        503=>"111110000",
        504=>"010110110",
        505=>"010000000",
        506=>"000111111",
        507=>"000000000",
        508=>"001011110",
        509=>"000101000",
        510=>"111111010",
        511=>"111010000",
        512=>"100010111",
        513=>"101000111",
        514=>"111100101",
        515=>"000000111",
        516=>"110110010",
        517=>"111011111",
        518=>"111111111",
        519=>"111111000",
        520=>"110010100",
        521=>"010000000",
        522=>"000000000",
        523=>"010000001",
        524=>"111101101",
        525=>"100100110",
        526=>"000011000",
        527=>"001001100",
        528=>"000000001",
        529=>"000000100",
        530=>"100110010",
        531=>"011001010",
        532=>"000001111",
        533=>"000010000",
        534=>"010011000",
        535=>"000010000",
        536=>"001011011",
        537=>"000011110",
        538=>"000111010",
        539=>"101011011",
        540=>"011101111",
        541=>"000110000",
        542=>"001110010",
        543=>"000000000",
        544=>"000101111",
        545=>"000100001",
        546=>"100110011",
        547=>"111000000",
        548=>"010000000",
        549=>"000000000",
        550=>"111010000",
        551=>"110000100",
        552=>"100111111",
        553=>"000000001",
        554=>"111110011",
        555=>"000001111",
        556=>"110110110",
        557=>"011000000",
        558=>"000111111",
        559=>"111111000",
        560=>"000101111",
        561=>"110000000",
        562=>"110110111",
        563=>"010011000",
        564=>"000011000",
        565=>"000000000",
        566=>"000000111",
        567=>"110000000",
        568=>"110000000",
        569=>"000100101",
        570=>"011000000",
        571=>"010000111",
        572=>"010111111",
        573=>"111111010",
        574=>"110110110",
        575=>"000000110",
        576=>"000001011",
        577=>"100000000",
        578=>"011000000",
        579=>"001010111",
        580=>"011111111",
        581=>"110100100",
        582=>"010010010",
        583=>"000111111",
        584=>"000000010",
        585=>"100100111",
        586=>"010111111",
        587=>"000010000",
        588=>"000010100",
        589=>"000001000",
        590=>"111111100",
        591=>"111000001",
        592=>"000001101",
        593=>"111011000",
        594=>"100101110",
        595=>"001000000",
        596=>"010011001",
        597=>"000100110",
        598=>"111111100",
        599=>"111000101",
        600=>"001001000",
        601=>"110000010",
        602=>"001111010",
        603=>"111100000",
        604=>"100100111",
        605=>"000100000",
        606=>"110110000",
        607=>"110111111",
        608=>"011100011",
        609=>"000000001",
        610=>"101000111",
        611=>"111111000",
        612=>"110011000",
        613=>"010011001",
        614=>"111011011",
        615=>"001111111",
        616=>"011000100",
        617=>"111111101",
        618=>"000001010",
        619=>"000111111",
        620=>"011000000",
        621=>"110111111",
        622=>"100100110",
        623=>"011110010",
        624=>"000000000",
        625=>"111011000",
        626=>"001100011",
        627=>"101100101",
        628=>"000000111",
        629=>"111011000",
        630=>"101111111",
        631=>"011011010",
        632=>"000111010",
        633=>"000001010",
        634=>"010010001",
        635=>"000010000",
        636=>"110010010",
        637=>"010000110",
        638=>"111111111",
        639=>"010011111",
        640=>"111011000",
        641=>"011010011",
        642=>"101100111",
        643=>"000000000",
        644=>"001111111",
        645=>"010011111",
        646=>"101001000",
        647=>"100000100",
        648=>"011111101",
        649=>"010111110",
        650=>"010100101",
        651=>"011101100",
        652=>"101001000",
        653=>"111111110",
        654=>"001011011",
        655=>"100100100",
        656=>"111001100",
        657=>"111111111",
        658=>"100100100",
        659=>"110000101",
        660=>"111000000",
        661=>"010000000",
        662=>"000000000",
        663=>"000010111",
        664=>"000001000",
        665=>"111101001",
        666=>"100100110",
        667=>"000110111",
        668=>"010111010",
        669=>"000001011",
        670=>"111100111",
        671=>"100001010",
        672=>"000000000",
        673=>"001111011",
        674=>"000001100",
        675=>"010000101",
        676=>"000111111",
        677=>"111000000",
        678=>"111101101",
        679=>"100100000",
        680=>"000000000",
        681=>"110110000",
        682=>"100100111",
        683=>"111110110",
        684=>"011011111",
        685=>"000010010",
        686=>"111011001",
        687=>"111101111",
        688=>"000111000",
        689=>"101000100",
        690=>"010101010",
        691=>"100100111",
        692=>"000110110",
        693=>"010111010",
        694=>"001111000",
        695=>"000011010",
        696=>"000100100",
        697=>"010100101",
        698=>"110101101",
        699=>"010011010",
        700=>"111100000",
        701=>"111101101",
        702=>"000001101",
        703=>"011111100",
        704=>"111000000",
        705=>"111100101",
        706=>"000010010",
        707=>"000010010",
        708=>"011101111",
        709=>"111100000",
        710=>"000010000",
        711=>"111110000",
        712=>"111100101",
        713=>"010111011",
        714=>"011011000",
        715=>"111000000",
        716=>"000000010",
        717=>"000000000",
        718=>"000000001",
        719=>"000000101",
        720=>"000000000",
        721=>"000100101",
        722=>"000000000",
        723=>"001000011",
        724=>"011001001",
        725=>"101010000",
        726=>"000111011",
        727=>"000111111",
        728=>"001011011",
        729=>"111111111",
        730=>"111110101",
        731=>"100000100",
        732=>"000001001",
        733=>"011001011",
        734=>"100000001",
        735=>"000000000",
        736=>"010011011",
        737=>"101011011",
        738=>"111101101",
        739=>"000011011",
        740=>"000000000",
        741=>"101100110",
        742=>"111100101",
        743=>"111011001",
        744=>"110111111",
        745=>"010111100",
        746=>"101110000",
        747=>"111011010",
        748=>"111111101",
        749=>"100000000",
        750=>"101100000",
        751=>"100110110",
        752=>"000000000",
        753=>"111001101",
        754=>"000000000",
        755=>"000110110",
        756=>"111101111",
        757=>"000100000",
        758=>"100000000",
        759=>"110000111",
        760=>"000100111",
        761=>"000000001",
        762=>"000100000",
        763=>"111000000",
        764=>"011001110",
        765=>"110111100",
        766=>"000000100",
        767=>"100111011",
        768=>"011001111",
        769=>"111100100",
        770=>"011011011",
        771=>"001001000",
        772=>"000001000",
        773=>"011011011",
        774=>"000001011",
        775=>"110110100",
        776=>"101111101",
        777=>"000001000",
        778=>"110010101",
        779=>"011111100",
        780=>"000011111",
        781=>"100101110",
        782=>"000000000",
        783=>"100100100",
        784=>"000011011",
        785=>"110110110",
        786=>"100001101",
        787=>"110100000",
        788=>"000000001",
        789=>"001110101",
        790=>"001000000",
        791=>"110110010",
        792=>"000000110",
        793=>"001001010",
        794=>"100001101",
        795=>"100111111",
        796=>"010111111",
        797=>"000000000",
        798=>"111011101",
        799=>"110110100",
        800=>"000001101",
        801=>"100100100",
        802=>"000111111",
        803=>"000000000",
        804=>"100001010",
        805=>"110100110",
        806=>"010111111",
        807=>"001001011",
        808=>"100100100",
        809=>"110000010",
        810=>"000000000",
        811=>"000001001",
        812=>"110111001",
        813=>"110100110",
        814=>"001111101",
        815=>"111111101",
        816=>"100111111",
        817=>"001001110",
        818=>"001011010",
        819=>"000001111",
        820=>"100111111",
        821=>"000000001",
        822=>"010110000",
        823=>"001001011",
        824=>"110111111",
        825=>"010011000",
        826=>"001011111",
        827=>"001100000",
        828=>"110100100",
        829=>"000000000",
        830=>"100100000",
        831=>"101111011",
        832=>"111111111",
        833=>"010000111",
        834=>"101000000",
        835=>"010010001",
        836=>"001011011",
        837=>"000101011",
        838=>"100100101",
        839=>"110111110",
        840=>"011000000",
        841=>"000000001",
        842=>"100000001",
        843=>"001100110",
        844=>"101111101",
        845=>"100000100",
        846=>"100100101",
        847=>"001011001",
        848=>"010100110",
        849=>"011000011",
        850=>"110000101",
        851=>"011011001",
        852=>"001011111",
        853=>"011110000",
        854=>"000000101",
        855=>"011000000",
        856=>"001111001",
        857=>"011101000",
        858=>"111111011",
        859=>"001001000",
        860=>"000001101",
        861=>"011111111",
        862=>"111101101",
        863=>"011000010",
        864=>"000000000",
        865=>"111110010",
        866=>"111110011",
        867=>"111011010",
        868=>"110110100",
        869=>"000001111",
        870=>"000001111",
        871=>"011110100",
        872=>"000001011",
        873=>"101000100",
        874=>"100000001",
        875=>"111111111",
        876=>"001001110",
        877=>"110100100",
        878=>"110011001",
        879=>"001001001",
        880=>"011011011",
        881=>"101011011",
        882=>"100001001",
        883=>"001011011",
        884=>"111100111",
        885=>"010011010",
        886=>"100110100",
        887=>"000001101",
        888=>"000001111",
        889=>"100110110",
        890=>"110110000",
        891=>"110100100",
        892=>"100000110",
        893=>"110010000",
        894=>"110000000",
        895=>"110000000",
        896=>"111111111",
        897=>"001100100",
        898=>"001001001",
        899=>"110011100",
        900=>"111000000",
        901=>"010010100",
        902=>"111101001",
        903=>"100100110",
        904=>"111011111",
        905=>"000000000",
        906=>"000110100",
        907=>"111110000",
        908=>"011011011",
        909=>"000111100",
        910=>"110111111",
        911=>"100111111",
        912=>"000100101",
        913=>"110100000",
        914=>"111101000",
        915=>"011011011",
        916=>"100110110",
        917=>"001001000",
        918=>"011011111",
        919=>"110110010",
        920=>"001001001",
        921=>"100110000",
        922=>"100010001",
        923=>"111111111",
        924=>"101111101",
        925=>"111011001",
        926=>"111101000",
        927=>"110100100",
        928=>"001100100",
        929=>"111110000",
        930=>"001001010",
        931=>"100010000",
        932=>"110110000",
        933=>"000001001",
        934=>"101100110",
        935=>"011011000",
        936=>"010000000",
        937=>"100110010",
        938=>"101011001",
        939=>"111011001",
        940=>"110100100",
        941=>"101100100",
        942=>"100100100",
        943=>"001011011",
        944=>"100110001",
        945=>"001001111",
        946=>"111000000",
        947=>"111111011",
        948=>"011001001",
        949=>"000000001",
        950=>"100110110",
        951=>"001011011",
        952=>"111111111",
        953=>"100110100",
        954=>"111111111",
        955=>"111001001",
        956=>"011001001",
        957=>"110100000",
        958=>"000000000",
        959=>"100110010",
        960=>"010111111",
        961=>"110100000",
        962=>"100100110",
        963=>"010010100",
        964=>"100011111",
        965=>"100000101",
        966=>"100101000",
        967=>"100110110",
        968=>"110110000",
        969=>"001011001",
        970=>"100100100",
        971=>"000001001",
        972=>"100100101",
        973=>"000010001",
        974=>"100110100",
        975=>"001011011",
        976=>"100100100",
        977=>"011011011",
        978=>"100000101",
        979=>"100001111",
        980=>"111110110",
        981=>"000001011",
        982=>"111111111",
        983=>"001001100",
        984=>"010111101",
        985=>"100000000",
        986=>"111010001",
        987=>"111111111",
        988=>"111011001",
        989=>"111101110",
        990=>"111011001",
        991=>"100001011",
        992=>"000000000",
        993=>"100000000",
        994=>"001010001",
        995=>"001111000",
        996=>"100000110",
        997=>"110011000",
        998=>"011011001",
        999=>"110110101",
        1000=>"100100110",
        1001=>"001000001",
        1002=>"110111001",
        1003=>"100100100",
        1004=>"011001001",
        1005=>"000000110",
        1006=>"100000100",
        1007=>"000000000",
        1008=>"111011011",
        1009=>"000000000",
        1010=>"111001000",
        1011=>"011011011",
        1012=>"000001011",
        1013=>"111110101",
        1014=>"100100100",
        1015=>"110111111",
        1016=>"000100100",
        1017=>"100100100",
        1018=>"111100100",
        1019=>"100100110",
        1020=>"110000000",
        1021=>"010110000",
        1022=>"000000010",
        1023=>"110011000",
        1024=>"000010011",
        1025=>"100100100",
        1026=>"110110100",
        1027=>"000001110",
        1028=>"111111111",
        1029=>"110110010",
        1030=>"000011011",
        1031=>"100101000",
        1032=>"101111101",
        1033=>"010001111",
        1034=>"011111111",
        1035=>"001001001",
        1036=>"001100100",
        1037=>"100111000",
        1038=>"111111001",
        1039=>"110110100",
        1040=>"111011011",
        1041=>"001011111",
        1042=>"000000000",
        1043=>"000000000",
        1044=>"100100000",
        1045=>"001001011",
        1046=>"000000010",
        1047=>"101001001",
        1048=>"101111111",
        1049=>"001101101",
        1050=>"001011101",
        1051=>"010011010",
        1052=>"000000101",
        1053=>"111111111",
        1054=>"000000000",
        1055=>"010001011",
        1056=>"101011111",
        1057=>"011011010",
        1058=>"101011001",
        1059=>"001001001",
        1060=>"010001011",
        1061=>"001001000",
        1062=>"000001001",
        1063=>"110110100",
        1064=>"001001011",
        1065=>"011011011",
        1066=>"111010111",
        1067=>"010010110",
        1068=>"101001100",
        1069=>"001001001",
        1070=>"001001011",
        1071=>"011011111",
        1072=>"000110110",
        1073=>"110100101",
        1074=>"001000100",
        1075=>"101001001",
        1076=>"000000000",
        1077=>"011001001",
        1078=>"110110100",
        1079=>"100100010",
        1080=>"011100011",
        1081=>"011011011",
        1082=>"101100110",
        1083=>"110111011",
        1084=>"001001001",
        1085=>"011000001",
        1086=>"001011101",
        1087=>"111100110",
        1088=>"010011110",
        1089=>"010000111",
        1090=>"001111000",
        1091=>"111001011",
        1092=>"010011001",
        1093=>"110111101",
        1094=>"100110100",
        1095=>"001001000",
        1096=>"001001110",
        1097=>"100100100",
        1098=>"000000000",
        1099=>"001001001",
        1100=>"010100100",
        1101=>"100000000",
        1102=>"000011001",
        1103=>"100100100",
        1104=>"110110101",
        1105=>"110100100",
        1106=>"001001001",
        1107=>"110110111",
        1108=>"001001001",
        1109=>"110100000",
        1110=>"001011011",
        1111=>"100110011",
        1112=>"001001001",
        1113=>"010010001",
        1114=>"001010100",
        1115=>"101001000",
        1116=>"000010000",
        1117=>"100100100",
        1118=>"011011011",
        1119=>"001001011",
        1120=>"011000001",
        1121=>"110110010",
        1122=>"100100100",
        1123=>"000100000",
        1124=>"011001001",
        1125=>"001001111",
        1126=>"100100000",
        1127=>"000111010",
        1128=>"110110011",
        1129=>"100100000",
        1130=>"101101010",
        1131=>"111100111",
        1132=>"111100110",
        1133=>"100000000",
        1134=>"100000001",
        1135=>"000000110",
        1136=>"011010001",
        1137=>"000100000",
        1138=>"010110110",
        1139=>"100100100",
        1140=>"001011011",
        1141=>"001001001",
        1142=>"011011011",
        1143=>"001011111",
        1144=>"001001010",
        1145=>"110001011",
        1146=>"111111001",
        1147=>"100001100",
        1148=>"000000000",
        1149=>"010000001",
        1150=>"001001101",
        1151=>"111011111",
        1152=>"111111111",
        1153=>"000111010",
        1154=>"111111100",
        1155=>"011011010",
        1156=>"001010111",
        1157=>"010000101",
        1158=>"111111111",
        1159=>"111100100",
        1160=>"001000000",
        1161=>"100000000",
        1162=>"111001000",
        1163=>"110100001",
        1164=>"010000100",
        1165=>"111110110",
        1166=>"111100111",
        1167=>"110000001",
        1168=>"111100100",
        1169=>"000110010",
        1170=>"111111001",
        1171=>"100001011",
        1172=>"111010010",
        1173=>"100000100",
        1174=>"000000100",
        1175=>"000000111",
        1176=>"101101100",
        1177=>"001000000",
        1178=>"001101101",
        1179=>"001110011",
        1180=>"101010000",
        1181=>"110110100",
        1182=>"101111101",
        1183=>"000000000",
        1184=>"110100000",
        1185=>"000010100",
        1186=>"000000000",
        1187=>"000000000",
        1188=>"000000000",
        1189=>"110110010",
        1190=>"010000010",
        1191=>"000000110",
        1192=>"001001000",
        1193=>"111101000",
        1194=>"101111101",
        1195=>"100101101",
        1196=>"111100000",
        1197=>"000000000",
        1198=>"000010010",
        1199=>"111111111",
        1200=>"110111010",
        1201=>"110010010",
        1202=>"111011000",
        1203=>"001000000",
        1204=>"101001100",
        1205=>"000000011",
        1206=>"000111111",
        1207=>"111000100",
        1208=>"011111111",
        1209=>"011101101",
        1210=>"011000101",
        1211=>"001000010",
        1212=>"100000000",
        1213=>"000010110",
        1214=>"100000100",
        1215=>"011010011",
        1216=>"000000000",
        1217=>"010110010",
        1218=>"110110000",
        1219=>"101000000",
        1220=>"000000000",
        1221=>"111111111",
        1222=>"111001000",
        1223=>"111111111",
        1224=>"110000001",
        1225=>"101100010",
        1226=>"011111111",
        1227=>"100111111",
        1228=>"000000000",
        1229=>"101100111",
        1230=>"000000000",
        1231=>"000000000",
        1232=>"000000000",
        1233=>"000011010",
        1234=>"110100100",
        1235=>"110111111",
        1236=>"111111111",
        1237=>"101000000",
        1238=>"111111111",
        1239=>"110000001",
        1240=>"111111111",
        1241=>"111010100",
        1242=>"000001001",
        1243=>"010000000",
        1244=>"001101001",
        1245=>"011000100",
        1246=>"100101100",
        1247=>"101111100",
        1248=>"110100100",
        1249=>"111001001",
        1250=>"000000010",
        1251=>"111111111",
        1252=>"111010000",
        1253=>"001011101",
        1254=>"000010010",
        1255=>"111101111",
        1256=>"110110000",
        1257=>"100100000",
        1258=>"111100110",
        1259=>"000000111",
        1260=>"101111010",
        1261=>"000000000",
        1262=>"101110100",
        1263=>"100001111",
        1264=>"000000000",
        1265=>"111101100",
        1266=>"000000010",
        1267=>"110101111",
        1268=>"111000000",
        1269=>"000000001",
        1270=>"000011111",
        1271=>"110110100",
        1272=>"111111100",
        1273=>"111011011",
        1274=>"011011010",
        1275=>"000000000",
        1276=>"000110100",
        1277=>"110110011",
        1278=>"000001001",
        1279=>"100011011",
        1280=>"010000010",
        1281=>"010110110",
        1282=>"011110111",
        1283=>"101001001",
        1284=>"111111000",
        1285=>"010110000",
        1286=>"111011110",
        1287=>"001000000",
        1288=>"010011001",
        1289=>"001000000",
        1290=>"010111111",
        1291=>"000000101",
        1292=>"000000000",
        1293=>"110110110",
        1294=>"111100110",
        1295=>"100000111",
        1296=>"111111111",
        1297=>"110111101",
        1298=>"101110111",
        1299=>"111000010",
        1300=>"000110011",
        1301=>"100001001",
        1302=>"011000001",
        1303=>"000000100",
        1304=>"111101111",
        1305=>"001011111",
        1306=>"001001000",
        1307=>"000000100",
        1308=>"110111110",
        1309=>"000111111",
        1310=>"010011101",
        1311=>"111111111",
        1312=>"110110111",
        1313=>"100011000",
        1314=>"011111101",
        1315=>"101001111",
        1316=>"011000000",
        1317=>"000111110",
        1318=>"110110101",
        1319=>"001000001",
        1320=>"111011011",
        1321=>"111111000",
        1322=>"111001001",
        1323=>"011001111",
        1324=>"111010010",
        1325=>"010000100",
        1326=>"000111111",
        1327=>"111111111",
        1328=>"000001000",
        1329=>"111010111",
        1330=>"010001000",
        1331=>"100000000",
        1332=>"000111000",
        1333=>"000000000",
        1334=>"000000000",
        1335=>"110111110",
        1336=>"110000000",
        1337=>"110111111",
        1338=>"000000000",
        1339=>"000110000",
        1340=>"111000001",
        1341=>"001000100",
        1342=>"000000001",
        1343=>"110110110",
        1344=>"010000000",
        1345=>"010010110",
        1346=>"010110110",
        1347=>"110000000",
        1348=>"001001011",
        1349=>"000010010",
        1350=>"110111110",
        1351=>"111011111",
        1352=>"111111111",
        1353=>"010111000",
        1354=>"000000000",
        1355=>"111000111",
        1356=>"001001000",
        1357=>"010011010",
        1358=>"001101111",
        1359=>"111011101",
        1360=>"110110010",
        1361=>"101001101",
        1362=>"000000000",
        1363=>"010000010",
        1364=>"010110111",
        1365=>"000000000",
        1366=>"101001001",
        1367=>"111111101",
        1368=>"011100000",
        1369=>"110100101",
        1370=>"000000000",
        1371=>"000000000",
        1372=>"111110111",
        1373=>"111111111",
        1374=>"101001101",
        1375=>"110110100",
        1376=>"001101001",
        1377=>"111001101",
        1378=>"111111111",
        1379=>"110110110",
        1380=>"111111111",
        1381=>"010010001",
        1382=>"001000101",
        1383=>"111011110",
        1384=>"100111010",
        1385=>"101101100",
        1386=>"101011110",
        1387=>"000010000",
        1388=>"001000000",
        1389=>"011001001",
        1390=>"110111110",
        1391=>"001101100",
        1392=>"001000001",
        1393=>"001101011",
        1394=>"001000001",
        1395=>"000111000",
        1396=>"111000000",
        1397=>"101000001",
        1398=>"111110000",
        1399=>"001001000",
        1400=>"111000110",
        1401=>"100000111",
        1402=>"100111110",
        1403=>"001000001",
        1404=>"001011001",
        1405=>"000000111",
        1406=>"011111000",
        1407=>"110111110",
        1408=>"100110010",
        1409=>"111101001",
        1410=>"111000001",
        1411=>"101101111",
        1412=>"000010100",
        1413=>"010111001",
        1414=>"000000000",
        1415=>"110001001",
        1416=>"011011101",
        1417=>"010100110",
        1418=>"110100101",
        1419=>"010010001",
        1420=>"111001000",
        1421=>"111111111",
        1422=>"000100000",
        1423=>"111100000",
        1424=>"101000000",
        1425=>"111101001",
        1426=>"000001101",
        1427=>"100100011",
        1428=>"000001111",
        1429=>"000001000",
        1430=>"011001000",
        1431=>"101111011",
        1432=>"001100110",
        1433=>"100100110",
        1434=>"001000100",
        1435=>"000000000",
        1436=>"001001101",
        1437=>"000000101",
        1438=>"011011111",
        1439=>"001010010",
        1440=>"000000100",
        1441=>"000000101",
        1442=>"000011011",
        1443=>"010110111",
        1444=>"000010111",
        1445=>"111101110",
        1446=>"110000000",
        1447=>"000001111",
        1448=>"010010011",
        1449=>"111110110",
        1450=>"111000000",
        1451=>"000000111",
        1452=>"010001011",
        1453=>"000010011",
        1454=>"010010100",
        1455=>"111111101",
        1456=>"111000101",
        1457=>"111001000",
        1458=>"011001101",
        1459=>"001010010",
        1460=>"000000101",
        1461=>"010111101",
        1462=>"111010001",
        1463=>"000010110",
        1464=>"101001001",
        1465=>"000011010",
        1466=>"110010111",
        1467=>"111001100",
        1468=>"111111000",
        1469=>"000010010",
        1470=>"000000000",
        1471=>"110111011",
        1472=>"111111011",
        1473=>"110000000",
        1474=>"111111111",
        1475=>"011011000",
        1476=>"000110101",
        1477=>"000010110",
        1478=>"001100100",
        1479=>"101000001",
        1480=>"101000000",
        1481=>"000110111",
        1482=>"110011011",
        1483=>"111101000",
        1484=>"111001000",
        1485=>"010111111",
        1486=>"000010010",
        1487=>"111001001",
        1488=>"001000011",
        1489=>"000000000",
        1490=>"000010111",
        1491=>"000000110",
        1492=>"000010011",
        1493=>"111001001",
        1494=>"110101000",
        1495=>"000111100",
        1496=>"000011111",
        1497=>"100110000",
        1498=>"100000010",
        1499=>"110001000",
        1500=>"000100101",
        1501=>"111011001",
        1502=>"111000001",
        1503=>"111111000",
        1504=>"000001101",
        1505=>"001000110",
        1506=>"111010000",
        1507=>"001000111",
        1508=>"110110000",
        1509=>"111001101",
        1510=>"010000000",
        1511=>"110100000",
        1512=>"111000001",
        1513=>"000101101",
        1514=>"000110111",
        1515=>"110111001",
        1516=>"011010001",
        1517=>"100110101",
        1518=>"000110110",
        1519=>"100011001",
        1520=>"101111000",
        1521=>"110110110",
        1522=>"111111000",
        1523=>"111001101",
        1524=>"000100000",
        1525=>"111101000",
        1526=>"000000000",
        1527=>"010100100",
        1528=>"111011000",
        1529=>"111010000",
        1530=>"111001000",
        1531=>"111101101",
        1532=>"011101100",
        1533=>"101111101",
        1534=>"010110111",
        1535=>"000010111",
        1536=>"101110111",
        1537=>"010111111",
        1538=>"000000000",
        1539=>"110101000",
        1540=>"001000000",
        1541=>"111111111",
        1542=>"010100111",
        1543=>"000001000",
        1544=>"111111101",
        1545=>"000111100",
        1546=>"100101110",
        1547=>"011111000",
        1548=>"110001001",
        1549=>"010111110",
        1550=>"100000100",
        1551=>"001111111",
        1552=>"111100100",
        1553=>"111010000",
        1554=>"001000000",
        1555=>"110010110",
        1556=>"010111000",
        1557=>"101111111",
        1558=>"000000001",
        1559=>"000000000",
        1560=>"000001001",
        1561=>"111111100",
        1562=>"000101100",
        1563=>"111111111",
        1564=>"111111110",
        1565=>"100100000",
        1566=>"101100111",
        1567=>"100001111",
        1568=>"011100000",
        1569=>"000000000",
        1570=>"000011000",
        1571=>"100000000",
        1572=>"011011111",
        1573=>"111111111",
        1574=>"011000000",
        1575=>"110000000",
        1576=>"000000000",
        1577=>"000000000",
        1578=>"111111111",
        1579=>"110100101",
        1580=>"101000100",
        1581=>"001000000",
        1582=>"001000110",
        1583=>"000000000",
        1584=>"111111111",
        1585=>"100101111",
        1586=>"011110110",
        1587=>"101001011",
        1588=>"000000000",
        1589=>"011001001",
        1590=>"111111110",
        1591=>"010011000",
        1592=>"111111111",
        1593=>"111111010",
        1594=>"111111001",
        1595=>"110111011",
        1596=>"000000000",
        1597=>"011111101",
        1598=>"110111011",
        1599=>"100101110",
        1600=>"111111101",
        1601=>"001010000",
        1602=>"000000001",
        1603=>"000100001",
        1604=>"111111111",
        1605=>"000010000",
        1606=>"000111010",
        1607=>"000000000",
        1608=>"001001001",
        1609=>"000000000",
        1610=>"011000100",
        1611=>"000000000",
        1612=>"001000100",
        1613=>"111111111",
        1614=>"111111111",
        1615=>"010110010",
        1616=>"011000000",
        1617=>"000000000",
        1618=>"000000100",
        1619=>"111111111",
        1620=>"000001000",
        1621=>"010100010",
        1622=>"111111111",
        1623=>"111111111",
        1624=>"000000100",
        1625=>"111101110",
        1626=>"001011001",
        1627=>"111111111",
        1628=>"100101101",
        1629=>"001001101",
        1630=>"001001001",
        1631=>"000000000",
        1632=>"111111111",
        1633=>"101101111",
        1634=>"111111111",
        1635=>"000001001",
        1636=>"000011110",
        1637=>"000000100",
        1638=>"100000101",
        1639=>"101100111",
        1640=>"011011000",
        1641=>"000100000",
        1642=>"100000001",
        1643=>"000000111",
        1644=>"111111101",
        1645=>"000110000",
        1646=>"001001001",
        1647=>"001001101",
        1648=>"000000000",
        1649=>"000000000",
        1650=>"010000111",
        1651=>"000111110",
        1652=>"011111000",
        1653=>"010000000",
        1654=>"001110011",
        1655=>"100111011",
        1656=>"011000100",
        1657=>"000000001",
        1658=>"101101100",
        1659=>"001111111",
        1660=>"110110111",
        1661=>"111111111",
        1662=>"000000000",
        1663=>"000011001",
        1664=>"111111111",
        1665=>"000100111",
        1666=>"000000000",
        1667=>"101101100",
        1668=>"001011011",
        1669=>"011101111",
        1670=>"000010011",
        1671=>"000100100",
        1672=>"111100101",
        1673=>"111100100",
        1674=>"000000010",
        1675=>"111001000",
        1676=>"101011000",
        1677=>"110111010",
        1678=>"000111111",
        1679=>"000110110",
        1680=>"110100011",
        1681=>"111000000",
        1682=>"001100100",
        1683=>"101111111",
        1684=>"000111010",
        1685=>"010010000",
        1686=>"010000011",
        1687=>"000010101",
        1688=>"100000000",
        1689=>"001011000",
        1690=>"100110010",
        1691=>"101111111",
        1692=>"100111110",
        1693=>"000000000",
        1694=>"001000000",
        1695=>"011111011",
        1696=>"110100000",
        1697=>"010111111",
        1698=>"100110010",
        1699=>"000000000",
        1700=>"011111111",
        1701=>"000010010",
        1702=>"111101100",
        1703=>"111111010",
        1704=>"000010111",
        1705=>"110110100",
        1706=>"111100110",
        1707=>"001001101",
        1708=>"101110111",
        1709=>"000111111",
        1710=>"111111111",
        1711=>"110101101",
        1712=>"111111111",
        1713=>"110111111",
        1714=>"101110111",
        1715=>"011000000",
        1716=>"000000000",
        1717=>"000000000",
        1718=>"010000010",
        1719=>"111000000",
        1720=>"111000100",
        1721=>"000000000",
        1722=>"011010000",
        1723=>"111111010",
        1724=>"010111111",
        1725=>"000000000",
        1726=>"100111111",
        1727=>"111111001",
        1728=>"010011111",
        1729=>"000000000",
        1730=>"000000111",
        1731=>"000111111",
        1732=>"110100011",
        1733=>"011011001",
        1734=>"000011010",
        1735=>"000010111",
        1736=>"001001100",
        1737=>"000000000",
        1738=>"000000111",
        1739=>"000111111",
        1740=>"111011111",
        1741=>"111111111",
        1742=>"000010000",
        1743=>"000000001",
        1744=>"010010010",
        1745=>"111100100",
        1746=>"000110000",
        1747=>"111100111",
        1748=>"010110100",
        1749=>"111000000",
        1750=>"000010001",
        1751=>"110111001",
        1752=>"110011011",
        1753=>"111001000",
        1754=>"000010101",
        1755=>"000000001",
        1756=>"111110100",
        1757=>"101011011",
        1758=>"000000000",
        1759=>"000000000",
        1760=>"011110111",
        1761=>"111111110",
        1762=>"010111011",
        1763=>"111111111",
        1764=>"010000000",
        1765=>"000011011",
        1766=>"011001001",
        1767=>"001000000",
        1768=>"011110000",
        1769=>"000000101",
        1770=>"010001001",
        1771=>"110000000",
        1772=>"001001111",
        1773=>"100001101",
        1774=>"111111111",
        1775=>"000001001",
        1776=>"000111010",
        1777=>"001000001",
        1778=>"100000000",
        1779=>"001000101",
        1780=>"000000001",
        1781=>"011000000",
        1782=>"000000000",
        1783=>"101001011",
        1784=>"111011000",
        1785=>"000010010",
        1786=>"110010011",
        1787=>"101101111",
        1788=>"100011001",
        1789=>"011011110",
        1790=>"000000000",
        1791=>"000000000",
        1792=>"000000000",
        1793=>"000000110",
        1794=>"000000000",
        1795=>"111111110",
        1796=>"000101110",
        1797=>"000000100",
        1798=>"010011011",
        1799=>"101101111",
        1800=>"111111000",
        1801=>"111110100",
        1802=>"100000000",
        1803=>"011001001",
        1804=>"001010000",
        1805=>"110110000",
        1806=>"001001101",
        1807=>"000011000",
        1808=>"011111010",
        1809=>"000101010",
        1810=>"100101111",
        1811=>"000100111",
        1812=>"010111000",
        1813=>"001000000",
        1814=>"100000111",
        1815=>"010111110",
        1816=>"011001111",
        1817=>"110100000",
        1818=>"101101111",
        1819=>"111111101",
        1820=>"111111111",
        1821=>"011000011",
        1822=>"100100110",
        1823=>"010111011",
        1824=>"000010000",
        1825=>"101110101",
        1826=>"011110110",
        1827=>"111000000",
        1828=>"001011010",
        1829=>"010001001",
        1830=>"001111110",
        1831=>"000000111",
        1832=>"000000000",
        1833=>"000010000",
        1834=>"000111111",
        1835=>"111100111",
        1836=>"000000111",
        1837=>"010011010",
        1838=>"000000111",
        1839=>"111111111",
        1840=>"011110110",
        1841=>"000000101",
        1842=>"001111111",
        1843=>"001001001",
        1844=>"011101111",
        1845=>"000000000",
        1846=>"000000001",
        1847=>"101101111",
        1848=>"100110000",
        1849=>"111101000",
        1850=>"101011011",
        1851=>"000010000",
        1852=>"000000111",
        1853=>"111001101",
        1854=>"001000110",
        1855=>"010100011",
        1856=>"110111111",
        1857=>"001101101",
        1858=>"011010111",
        1859=>"111010111",
        1860=>"011011000",
        1861=>"011011000",
        1862=>"000000000",
        1863=>"000000110",
        1864=>"001011001",
        1865=>"111000011",
        1866=>"111111110",
        1867=>"011111010",
        1868=>"000100000",
        1869=>"111011111",
        1870=>"111111000",
        1871=>"010010010",
        1872=>"000010111",
        1873=>"000000111",
        1874=>"101100101",
        1875=>"111000100",
        1876=>"010110010",
        1877=>"111000000",
        1878=>"000011011",
        1879=>"001001001",
        1880=>"001011111",
        1881=>"111100111",
        1882=>"001001001",
        1883=>"111111111",
        1884=>"110110111",
        1885=>"100001101",
        1886=>"101111111",
        1887=>"101000100",
        1888=>"111110000",
        1889=>"100100001",
        1890=>"000010000",
        1891=>"111111010",
        1892=>"000000000",
        1893=>"000000101",
        1894=>"000000110",
        1895=>"010000001",
        1896=>"110110110",
        1897=>"101001100",
        1898=>"110101101",
        1899=>"111111111",
        1900=>"010011000",
        1901=>"101001111",
        1902=>"110000000",
        1903=>"001101111",
        1904=>"100000000",
        1905=>"000000100",
        1906=>"000100111",
        1907=>"001000000",
        1908=>"000000000",
        1909=>"000000000",
        1910=>"000000000",
        1911=>"101111111",
        1912=>"111011111",
        1913=>"001001011",
        1914=>"000110111",
        1915=>"111111001",
        1916=>"000100110",
        1917=>"111110000",
        1918=>"000000000",
        1919=>"111111111",
        1920=>"010111100",
        1921=>"011111010",
        1922=>"110111110",
        1923=>"000000000",
        1924=>"000100100",
        1925=>"111111111",
        1926=>"111111111",
        1927=>"111111111",
        1928=>"100100000",
        1929=>"111110110",
        1930=>"000000000",
        1931=>"010000000",
        1932=>"100101100",
        1933=>"000000000",
        1934=>"001100101",
        1935=>"001011111",
        1936=>"110100111",
        1937=>"101011000",
        1938=>"000110110",
        1939=>"110001111",
        1940=>"111011011",
        1941=>"111011010",
        1942=>"101101111",
        1943=>"111011111",
        1944=>"100100000",
        1945=>"101000000",
        1946=>"110110110",
        1947=>"001111111",
        1948=>"111111111",
        1949=>"110010000",
        1950=>"000101110",
        1951=>"111011111",
        1952=>"000010011",
        1953=>"000100001",
        1954=>"000101100",
        1955=>"000000000",
        1956=>"011011111",
        1957=>"011011010",
        1958=>"111111111",
        1959=>"111010100",
        1960=>"000100100",
        1961=>"110010101",
        1962=>"000000100",
        1963=>"110101001",
        1964=>"101010111",
        1965=>"011011011",
        1966=>"001001111",
        1967=>"110111010",
        1968=>"010000000",
        1969=>"101100000",
        1970=>"110110111",
        1971=>"100111001",
        1972=>"100110000",
        1973=>"011111001",
        1974=>"111001001",
        1975=>"111011111",
        1976=>"011010000",
        1977=>"000010111",
        1978=>"001001000",
        1979=>"001001000",
        1980=>"111011111",
        1981=>"111111011",
        1982=>"111111111",
        1983=>"000011111",
        1984=>"111111010",
        1985=>"111011101",
        1986=>"000111011",
        1987=>"111111111",
        1988=>"100000110",
        1989=>"011101101",
        1990=>"000010000",
        1991=>"001011011",
        1992=>"101000111",
        1993=>"010000101",
        1994=>"000110111",
        1995=>"110111110",
        1996=>"000000010",
        1997=>"000000000",
        1998=>"001111111",
        1999=>"011011111",
        2000=>"100110011",
        2001=>"111111011",
        2002=>"000000000",
        2003=>"011111101",
        2004=>"111111111",
        2005=>"111111111",
        2006=>"011111111",
        2007=>"111111011",
        2008=>"000110100",
        2009=>"011000000",
        2010=>"000001000",
        2011=>"110110111",
        2012=>"110110000",
        2013=>"010001011",
        2014=>"001100000",
        2015=>"000000100",
        2016=>"110110111",
        2017=>"000100110",
        2018=>"101000000",
        2019=>"100110110",
        2020=>"111111101",
        2021=>"111011010",
        2022=>"111110111",
        2023=>"001101011",
        2024=>"011011001",
        2025=>"100111010",
        2026=>"100100100",
        2027=>"111011111",
        2028=>"010000101",
        2029=>"111010111",
        2030=>"010111011",
        2031=>"111111111",
        2032=>"000110011",
        2033=>"001011111",
        2034=>"111110000",
        2035=>"111001010",
        2036=>"000000001",
        2037=>"000011001",
        2038=>"001011000",
        2039=>"010000000",
        2040=>"001011011",
        2041=>"011000011",
        2042=>"111111111",
        2043=>"000000000",
        2044=>"110100100",
        2045=>"000000000",
        2046=>"111010011",
        2047=>"000001000",
        2048=>"111110010",
        2049=>"100100100",
        2050=>"011001001",
        2051=>"000111011",
        2052=>"000000100",
        2053=>"100110000",
        2054=>"000010010",
        2055=>"000101101",
        2056=>"000100000",
        2057=>"011110000",
        2058=>"111001011",
        2059=>"110100000",
        2060=>"100110110",
        2061=>"000110000",
        2062=>"101101100",
        2063=>"001001001",
        2064=>"100110110",
        2065=>"010001000",
        2066=>"101010001",
        2067=>"111011000",
        2068=>"001001001",
        2069=>"001001001",
        2070=>"010100110",
        2071=>"101101101",
        2072=>"110111101",
        2073=>"101111010",
        2074=>"010010010",
        2075=>"101110001",
        2076=>"110111000",
        2077=>"000000000",
        2078=>"100001011",
        2079=>"010011000",
        2080=>"010110110",
        2081=>"100100100",
        2082=>"010110000",
        2083=>"000001100",
        2084=>"000100011",
        2085=>"011001001",
        2086=>"100110100",
        2087=>"001011000",
        2088=>"100000000",
        2089=>"100001110",
        2090=>"100110110",
        2091=>"010111111",
        2092=>"110011011",
        2093=>"001001110",
        2094=>"100110111",
        2095=>"110100100",
        2096=>"100110110",
        2097=>"100100000",
        2098=>"010110110",
        2099=>"001011011",
        2100=>"110110110",
        2101=>"000010000",
        2102=>"010110110",
        2103=>"101001101",
        2104=>"110101100",
        2105=>"110000000",
        2106=>"000110110",
        2107=>"000000010",
        2108=>"111100000",
        2109=>"001001011",
        2110=>"111111011",
        2111=>"001001001",
        2112=>"000000000",
        2113=>"100100100",
        2114=>"100011011",
        2115=>"101001111",
        2116=>"100110010",
        2117=>"101100101",
        2118=>"001000001",
        2119=>"110100000",
        2120=>"000110110",
        2121=>"011000000",
        2122=>"001000100",
        2123=>"000000001",
        2124=>"110100000",
        2125=>"100110110",
        2126=>"000010101",
        2127=>"100100100",
        2128=>"100100100",
        2129=>"001001000",
        2130=>"001001001",
        2131=>"111110110",
        2132=>"001111001",
        2133=>"111001001",
        2134=>"000110100",
        2135=>"011000100",
        2136=>"111011001",
        2137=>"101110010",
        2138=>"100000101",
        2139=>"000100100",
        2140=>"000000000",
        2141=>"110101001",
        2142=>"110111011",
        2143=>"101100100",
        2144=>"101100011",
        2145=>"000000110",
        2146=>"011001001",
        2147=>"110100000",
        2148=>"110110000",
        2149=>"101100110",
        2150=>"111100100",
        2151=>"110000000",
        2152=>"100110100",
        2153=>"111000000",
        2154=>"011111111",
        2155=>"111100101",
        2156=>"001000001",
        2157=>"101001001",
        2158=>"111011011",
        2159=>"111110100",
        2160=>"011001001",
        2161=>"111000101",
        2162=>"100110110",
        2163=>"100100100",
        2164=>"011001000",
        2165=>"000100110",
        2166=>"111100100",
        2167=>"100110110",
        2168=>"110111011",
        2169=>"100100110",
        2170=>"100110100",
        2171=>"100110100",
        2172=>"110001100",
        2173=>"110111110",
        2174=>"111001101",
        2175=>"101011011",
        2176=>"110111111",
        2177=>"000000000",
        2178=>"001000011",
        2179=>"000000000",
        2180=>"100000100",
        2181=>"001100111",
        2182=>"011001011",
        2183=>"100101101",
        2184=>"110110110",
        2185=>"111111111",
        2186=>"111010001",
        2187=>"100100100",
        2188=>"111101000",
        2189=>"111101100",
        2190=>"100110010",
        2191=>"001001011",
        2192=>"110100100",
        2193=>"111000000",
        2194=>"101000001",
        2195=>"001001001",
        2196=>"101101000",
        2197=>"111101101",
        2198=>"000100101",
        2199=>"101000110",
        2200=>"100000000",
        2201=>"011011001",
        2202=>"010110011",
        2203=>"100000000",
        2204=>"010010111",
        2205=>"011000000",
        2206=>"101100100",
        2207=>"000001001",
        2208=>"111111101",
        2209=>"100000000",
        2210=>"011111010",
        2211=>"011001111",
        2212=>"001010111",
        2213=>"101101001",
        2214=>"000010110",
        2215=>"111110010",
        2216=>"111000000",
        2217=>"101101011",
        2218=>"000000000",
        2219=>"111000000",
        2220=>"110100001",
        2221=>"101001101",
        2222=>"111000110",
        2223=>"011000001",
        2224=>"100000000",
        2225=>"100111111",
        2226=>"100100000",
        2227=>"000000001",
        2228=>"100000000",
        2229=>"011000100",
        2230=>"100101111",
        2231=>"000010100",
        2232=>"000000000",
        2233=>"111100010",
        2234=>"110111111",
        2235=>"011010000",
        2236=>"001000111",
        2237=>"110000010",
        2238=>"000000000",
        2239=>"110001001",
        2240=>"110100100",
        2241=>"000100000",
        2242=>"101101000",
        2243=>"001000111",
        2244=>"111111110",
        2245=>"100101111",
        2246=>"111101100",
        2247=>"001010010",
        2248=>"011001001",
        2249=>"010000000",
        2250=>"101101000",
        2251=>"000000000",
        2252=>"111100010",
        2253=>"111101010",
        2254=>"000011111",
        2255=>"000110110",
        2256=>"000100000",
        2257=>"011001001",
        2258=>"100000010",
        2259=>"000111010",
        2260=>"010000001",
        2261=>"000100101",
        2262=>"000010000",
        2263=>"100100001",
        2264=>"001000100",
        2265=>"010111111",
        2266=>"000000000",
        2267=>"110110010",
        2268=>"101001001",
        2269=>"100100110",
        2270=>"001110111",
        2271=>"011100010",
        2272=>"011011011",
        2273=>"001000000",
        2274=>"011111111",
        2275=>"001010010",
        2276=>"101111000",
        2277=>"111101101",
        2278=>"110100100",
        2279=>"100101101",
        2280=>"001001001",
        2281=>"001010001",
        2282=>"111000000",
        2283=>"000000000",
        2284=>"001000101",
        2285=>"111100111",
        2286=>"111110111",
        2287=>"001011011",
        2288=>"100101111",
        2289=>"000000111",
        2290=>"111010000",
        2291=>"100000111",
        2292=>"111111011",
        2293=>"000011000",
        2294=>"000100001",
        2295=>"001001000",
        2296=>"000100110",
        2297=>"000000000",
        2298=>"100100100",
        2299=>"000001001",
        2300=>"011011111",
        2301=>"010010111",
        2302=>"101111111",
        2303=>"010011011",
        2304=>"001000000",
        2305=>"000011111",
        2306=>"111100111",
        2307=>"000000000",
        2308=>"001011000",
        2309=>"010110110",
        2310=>"010010000",
        2311=>"010111110",
        2312=>"001011001",
        2313=>"110110111",
        2314=>"010111110",
        2315=>"010001000",
        2316=>"111111111",
        2317=>"010111010",
        2318=>"000000001",
        2319=>"110100111",
        2320=>"010111111",
        2321=>"101000001",
        2322=>"100100111",
        2323=>"100110000",
        2324=>"110111000",
        2325=>"110110101",
        2326=>"111000011",
        2327=>"110000101",
        2328=>"010110100",
        2329=>"010110001",
        2330=>"000101101",
        2331=>"101011111",
        2332=>"000000000",
        2333=>"000100000",
        2334=>"001011000",
        2335=>"111000000",
        2336=>"110110000",
        2337=>"000000001",
        2338=>"011011100",
        2339=>"110100110",
        2340=>"101100101",
        2341=>"110110000",
        2342=>"111011111",
        2343=>"111111100",
        2344=>"000101001",
        2345=>"110101000",
        2346=>"111111111",
        2347=>"001101101",
        2348=>"011001100",
        2349=>"111010000",
        2350=>"101001000",
        2351=>"001000000",
        2352=>"110000111",
        2353=>"011010100",
        2354=>"001000101",
        2355=>"000100000",
        2356=>"100101100",
        2357=>"110111111",
        2358=>"111111111",
        2359=>"000111111",
        2360=>"000000000",
        2361=>"100010011",
        2362=>"011011100",
        2363=>"100101000",
        2364=>"000000000",
        2365=>"001000110",
        2366=>"110011111",
        2367=>"010111111",
        2368=>"001010000",
        2369=>"100000000",
        2370=>"000001111",
        2371=>"101000000",
        2372=>"111001011",
        2373=>"100000001",
        2374=>"000110011",
        2375=>"111000000",
        2376=>"010111111",
        2377=>"000000000",
        2378=>"111011000",
        2379=>"100000000",
        2380=>"000001101",
        2381=>"000000000",
        2382=>"111100001",
        2383=>"001001111",
        2384=>"010001100",
        2385=>"000010000",
        2386=>"000100000",
        2387=>"000010101",
        2388=>"000000100",
        2389=>"000101101",
        2390=>"000010110",
        2391=>"010110010",
        2392=>"011001100",
        2393=>"111111011",
        2394=>"001101111",
        2395=>"001000001",
        2396=>"100111111",
        2397=>"001111110",
        2398=>"011001111",
        2399=>"001000101",
        2400=>"000110100",
        2401=>"000001001",
        2402=>"101111001",
        2403=>"000000000",
        2404=>"001010110",
        2405=>"000010010",
        2406=>"001010100",
        2407=>"111111011",
        2408=>"010111111",
        2409=>"100100101",
        2410=>"100111010",
        2411=>"000110111",
        2412=>"000000000",
        2413=>"000000000",
        2414=>"111110100",
        2415=>"000100000",
        2416=>"101000001",
        2417=>"111001000",
        2418=>"010111111",
        2419=>"000010000",
        2420=>"101001111",
        2421=>"111110111",
        2422=>"111010000",
        2423=>"000100001",
        2424=>"001000100",
        2425=>"000000000",
        2426=>"000011011",
        2427=>"010111111",
        2428=>"110101111",
        2429=>"110000000",
        2430=>"010000000",
        2431=>"110101001",
        2432=>"001001001",
        2433=>"111010000",
        2434=>"111100100",
        2435=>"010000001",
        2436=>"100110100",
        2437=>"101111010",
        2438=>"001000000",
        2439=>"000110111",
        2440=>"111011111",
        2441=>"001100110",
        2442=>"000110000",
        2443=>"110111101",
        2444=>"001111101",
        2445=>"010000010",
        2446=>"011001010",
        2447=>"011011011",
        2448=>"000100000",
        2449=>"111010000",
        2450=>"000100001",
        2451=>"001001011",
        2452=>"001000100",
        2453=>"100101011",
        2454=>"111110111",
        2455=>"000111111",
        2456=>"001010000",
        2457=>"011111101",
        2458=>"000010000",
        2459=>"000001011",
        2460=>"111011000",
        2461=>"001011011",
        2462=>"100100000",
        2463=>"100111111",
        2464=>"001010000",
        2465=>"011000000",
        2466=>"110110100",
        2467=>"111111111",
        2468=>"000011010",
        2469=>"100110010",
        2470=>"111111111",
        2471=>"111101101",
        2472=>"101111110",
        2473=>"011010001",
        2474=>"011011000",
        2475=>"001001001",
        2476=>"100110110",
        2477=>"000111111",
        2478=>"000000110",
        2479=>"111000000",
        2480=>"000011111",
        2481=>"111110110",
        2482=>"010110110",
        2483=>"001001011",
        2484=>"000001001",
        2485=>"110111110",
        2486=>"100010110",
        2487=>"111000010",
        2488=>"010010000",
        2489=>"100110010",
        2490=>"000101001",
        2491=>"000000000",
        2492=>"011000000",
        2493=>"111111111",
        2494=>"001001100",
        2495=>"101111110",
        2496=>"101011000",
        2497=>"010000101",
        2498=>"000011011",
        2499=>"100101010",
        2500=>"100111111",
        2501=>"000001111",
        2502=>"000010110",
        2503=>"011100010",
        2504=>"000001000",
        2505=>"111010000",
        2506=>"110110110",
        2507=>"101111000",
        2508=>"010000011",
        2509=>"000010000",
        2510=>"000110111",
        2511=>"111000001",
        2512=>"000111111",
        2513=>"001001011",
        2514=>"111000100",
        2515=>"111111111",
        2516=>"111100111",
        2517=>"111001000",
        2518=>"000111111",
        2519=>"100001100",
        2520=>"110010100",
        2521=>"001111110",
        2522=>"110110001",
        2523=>"111110010",
        2524=>"111001000",
        2525=>"100100100",
        2526=>"110010000",
        2527=>"010000001",
        2528=>"110110110",
        2529=>"100110110",
        2530=>"000111111",
        2531=>"101111000",
        2532=>"101110111",
        2533=>"000111100",
        2534=>"100100100",
        2535=>"000011111",
        2536=>"101011001",
        2537=>"111111000",
        2538=>"011011001",
        2539=>"101011110",
        2540=>"001000000",
        2541=>"111110000",
        2542=>"000001100",
        2543=>"110110000",
        2544=>"000010000",
        2545=>"100100111",
        2546=>"001101000",
        2547=>"111000000",
        2548=>"010010011",
        2549=>"000000000",
        2550=>"110001000",
        2551=>"001001011",
        2552=>"100110010",
        2553=>"110110100",
        2554=>"001101000",
        2555=>"101010101",
        2556=>"011100100",
        2557=>"010110111",
        2558=>"000000000",
        2559=>"011011011",
        2560=>"101001111",
        2561=>"110110010",
        2562=>"010110111",
        2563=>"111111111",
        2564=>"101100100",
        2565=>"011001011",
        2566=>"111111010",
        2567=>"110111100",
        2568=>"011000011",
        2569=>"100000100",
        2570=>"111000011",
        2571=>"100100000",
        2572=>"011001001",
        2573=>"110100100",
        2574=>"000000001",
        2575=>"011011011",
        2576=>"100100100",
        2577=>"110110010",
        2578=>"001001000",
        2579=>"001010011",
        2580=>"001001000",
        2581=>"111000001",
        2582=>"000001011",
        2583=>"000110110",
        2584=>"100001000",
        2585=>"001000000",
        2586=>"011001101",
        2587=>"110100101",
        2588=>"011101001",
        2589=>"000000100",
        2590=>"000100100",
        2591=>"100111110",
        2592=>"101110110",
        2593=>"100100000",
        2594=>"000000001",
        2595=>"001111011",
        2596=>"111111111",
        2597=>"000111001",
        2598=>"100110100",
        2599=>"001000001",
        2600=>"101111000",
        2601=>"011111111",
        2602=>"011011011",
        2603=>"101000101",
        2604=>"000100100",
        2605=>"101110110",
        2606=>"011110110",
        2607=>"111111101",
        2608=>"000111011",
        2609=>"000110011",
        2610=>"100000000",
        2611=>"001001001",
        2612=>"011001001",
        2613=>"000000001",
        2614=>"010110111",
        2615=>"111111011",
        2616=>"010011011",
        2617=>"001001101",
        2618=>"000001000",
        2619=>"000000001",
        2620=>"000111101",
        2621=>"000000010",
        2622=>"011001110",
        2623=>"011101100",
        2624=>"100001101",
        2625=>"100110111",
        2626=>"111111000",
        2627=>"010000000",
        2628=>"001001000",
        2629=>"010011000",
        2630=>"101011100",
        2631=>"111111110",
        2632=>"011001001",
        2633=>"001001000",
        2634=>"011111110",
        2635=>"000000111",
        2636=>"111111111",
        2637=>"000000010",
        2638=>"111111111",
        2639=>"000000011",
        2640=>"000000010",
        2641=>"111000001",
        2642=>"101100111",
        2643=>"111111011",
        2644=>"110111111",
        2645=>"111110000",
        2646=>"111101111",
        2647=>"000000101",
        2648=>"100100011",
        2649=>"000000000",
        2650=>"011111111",
        2651=>"000000000",
        2652=>"001001001",
        2653=>"100100100",
        2654=>"100101101",
        2655=>"001111000",
        2656=>"100100000",
        2657=>"001001011",
        2658=>"110110010",
        2659=>"001011101",
        2660=>"101111111",
        2661=>"110000000",
        2662=>"011001111",
        2663=>"001111011",
        2664=>"011011001",
        2665=>"110000000",
        2666=>"001001000",
        2667=>"000111111",
        2668=>"101110000",
        2669=>"011010011",
        2670=>"000001000",
        2671=>"101000000",
        2672=>"011001001",
        2673=>"100100110",
        2674=>"101100110",
        2675=>"001001001",
        2676=>"010111111",
        2677=>"011000010",
        2678=>"000110111",
        2679=>"011011001",
        2680=>"111110110",
        2681=>"011111111",
        2682=>"110100100",
        2683=>"110110100",
        2684=>"100100110",
        2685=>"011010000",
        2686=>"100100000",
        2687=>"000100110",
        2688=>"000000000",
        2689=>"000000000",
        2690=>"001111011",
        2691=>"000011111",
        2692=>"000000000",
        2693=>"010000100",
        2694=>"000000000",
        2695=>"000010110",
        2696=>"011000000",
        2697=>"000000000",
        2698=>"111101111",
        2699=>"101011011",
        2700=>"000000000",
        2701=>"000010000",
        2702=>"000000000",
        2703=>"111111001",
        2704=>"101101001",
        2705=>"000000000",
        2706=>"000000000",
        2707=>"001001001",
        2708=>"100011000",
        2709=>"111010110",
        2710=>"111011111",
        2711=>"101101110",
        2712=>"000000000",
        2713=>"000101101",
        2714=>"000000000",
        2715=>"111110110",
        2716=>"000000000",
        2717=>"000000000",
        2718=>"000000000",
        2719=>"111111111",
        2720=>"000011001",
        2721=>"001000000",
        2722=>"000000000",
        2723=>"000111111",
        2724=>"111110111",
        2725=>"110111001",
        2726=>"101101101",
        2727=>"000111111",
        2728=>"111111111",
        2729=>"111111011",
        2730=>"110110100",
        2731=>"000000000",
        2732=>"110011111",
        2733=>"111111111",
        2734=>"111111111",
        2735=>"111111001",
        2736=>"101101111",
        2737=>"111111111",
        2738=>"110111111",
        2739=>"101001110",
        2740=>"000000000",
        2741=>"000000000",
        2742=>"000000000",
        2743=>"010000000",
        2744=>"100110100",
        2745=>"111111111",
        2746=>"000010011",
        2747=>"111111111",
        2748=>"000000111",
        2749=>"000010000",
        2750=>"101011010",
        2751=>"010111101",
        2752=>"111101100",
        2753=>"001000111",
        2754=>"111111101",
        2755=>"000000000",
        2756=>"000000010",
        2757=>"000000000",
        2758=>"000000011",
        2759=>"111111111",
        2760=>"101011111",
        2761=>"000000000",
        2762=>"101111111",
        2763=>"100000000",
        2764=>"111111101",
        2765=>"111111001",
        2766=>"111111110",
        2767=>"001011000",
        2768=>"101111000",
        2769=>"000000010",
        2770=>"000000000",
        2771=>"010000000",
        2772=>"000000000",
        2773=>"001111001",
        2774=>"000000000",
        2775=>"010111110",
        2776=>"000000000",
        2777=>"000110100",
        2778=>"000000000",
        2779=>"111111000",
        2780=>"000000000",
        2781=>"110000100",
        2782=>"000000000",
        2783=>"111001111",
        2784=>"000000001",
        2785=>"100111001",
        2786=>"111111111",
        2787=>"000111100",
        2788=>"001111111",
        2789=>"000010010",
        2790=>"010000111",
        2791=>"111111111",
        2792=>"000000011",
        2793=>"000000000",
        2794=>"000000000",
        2795=>"010001111",
        2796=>"000000000",
        2797=>"111010011",
        2798=>"111000000",
        2799=>"000000000",
        2800=>"110000101",
        2801=>"000111110",
        2802=>"000000000",
        2803=>"010000000",
        2804=>"111111000",
        2805=>"000000110",
        2806=>"000110000",
        2807=>"111111110",
        2808=>"111111111",
        2809=>"111111111",
        2810=>"100000000",
        2811=>"000000101",
        2812=>"000000000",
        2813=>"111111111",
        2814=>"010000010",
        2815=>"000010001",
        2816=>"000100001",
        2817=>"101101101",
        2818=>"001111110",
        2819=>"000010000",
        2820=>"000100111",
        2821=>"111111101",
        2822=>"010000010",
        2823=>"001101110",
        2824=>"001111001",
        2825=>"110110001",
        2826=>"111100101",
        2827=>"111111001",
        2828=>"000110100",
        2829=>"111111010",
        2830=>"010111111",
        2831=>"000000011",
        2832=>"111111111",
        2833=>"000000001",
        2834=>"000111111",
        2835=>"110111111",
        2836=>"100000000",
        2837=>"000000000",
        2838=>"101000000",
        2839=>"111011111",
        2840=>"000111000",
        2841=>"110000000",
        2842=>"101111111",
        2843=>"000011111",
        2844=>"100001100",
        2845=>"100111001",
        2846=>"001111100",
        2847=>"111111111",
        2848=>"000110001",
        2849=>"110110101",
        2850=>"100101100",
        2851=>"010111111",
        2852=>"000010000",
        2853=>"000110010",
        2854=>"011011011",
        2855=>"011000000",
        2856=>"010000000",
        2857=>"011001111",
        2858=>"011011100",
        2859=>"000110110",
        2860=>"001001000",
        2861=>"010011011",
        2862=>"001111111",
        2863=>"010111111",
        2864=>"000000111",
        2865=>"011001010",
        2866=>"010111101",
        2867=>"110010000",
        2868=>"000000000",
        2869=>"000000000",
        2870=>"101101111",
        2871=>"100000000",
        2872=>"100100001",
        2873=>"110010010",
        2874=>"010111111",
        2875=>"100000000",
        2876=>"000000000",
        2877=>"000000101",
        2878=>"010010111",
        2879=>"011111000",
        2880=>"000000101",
        2881=>"010010000",
        2882=>"000000000",
        2883=>"111111100",
        2884=>"111111111",
        2885=>"000111011",
        2886=>"000000000",
        2887=>"011011111",
        2888=>"110111111",
        2889=>"001000000",
        2890=>"111011000",
        2891=>"111101101",
        2892=>"010110110",
        2893=>"000000000",
        2894=>"010111110",
        2895=>"000000000",
        2896=>"001111111",
        2897=>"000001010",
        2898=>"000000000",
        2899=>"011111010",
        2900=>"011111100",
        2901=>"000000001",
        2902=>"100011111",
        2903=>"001001000",
        2904=>"100111100",
        2905=>"111111101",
        2906=>"000011001",
        2907=>"010110000",
        2908=>"000001011",
        2909=>"001001110",
        2910=>"100001000",
        2911=>"101101111",
        2912=>"010100100",
        2913=>"000011000",
        2914=>"111111111",
        2915=>"111111111",
        2916=>"111101110",
        2917=>"001111010",
        2918=>"001100010",
        2919=>"000000000",
        2920=>"110011011",
        2921=>"101000000",
        2922=>"000101101",
        2923=>"111110000",
        2924=>"100100100",
        2925=>"011000000",
        2926=>"010101110",
        2927=>"101111111",
        2928=>"010010110",
        2929=>"000011100",
        2930=>"111110101",
        2931=>"000000011",
        2932=>"000000000",
        2933=>"000000000",
        2934=>"000100000",
        2935=>"010111001",
        2936=>"000000110",
        2937=>"000010011",
        2938=>"100110010",
        2939=>"000000100",
        2940=>"000111001",
        2941=>"111011111",
        2942=>"010111101",
        2943=>"101111111",
        2944=>"010110010",
        2945=>"001001011",
        2946=>"110110000",
        2947=>"110000000",
        2948=>"011000000",
        2949=>"101001111",
        2950=>"100000100",
        2951=>"001001111",
        2952=>"110100000",
        2953=>"000001001",
        2954=>"001001001",
        2955=>"011001011",
        2956=>"000000110",
        2957=>"110110110",
        2958=>"101011010",
        2959=>"011001011",
        2960=>"110100100",
        2961=>"000001011",
        2962=>"111010010",
        2963=>"111111111",
        2964=>"111111111",
        2965=>"000001010",
        2966=>"000000000",
        2967=>"001000100",
        2968=>"111110100",
        2969=>"000001000",
        2970=>"000000001",
        2971=>"111111110",
        2972=>"111001111",
        2973=>"011111011",
        2974=>"001100100",
        2975=>"100100100",
        2976=>"110011110",
        2977=>"101101110",
        2978=>"100111111",
        2979=>"001111101",
        2980=>"110110100",
        2981=>"011001101",
        2982=>"011010111",
        2983=>"110010000",
        2984=>"001011111",
        2985=>"011110110",
        2986=>"011010110",
        2987=>"111010110",
        2988=>"111110010",
        2989=>"110110100",
        2990=>"100110110",
        2991=>"011011111",
        2992=>"110100100",
        2993=>"000100001",
        2994=>"011011001",
        2995=>"110110110",
        2996=>"111110111",
        2997=>"011011010",
        2998=>"000001011",
        2999=>"110000100",
        3000=>"101001000",
        3001=>"111111100",
        3002=>"000001011",
        3003=>"001010010",
        3004=>"001001011",
        3005=>"110100110",
        3006=>"100000010",
        3007=>"001001100",
        3008=>"001001111",
        3009=>"010100001",
        3010=>"001001111",
        3011=>"001001011",
        3012=>"111110110",
        3013=>"111110100",
        3014=>"100000110",
        3015=>"001011111",
        3016=>"000010110",
        3017=>"011001011",
        3018=>"110110100",
        3019=>"000001011",
        3020=>"110000111",
        3021=>"110110000",
        3022=>"110100100",
        3023=>"110100000",
        3024=>"110100000",
        3025=>"001001011",
        3026=>"001001111",
        3027=>"111011101",
        3028=>"100100100",
        3029=>"001001011",
        3030=>"110110100",
        3031=>"110110100",
        3032=>"001111111",
        3033=>"110110000",
        3034=>"011010110",
        3035=>"100100100",
        3036=>"100110110",
        3037=>"000001101",
        3038=>"011001010",
        3039=>"111101111",
        3040=>"111111011",
        3041=>"110110000",
        3042=>"110110000",
        3043=>"100000000",
        3044=>"100000000",
        3045=>"000001011",
        3046=>"001001011",
        3047=>"000011111",
        3048=>"000001001",
        3049=>"000000001",
        3050=>"011010010",
        3051=>"000101000",
        3052=>"110010010",
        3053=>"011011111",
        3054=>"010011110",
        3055=>"110000100",
        3056=>"100001000",
        3057=>"000001111",
        3058=>"000001010",
        3059=>"001001111",
        3060=>"010000011",
        3061=>"011001111",
        3062=>"011011000",
        3063=>"101111101",
        3064=>"101011110",
        3065=>"001001001",
        3066=>"000000010",
        3067=>"110110110",
        3068=>"000000001",
        3069=>"101101101",
        3070=>"011011011",
        3071=>"011110100",
        3072=>"000000000",
        3073=>"111001011",
        3074=>"000000000",
        3075=>"111111100",
        3076=>"001100100",
        3077=>"100100010",
        3078=>"110111111",
        3079=>"101101101",
        3080=>"011001001",
        3081=>"011111100",
        3082=>"100111010",
        3083=>"011000000",
        3084=>"000010001",
        3085=>"111101010",
        3086=>"000010001",
        3087=>"100001011",
        3088=>"000111111",
        3089=>"000001000",
        3090=>"001100000",
        3091=>"100001011",
        3092=>"000111010",
        3093=>"111101000",
        3094=>"101101100",
        3095=>"111010101",
        3096=>"000001101",
        3097=>"100100001",
        3098=>"100101111",
        3099=>"010011001",
        3100=>"000010110",
        3101=>"100100100",
        3102=>"000000100",
        3103=>"000010000",
        3104=>"000101000",
        3105=>"100110100",
        3106=>"001001100",
        3107=>"000000011",
        3108=>"010111000",
        3109=>"011111111",
        3110=>"100100111",
        3111=>"111101010",
        3112=>"111000000",
        3113=>"110110000",
        3114=>"000001100",
        3115=>"110101001",
        3116=>"011000100",
        3117=>"000011111",
        3118=>"000010111",
        3119=>"111000010",
        3120=>"010100001",
        3121=>"111101111",
        3122=>"001100111",
        3123=>"000100000",
        3124=>"000011111",
        3125=>"000110001",
        3126=>"010111011",
        3127=>"000010110",
        3128=>"100000000",
        3129=>"000000100",
        3130=>"011001001",
        3131=>"000000101",
        3132=>"000000000",
        3133=>"100000001",
        3134=>"110110100",
        3135=>"000011000",
        3136=>"100111000",
        3137=>"000001101",
        3138=>"010111111",
        3139=>"011010101",
        3140=>"110110000",
        3141=>"011011001",
        3142=>"010110010",
        3143=>"001000010",
        3144=>"000100001",
        3145=>"110101000",
        3146=>"111011000",
        3147=>"000000001",
        3148=>"111111000",
        3149=>"110100101",
        3150=>"111111111",
        3151=>"111101101",
        3152=>"000011001",
        3153=>"111100111",
        3154=>"100101111",
        3155=>"000000110",
        3156=>"100110100",
        3157=>"101000111",
        3158=>"000101101",
        3159=>"100000101",
        3160=>"000011000",
        3161=>"001000110",
        3162=>"000001001",
        3163=>"000000100",
        3164=>"100001000",
        3165=>"011001000",
        3166=>"101100101",
        3167=>"011111011",
        3168=>"110110100",
        3169=>"011011101",
        3170=>"111000010",
        3171=>"010111010",
        3172=>"010001001",
        3173=>"100101111",
        3174=>"001001101",
        3175=>"111100001",
        3176=>"000011111",
        3177=>"100000100",
        3178=>"110111001",
        3179=>"010100110",
        3180=>"010000000",
        3181=>"111000111",
        3182=>"100000100",
        3183=>"011111001",
        3184=>"010010000",
        3185=>"111010111",
        3186=>"001000001",
        3187=>"111000101",
        3188=>"100000111",
        3189=>"000000011",
        3190=>"000101000",
        3191=>"101001110",
        3192=>"000000111",
        3193=>"110000000",
        3194=>"000110111",
        3195=>"000000111",
        3196=>"000100100",
        3197=>"110100111",
        3198=>"001000111",
        3199=>"110101010",
        3200=>"011000010",
        3201=>"100010010",
        3202=>"100101111",
        3203=>"011101000",
        3204=>"000000100",
        3205=>"100111000",
        3206=>"101000101",
        3207=>"000000001",
        3208=>"100000000",
        3209=>"000101000",
        3210=>"101101011",
        3211=>"010000110",
        3212=>"000000000",
        3213=>"110110111",
        3214=>"011001011",
        3215=>"000100011",
        3216=>"011011000",
        3217=>"011010000",
        3218=>"111000000",
        3219=>"001000000",
        3220=>"000010010",
        3221=>"100000110",
        3222=>"000000000",
        3223=>"000111111",
        3224=>"111000000",
        3225=>"010000001",
        3226=>"110110000",
        3227=>"111110000",
        3228=>"100000011",
        3229=>"001001000",
        3230=>"101001100",
        3231=>"111111111",
        3232=>"100111000",
        3233=>"110001001",
        3234=>"011101100",
        3235=>"111000000",
        3236=>"000100000",
        3237=>"111110010",
        3238=>"000111010",
        3239=>"010010000",
        3240=>"000110101",
        3241=>"000000001",
        3242=>"001000000",
        3243=>"001001001",
        3244=>"111010000",
        3245=>"000000101",
        3246=>"111111000",
        3247=>"000101111",
        3248=>"010000000",
        3249=>"001011011",
        3250=>"101111000",
        3251=>"010100000",
        3252=>"010111110",
        3253=>"000100000",
        3254=>"100000000",
        3255=>"000000111",
        3256=>"000100111",
        3257=>"001011110",
        3258=>"010001000",
        3259=>"000011000",
        3260=>"101110110",
        3261=>"001000001",
        3262=>"111011001",
        3263=>"010000100",
        3264=>"101111000",
        3265=>"000000000",
        3266=>"000111010",
        3267=>"000000101",
        3268=>"000000000",
        3269=>"111000100",
        3270=>"110000000",
        3271=>"000000000",
        3272=>"010010000",
        3273=>"010110000",
        3274=>"100100110",
        3275=>"101000000",
        3276=>"011101111",
        3277=>"111011000",
        3278=>"000000000",
        3279=>"000101111",
        3280=>"001010000",
        3281=>"000000101",
        3282=>"101000000",
        3283=>"010100111",
        3284=>"111000101",
        3285=>"010010000",
        3286=>"111100100",
        3287=>"000001011",
        3288=>"100000000",
        3289=>"111000000",
        3290=>"111111100",
        3291=>"000110010",
        3292=>"111100101",
        3293=>"110000000",
        3294=>"100011110",
        3295=>"000101011",
        3296=>"011001000",
        3297=>"010000100",
        3298=>"000010111",
        3299=>"000001001",
        3300=>"111000000",
        3301=>"000100101",
        3302=>"000000100",
        3303=>"001101011",
        3304=>"100011000",
        3305=>"100100010",
        3306=>"111000001",
        3307=>"110111101",
        3308=>"000101101",
        3309=>"010001000",
        3310=>"010110110",
        3311=>"110100100",
        3312=>"101000101",
        3313=>"111111110",
        3314=>"101111000",
        3315=>"000111111",
        3316=>"101010010",
        3317=>"000010111",
        3318=>"000010000",
        3319=>"111110000",
        3320=>"000000110",
        3321=>"110101100",
        3322=>"000100001",
        3323=>"000101011",
        3324=>"110111000",
        3325=>"001111111",
        3326=>"011100101",
        3327=>"010111111",
        3328=>"001111011",
        3329=>"000000100",
        3330=>"000000100",
        3331=>"111111111",
        3332=>"111111111",
        3333=>"011010101",
        3334=>"111111011",
        3335=>"001101111",
        3336=>"111100101",
        3337=>"111111110",
        3338=>"111111111",
        3339=>"011000000",
        3340=>"101011011",
        3341=>"110110111",
        3342=>"000000100",
        3343=>"100001001",
        3344=>"111101000",
        3345=>"000000000",
        3346=>"111011011",
        3347=>"001111001",
        3348=>"000000000",
        3349=>"000000000",
        3350=>"100100100",
        3351=>"000010010",
        3352=>"100100100",
        3353=>"001011000",
        3354=>"111101101",
        3355=>"111011111",
        3356=>"111011110",
        3357=>"001100011",
        3358=>"001111100",
        3359=>"111110111",
        3360=>"000001010",
        3361=>"111100000",
        3362=>"001001011",
        3363=>"000001011",
        3364=>"111000000",
        3365=>"111001000",
        3366=>"111101001",
        3367=>"000111100",
        3368=>"111011110",
        3369=>"111111111",
        3370=>"000001000",
        3371=>"000000000",
        3372=>"000000000",
        3373=>"010010000",
        3374=>"011111000",
        3375=>"000111011",
        3376=>"000111010",
        3377=>"010000000",
        3378=>"000000000",
        3379=>"011011011",
        3380=>"111101101",
        3381=>"111011000",
        3382=>"111010011",
        3383=>"111111000",
        3384=>"111111111",
        3385=>"001111111",
        3386=>"010111011",
        3387=>"111010000",
        3388=>"000000101",
        3389=>"000000000",
        3390=>"111110110",
        3391=>"000000000",
        3392=>"101111111",
        3393=>"000000000",
        3394=>"111011000",
        3395=>"010110101",
        3396=>"111111111",
        3397=>"011011100",
        3398=>"111110000",
        3399=>"000010001",
        3400=>"111111011",
        3401=>"111111010",
        3402=>"001000100",
        3403=>"000000000",
        3404=>"001000000",
        3405=>"000000000",
        3406=>"010111011",
        3407=>"110111010",
        3408=>"000001101",
        3409=>"000101111",
        3410=>"101100110",
        3411=>"111111011",
        3412=>"100110000",
        3413=>"111111111",
        3414=>"110110010",
        3415=>"010000000",
        3416=>"111101110",
        3417=>"110011000",
        3418=>"111011011",
        3419=>"100100011",
        3420=>"000000001",
        3421=>"111111100",
        3422=>"000000000",
        3423=>"010001001",
        3424=>"000110000",
        3425=>"000100000",
        3426=>"000000110",
        3427=>"010101000",
        3428=>"000010100",
        3429=>"011001001",
        3430=>"111011111",
        3431=>"000000000",
        3432=>"111011001",
        3433=>"001000101",
        3434=>"100001011",
        3435=>"111111001",
        3436=>"111000000",
        3437=>"001001000",
        3438=>"000000000",
        3439=>"000010001",
        3440=>"110111111",
        3441=>"110111110",
        3442=>"010111000",
        3443=>"101001001",
        3444=>"000111000",
        3445=>"000001000",
        3446=>"110111000",
        3447=>"000001001",
        3448=>"000001000",
        3449=>"000111000",
        3450=>"011110000",
        3451=>"010000000",
        3452=>"100110100",
        3453=>"111000011",
        3454=>"010000000",
        3455=>"111100100",
        3456=>"101101111",
        3457=>"010011111",
        3458=>"000000000",
        3459=>"101111010",
        3460=>"100111111",
        3461=>"000000000",
        3462=>"111100111",
        3463=>"000000000",
        3464=>"000001000",
        3465=>"000000000",
        3466=>"111111111",
        3467=>"000000000",
        3468=>"111111101",
        3469=>"011000000",
        3470=>"001001000",
        3471=>"011000000",
        3472=>"001001101",
        3473=>"111011001",
        3474=>"000000001",
        3475=>"000000101",
        3476=>"000110110",
        3477=>"000011000",
        3478=>"101001001",
        3479=>"000111000",
        3480=>"000000100",
        3481=>"000001001",
        3482=>"000100110",
        3483=>"000110000",
        3484=>"110111111",
        3485=>"101101111",
        3486=>"111000000",
        3487=>"111111111",
        3488=>"000000010",
        3489=>"111101111",
        3490=>"000100000",
        3491=>"000000000",
        3492=>"111010000",
        3493=>"001110110",
        3494=>"111000100",
        3495=>"000110010",
        3496=>"000111001",
        3497=>"001111111",
        3498=>"000110101",
        3499=>"001001001",
        3500=>"111101110",
        3501=>"111111111",
        3502=>"001111111",
        3503=>"111111010",
        3504=>"111111111",
        3505=>"111011000",
        3506=>"000001000",
        3507=>"111111001",
        3508=>"101111111",
        3509=>"000101111",
        3510=>"000000000",
        3511=>"000000000",
        3512=>"000111111",
        3513=>"000000000",
        3514=>"000000000",
        3515=>"110111111",
        3516=>"111000001",
        3517=>"000000000",
        3518=>"010010000",
        3519=>"010111010",
        3520=>"110101111",
        3521=>"110110111",
        3522=>"101111010",
        3523=>"111111010",
        3524=>"101011001",
        3525=>"010000000",
        3526=>"000001000",
        3527=>"101111111",
        3528=>"000000100",
        3529=>"011100111",
        3530=>"100110111",
        3531=>"101100101",
        3532=>"111111111",
        3533=>"000000111",
        3534=>"111111111",
        3535=>"110010010",
        3536=>"011111000",
        3537=>"000001001",
        3538=>"000000111",
        3539=>"010111111",
        3540=>"101000000",
        3541=>"010101000",
        3542=>"000001000",
        3543=>"000000000",
        3544=>"001110110",
        3545=>"000000010",
        3546=>"000000000",
        3547=>"000100100",
        3548=>"100101101",
        3549=>"010010000",
        3550=>"110010111",
        3551=>"111111111",
        3552=>"000000001",
        3553=>"111111111",
        3554=>"111000010",
        3555=>"111111111",
        3556=>"000000000",
        3557=>"000111000",
        3558=>"000000110",
        3559=>"101111101",
        3560=>"111111111",
        3561=>"000101101",
        3562=>"000001001",
        3563=>"111111000",
        3564=>"101001111",
        3565=>"111000111",
        3566=>"001100011",
        3567=>"000000000",
        3568=>"111111000",
        3569=>"000100010",
        3570=>"000000110",
        3571=>"000111111",
        3572=>"010000000",
        3573=>"001000100",
        3574=>"000000000",
        3575=>"001000000",
        3576=>"000111110",
        3577=>"000010010",
        3578=>"111111111",
        3579=>"000000000",
        3580=>"000000000",
        3581=>"000001011",
        3582=>"000101000",
        3583=>"110111100",
        3584=>"111111000",
        3585=>"000001111",
        3586=>"111111000",
        3587=>"111111100",
        3588=>"000000000",
        3589=>"111101011",
        3590=>"001101100",
        3591=>"000100101",
        3592=>"011011010",
        3593=>"000100111",
        3594=>"000000000",
        3595=>"001100000",
        3596=>"101000010",
        3597=>"110111000",
        3598=>"100000000",
        3599=>"100001000",
        3600=>"111110000",
        3601=>"000000110",
        3602=>"011111000",
        3603=>"110111010",
        3604=>"111110000",
        3605=>"100110110",
        3606=>"001101101",
        3607=>"010000001",
        3608=>"010110000",
        3609=>"000010010",
        3610=>"011111000",
        3611=>"011000100",
        3612=>"000000101",
        3613=>"011111010",
        3614=>"111001000",
        3615=>"111111011",
        3616=>"110100000",
        3617=>"100011001",
        3618=>"110010000",
        3619=>"111011111",
        3620=>"000111111",
        3621=>"011111010",
        3622=>"110000000",
        3623=>"110110000",
        3624=>"100011110",
        3625=>"011111111",
        3626=>"111111010",
        3627=>"101011011",
        3628=>"000110111",
        3629=>"011111101",
        3630=>"000001011",
        3631=>"000000000",
        3632=>"001110010",
        3633=>"111111000",
        3634=>"001111000",
        3635=>"000000000",
        3636=>"001011000",
        3637=>"110110110",
        3638=>"001101101",
        3639=>"010000000",
        3640=>"000011010",
        3641=>"000000111",
        3642=>"110001111",
        3643=>"000000110",
        3644=>"011111111",
        3645=>"110000111",
        3646=>"110110000",
        3647=>"111111000",
        3648=>"001011000",
        3649=>"100110000",
        3650=>"000100111",
        3651=>"000000001",
        3652=>"111110000",
        3653=>"010010001",
        3654=>"001000000",
        3655=>"111110100",
        3656=>"000000000",
        3657=>"000001111",
        3658=>"011001000",
        3659=>"000111000",
        3660=>"000001111",
        3661=>"000001111",
        3662=>"011001000",
        3663=>"110110000",
        3664=>"000011000",
        3665=>"011000011",
        3666=>"100100000",
        3667=>"000000000",
        3668=>"010010000",
        3669=>"011000100",
        3670=>"111111110",
        3671=>"000000111",
        3672=>"110110110",
        3673=>"100001101",
        3674=>"001000010",
        3675=>"100000101",
        3676=>"001011110",
        3677=>"110100100",
        3678=>"011110000",
        3679=>"000001111",
        3680=>"110000000",
        3681=>"111110000",
        3682=>"010010100",
        3683=>"001010010",
        3684=>"110110001",
        3685=>"110110000",
        3686=>"110100000",
        3687=>"000000000",
        3688=>"000000000",
        3689=>"000000000",
        3690=>"110100000",
        3691=>"110111111",
        3692=>"101011000",
        3693=>"001000100",
        3694=>"000001010",
        3695=>"011100000",
        3696=>"111001000",
        3697=>"101101010",
        3698=>"001000111",
        3699=>"101001001",
        3700=>"010000010",
        3701=>"100101100",
        3702=>"000001111",
        3703=>"111110110",
        3704=>"100111111",
        3705=>"100111110",
        3706=>"000100010",
        3707=>"001000000",
        3708=>"000001000",
        3709=>"011001100",
        3710=>"000010000",
        3711=>"110110010",
        3712=>"111111000",
        3713=>"000111000",
        3714=>"000000001",
        3715=>"101111111",
        3716=>"111111110",
        3717=>"110110110",
        3718=>"101001011",
        3719=>"111000111",
        3720=>"001111100",
        3721=>"001011110",
        3722=>"110111100",
        3723=>"101100000",
        3724=>"000000101",
        3725=>"000110110",
        3726=>"101000000",
        3727=>"111001111",
        3728=>"001100100",
        3729=>"010111111",
        3730=>"011011011",
        3731=>"111110100",
        3732=>"100110100",
        3733=>"000000000",
        3734=>"010000001",
        3735=>"111110111",
        3736=>"111110110",
        3737=>"000001000",
        3738=>"101000001",
        3739=>"000101110",
        3740=>"111111111",
        3741=>"101111111",
        3742=>"000100100",
        3743=>"111110010",
        3744=>"011000000",
        3745=>"000000000",
        3746=>"001100000",
        3747=>"000000101",
        3748=>"111111111",
        3749=>"001110111",
        3750=>"000100110",
        3751=>"111000111",
        3752=>"100100000",
        3753=>"011111111",
        3754=>"000000001",
        3755=>"010000100",
        3756=>"111001001",
        3757=>"110111110",
        3758=>"111000111",
        3759=>"111111111",
        3760=>"000111111",
        3761=>"000000001",
        3762=>"001100110",
        3763=>"001000000",
        3764=>"000010110",
        3765=>"000000011",
        3766=>"000011011",
        3767=>"000000001",
        3768=>"101000000",
        3769=>"111111000",
        3770=>"111110110",
        3771=>"111111010",
        3772=>"000000000",
        3773=>"000000100",
        3774=>"100011011",
        3775=>"000000100",
        3776=>"000000110",
        3777=>"101000001",
        3778=>"110111111",
        3779=>"111111110",
        3780=>"111110000",
        3781=>"110110001",
        3782=>"000001000",
        3783=>"111000101",
        3784=>"111011011",
        3785=>"001011000",
        3786=>"100110100",
        3787=>"000000111",
        3788=>"111111111",
        3789=>"111001011",
        3790=>"110111100",
        3791=>"110111000",
        3792=>"000000111",
        3793=>"000101111",
        3794=>"100000000",
        3795=>"000000000",
        3796=>"010111100",
        3797=>"000000111",
        3798=>"011111001",
        3799=>"010001000",
        3800=>"010110110",
        3801=>"111010000",
        3802=>"001000111",
        3803=>"010111111",
        3804=>"000000001",
        3805=>"111100000",
        3806=>"000000000",
        3807=>"101000000",
        3808=>"000101100",
        3809=>"001011000",
        3810=>"111111010",
        3811=>"000111111",
        3812=>"110111010",
        3813=>"001010011",
        3814=>"001101111",
        3815=>"111111100",
        3816=>"001000001",
        3817=>"001000000",
        3818=>"001111001",
        3819=>"010000011",
        3820=>"101011000",
        3821=>"100000111",
        3822=>"000000000",
        3823=>"111110011",
        3824=>"111110100",
        3825=>"000100100",
        3826=>"111000001",
        3827=>"000111111",
        3828=>"000000001",
        3829=>"000000000",
        3830=>"111000000",
        3831=>"110000011",
        3832=>"000110001",
        3833=>"001000110",
        3834=>"010000001",
        3835=>"111110000",
        3836=>"100001101",
        3837=>"100111011",
        3838=>"000000000",
        3839=>"001000100",
        3840=>"011000000",
        3841=>"111000000",
        3842=>"111101000",
        3843=>"111111000",
        3844=>"000010100",
        3845=>"000010110",
        3846=>"111100100",
        3847=>"000110111",
        3848=>"111011100",
        3849=>"000010011",
        3850=>"010000100",
        3851=>"100011001",
        3852=>"110000011",
        3853=>"110111000",
        3854=>"000000110",
        3855=>"111000000",
        3856=>"111001000",
        3857=>"100000010",
        3858=>"000000110",
        3859=>"000000000",
        3860=>"000110111",
        3861=>"000000111",
        3862=>"011000111",
        3863=>"000111000",
        3864=>"000010001",
        3865=>"111110100",
        3866=>"000000111",
        3867=>"111101111",
        3868=>"000110100",
        3869=>"000000110",
        3870=>"111111101",
        3871=>"011000111",
        3872=>"111110000",
        3873=>"000000001",
        3874=>"111100001",
        3875=>"000111101",
        3876=>"011000000",
        3877=>"111100000",
        3878=>"111000100",
        3879=>"110101000",
        3880=>"000000000",
        3881=>"110111110",
        3882=>"111001110",
        3883=>"100000101",
        3884=>"100010101",
        3885=>"000101111",
        3886=>"110010101",
        3887=>"111101000",
        3888=>"001000010",
        3889=>"110000000",
        3890=>"110110001",
        3891=>"001000000",
        3892=>"100000111",
        3893=>"000000100",
        3894=>"000111000",
        3895=>"111000111",
        3896=>"001110101",
        3897=>"000000001",
        3898=>"001011001",
        3899=>"111001000",
        3900=>"000000111",
        3901=>"111010000",
        3902=>"111111010",
        3903=>"011001000",
        3904=>"111010010",
        3905=>"111111111",
        3906=>"000110111",
        3907=>"111110000",
        3908=>"111000000",
        3909=>"011000100",
        3910=>"000000110",
        3911=>"111101000",
        3912=>"100110000",
        3913=>"111000111",
        3914=>"000000000",
        3915=>"000010111",
        3916=>"000000111",
        3917=>"011101111",
        3918=>"000100011",
        3919=>"111001000",
        3920=>"111101000",
        3921=>"000000110",
        3922=>"000000111",
        3923=>"010000111",
        3924=>"101000000",
        3925=>"000000010",
        3926=>"010001010",
        3927=>"111000110",
        3928=>"001011011",
        3929=>"001111111",
        3930=>"000000000",
        3931=>"111001000",
        3932=>"001011110",
        3933=>"000011011",
        3934=>"111001001",
        3935=>"101101111",
        3936=>"110000000",
        3937=>"110000000",
        3938=>"111111000",
        3939=>"000000111",
        3940=>"111111111",
        3941=>"001000000",
        3942=>"000000110",
        3943=>"110000000",
        3944=>"001000000",
        3945=>"100010100",
        3946=>"000101100",
        3947=>"111111111",
        3948=>"111000000",
        3949=>"000000111",
        3950=>"001001111",
        3951=>"000010011",
        3952=>"000000010",
        3953=>"101111110",
        3954=>"001100010",
        3955=>"010111111",
        3956=>"111001000",
        3957=>"100110100",
        3958=>"111000000",
        3959=>"010111110",
        3960=>"000110111",
        3961=>"000111010",
        3962=>"100000000",
        3963=>"100111111",
        3964=>"011000100",
        3965=>"111111000",
        3966=>"000000111",
        3967=>"111111101",
        3968=>"111111011",
        3969=>"111111111",
        3970=>"111111010",
        3971=>"001101000",
        3972=>"010001000",
        3973=>"000000000",
        3974=>"111010011",
        3975=>"111111111",
        3976=>"001000001",
        3977=>"000000001",
        3978=>"001000000",
        3979=>"000000100",
        3980=>"111111011",
        3981=>"000100000",
        3982=>"111100101",
        3983=>"000010000",
        3984=>"001101000",
        3985=>"010000010",
        3986=>"111111000",
        3987=>"110100100",
        3988=>"101000111",
        3989=>"111111111",
        3990=>"011111111",
        3991=>"111001100",
        3992=>"001011000",
        3993=>"101001011",
        3994=>"111111111",
        3995=>"100100100",
        3996=>"000000000",
        3997=>"111001001",
        3998=>"110110110",
        3999=>"011111111",
        4000=>"111101000",
        4001=>"110100100",
        4002=>"110101100",
        4003=>"000011011",
        4004=>"111010000",
        4005=>"000111110",
        4006=>"111110110",
        4007=>"110111010",
        4008=>"000001000",
        4009=>"010111111",
        4010=>"101101000",
        4011=>"111100100",
        4012=>"000101111",
        4013=>"000011111",
        4014=>"110101101",
        4015=>"110111111",
        4016=>"000000110",
        4017=>"010011010",
        4018=>"000000000",
        4019=>"010111111",
        4020=>"101100000",
        4021=>"001000000",
        4022=>"000000000",
        4023=>"111111110",
        4024=>"110111111",
        4025=>"111001000",
        4026=>"000100010",
        4027=>"110011000",
        4028=>"001111110",
        4029=>"000001101",
        4030=>"001001000",
        4031=>"011111111",
        4032=>"000100000",
        4033=>"001111111",
        4034=>"000000111",
        4035=>"001111111",
        4036=>"111111011",
        4037=>"100111110",
        4038=>"000001001",
        4039=>"111000010",
        4040=>"111101001",
        4041=>"000010010",
        4042=>"001000110",
        4043=>"011001001",
        4044=>"111100010",
        4045=>"000000000",
        4046=>"111111111",
        4047=>"011011001",
        4048=>"011111111",
        4049=>"111111111",
        4050=>"111101100",
        4051=>"000000000",
        4052=>"011011001",
        4053=>"111111111",
        4054=>"001001001",
        4055=>"101000000",
        4056=>"100110110",
        4057=>"000000111",
        4058=>"111111111",
        4059=>"110111011",
        4060=>"101001011",
        4061=>"011011111",
        4062=>"101000000",
        4063=>"110110000",
        4064=>"101000000",
        4065=>"000100000",
        4066=>"010111010",
        4067=>"000000000",
        4068=>"101111111",
        4069=>"111111111",
        4070=>"111111111",
        4071=>"111101111",
        4072=>"111111111",
        4073=>"000011010",
        4074=>"111100000",
        4075=>"000000000",
        4076=>"111111111",
        4077=>"000111000",
        4078=>"001000000",
        4079=>"111101101",
        4080=>"010111111",
        4081=>"000100111",
        4082=>"000000000",
        4083=>"000010011",
        4084=>"110110111",
        4085=>"111011000",
        4086=>"101100111",
        4087=>"001101000",
        4088=>"000100111",
        4089=>"111011100",
        4090=>"011111111",
        4091=>"001000000",
        4092=>"111111111",
        4093=>"000000110",
        4094=>"100111010",
        4095=>"000000000",
        4096=>"000000100",
        4097=>"011001111",
        4098=>"001001111",
        4099=>"110111110",
        4100=>"110000000",
        4101=>"110000100",
        4102=>"000000000",
        4103=>"001101110",
        4104=>"000111000",
        4105=>"110110010",
        4106=>"010001010",
        4107=>"110100000",
        4108=>"110000000",
        4109=>"101101100",
        4110=>"100111111",
        4111=>"001111111",
        4112=>"110100000",
        4113=>"011000100",
        4114=>"110011100",
        4115=>"001000101",
        4116=>"011000000",
        4117=>"000001010",
        4118=>"000001001",
        4119=>"011110011",
        4120=>"100011101",
        4121=>"000100010",
        4122=>"000001000",
        4123=>"000110010",
        4124=>"000110100",
        4125=>"000110101",
        4126=>"111111001",
        4127=>"111111110",
        4128=>"100100110",
        4129=>"100111011",
        4130=>"111001100",
        4131=>"000000110",
        4132=>"110110000",
        4133=>"111000010",
        4134=>"011001011",
        4135=>"110011011",
        4136=>"100100000",
        4137=>"000000110",
        4138=>"100110111",
        4139=>"000110100",
        4140=>"110100110",
        4141=>"001101110",
        4142=>"000100010",
        4143=>"011111010",
        4144=>"000110000",
        4145=>"111001011",
        4146=>"111100100",
        4147=>"000010011",
        4148=>"100110100",
        4149=>"110110100",
        4150=>"001100001",
        4151=>"001001000",
        4152=>"001000001",
        4153=>"110110110",
        4154=>"000000000",
        4155=>"011001111",
        4156=>"011001010",
        4157=>"110010000",
        4158=>"110110000",
        4159=>"110110100",
        4160=>"110110100",
        4161=>"111100000",
        4162=>"100100100",
        4163=>"000001001",
        4164=>"110000001",
        4165=>"111111111",
        4166=>"000001000",
        4167=>"110110010",
        4168=>"100100100",
        4169=>"000001001",
        4170=>"100000100",
        4171=>"110111111",
        4172=>"001100100",
        4173=>"111111100",
        4174=>"111110100",
        4175=>"001011011",
        4176=>"101100011",
        4177=>"001001111",
        4178=>"000000000",
        4179=>"100110010",
        4180=>"111000000",
        4181=>"001001111",
        4182=>"000100010",
        4183=>"110000010",
        4184=>"111101100",
        4185=>"011110001",
        4186=>"001001101",
        4187=>"111001000",
        4188=>"000001001",
        4189=>"111111000",
        4190=>"100101000",
        4191=>"011010111",
        4192=>"110000000",
        4193=>"001001000",
        4194=>"001101111",
        4195=>"100110111",
        4196=>"100100000",
        4197=>"110110100",
        4198=>"110001000",
        4199=>"110110110",
        4200=>"111101001",
        4201=>"100001011",
        4202=>"000111110",
        4203=>"111100011",
        4204=>"000001000",
        4205=>"100001010",
        4206=>"100100110",
        4207=>"110000000",
        4208=>"011001111",
        4209=>"001101100",
        4210=>"110000100",
        4211=>"000010111",
        4212=>"111001111",
        4213=>"000100000",
        4214=>"000100110",
        4215=>"100100111",
        4216=>"100000000",
        4217=>"010100110",
        4218=>"001100111",
        4219=>"010110110",
        4220=>"001001000",
        4221=>"110110110",
        4222=>"100001011",
        4223=>"000010110",
        4224=>"000000100",
        4225=>"000010111",
        4226=>"001000111",
        4227=>"111010000",
        4228=>"001010111",
        4229=>"100010001",
        4230=>"001100011",
        4231=>"000110010",
        4232=>"100111111",
        4233=>"001001000",
        4234=>"101100000",
        4235=>"000000000",
        4236=>"111100000",
        4237=>"110010110",
        4238=>"110100110",
        4239=>"000010110",
        4240=>"111000000",
        4241=>"000011000",
        4242=>"000000000",
        4243=>"010110111",
        4244=>"010100000",
        4245=>"010000000",
        4246=>"000000100",
        4247=>"000111111",
        4248=>"100001010",
        4249=>"110000000",
        4250=>"000000011",
        4251=>"000001000",
        4252=>"101101011",
        4253=>"000000000",
        4254=>"000001100",
        4255=>"000011111",
        4256=>"110111111",
        4257=>"000100101",
        4258=>"011001110",
        4259=>"100111101",
        4260=>"111111101",
        4261=>"000101111",
        4262=>"010110000",
        4263=>"111000000",
        4264=>"000011010",
        4265=>"000111111",
        4266=>"111010001",
        4267=>"010000000",
        4268=>"000000110",
        4269=>"001010000",
        4270=>"010000001",
        4271=>"111011111",
        4272=>"010000110",
        4273=>"111010000",
        4274=>"110000000",
        4275=>"110101000",
        4276=>"000011011",
        4277=>"000100000",
        4278=>"000000111",
        4279=>"111111101",
        4280=>"000111111",
        4281=>"000111111",
        4282=>"010110000",
        4283=>"010011010",
        4284=>"010010010",
        4285=>"010000000",
        4286=>"000000000",
        4287=>"000101111",
        4288=>"000000001",
        4289=>"000011001",
        4290=>"010101111",
        4291=>"101000000",
        4292=>"111000000",
        4293=>"111011001",
        4294=>"110111001",
        4295=>"010111110",
        4296=>"111110000",
        4297=>"111101101",
        4298=>"000010110",
        4299=>"000110111",
        4300=>"110010010",
        4301=>"000000101",
        4302=>"000010010",
        4303=>"101010010",
        4304=>"111010000",
        4305=>"111100000",
        4306=>"000111100",
        4307=>"010100111",
        4308=>"111100110",
        4309=>"111000000",
        4310=>"110001000",
        4311=>"100111111",
        4312=>"011011110",
        4313=>"010000000",
        4314=>"000110111",
        4315=>"110000101",
        4316=>"100000001",
        4317=>"000001111",
        4318=>"100001110",
        4319=>"000010111",
        4320=>"000101111",
        4321=>"111100000",
        4322=>"111111100",
        4323=>"000000101",
        4324=>"001001110",
        4325=>"100111010",
        4326=>"111001000",
        4327=>"000010111",
        4328=>"010011111",
        4329=>"001001011",
        4330=>"000000100",
        4331=>"000101001",
        4332=>"101000101",
        4333=>"100101010",
        4334=>"110111111",
        4335=>"001001101",
        4336=>"111000000",
        4337=>"000000111",
        4338=>"101000000",
        4339=>"111000000",
        4340=>"111101001",
        4341=>"100000000",
        4342=>"000010010",
        4343=>"011010000",
        4344=>"000010110",
        4345=>"000011111",
        4346=>"000110111",
        4347=>"000110111",
        4348=>"100111111",
        4349=>"000100001",
        4350=>"111100010",
        4351=>"010100000",
        4352=>"101010111",
        4353=>"001000111",
        4354=>"000000100",
        4355=>"000011111",
        4356=>"111111111",
        4357=>"111000100",
        4358=>"000000000",
        4359=>"001001001",
        4360=>"101001000",
        4361=>"110110010",
        4362=>"010110000",
        4363=>"011001100",
        4364=>"001000000",
        4365=>"111111111",
        4366=>"010011101",
        4367=>"000001001",
        4368=>"000001011",
        4369=>"001000000",
        4370=>"000101111",
        4371=>"101101100",
        4372=>"010010010",
        4373=>"101000010",
        4374=>"101000101",
        4375=>"010010111",
        4376=>"000001111",
        4377=>"110100001",
        4378=>"110100111",
        4379=>"001001110",
        4380=>"000000011",
        4381=>"100100101",
        4382=>"111111110",
        4383=>"101111111",
        4384=>"000000000",
        4385=>"111100011",
        4386=>"010001000",
        4387=>"111111011",
        4388=>"111111110",
        4389=>"110111110",
        4390=>"000111111",
        4391=>"001000010",
        4392=>"000000000",
        4393=>"110000011",
        4394=>"001000001",
        4395=>"011001100",
        4396=>"101110110",
        4397=>"011111011",
        4398=>"000010010",
        4399=>"000001101",
        4400=>"000010010",
        4401=>"001001111",
        4402=>"000110111",
        4403=>"000011010",
        4404=>"000100100",
        4405=>"111101000",
        4406=>"111100100",
        4407=>"110010000",
        4408=>"011000001",
        4409=>"111000111",
        4410=>"111011001",
        4411=>"101101111",
        4412=>"101000100",
        4413=>"000010000",
        4414=>"110111011",
        4415=>"010011011",
        4416=>"000101101",
        4417=>"000000000",
        4418=>"111111111",
        4419=>"000000000",
        4420=>"111111000",
        4421=>"111110011",
        4422=>"110110000",
        4423=>"001000000",
        4424=>"000010011",
        4425=>"000010010",
        4426=>"000000010",
        4427=>"010001111",
        4428=>"000000000",
        4429=>"111111000",
        4430=>"010110110",
        4431=>"101001111",
        4432=>"000111101",
        4433=>"101000001",
        4434=>"000000111",
        4435=>"111001100",
        4436=>"011011100",
        4437=>"101001101",
        4438=>"100111000",
        4439=>"111010000",
        4440=>"011111110",
        4441=>"011010000",
        4442=>"111001111",
        4443=>"011110000",
        4444=>"101101011",
        4445=>"000000001",
        4446=>"000000111",
        4447=>"000000000",
        4448=>"001010011",
        4449=>"100100110",
        4450=>"000000000",
        4451=>"010010000",
        4452=>"000000010",
        4453=>"000000010",
        4454=>"100000100",
        4455=>"001101111",
        4456=>"001001001",
        4457=>"111100100",
        4458=>"100001111",
        4459=>"010000001",
        4460=>"111001111",
        4461=>"111101000",
        4462=>"111111111",
        4463=>"111111101",
        4464=>"011010000",
        4465=>"001110110",
        4466=>"101000000",
        4467=>"011000101",
        4468=>"111111101",
        4469=>"001000000",
        4470=>"101111111",
        4471=>"000011010",
        4472=>"000000000",
        4473=>"110100001",
        4474=>"100100100",
        4475=>"100001001",
        4476=>"000101111",
        4477=>"010100101",
        4478=>"010000000",
        4479=>"010111110",
        4480=>"000111110",
        4481=>"111001111",
        4482=>"101100111",
        4483=>"111101111",
        4484=>"011100000",
        4485=>"010000100",
        4486=>"110010101",
        4487=>"101101000",
        4488=>"000001001",
        4489=>"111110000",
        4490=>"111100010",
        4491=>"011100010",
        4492=>"111101111",
        4493=>"111000111",
        4494=>"011011001",
        4495=>"000010010",
        4496=>"101000111",
        4497=>"101111111",
        4498=>"110100100",
        4499=>"001001010",
        4500=>"010010000",
        4501=>"000000000",
        4502=>"000101110",
        4503=>"111010010",
        4504=>"100001000",
        4505=>"110000010",
        4506=>"110111001",
        4507=>"011011000",
        4508=>"111010001",
        4509=>"011001000",
        4510=>"111111100",
        4511=>"101111000",
        4512=>"111100000",
        4513=>"111011011",
        4514=>"010100000",
        4515=>"010010000",
        4516=>"000010010",
        4517=>"110111111",
        4518=>"111111111",
        4519=>"010000111",
        4520=>"000010111",
        4521=>"101011001",
        4522=>"000000000",
        4523=>"111000100",
        4524=>"100010000",
        4525=>"101000111",
        4526=>"000000000",
        4527=>"101111111",
        4528=>"000100100",
        4529=>"000100110",
        4530=>"100100000",
        4531=>"000010000",
        4532=>"110100000",
        4533=>"110000001",
        4534=>"110000000",
        4535=>"000000100",
        4536=>"011010011",
        4537=>"000010110",
        4538=>"010010101",
        4539=>"110000111",
        4540=>"000111111",
        4541=>"000100111",
        4542=>"110110000",
        4543=>"011001000",
        4544=>"111000110",
        4545=>"001111000",
        4546=>"010010000",
        4547=>"001000111",
        4548=>"100001010",
        4549=>"101001011",
        4550=>"000000000",
        4551=>"010000000",
        4552=>"111001100",
        4553=>"010000100",
        4554=>"111110010",
        4555=>"100111010",
        4556=>"111101000",
        4557=>"000001111",
        4558=>"111010000",
        4559=>"000111111",
        4560=>"100101111",
        4561=>"001001110",
        4562=>"000000000",
        4563=>"011111010",
        4564=>"100100011",
        4565=>"001001111",
        4566=>"000011001",
        4567=>"111110000",
        4568=>"111100000",
        4569=>"111111011",
        4570=>"111101100",
        4571=>"100110111",
        4572=>"011000000",
        4573=>"100110001",
        4574=>"111100110",
        4575=>"000000111",
        4576=>"011000000",
        4577=>"100100111",
        4578=>"000100111",
        4579=>"010010111",
        4580=>"010010000",
        4581=>"110000000",
        4582=>"011101011",
        4583=>"011000000",
        4584=>"111000111",
        4585=>"110101011",
        4586=>"101001001",
        4587=>"000011001",
        4588=>"101101111",
        4589=>"000011010",
        4590=>"110010001",
        4591=>"100110000",
        4592=>"001111000",
        4593=>"011110100",
        4594=>"110101100",
        4595=>"011011000",
        4596=>"111111111",
        4597=>"101101000",
        4598=>"111101100",
        4599=>"101001001",
        4600=>"010110110",
        4601=>"101101101",
        4602=>"111100101",
        4603=>"001000001",
        4604=>"101001000",
        4605=>"110110001",
        4606=>"111111111",
        4607=>"011011000",
        4608=>"000000011",
        4609=>"111100000",
        4610=>"101010100",
        4611=>"000010010",
        4612=>"000100110",
        4613=>"100000010",
        4614=>"010101010",
        4615=>"101101101",
        4616=>"100111111",
        4617=>"001011011",
        4618=>"111111000",
        4619=>"110111000",
        4620=>"000110111",
        4621=>"111110110",
        4622=>"011101111",
        4623=>"111100000",
        4624=>"000011011",
        4625=>"000000000",
        4626=>"110001001",
        4627=>"001000000",
        4628=>"111000000",
        4629=>"110000000",
        4630=>"000000000",
        4631=>"111111010",
        4632=>"001100010",
        4633=>"011110011",
        4634=>"110111100",
        4635=>"011000000",
        4636=>"111111010",
        4637=>"000001001",
        4638=>"001101000",
        4639=>"000100010",
        4640=>"001101000",
        4641=>"000101110",
        4642=>"100100100",
        4643=>"101111111",
        4644=>"101011111",
        4645=>"111000000",
        4646=>"111011010",
        4647=>"000000111",
        4648=>"011111111",
        4649=>"000001011",
        4650=>"110101111",
        4651=>"100001001",
        4652=>"000000000",
        4653=>"000000111",
        4654=>"000010010",
        4655=>"000010111",
        4656=>"000111111",
        4657=>"000010111",
        4658=>"000101101",
        4659=>"000100111",
        4660=>"000100111",
        4661=>"000000000",
        4662=>"110000000",
        4663=>"110001001",
        4664=>"101111010",
        4665=>"001110010",
        4666=>"100111011",
        4667=>"001001111",
        4668=>"000000111",
        4669=>"000111111",
        4670=>"100100100",
        4671=>"111100000",
        4672=>"111000000",
        4673=>"010000011",
        4674=>"111111010",
        4675=>"111111000",
        4676=>"111111111",
        4677=>"000011011",
        4678=>"111111100",
        4679=>"010011001",
        4680=>"001010001",
        4681=>"111100000",
        4682=>"101000011",
        4683=>"000000010",
        4684=>"111000110",
        4685=>"100111111",
        4686=>"001101111",
        4687=>"000010111",
        4688=>"000001111",
        4689=>"000000111",
        4690=>"011010011",
        4691=>"100100010",
        4692=>"000111110",
        4693=>"111000011",
        4694=>"000011001",
        4695=>"001111010",
        4696=>"101110111",
        4697=>"011111000",
        4698=>"111101001",
        4699=>"111000000",
        4700=>"011110100",
        4701=>"100011010",
        4702=>"111100100",
        4703=>"000111001",
        4704=>"001100010",
        4705=>"000110111",
        4706=>"000111111",
        4707=>"000000000",
        4708=>"111011010",
        4709=>"101000000",
        4710=>"000000001",
        4711=>"000000101",
        4712=>"001100100",
        4713=>"111000000",
        4714=>"011110100",
        4715=>"111000000",
        4716=>"000101100",
        4717=>"000011011",
        4718=>"011000000",
        4719=>"001100011",
        4720=>"000000111",
        4721=>"101000000",
        4722=>"000100100",
        4723=>"100000011",
        4724=>"111101000",
        4725=>"000000111",
        4726=>"001100001",
        4727=>"000001111",
        4728=>"111111000",
        4729=>"000011011",
        4730=>"010000001",
        4731=>"000111111",
        4732=>"110101110",
        4733=>"111001000",
        4734=>"111111110",
        4735=>"010000001",
        4736=>"111011110",
        4737=>"000001011",
        4738=>"110110110",
        4739=>"001111100",
        4740=>"000100011",
        4741=>"001001001",
        4742=>"111111110",
        4743=>"100100100",
        4744=>"000001001",
        4745=>"001011011",
        4746=>"110101001",
        4747=>"000000110",
        4748=>"111110110",
        4749=>"101101101",
        4750=>"000000000",
        4751=>"111110000",
        4752=>"111111111",
        4753=>"001011011",
        4754=>"001001110",
        4755=>"111111000",
        4756=>"001001001",
        4757=>"001100001",
        4758=>"001011011",
        4759=>"011001011",
        4760=>"100100001",
        4761=>"111100001",
        4762=>"100110111",
        4763=>"000000000",
        4764=>"000001001",
        4765=>"110110010",
        4766=>"000000000",
        4767=>"000011001",
        4768=>"111110110",
        4769=>"011000000",
        4770=>"010110010",
        4771=>"001001000",
        4772=>"001011001",
        4773=>"001001001",
        4774=>"000001111",
        4775=>"110110110",
        4776=>"000000000",
        4777=>"111111101",
        4778=>"111001011",
        4779=>"000000000",
        4780=>"111001011",
        4781=>"101111101",
        4782=>"001001001",
        4783=>"000110010",
        4784=>"001000000",
        4785=>"110110110",
        4786=>"101101111",
        4787=>"111000001",
        4788=>"100101010",
        4789=>"001001001",
        4790=>"011001001",
        4791=>"100100000",
        4792=>"110010000",
        4793=>"001001001",
        4794=>"000000000",
        4795=>"111111110",
        4796=>"100110111",
        4797=>"011001011",
        4798=>"111001011",
        4799=>"001000001",
        4800=>"000001000",
        4801=>"110111001",
        4802=>"001001001",
        4803=>"000000000",
        4804=>"000001011",
        4805=>"100000110",
        4806=>"001001000",
        4807=>"001001000",
        4808=>"000011001",
        4809=>"110110111",
        4810=>"111100111",
        4811=>"011011011",
        4812=>"011011011",
        4813=>"001001001",
        4814=>"111001001",
        4815=>"010110110",
        4816=>"111010001",
        4817=>"110110100",
        4818=>"000001001",
        4819=>"000000000",
        4820=>"111100101",
        4821=>"111100110",
        4822=>"010010001",
        4823=>"001000001",
        4824=>"000000000",
        4825=>"000001011",
        4826=>"100100110",
        4827=>"000111111",
        4828=>"110101010",
        4829=>"000000010",
        4830=>"111110110",
        4831=>"110110110",
        4832=>"110001011",
        4833=>"101010110",
        4834=>"110110100",
        4835=>"001001011",
        4836=>"101001001",
        4837=>"010010001",
        4838=>"110110110",
        4839=>"110110100",
        4840=>"110110111",
        4841=>"111111011",
        4842=>"110110100",
        4843=>"001001011",
        4844=>"110110000",
        4845=>"010111111",
        4846=>"001001011",
        4847=>"001001111",
        4848=>"111110110",
        4849=>"000000000",
        4850=>"011011010",
        4851=>"000001000",
        4852=>"000110110",
        4853=>"011110110",
        4854=>"001001001",
        4855=>"011111001",
        4856=>"111000000",
        4857=>"011111001",
        4858=>"111000101",
        4859=>"011001001",
        4860=>"000000001",
        4861=>"000001001",
        4862=>"001110100",
        4863=>"100100111",
        4864=>"000100010",
        4865=>"101100100",
        4866=>"111111101",
        4867=>"001111100",
        4868=>"011111101",
        4869=>"011011000",
        4870=>"101011000",
        4871=>"111100100",
        4872=>"000111111",
        4873=>"110000011",
        4874=>"011100100",
        4875=>"111000001",
        4876=>"100100111",
        4877=>"000111111",
        4878=>"000011001",
        4879=>"111000011",
        4880=>"001100110",
        4881=>"111100100",
        4882=>"001111011",
        4883=>"110000010",
        4884=>"110000111",
        4885=>"000000100",
        4886=>"000000100",
        4887=>"100100101",
        4888=>"100100010",
        4889=>"110110110",
        4890=>"100100111",
        4891=>"001100101",
        4892=>"111011111",
        4893=>"110111110",
        4894=>"000000001",
        4895=>"011011100",
        4896=>"011000111",
        4897=>"110110111",
        4898=>"100100001",
        4899=>"000100100",
        4900=>"011011100",
        4901=>"100100101",
        4902=>"100100101",
        4903=>"100111110",
        4904=>"111000101",
        4905=>"110011110",
        4906=>"110101100",
        4907=>"110101001",
        4908=>"101101001",
        4909=>"111100100",
        4910=>"011000111",
        4911=>"111000100",
        4912=>"011000110",
        4913=>"101000000",
        4914=>"111101111",
        4915=>"001011011",
        4916=>"011101010",
        4917=>"000100111",
        4918=>"111100100",
        4919=>"010011011",
        4920=>"111100100",
        4921=>"100000000",
        4922=>"001000000",
        4923=>"010000000",
        4924=>"111000100",
        4925=>"100011100",
        4926=>"110110110",
        4927=>"100100011",
        4928=>"111111111",
        4929=>"111000100",
        4930=>"111100000",
        4931=>"111100000",
        4932=>"000110000",
        4933=>"000001110",
        4934=>"010011010",
        4935=>"011000111",
        4936=>"110000001",
        4937=>"100111100",
        4938=>"001110000",
        4939=>"000100100",
        4940=>"011000100",
        4941=>"000011010",
        4942=>"011011000",
        4943=>"000000000",
        4944=>"100011100",
        4945=>"100100100",
        4946=>"011010010",
        4947=>"011011111",
        4948=>"000010011",
        4949=>"111010000",
        4950=>"110101000",
        4951=>"010111110",
        4952=>"011111101",
        4953=>"000011011",
        4954=>"000001011",
        4955=>"000010011",
        4956=>"110110100",
        4957=>"001000000",
        4958=>"100001011",
        4959=>"000000000",
        4960=>"101111011",
        4961=>"010011101",
        4962=>"000011000",
        4963=>"000000100",
        4964=>"111101100",
        4965=>"100100100",
        4966=>"000000100",
        4967=>"010110100",
        4968=>"100000001",
        4969=>"111100110",
        4970=>"100100001",
        4971=>"101000000",
        4972=>"000000000",
        4973=>"010100101",
        4974=>"110100010",
        4975=>"000110110",
        4976=>"011010000",
        4977=>"000000001",
        4978=>"100000111",
        4979=>"101100100",
        4980=>"000000000",
        4981=>"000000111",
        4982=>"111100001",
        4983=>"101100111",
        4984=>"011001101",
        4985=>"011111100",
        4986=>"100000101",
        4987=>"100000101",
        4988=>"100010010",
        4989=>"101000011",
        4990=>"110111000",
        4991=>"110111111",
        4992=>"010010110",
        4993=>"000000000",
        4994=>"110010000",
        4995=>"000000100",
        4996=>"001001001",
        4997=>"001000000",
        4998=>"000000000",
        4999=>"000010101",
        5000=>"100001000",
        5001=>"111100100",
        5002=>"111111110",
        5003=>"011001100",
        5004=>"010010000",
        5005=>"010111010",
        5006=>"011100001",
        5007=>"110110011",
        5008=>"111111110",
        5009=>"000000000",
        5010=>"100100000",
        5011=>"010000000",
        5012=>"110010000",
        5013=>"001001010",
        5014=>"000000001",
        5015=>"000101111",
        5016=>"011011011",
        5017=>"110100000",
        5018=>"101101100",
        5019=>"011011010",
        5020=>"111111111",
        5021=>"110110100",
        5022=>"101110111",
        5023=>"100011011",
        5024=>"001001000",
        5025=>"111111101",
        5026=>"011001001",
        5027=>"010111110",
        5028=>"010111110",
        5029=>"001000011",
        5030=>"110110010",
        5031=>"011111111",
        5032=>"111000100",
        5033=>"111011011",
        5034=>"000101011",
        5035=>"100110100",
        5036=>"111001000",
        5037=>"101010000",
        5038=>"101111111",
        5039=>"111111010",
        5040=>"110111110",
        5041=>"000000000",
        5042=>"000100110",
        5043=>"000011011",
        5044=>"111001100",
        5045=>"000000100",
        5046=>"100100000",
        5047=>"000000111",
        5048=>"000000000",
        5049=>"111111001",
        5050=>"111011001",
        5051=>"000000000",
        5052=>"001000000",
        5053=>"000000001",
        5054=>"110110010",
        5055=>"000000011",
        5056=>"010010010",
        5057=>"111111111",
        5058=>"111000101",
        5059=>"110110100",
        5060=>"111110000",
        5061=>"110110110",
        5062=>"010111110",
        5063=>"111111111",
        5064=>"110111101",
        5065=>"111000111",
        5066=>"100110010",
        5067=>"000000101",
        5068=>"111111110",
        5069=>"000101111",
        5070=>"000000111",
        5071=>"000000001",
        5072=>"000010110",
        5073=>"010010000",
        5074=>"000000000",
        5075=>"111101010",
        5076=>"011111111",
        5077=>"000001101",
        5078=>"000010010",
        5079=>"111111101",
        5080=>"101101111",
        5081=>"000000100",
        5082=>"001001011",
        5083=>"111100111",
        5084=>"001011110",
        5085=>"000011001",
        5086=>"001001101",
        5087=>"000000000",
        5088=>"001101011",
        5089=>"110110110",
        5090=>"000000000",
        5091=>"000000000",
        5092=>"000010010",
        5093=>"111010000",
        5094=>"100011000",
        5095=>"010000000",
        5096=>"001010000",
        5097=>"101000101",
        5098=>"000011011",
        5099=>"001101111",
        5100=>"111010000",
        5101=>"001000000",
        5102=>"111001001",
        5103=>"011011001",
        5104=>"010010000",
        5105=>"000001001",
        5106=>"111111011",
        5107=>"001000111",
        5108=>"000000001",
        5109=>"001000000",
        5110=>"000000111",
        5111=>"000001011",
        5112=>"011010000",
        5113=>"101101111",
        5114=>"000000000",
        5115=>"111111111",
        5116=>"100100110",
        5117=>"111101100",
        5118=>"001001111",
        5119=>"110111011",
        5120=>"000111111",
        5121=>"010000000",
        5122=>"010111110",
        5123=>"000111111",
        5124=>"001001111",
        5125=>"111111010",
        5126=>"001111111",
        5127=>"111000000",
        5128=>"000100001",
        5129=>"111011011",
        5130=>"011100111",
        5131=>"101000000",
        5132=>"000000111",
        5133=>"110010000",
        5134=>"110111111",
        5135=>"111000000",
        5136=>"000111100",
        5137=>"110000111",
        5138=>"000111111",
        5139=>"010001011",
        5140=>"000000111",
        5141=>"100000000",
        5142=>"111000000",
        5143=>"111000011",
        5144=>"000001111",
        5145=>"000000101",
        5146=>"100111111",
        5147=>"100011000",
        5148=>"111110111",
        5149=>"001111111",
        5150=>"100100011",
        5151=>"111111011",
        5152=>"000101111",
        5153=>"100100101",
        5154=>"000111111",
        5155=>"111000011",
        5156=>"110111000",
        5157=>"110111111",
        5158=>"011001000",
        5159=>"000100111",
        5160=>"000001101",
        5161=>"111001001",
        5162=>"000000000",
        5163=>"100001101",
        5164=>"111000000",
        5165=>"111000000",
        5166=>"000000000",
        5167=>"111000111",
        5168=>"111011000",
        5169=>"000000011",
        5170=>"100111100",
        5171=>"100111111",
        5172=>"100111101",
        5173=>"111000000",
        5174=>"111110000",
        5175=>"000000111",
        5176=>"010000000",
        5177=>"000000000",
        5178=>"101100000",
        5179=>"000000111",
        5180=>"000111101",
        5181=>"000111111",
        5182=>"011101000",
        5183=>"110010010",
        5184=>"110110100",
        5185=>"000000111",
        5186=>"111000001",
        5187=>"000000000",
        5188=>"000010111",
        5189=>"000111000",
        5190=>"111001000",
        5191=>"111000000",
        5192=>"000000111",
        5193=>"000111111",
        5194=>"111000000",
        5195=>"000100111",
        5196=>"110000000",
        5197=>"110011111",
        5198=>"111000001",
        5199=>"000110110",
        5200=>"111111000",
        5201=>"000001111",
        5202=>"000000100",
        5203=>"101000000",
        5204=>"000111100",
        5205=>"011000000",
        5206=>"000000011",
        5207=>"000101000",
        5208=>"000000111",
        5209=>"001101111",
        5210=>"000111111",
        5211=>"010010000",
        5212=>"000101111",
        5213=>"111000000",
        5214=>"000110111",
        5215=>"111101000",
        5216=>"001101110",
        5217=>"001111001",
        5218=>"111011111",
        5219=>"000000010",
        5220=>"011000000",
        5221=>"000100101",
        5222=>"000100111",
        5223=>"111111000",
        5224=>"001000001",
        5225=>"000000100",
        5226=>"000100111",
        5227=>"110000000",
        5228=>"000111101",
        5229=>"000001001",
        5230=>"111000111",
        5231=>"000001111",
        5232=>"011000101",
        5233=>"111111110",
        5234=>"000000000",
        5235=>"000000111",
        5236=>"011010010",
        5237=>"000000111",
        5238=>"111111001",
        5239=>"101011001",
        5240=>"111000000",
        5241=>"111111110",
        5242=>"100001000",
        5243=>"111111000",
        5244=>"000100111",
        5245=>"000000010",
        5246=>"010010111",
        5247=>"100111010",
        5248=>"101011111",
        5249=>"000000111",
        5250=>"111010000",
        5251=>"000100010",
        5252=>"000101111",
        5253=>"011000000",
        5254=>"010101010",
        5255=>"111000000",
        5256=>"011100100",
        5257=>"000000100",
        5258=>"000101111",
        5259=>"001001001",
        5260=>"001001011",
        5261=>"110110010",
        5262=>"111010000",
        5263=>"011011000",
        5264=>"100110000",
        5265=>"011010010",
        5266=>"000101111",
        5267=>"000001011",
        5268=>"101000111",
        5269=>"001000000",
        5270=>"111101000",
        5271=>"000000000",
        5272=>"001001111",
        5273=>"000100101",
        5274=>"001100111",
        5275=>"011011001",
        5276=>"000000101",
        5277=>"100100000",
        5278=>"100100111",
        5279=>"101111001",
        5280=>"101101111",
        5281=>"100100110",
        5282=>"100100001",
        5283=>"010000000",
        5284=>"101010000",
        5285=>"111000000",
        5286=>"111110000",
        5287=>"101000010",
        5288=>"000101100",
        5289=>"101111011",
        5290=>"001101111",
        5291=>"000001101",
        5292=>"111111101",
        5293=>"111000101",
        5294=>"100110111",
        5295=>"111111000",
        5296=>"110100010",
        5297=>"110000000",
        5298=>"000111111",
        5299=>"111001010",
        5300=>"001001111",
        5301=>"000001111",
        5302=>"100101111",
        5303=>"001100101",
        5304=>"000000100",
        5305=>"111001000",
        5306=>"000000011",
        5307=>"000001101",
        5308=>"000000100",
        5309=>"111110000",
        5310=>"111110100",
        5311=>"100100000",
        5312=>"000101111",
        5313=>"111000000",
        5314=>"001010010",
        5315=>"010000000",
        5316=>"011111000",
        5317=>"100110011",
        5318=>"111000111",
        5319=>"001101101",
        5320=>"001001111",
        5321=>"000000111",
        5322=>"100100100",
        5323=>"000000100",
        5324=>"111111010",
        5325=>"000111101",
        5326=>"111010000",
        5327=>"111010000",
        5328=>"000100000",
        5329=>"011000100",
        5330=>"100000111",
        5331=>"110100110",
        5332=>"011111110",
        5333=>"000000000",
        5334=>"111101000",
        5335=>"111010000",
        5336=>"000100111",
        5337=>"000000000",
        5338=>"001001011",
        5339=>"011110010",
        5340=>"000101100",
        5341=>"100100110",
        5342=>"000100001",
        5343=>"100110000",
        5344=>"110110000",
        5345=>"111001000",
        5346=>"111111010",
        5347=>"001111010",
        5348=>"111111000",
        5349=>"111000101",
        5350=>"100000001",
        5351=>"011111100",
        5352=>"000000001",
        5353=>"000000101",
        5354=>"000001110",
        5355=>"010111111",
        5356=>"010000111",
        5357=>"011000101",
        5358=>"000000001",
        5359=>"111011001",
        5360=>"000111000",
        5361=>"100101101",
        5362=>"000000111",
        5363=>"000000100",
        5364=>"010011100",
        5365=>"111000000",
        5366=>"000011001",
        5367=>"010111111",
        5368=>"111101000",
        5369=>"000100111",
        5370=>"001001101",
        5371=>"000001101",
        5372=>"100110111",
        5373=>"000110000",
        5374=>"000101111",
        5375=>"001111011",
        5376=>"101111000",
        5377=>"001000100",
        5378=>"111111000",
        5379=>"000000100",
        5380=>"011011111",
        5381=>"001001111",
        5382=>"000101000",
        5383=>"000000000",
        5384=>"100101111",
        5385=>"010000001",
        5386=>"111110110",
        5387=>"001001000",
        5388=>"000000001",
        5389=>"110111110",
        5390=>"000100000",
        5391=>"110110001",
        5392=>"110111111",
        5393=>"000000000",
        5394=>"111011100",
        5395=>"110110101",
        5396=>"010000000",
        5397=>"000111000",
        5398=>"000000000",
        5399=>"011111000",
        5400=>"110100101",
        5401=>"100101101",
        5402=>"010001101",
        5403=>"000000011",
        5404=>"000001111",
        5405=>"100100000",
        5406=>"110000101",
        5407=>"010010110",
        5408=>"000000111",
        5409=>"001000100",
        5410=>"001001100",
        5411=>"000101110",
        5412=>"010011000",
        5413=>"011000000",
        5414=>"000000000",
        5415=>"111110010",
        5416=>"110000000",
        5417=>"000011111",
        5418=>"001000001",
        5419=>"000000000",
        5420=>"011001000",
        5421=>"000111000",
        5422=>"000000100",
        5423=>"000000000",
        5424=>"101111010",
        5425=>"110110000",
        5426=>"000100001",
        5427=>"100100001",
        5428=>"000100101",
        5429=>"101001101",
        5430=>"111111111",
        5431=>"000000010",
        5432=>"000111011",
        5433=>"000101000",
        5434=>"010000000",
        5435=>"000001101",
        5436=>"111111111",
        5437=>"000000111",
        5438=>"000000110",
        5439=>"101101011",
        5440=>"110110100",
        5441=>"000000000",
        5442=>"101111111",
        5443=>"101000000",
        5444=>"110011010",
        5445=>"000110100",
        5446=>"011101111",
        5447=>"000000000",
        5448=>"011100001",
        5449=>"001111110",
        5450=>"000000110",
        5451=>"000000000",
        5452=>"000000111",
        5453=>"110111010",
        5454=>"010110110",
        5455=>"000110010",
        5456=>"011111111",
        5457=>"000000000",
        5458=>"000010010",
        5459=>"000000100",
        5460=>"000010000",
        5461=>"000000000",
        5462=>"000000000",
        5463=>"111001001",
        5464=>"001110110",
        5465=>"111010011",
        5466=>"000000110",
        5467=>"000000000",
        5468=>"100100110",
        5469=>"000010110",
        5470=>"111111101",
        5471=>"111101111",
        5472=>"010010010",
        5473=>"101111110",
        5474=>"111111111",
        5475=>"000000000",
        5476=>"000000000",
        5477=>"000010011",
        5478=>"000000000",
        5479=>"011000001",
        5480=>"000000000",
        5481=>"011000010",
        5482=>"000011011",
        5483=>"010000101",
        5484=>"010111011",
        5485=>"111111111",
        5486=>"111000111",
        5487=>"000001001",
        5488=>"111111110",
        5489=>"111100110",
        5490=>"111101101",
        5491=>"000000111",
        5492=>"111111000",
        5493=>"000000001",
        5494=>"101000100",
        5495=>"000000000",
        5496=>"011001000",
        5497=>"100000000",
        5498=>"000001001",
        5499=>"001101100",
        5500=>"011111111",
        5501=>"011010100",
        5502=>"111110010",
        5503=>"010000010",
        5504=>"010011011",
        5505=>"011011011",
        5506=>"010100110",
        5507=>"111100010",
        5508=>"110111111",
        5509=>"111101100",
        5510=>"001000010",
        5511=>"111111000",
        5512=>"000010100",
        5513=>"000000000",
        5514=>"101000001",
        5515=>"111011001",
        5516=>"111110101",
        5517=>"000010110",
        5518=>"000000000",
        5519=>"111110100",
        5520=>"000111010",
        5521=>"100101001",
        5522=>"000111111",
        5523=>"011111111",
        5524=>"100100111",
        5525=>"111111111",
        5526=>"101101101",
        5527=>"000000000",
        5528=>"010110111",
        5529=>"111110101",
        5530=>"110110111",
        5531=>"000000000",
        5532=>"111101111",
        5533=>"001011111",
        5534=>"010001001",
        5535=>"100111101",
        5536=>"101111111",
        5537=>"000000110",
        5538=>"011111001",
        5539=>"000000000",
        5540=>"000000000",
        5541=>"111101111",
        5542=>"111001101",
        5543=>"110111110",
        5544=>"111111001",
        5545=>"110111100",
        5546=>"011011010",
        5547=>"001011110",
        5548=>"110111011",
        5549=>"111010000",
        5550=>"000100100",
        5551=>"110101111",
        5552=>"010000000",
        5553=>"000000111",
        5554=>"100111101",
        5555=>"110110100",
        5556=>"010111111",
        5557=>"000000000",
        5558=>"000010110",
        5559=>"101111001",
        5560=>"000000010",
        5561=>"100111111",
        5562=>"000000000",
        5563=>"000010111",
        5564=>"000001111",
        5565=>"000010000",
        5566=>"000000000",
        5567=>"100000100",
        5568=>"110010000",
        5569=>"011111111",
        5570=>"111111101",
        5571=>"000010000",
        5572=>"111011101",
        5573=>"100110110",
        5574=>"011111110",
        5575=>"111011000",
        5576=>"111111011",
        5577=>"010010010",
        5578=>"111111011",
        5579=>"000000000",
        5580=>"100111110",
        5581=>"000010010",
        5582=>"000111100",
        5583=>"101101100",
        5584=>"100111101",
        5585=>"011011110",
        5586=>"000011110",
        5587=>"110100110",
        5588=>"001001011",
        5589=>"111000000",
        5590=>"000000000",
        5591=>"000000100",
        5592=>"011011011",
        5593=>"000000000",
        5594=>"011011111",
        5595=>"100000001",
        5596=>"001010111",
        5597=>"111110111",
        5598=>"011111111",
        5599=>"001111100",
        5600=>"000010000",
        5601=>"110001001",
        5602=>"111100110",
        5603=>"010101111",
        5604=>"111111000",
        5605=>"010011011",
        5606=>"110111011",
        5607=>"101000100",
        5608=>"111111111",
        5609=>"011000111",
        5610=>"000111110",
        5611=>"000000000",
        5612=>"111010010",
        5613=>"000001111",
        5614=>"000000000",
        5615=>"000000000",
        5616=>"101111111",
        5617=>"111111111",
        5618=>"010111011",
        5619=>"101100101",
        5620=>"000011111",
        5621=>"111011101",
        5622=>"111111101",
        5623=>"001111100",
        5624=>"010111000",
        5625=>"010010000",
        5626=>"111111111",
        5627=>"111111010",
        5628=>"011000011",
        5629=>"000000000",
        5630=>"101101000",
        5631=>"101101110",
        5632=>"111111111",
        5633=>"001000001",
        5634=>"000100111",
        5635=>"101110111",
        5636=>"101101111",
        5637=>"111111000",
        5638=>"000100110",
        5639=>"010100101",
        5640=>"101101010",
        5641=>"011001110",
        5642=>"101101000",
        5643=>"011000100",
        5644=>"100000000",
        5645=>"111111000",
        5646=>"001101111",
        5647=>"110000001",
        5648=>"000000100",
        5649=>"110000101",
        5650=>"100100110",
        5651=>"111100111",
        5652=>"101001101",
        5653=>"000001000",
        5654=>"000000000",
        5655=>"000000110",
        5656=>"000000110",
        5657=>"110100111",
        5658=>"001110111",
        5659=>"000100111",
        5660=>"111000000",
        5661=>"000011110",
        5662=>"001001000",
        5663=>"011101111",
        5664=>"000101101",
        5665=>"101101110",
        5666=>"011101111",
        5667=>"010110110",
        5668=>"111111111",
        5669=>"001001100",
        5670=>"000110111",
        5671=>"000000101",
        5672=>"010000000",
        5673=>"000111111",
        5674=>"000000111",
        5675=>"100110010",
        5676=>"001011010",
        5677=>"000000111",
        5678=>"110000000",
        5679=>"000100111",
        5680=>"000111111",
        5681=>"000000000",
        5682=>"001000110",
        5683=>"000001001",
        5684=>"001110011",
        5685=>"111111000",
        5686=>"000010000",
        5687=>"010110000",
        5688=>"100100111",
        5689=>"101011010",
        5690=>"110100011",
        5691=>"000111110",
        5692=>"000100101",
        5693=>"000000110",
        5694=>"001011110",
        5695=>"011011010",
        5696=>"101111001",
        5697=>"000000110",
        5698=>"010010111",
        5699=>"000000000",
        5700=>"101101101",
        5701=>"100110111",
        5702=>"010110110",
        5703=>"111000000",
        5704=>"000000000",
        5705=>"110111000",
        5706=>"010000001",
        5707=>"001000001",
        5708=>"000100011",
        5709=>"000100000",
        5710=>"010111101",
        5711=>"010110000",
        5712=>"010000111",
        5713=>"000000100",
        5714=>"010000000",
        5715=>"111111010",
        5716=>"000111111",
        5717=>"000000000",
        5718=>"000100111",
        5719=>"111111100",
        5720=>"111111111",
        5721=>"110101000",
        5722=>"000111111",
        5723=>"100000001",
        5724=>"101111010",
        5725=>"001000000",
        5726=>"100001111",
        5727=>"010000000",
        5728=>"101001010",
        5729=>"000110100",
        5730=>"011001000",
        5731=>"000001111",
        5732=>"010000111",
        5733=>"001100110",
        5734=>"000000001",
        5735=>"010010000",
        5736=>"100000001",
        5737=>"111100100",
        5738=>"100101111",
        5739=>"111000000",
        5740=>"001101000",
        5741=>"000111000",
        5742=>"110111001",
        5743=>"100100110",
        5744=>"010010000",
        5745=>"111100000",
        5746=>"000000100",
        5747=>"000000000",
        5748=>"010111111",
        5749=>"000000000",
        5750=>"101111000",
        5751=>"100100001",
        5752=>"000000111",
        5753=>"111000110",
        5754=>"011000101",
        5755=>"001000000",
        5756=>"000101111",
        5757=>"110010010",
        5758=>"010110101",
        5759=>"101110010",
        5760=>"000000000",
        5761=>"000111111",
        5762=>"111000000",
        5763=>"011011111",
        5764=>"001000000",
        5765=>"000110111",
        5766=>"000000000",
        5767=>"110000000",
        5768=>"001001011",
        5769=>"011000111",
        5770=>"001000000",
        5771=>"001000100",
        5772=>"001000001",
        5773=>"000111110",
        5774=>"000001001",
        5775=>"110111111",
        5776=>"011010111",
        5777=>"100111010",
        5778=>"001001101",
        5779=>"100100100",
        5780=>"111111000",
        5781=>"000100111",
        5782=>"101000001",
        5783=>"000000000",
        5784=>"101100101",
        5785=>"000000001",
        5786=>"001001101",
        5787=>"011111110",
        5788=>"000000000",
        5789=>"111101101",
        5790=>"001000000",
        5791=>"000000000",
        5792=>"101100011",
        5793=>"111100100",
        5794=>"001011100",
        5795=>"111111111",
        5796=>"100000111",
        5797=>"111000000",
        5798=>"000111111",
        5799=>"011101101",
        5800=>"011000000",
        5801=>"000000001",
        5802=>"001111110",
        5803=>"101101101",
        5804=>"001001100",
        5805=>"111101000",
        5806=>"101000000",
        5807=>"111010111",
        5808=>"011111011",
        5809=>"011110110",
        5810=>"011010010",
        5811=>"000000000",
        5812=>"101101101",
        5813=>"010000000",
        5814=>"111000000",
        5815=>"000100001",
        5816=>"000000000",
        5817=>"001000000",
        5818=>"110000011",
        5819=>"000000000",
        5820=>"000010111",
        5821=>"011011101",
        5822=>"110111111",
        5823=>"101000000",
        5824=>"000100100",
        5825=>"001000000",
        5826=>"111001001",
        5827=>"000011000",
        5828=>"000000000",
        5829=>"111111111",
        5830=>"111100000",
        5831=>"000000000",
        5832=>"110110011",
        5833=>"000111111",
        5834=>"111000100",
        5835=>"000111111",
        5836=>"111111100",
        5837=>"011011000",
        5838=>"000000000",
        5839=>"010111010",
        5840=>"111101111",
        5841=>"110101011",
        5842=>"000111111",
        5843=>"001000000",
        5844=>"111111111",
        5845=>"010111010",
        5846=>"111111101",
        5847=>"000000000",
        5848=>"000000100",
        5849=>"001101110",
        5850=>"000000001",
        5851=>"010110010",
        5852=>"100101111",
        5853=>"011001011",
        5854=>"000110110",
        5855=>"000000000",
        5856=>"100110111",
        5857=>"110011011",
        5858=>"111111111",
        5859=>"111111000",
        5860=>"111000000",
        5861=>"001000111",
        5862=>"011111110",
        5863=>"101000000",
        5864=>"001000000",
        5865=>"110110111",
        5866=>"100100001",
        5867=>"000000000",
        5868=>"011010111",
        5869=>"111111111",
        5870=>"000000000",
        5871=>"101100000",
        5872=>"111001010",
        5873=>"000000000",
        5874=>"000000000",
        5875=>"101000000",
        5876=>"000111111",
        5877=>"001000001",
        5878=>"000000011",
        5879=>"000010010",
        5880=>"111001100",
        5881=>"111000000",
        5882=>"100000001",
        5883=>"000000010",
        5884=>"000100100",
        5885=>"111111111",
        5886=>"100000000",
        5887=>"110110110",
        5888=>"011011111",
        5889=>"101100000",
        5890=>"000010000",
        5891=>"000110000",
        5892=>"001011110",
        5893=>"010111000",
        5894=>"011010000",
        5895=>"100101001",
        5896=>"010110111",
        5897=>"100000000",
        5898=>"100110100",
        5899=>"011111111",
        5900=>"001011000",
        5901=>"001010001",
        5902=>"011111110",
        5903=>"100100101",
        5904=>"000000001",
        5905=>"100001011",
        5906=>"100110100",
        5907=>"011010110",
        5908=>"001010010",
        5909=>"011101100",
        5910=>"000000000",
        5911=>"001001011",
        5912=>"111110100",
        5913=>"001000000",
        5914=>"000000110",
        5915=>"000000000",
        5916=>"110011110",
        5917=>"001010110",
        5918=>"000110110",
        5919=>"010100000",
        5920=>"011110110",
        5921=>"010010100",
        5922=>"000000000",
        5923=>"010101100",
        5924=>"001011011",
        5925=>"010010011",
        5926=>"000001001",
        5927=>"001011110",
        5928=>"011011001",
        5929=>"011010110",
        5930=>"011111111",
        5931=>"011110110",
        5932=>"000001000",
        5933=>"100100001",
        5934=>"000110100",
        5935=>"010011010",
        5936=>"011111000",
        5937=>"100101000",
        5938=>"011011011",
        5939=>"011010110",
        5940=>"010010100",
        5941=>"001100100",
        5942=>"011010000",
        5943=>"100101110",
        5944=>"100101011",
        5945=>"010110100",
        5946=>"000001010",
        5947=>"000101001",
        5948=>"111101001",
        5949=>"000000010",
        5950=>"011111000",
        5951=>"011011011",
        5952=>"011011000",
        5953=>"100100000",
        5954=>"001010000",
        5955=>"100111110",
        5956=>"011010000",
        5957=>"011011010",
        5958=>"001011110",
        5959=>"111011011",
        5960=>"011011010",
        5961=>"001000011",
        5962=>"000001001",
        5963=>"000101001",
        5964=>"100000000",
        5965=>"100100100",
        5966=>"000000000",
        5967=>"100001001",
        5968=>"001001001",
        5969=>"011010000",
        5970=>"101100100",
        5971=>"111111111",
        5972=>"001010100",
        5973=>"100000001",
        5974=>"011011011",
        5975=>"110101010",
        5976=>"000000100",
        5977=>"010000011",
        5978=>"001101111",
        5979=>"000001000",
        5980=>"011110110",
        5981=>"100001001",
        5982=>"000000011",
        5983=>"110101001",
        5984=>"011010011",
        5985=>"000001000",
        5986=>"101111010",
        5987=>"001010110",
        5988=>"001001000",
        5989=>"100001000",
        5990=>"100101001",
        5991=>"010011110",
        5992=>"100101001",
        5993=>"010110100",
        5994=>"011010110",
        5995=>"101000010",
        5996=>"110101101",
        5997=>"100101001",
        5998=>"100111010",
        5999=>"111110100",
        6000=>"100001001",
        6001=>"001001011",
        6002=>"010011000",
        6003=>"011011110",
        6004=>"000101110",
        6005=>"000100000",
        6006=>"011101101",
        6007=>"100000001",
        6008=>"000001000",
        6009=>"011111101",
        6010=>"010010110",
        6011=>"110100011",
        6012=>"000000100",
        6013=>"101111100",
        6014=>"100101000",
        6015=>"111111110",
        6016=>"110111111",
        6017=>"101100100",
        6018=>"000011000",
        6019=>"000111011",
        6020=>"000000001",
        6021=>"000011111",
        6022=>"111111010",
        6023=>"000000100",
        6024=>"100101111",
        6025=>"001001001",
        6026=>"111100000",
        6027=>"101101000",
        6028=>"000000000",
        6029=>"111101111",
        6030=>"110110001",
        6031=>"000010111",
        6032=>"100000100",
        6033=>"000111011",
        6034=>"110101101",
        6035=>"000100100",
        6036=>"010110000",
        6037=>"100000001",
        6038=>"011100000",
        6039=>"111111100",
        6040=>"100101111",
        6041=>"110100000",
        6042=>"100101101",
        6043=>"111100001",
        6044=>"001110011",
        6045=>"000111111",
        6046=>"001100001",
        6047=>"000010000",
        6048=>"110000100",
        6049=>"100100100",
        6050=>"010001100",
        6051=>"011000000",
        6052=>"111111001",
        6053=>"010111111",
        6054=>"111111111",
        6055=>"000011111",
        6056=>"111111111",
        6057=>"111000111",
        6058=>"101000001",
        6059=>"000101101",
        6060=>"011101010",
        6061=>"000000100",
        6062=>"111111111",
        6063=>"111111111",
        6064=>"100100100",
        6065=>"000000100",
        6066=>"110000000",
        6067=>"000011000",
        6068=>"000100101",
        6069=>"011001111",
        6070=>"100100101",
        6071=>"000111110",
        6072=>"111101000",
        6073=>"111001000",
        6074=>"100100100",
        6075=>"110000000",
        6076=>"100000000",
        6077=>"100111010",
        6078=>"111001100",
        6079=>"111000010",
        6080=>"101100111",
        6081=>"000000000",
        6082=>"010111000",
        6083=>"101001101",
        6084=>"101111000",
        6085=>"000101011",
        6086=>"100111110",
        6087=>"000010011",
        6088=>"001000001",
        6089=>"010111111",
        6090=>"111101111",
        6091=>"011101101",
        6092=>"011000000",
        6093=>"111100010",
        6094=>"110001000",
        6095=>"000011110",
        6096=>"011000100",
        6097=>"001111101",
        6098=>"100000110",
        6099=>"100011111",
        6100=>"100100110",
        6101=>"000000001",
        6102=>"111000000",
        6103=>"000011111",
        6104=>"111101110",
        6105=>"000000111",
        6106=>"001001001",
        6107=>"000010111",
        6108=>"100001000",
        6109=>"000011001",
        6110=>"100100110",
        6111=>"000000000",
        6112=>"111101110",
        6113=>"000100001",
        6114=>"000010101",
        6115=>"011111010",
        6116=>"010001110",
        6117=>"101000101",
        6118=>"100000000",
        6119=>"010100111",
        6120=>"000001000",
        6121=>"100000000",
        6122=>"000100101",
        6123=>"111010111",
        6124=>"000100000",
        6125=>"000010111",
        6126=>"111101011",
        6127=>"011011111",
        6128=>"000011000",
        6129=>"000000000",
        6130=>"100000000",
        6131=>"111111111",
        6132=>"000001001",
        6133=>"000000000",
        6134=>"000000010",
        6135=>"100000000",
        6136=>"011000011",
        6137=>"010000100",
        6138=>"000100000",
        6139=>"000000000",
        6140=>"000100100",
        6141=>"111011010",
        6142=>"111101100",
        6143=>"010111111",
        6144=>"011111011",
        6145=>"000000000",
        6146=>"001000000",
        6147=>"100001000",
        6148=>"001001100",
        6149=>"111111100",
        6150=>"010111110",
        6151=>"000111101",
        6152=>"110110001",
        6153=>"001100100",
        6154=>"010110110",
        6155=>"001001001",
        6156=>"001000001",
        6157=>"111111111",
        6158=>"100001001",
        6159=>"110010010",
        6160=>"100100001",
        6161=>"000000100",
        6162=>"000001001",
        6163=>"100100001",
        6164=>"011111011",
        6165=>"100000000",
        6166=>"100100000",
        6167=>"101010111",
        6168=>"100101101",
        6169=>"000000000",
        6170=>"000011100",
        6171=>"001001011",
        6172=>"000000010",
        6173=>"100100001",
        6174=>"001001010",
        6175=>"110011001",
        6176=>"001100110",
        6177=>"101100001",
        6178=>"101010100",
        6179=>"000010010",
        6180=>"111111000",
        6181=>"111101101",
        6182=>"111010110",
        6183=>"111010000",
        6184=>"110010100",
        6185=>"110110111",
        6186=>"000000110",
        6187=>"100101001",
        6188=>"011110100",
        6189=>"011111010",
        6190=>"101110110",
        6191=>"000101101",
        6192=>"000111111",
        6193=>"000000100",
        6194=>"101100100",
        6195=>"100100011",
        6196=>"000101111",
        6197=>"111011110",
        6198=>"000100100",
        6199=>"001010010",
        6200=>"111101110",
        6201=>"101000000",
        6202=>"000001001",
        6203=>"000001111",
        6204=>"010111000",
        6205=>"100100011",
        6206=>"000100101",
        6207=>"000001011",
        6208=>"111110000",
        6209=>"000010000",
        6210=>"010000010",
        6211=>"111010000",
        6212=>"101001001",
        6213=>"100111111",
        6214=>"011011110",
        6215=>"101011000",
        6216=>"001001100",
        6217=>"000110011",
        6218=>"011000110",
        6219=>"000001000",
        6220=>"111010110",
        6221=>"010110000",
        6222=>"110110111",
        6223=>"100011001",
        6224=>"010000011",
        6225=>"100110011",
        6226=>"011011100",
        6227=>"000011001",
        6228=>"001101110",
        6229=>"111000111",
        6230=>"001000111",
        6231=>"101101101",
        6232=>"001101110",
        6233=>"101101111",
        6234=>"000010001",
        6235=>"111110110",
        6236=>"101101001",
        6237=>"001010100",
        6238=>"001100001",
        6239=>"111111111",
        6240=>"011011001",
        6241=>"001100110",
        6242=>"111111000",
        6243=>"110111000",
        6244=>"010010010",
        6245=>"000110111",
        6246=>"001000100",
        6247=>"110010100",
        6248=>"000000001",
        6249=>"000000010",
        6250=>"100101001",
        6251=>"111000111",
        6252=>"000101001",
        6253=>"000000110",
        6254=>"100110101",
        6255=>"001101101",
        6256=>"000010100",
        6257=>"000010110",
        6258=>"011000000",
        6259=>"101111100",
        6260=>"110010010",
        6261=>"000000000",
        6262=>"100100010",
        6263=>"101001011",
        6264=>"011010110",
        6265=>"010000000",
        6266=>"000000000",
        6267=>"000101101",
        6268=>"011000000",
        6269=>"111110110",
        6270=>"000010110",
        6271=>"010011011",
        6272=>"100100110",
        6273=>"011010000",
        6274=>"111100000",
        6275=>"101011001",
        6276=>"100110100",
        6277=>"111111000",
        6278=>"110110100",
        6279=>"000001110",
        6280=>"110010111",
        6281=>"000000001",
        6282=>"011011001",
        6283=>"100001001",
        6284=>"110000001",
        6285=>"111100010",
        6286=>"110100000",
        6287=>"001001000",
        6288=>"000111001",
        6289=>"001001001",
        6290=>"010110101",
        6291=>"111000000",
        6292=>"000100101",
        6293=>"011100000",
        6294=>"100000000",
        6295=>"001011111",
        6296=>"111110100",
        6297=>"001000000",
        6298=>"110110000",
        6299=>"110000100",
        6300=>"011011110",
        6301=>"010010000",
        6302=>"011100001",
        6303=>"001011110",
        6304=>"000001000",
        6305=>"011000000",
        6306=>"110111111",
        6307=>"000011011",
        6308=>"110110011",
        6309=>"000011011",
        6310=>"001011110",
        6311=>"110100000",
        6312=>"001011011",
        6313=>"001001000",
        6314=>"010111110",
        6315=>"110110000",
        6316=>"000111111",
        6317=>"001001011",
        6318=>"000000000",
        6319=>"101101000",
        6320=>"100011111",
        6321=>"000100100",
        6322=>"000010111",
        6323=>"110100110",
        6324=>"010000111",
        6325=>"001001001",
        6326=>"000001011",
        6327=>"000100100",
        6328=>"001001011",
        6329=>"010001110",
        6330=>"110101011",
        6331=>"000000000",
        6332=>"000010000",
        6333=>"000000000",
        6334=>"011111110",
        6335=>"110101100",
        6336=>"011001101",
        6337=>"011011100",
        6338=>"001001011",
        6339=>"011111100",
        6340=>"111111111",
        6341=>"110100100",
        6342=>"000100111",
        6343=>"001011010",
        6344=>"001001001",
        6345=>"000000000",
        6346=>"001011111",
        6347=>"000110100",
        6348=>"001001111",
        6349=>"111110111",
        6350=>"001011111",
        6351=>"100100110",
        6352=>"001001010",
        6353=>"110100101",
        6354=>"000000111",
        6355=>"110100000",
        6356=>"100110111",
        6357=>"001101110",
        6358=>"100110110",
        6359=>"100110110",
        6360=>"011110101",
        6361=>"100000010",
        6362=>"111111100",
        6363=>"001000000",
        6364=>"110100000",
        6365=>"101111111",
        6366=>"011111100",
        6367=>"100000011",
        6368=>"000111110",
        6369=>"001000110",
        6370=>"101111111",
        6371=>"011010000",
        6372=>"001011010",
        6373=>"010000000",
        6374=>"000100000",
        6375=>"000001011",
        6376=>"110011011",
        6377=>"000000000",
        6378=>"011110000",
        6379=>"000001110",
        6380=>"010100000",
        6381=>"100100011",
        6382=>"011010000",
        6383=>"100111110",
        6384=>"101100111",
        6385=>"100000110",
        6386=>"110100000",
        6387=>"000010001",
        6388=>"111101110",
        6389=>"011101001",
        6390=>"001001001",
        6391=>"000000000",
        6392=>"000111111",
        6393=>"011011011",
        6394=>"000001011",
        6395=>"000001011",
        6396=>"001110100",
        6397=>"001011110",
        6398=>"000110111",
        6399=>"000110110",
        6400=>"001111011",
        6401=>"000110000",
        6402=>"010011000",
        6403=>"111111111",
        6404=>"001110111",
        6405=>"100000000",
        6406=>"000000000",
        6407=>"011111111",
        6408=>"111111110",
        6409=>"000000000",
        6410=>"001000001",
        6411=>"000110111",
        6412=>"111111000",
        6413=>"010010111",
        6414=>"111110110",
        6415=>"000110000",
        6416=>"000110110",
        6417=>"000000000",
        6418=>"110110011",
        6419=>"100111110",
        6420=>"110100100",
        6421=>"000010000",
        6422=>"000000000",
        6423=>"001000000",
        6424=>"111001101",
        6425=>"000101110",
        6426=>"011011001",
        6427=>"100110000",
        6428=>"000000001",
        6429=>"000001010",
        6430=>"110110110",
        6431=>"111111111",
        6432=>"111111110",
        6433=>"011010000",
        6434=>"000010011",
        6435=>"101000000",
        6436=>"000100111",
        6437=>"000110110",
        6438=>"111011000",
        6439=>"000000000",
        6440=>"000000101",
        6441=>"111001101",
        6442=>"001011111",
        6443=>"110110110",
        6444=>"000000100",
        6445=>"000010001",
        6446=>"111111000",
        6447=>"000110110",
        6448=>"000100100",
        6449=>"110110110",
        6450=>"010111111",
        6451=>"100100100",
        6452=>"000011000",
        6453=>"000000000",
        6454=>"110000000",
        6455=>"111111110",
        6456=>"000000000",
        6457=>"011001000",
        6458=>"000000000",
        6459=>"011000000",
        6460=>"000000000",
        6461=>"101001101",
        6462=>"011011000",
        6463=>"111001001",
        6464=>"000000000",
        6465=>"000010000",
        6466=>"111110101",
        6467=>"000001101",
        6468=>"000000110",
        6469=>"110100111",
        6470=>"000000000",
        6471=>"000000001",
        6472=>"000000001",
        6473=>"100100111",
        6474=>"111001001",
        6475=>"000000000",
        6476=>"000000000",
        6477=>"101001101",
        6478=>"000000100",
        6479=>"000000000",
        6480=>"011010111",
        6481=>"000100000",
        6482=>"101101000",
        6483=>"111111111",
        6484=>"111001111",
        6485=>"111111100",
        6486=>"000000001",
        6487=>"001100000",
        6488=>"011001111",
        6489=>"010111111",
        6490=>"110111101",
        6491=>"000000000",
        6492=>"001011011",
        6493=>"000010000",
        6494=>"111111111",
        6495=>"011110111",
        6496=>"000110010",
        6497=>"111000001",
        6498=>"010000000",
        6499=>"110111111",
        6500=>"100101001",
        6501=>"000111000",
        6502=>"011101010",
        6503=>"010000000",
        6504=>"101100101",
        6505=>"010111111",
        6506=>"110110100",
        6507=>"000111100",
        6508=>"111111101",
        6509=>"111111101",
        6510=>"110110110",
        6511=>"111011111",
        6512=>"011010011",
        6513=>"111111101",
        6514=>"101111111",
        6515=>"011111011",
        6516=>"000101111",
        6517=>"000100110",
        6518=>"000001000",
        6519=>"010010111",
        6520=>"000100111",
        6521=>"110101111",
        6522=>"001011100",
        6523=>"111111111",
        6524=>"101001101",
        6525=>"000100000",
        6526=>"001000111",
        6527=>"101111111",
        6528=>"011010011",
        6529=>"011100111",
        6530=>"100111111",
        6531=>"100100100",
        6532=>"110111011",
        6533=>"000000000",
        6534=>"111011011",
        6535=>"100110111",
        6536=>"100011001",
        6537=>"011011111",
        6538=>"100101110",
        6539=>"000100111",
        6540=>"101001001",
        6541=>"000010000",
        6542=>"000000000",
        6543=>"000100100",
        6544=>"011011000",
        6545=>"110100111",
        6546=>"110110111",
        6547=>"000110000",
        6548=>"011001001",
        6549=>"000010010",
        6550=>"000000000",
        6551=>"001011011",
        6552=>"110111010",
        6553=>"000000000",
        6554=>"110110010",
        6555=>"000001000",
        6556=>"110111111",
        6557=>"010010000",
        6558=>"110010001",
        6559=>"101111111",
        6560=>"100110010",
        6561=>"001011001",
        6562=>"100100110",
        6563=>"001011011",
        6564=>"001000010",
        6565=>"011111101",
        6566=>"011011000",
        6567=>"011011001",
        6568=>"000110110",
        6569=>"000000001",
        6570=>"100000000",
        6571=>"000110011",
        6572=>"111011011",
        6573=>"011011001",
        6574=>"101011001",
        6575=>"100110110",
        6576=>"001001000",
        6577=>"000110111",
        6578=>"101111001",
        6579=>"000001000",
        6580=>"111110000",
        6581=>"011011001",
        6582=>"001000100",
        6583=>"111011110",
        6584=>"000000110",
        6585=>"111111011",
        6586=>"000000100",
        6587=>"011101111",
        6588=>"110110110",
        6589=>"000000001",
        6590=>"100111111",
        6591=>"100000000",
        6592=>"000000100",
        6593=>"001011111",
        6594=>"001000000",
        6595=>"000001000",
        6596=>"110011001",
        6597=>"101001011",
        6598=>"011111000",
        6599=>"001001001",
        6600=>"001000000",
        6601=>"111010000",
        6602=>"110111011",
        6603=>"000000000",
        6604=>"100100111",
        6605=>"111011101",
        6606=>"100001000",
        6607=>"001101100",
        6608=>"001001001",
        6609=>"000100110",
        6610=>"110011001",
        6611=>"000111000",
        6612=>"111001000",
        6613=>"011101100",
        6614=>"011010000",
        6615=>"111011001",
        6616=>"100110100",
        6617=>"001000000",
        6618=>"100101000",
        6619=>"111111100",
        6620=>"100010000",
        6621=>"000110011",
        6622=>"100100100",
        6623=>"000111111",
        6624=>"011000000",
        6625=>"111110111",
        6626=>"010001101",
        6627=>"110110111",
        6628=>"000011001",
        6629=>"010110100",
        6630=>"100000001",
        6631=>"000010001",
        6632=>"000100110",
        6633=>"100100110",
        6634=>"110010000",
        6635=>"101100000",
        6636=>"100100110",
        6637=>"000111110",
        6638=>"111010000",
        6639=>"110111111",
        6640=>"001100110",
        6641=>"000000111",
        6642=>"011101001",
        6643=>"100100110",
        6644=>"000111000",
        6645=>"010001101",
        6646=>"000001001",
        6647=>"000001000",
        6648=>"110111011",
        6649=>"000000011",
        6650=>"011001000",
        6651=>"000111011",
        6652=>"111111111",
        6653=>"111111011",
        6654=>"001110110",
        6655=>"100000000",
        6656=>"100000000",
        6657=>"001011000",
        6658=>"001001001",
        6659=>"000101100",
        6660=>"100110000",
        6661=>"100100110",
        6662=>"110010110",
        6663=>"011011011",
        6664=>"100100100",
        6665=>"010011100",
        6666=>"111001011",
        6667=>"001011111",
        6668=>"011011011",
        6669=>"001100001",
        6670=>"100110010",
        6671=>"011001001",
        6672=>"001001011",
        6673=>"000001000",
        6674=>"100100000",
        6675=>"001001001",
        6676=>"100110100",
        6677=>"011011001",
        6678=>"011011011",
        6679=>"011110100",
        6680=>"000100110",
        6681=>"010000110",
        6682=>"001001001",
        6683=>"100010110",
        6684=>"100100100",
        6685=>"100100000",
        6686=>"110110100",
        6687=>"100110000",
        6688=>"000001011",
        6689=>"100000010",
        6690=>"001110110",
        6691=>"100100000",
        6692=>"100100110",
        6693=>"111111100",
        6694=>"001001101",
        6695=>"011110011",
        6696=>"101010000",
        6697=>"100100011",
        6698=>"001001000",
        6699=>"100110000",
        6700=>"011101111",
        6701=>"110111011",
        6702=>"100100110",
        6703=>"111001001",
        6704=>"001011110",
        6705=>"011001011",
        6706=>"100000111",
        6707=>"010110100",
        6708=>"001101101",
        6709=>"000000000",
        6710=>"110011011",
        6711=>"110100100",
        6712=>"011011111",
        6713=>"100110100",
        6714=>"110110110",
        6715=>"000011111",
        6716=>"001011011",
        6717=>"100100110",
        6718=>"000000011",
        6719=>"100100000",
        6720=>"100000000",
        6721=>"011011010",
        6722=>"101100100",
        6723=>"110100000",
        6724=>"110110110",
        6725=>"101100000",
        6726=>"100100100",
        6727=>"011011110",
        6728=>"011011011",
        6729=>"100100100",
        6730=>"101101100",
        6731=>"001001001",
        6732=>"001011011",
        6733=>"110100100",
        6734=>"100110100",
        6735=>"010001101",
        6736=>"001011001",
        6737=>"011011001",
        6738=>"000100110",
        6739=>"110111110",
        6740=>"000101101",
        6741=>"011011011",
        6742=>"110010100",
        6743=>"001000000",
        6744=>"110110111",
        6745=>"100010100",
        6746=>"001111001",
        6747=>"100100100",
        6748=>"000000000",
        6749=>"000001111",
        6750=>"000000100",
        6751=>"111001000",
        6752=>"111111110",
        6753=>"011000100",
        6754=>"001111111",
        6755=>"100100100",
        6756=>"011011110",
        6757=>"011011001",
        6758=>"011001001",
        6759=>"111011111",
        6760=>"011011011",
        6761=>"010000000",
        6762=>"100100100",
        6763=>"110000011",
        6764=>"100001001",
        6765=>"100001001",
        6766=>"100100100",
        6767=>"000000000",
        6768=>"101001011",
        6769=>"110010110",
        6770=>"001011011",
        6771=>"011000100",
        6772=>"100100110",
        6773=>"001001011",
        6774=>"010011010",
        6775=>"110000101",
        6776=>"111001011",
        6777=>"011011011",
        6778=>"001011011",
        6779=>"011011001",
        6780=>"101001101",
        6781=>"000010110",
        6782=>"100100000",
        6783=>"100110100",
        6784=>"001100100",
        6785=>"111000101",
        6786=>"000001111",
        6787=>"110111111",
        6788=>"000001100",
        6789=>"000010010",
        6790=>"000110110",
        6791=>"101001001",
        6792=>"000000001",
        6793=>"110000000",
        6794=>"010000000",
        6795=>"001011001",
        6796=>"011001000",
        6797=>"111000001",
        6798=>"100110011",
        6799=>"001100110",
        6800=>"101111110",
        6801=>"111000111",
        6802=>"111111101",
        6803=>"000100001",
        6804=>"000010111",
        6805=>"001000000",
        6806=>"101000000",
        6807=>"100000110",
        6808=>"110001000",
        6809=>"011100001",
        6810=>"111101101",
        6811=>"011000100",
        6812=>"000000111",
        6813=>"100100001",
        6814=>"000010110",
        6815=>"011011100",
        6816=>"111101100",
        6817=>"100100100",
        6818=>"110011001",
        6819=>"001001101",
        6820=>"011111011",
        6821=>"111111111",
        6822=>"011111111",
        6823=>"000100110",
        6824=>"110010001",
        6825=>"100101111",
        6826=>"010100000",
        6827=>"111110001",
        6828=>"111111000",
        6829=>"011110100",
        6830=>"110000000",
        6831=>"111111111",
        6832=>"010001010",
        6833=>"111010000",
        6834=>"111001100",
        6835=>"101100010",
        6836=>"011001001",
        6837=>"111110010",
        6838=>"111100000",
        6839=>"000000110",
        6840=>"000000000",
        6841=>"100000110",
        6842=>"000110000",
        6843=>"111111111",
        6844=>"111101001",
        6845=>"101010010",
        6846=>"000000001",
        6847=>"010110100",
        6848=>"000000101",
        6849=>"000011111",
        6850=>"110000000",
        6851=>"111001001",
        6852=>"001111111",
        6853=>"111111111",
        6854=>"000000000",
        6855=>"100000001",
        6856=>"100111111",
        6857=>"111001001",
        6858=>"110101111",
        6859=>"111101001",
        6860=>"100110101",
        6861=>"101000000",
        6862=>"110111111",
        6863=>"000001111",
        6864=>"111001001",
        6865=>"111101001",
        6866=>"110000000",
        6867=>"000111111",
        6868=>"101111111",
        6869=>"001000000",
        6870=>"101001000",
        6871=>"000110110",
        6872=>"010111111",
        6873=>"111000110",
        6874=>"111011011",
        6875=>"010000110",
        6876=>"100110111",
        6877=>"001010110",
        6878=>"110011111",
        6879=>"000000010",
        6880=>"000011011",
        6881=>"100001101",
        6882=>"111001001",
        6883=>"111001101",
        6884=>"000000101",
        6885=>"010101101",
        6886=>"111001101",
        6887=>"111010101",
        6888=>"011000011",
        6889=>"000000011",
        6890=>"110110111",
        6891=>"010110000",
        6892=>"000000101",
        6893=>"011000000",
        6894=>"100110100",
        6895=>"000000100",
        6896=>"000110110",
        6897=>"111010101",
        6898=>"111110110",
        6899=>"000000000",
        6900=>"111000000",
        6901=>"000010101",
        6902=>"111000000",
        6903=>"111001011",
        6904=>"000011001",
        6905=>"111110101",
        6906=>"110111101",
        6907=>"000001000",
        6908=>"001101111",
        6909=>"101101011",
        6910=>"111001000",
        6911=>"100100111",
        6912=>"101001101",
        6913=>"000011000",
        6914=>"001111111",
        6915=>"111001001",
        6916=>"011000100",
        6917=>"110000000",
        6918=>"111110001",
        6919=>"001101000",
        6920=>"110001011",
        6921=>"101011000",
        6922=>"001000110",
        6923=>"000001100",
        6924=>"000000100",
        6925=>"111111000",
        6926=>"110001001",
        6927=>"000110111",
        6928=>"001100110",
        6929=>"000001000",
        6930=>"011011001",
        6931=>"000011011",
        6932=>"001010001",
        6933=>"110000000",
        6934=>"000011110",
        6935=>"110100000",
        6936=>"000001010",
        6937=>"001001010",
        6938=>"000001011",
        6939=>"011110011",
        6940=>"100000000",
        6941=>"110010000",
        6942=>"111000000",
        6943=>"111111100",
        6944=>"010111111",
        6945=>"101111111",
        6946=>"001111111",
        6947=>"001100001",
        6948=>"011110000",
        6949=>"000100000",
        6950=>"001111111",
        6951=>"011111111",
        6952=>"001001011",
        6953=>"000100000",
        6954=>"001100001",
        6955=>"101101001",
        6956=>"011111110",
        6957=>"100000000",
        6958=>"110000000",
        6959=>"100000011",
        6960=>"001101101",
        6961=>"001001001",
        6962=>"110111010",
        6963=>"101000000",
        6964=>"111001011",
        6965=>"100000000",
        6966=>"100110110",
        6967=>"001001000",
        6968=>"110110110",
        6969=>"110100100",
        6970=>"110001000",
        6971=>"000001011",
        6972=>"000000000",
        6973=>"000110011",
        6974=>"100001110",
        6975=>"111000100",
        6976=>"000001111",
        6977=>"001001001",
        6978=>"100000110",
        6979=>"110100001",
        6980=>"000010010",
        6981=>"000011111",
        6982=>"111100111",
        6983=>"000110110",
        6984=>"100011011",
        6985=>"111101000",
        6986=>"011000110",
        6987=>"001011011",
        6988=>"000111001",
        6989=>"001010110",
        6990=>"010110111",
        6991=>"001011111",
        6992=>"001011111",
        6993=>"000011110",
        6994=>"111000000",
        6995=>"111100000",
        6996=>"011111011",
        6997=>"000001111",
        6998=>"110110001",
        6999=>"110100000",
        7000=>"001111111",
        7001=>"100010010",
        7002=>"000000001",
        7003=>"001011111",
        7004=>"010010110",
        7005=>"111000100",
        7006=>"000010111",
        7007=>"001000110",
        7008=>"110010000",
        7009=>"000000001",
        7010=>"111111111",
        7011=>"000000111",
        7012=>"111001111",
        7013=>"100110000",
        7014=>"011101101",
        7015=>"110110100",
        7016=>"000001110",
        7017=>"001000101",
        7018=>"100001010",
        7019=>"100000000",
        7020=>"001011111",
        7021=>"101111111",
        7022=>"100110000",
        7023=>"110100000",
        7024=>"000011011",
        7025=>"011111110",
        7026=>"100111100",
        7027=>"100001000",
        7028=>"001100111",
        7029=>"111100011",
        7030=>"100011011",
        7031=>"111111100",
        7032=>"000111111",
        7033=>"100100000",
        7034=>"001111110",
        7035=>"000111111",
        7036=>"000000100",
        7037=>"000000000",
        7038=>"000011111",
        7039=>"011001001",
        7040=>"010111110",
        7041=>"111000000",
        7042=>"110010101",
        7043=>"000010011",
        7044=>"001101100",
        7045=>"100110111",
        7046=>"100110001",
        7047=>"000000010",
        7048=>"111011000",
        7049=>"111110100",
        7050=>"000100000",
        7051=>"011011001",
        7052=>"001000000",
        7053=>"010111110",
        7054=>"000000000",
        7055=>"000000011",
        7056=>"011000100",
        7057=>"101001001",
        7058=>"101110010",
        7059=>"100100000",
        7060=>"000111001",
        7061=>"000000000",
        7062=>"000000000",
        7063=>"011000010",
        7064=>"011011001",
        7065=>"110100001",
        7066=>"011101101",
        7067=>"001000001",
        7068=>"110111111",
        7069=>"000110101",
        7070=>"000001101",
        7071=>"010110110",
        7072=>"111000000",
        7073=>"110111101",
        7074=>"011111100",
        7075=>"011101001",
        7076=>"111011001",
        7077=>"001010000",
        7078=>"000111110",
        7079=>"001101001",
        7080=>"001100100",
        7081=>"110100001",
        7082=>"000000101",
        7083=>"100100011",
        7084=>"011000111",
        7085=>"010111010",
        7086=>"101000111",
        7087=>"111001011",
        7088=>"110000000",
        7089=>"001000000",
        7090=>"001000100",
        7091=>"001010011",
        7092=>"011001101",
        7093=>"000101000",
        7094=>"110000010",
        7095=>"000110010",
        7096=>"110010011",
        7097=>"001001111",
        7098=>"111011001",
        7099=>"111110010",
        7100=>"101000000",
        7101=>"000000110",
        7102=>"000000101",
        7103=>"000111100",
        7104=>"000101000",
        7105=>"000100010",
        7106=>"111110000",
        7107=>"001110110",
        7108=>"001000000",
        7109=>"011110100",
        7110=>"000110111",
        7111=>"110000010",
        7112=>"110000001",
        7113=>"001001101",
        7114=>"111011100",
        7115=>"000000001",
        7116=>"001010000",
        7117=>"000100111",
        7118=>"000010010",
        7119=>"111101111",
        7120=>"000011000",
        7121=>"000000001",
        7122=>"000000111",
        7123=>"111010111",
        7124=>"000010011",
        7125=>"110010000",
        7126=>"000000111",
        7127=>"101111111",
        7128=>"011011100",
        7129=>"111010000",
        7130=>"111001011",
        7131=>"000000001",
        7132=>"001011011",
        7133=>"011011100",
        7134=>"001101111",
        7135=>"000000111",
        7136=>"000100110",
        7137=>"100000001",
        7138=>"000001000",
        7139=>"110111000",
        7140=>"010010111",
        7141=>"101000111",
        7142=>"000000100",
        7143=>"111000011",
        7144=>"010010000",
        7145=>"100100100",
        7146=>"000100100",
        7147=>"000010111",
        7148=>"001000000",
        7149=>"001001101",
        7150=>"000011111",
        7151=>"000000000",
        7152=>"110010000",
        7153=>"001000010",
        7154=>"101101001",
        7155=>"011110100",
        7156=>"111000101",
        7157=>"000000010",
        7158=>"110000000",
        7159=>"000000001",
        7160=>"011111110",
        7161=>"110010010",
        7162=>"100000000",
        7163=>"000000111",
        7164=>"000111100",
        7165=>"011000000",
        7166=>"111101101",
        7167=>"100111111",
        7168=>"111011011",
        7169=>"001010000",
        7170=>"011111011",
        7171=>"111110101",
        7172=>"111110000",
        7173=>"100101101",
        7174=>"011111100",
        7175=>"000001001",
        7176=>"010000110",
        7177=>"000000001",
        7178=>"000011010",
        7179=>"000011011",
        7180=>"100100110",
        7181=>"111100000",
        7182=>"100100111",
        7183=>"000101111",
        7184=>"111000000",
        7185=>"011111010",
        7186=>"011010010",
        7187=>"000011111",
        7188=>"011010011",
        7189=>"111001100",
        7190=>"111011011",
        7191=>"001000001",
        7192=>"110000010",
        7193=>"000000100",
        7194=>"111111000",
        7195=>"111111111",
        7196=>"111111111",
        7197=>"110111110",
        7198=>"010111100",
        7199=>"000001001",
        7200=>"110100010",
        7201=>"000000000",
        7202=>"111100000",
        7203=>"000000100",
        7204=>"100000000",
        7205=>"111100001",
        7206=>"111111101",
        7207=>"110110000",
        7208=>"111100001",
        7209=>"001011111",
        7210=>"000000000",
        7211=>"100100010",
        7212=>"110000001",
        7213=>"010010010",
        7214=>"010000010",
        7215=>"111011011",
        7216=>"111001010",
        7217=>"111000000",
        7218=>"000000111",
        7219=>"111001111",
        7220=>"110011111",
        7221=>"001000000",
        7222=>"001000000",
        7223=>"100110100",
        7224=>"011011001",
        7225=>"111000000",
        7226=>"111111100",
        7227=>"100101111",
        7228=>"101011011",
        7229=>"000000100",
        7230=>"000000001",
        7231=>"100110000",
        7232=>"111101110",
        7233=>"000100101",
        7234=>"111001101",
        7235=>"100000001",
        7236=>"100100010",
        7237=>"100101111",
        7238=>"110010110",
        7239=>"011000001",
        7240=>"000000111",
        7241=>"010111000",
        7242=>"010000000",
        7243=>"000000000",
        7244=>"110100101",
        7245=>"000100100",
        7246=>"110110011",
        7247=>"000000101",
        7248=>"011000000",
        7249=>"000110111",
        7250=>"100000100",
        7251=>"010010111",
        7252=>"011010000",
        7253=>"101001001",
        7254=>"110010000",
        7255=>"000101001",
        7256=>"110110100",
        7257=>"001101010",
        7258=>"000111111",
        7259=>"011010011",
        7260=>"000011111",
        7261=>"111110000",
        7262=>"001011011",
        7263=>"001110111",
        7264=>"010110001",
        7265=>"100001100",
        7266=>"011111111",
        7267=>"110110011",
        7268=>"100000101",
        7269=>"000000100",
        7270=>"111100000",
        7271=>"100000011",
        7272=>"111100000",
        7273=>"000100110",
        7274=>"101010110",
        7275=>"000000110",
        7276=>"000111101",
        7277=>"100100111",
        7278=>"110100111",
        7279=>"010111110",
        7280=>"101000111",
        7281=>"100110111",
        7282=>"111010000",
        7283=>"011000010",
        7284=>"011000111",
        7285=>"000101000",
        7286=>"010011111",
        7287=>"111101000",
        7288=>"111100000",
        7289=>"101001001",
        7290=>"000010110",
        7291=>"110001001",
        7292=>"111111000",
        7293=>"000000111",
        7294=>"010110101",
        7295=>"000111111",
        7296=>"111110101",
        7297=>"001011011",
        7298=>"110100110",
        7299=>"110110001",
        7300=>"101111001",
        7301=>"111100101",
        7302=>"110110100",
        7303=>"011011001",
        7304=>"000000000",
        7305=>"111110100",
        7306=>"011000011",
        7307=>"010110010",
        7308=>"110100100",
        7309=>"001000001",
        7310=>"100000100",
        7311=>"011001001",
        7312=>"110110100",
        7313=>"001010110",
        7314=>"101100000",
        7315=>"110000010",
        7316=>"100100010",
        7317=>"111100110",
        7318=>"000100100",
        7319=>"011011001",
        7320=>"100100000",
        7321=>"111001110",
        7322=>"110000011",
        7323=>"110110000",
        7324=>"000010010",
        7325=>"110100101",
        7326=>"110100000",
        7327=>"011111011",
        7328=>"100001011",
        7329=>"100101010",
        7330=>"111000000",
        7331=>"110111110",
        7332=>"111011011",
        7333=>"100110101",
        7334=>"111111001",
        7335=>"100100110",
        7336=>"110111000",
        7337=>"100110011",
        7338=>"100100110",
        7339=>"100100100",
        7340=>"111111100",
        7341=>"000111111",
        7342=>"100110110",
        7343=>"100111111",
        7344=>"000110110",
        7345=>"100111110",
        7346=>"110110110",
        7347=>"110100000",
        7348=>"100000000",
        7349=>"100100000",
        7350=>"000001000",
        7351=>"100101111",
        7352=>"000000000",
        7353=>"100110100",
        7354=>"001001011",
        7355=>"011000000",
        7356=>"110111111",
        7357=>"100000100",
        7358=>"111100111",
        7359=>"011011001",
        7360=>"000000000",
        7361=>"110000011",
        7362=>"111111000",
        7363=>"000011000",
        7364=>"110110100",
        7365=>"101110100",
        7366=>"000000000",
        7367=>"011011001",
        7368=>"000001111",
        7369=>"100100011",
        7370=>"010111011",
        7371=>"100100100",
        7372=>"011000011",
        7373=>"110001000",
        7374=>"111011000",
        7375=>"100100110",
        7376=>"010010010",
        7377=>"110100110",
        7378=>"000100110",
        7379=>"000100111",
        7380=>"100100000",
        7381=>"010010010",
        7382=>"100110000",
        7383=>"111101011",
        7384=>"110100000",
        7385=>"011000011",
        7386=>"001001001",
        7387=>"010110110",
        7388=>"000000000",
        7389=>"000110110",
        7390=>"000100000",
        7391=>"010000110",
        7392=>"111111111",
        7393=>"100110100",
        7394=>"010011010",
        7395=>"100110110",
        7396=>"111111010",
        7397=>"110100100",
        7398=>"110100000",
        7399=>"110101110",
        7400=>"111001000",
        7401=>"010010111",
        7402=>"100000100",
        7403=>"000110001",
        7404=>"110100001",
        7405=>"001011101",
        7406=>"100100000",
        7407=>"111100000",
        7408=>"110110100",
        7409=>"110111111",
        7410=>"000000111",
        7411=>"000100100",
        7412=>"011001111",
        7413=>"101001000",
        7414=>"000001010",
        7415=>"110100100",
        7416=>"110011000",
        7417=>"001011011",
        7418=>"010110111",
        7419=>"011011011",
        7420=>"111111111",
        7421=>"000000000",
        7422=>"011010001",
        7423=>"001001000",
        7424=>"011000110",
        7425=>"000000111",
        7426=>"011101101",
        7427=>"011111101",
        7428=>"010000000",
        7429=>"010111000",
        7430=>"001111111",
        7431=>"111000000",
        7432=>"001110000",
        7433=>"111111101",
        7434=>"010000110",
        7435=>"100100110",
        7436=>"111000000",
        7437=>"010100111",
        7438=>"110101001",
        7439=>"011000101",
        7440=>"111111000",
        7441=>"000111111",
        7442=>"111111101",
        7443=>"000000011",
        7444=>"001011111",
        7445=>"010000010",
        7446=>"000101000",
        7447=>"100000000",
        7448=>"111011111",
        7449=>"111001000",
        7450=>"001111111",
        7451=>"000000000",
        7452=>"110111111",
        7453=>"110000000",
        7454=>"110011111",
        7455=>"111111111",
        7456=>"111111000",
        7457=>"111111011",
        7458=>"111101000",
        7459=>"100000000",
        7460=>"111111000",
        7461=>"011000000",
        7462=>"000111001",
        7463=>"000111111",
        7464=>"110101101",
        7465=>"111010110",
        7466=>"001011111",
        7467=>"001101001",
        7468=>"100000000",
        7469=>"011011000",
        7470=>"111000000",
        7471=>"010101110",
        7472=>"010000111",
        7473=>"111100100",
        7474=>"100100100",
        7475=>"111110000",
        7476=>"111011000",
        7477=>"111000110",
        7478=>"010000101",
        7479=>"111111100",
        7480=>"000001101",
        7481=>"100000010",
        7482=>"111111111",
        7483=>"000000011",
        7484=>"000000111",
        7485=>"110100000",
        7486=>"000001000",
        7487=>"011010111",
        7488=>"100010010",
        7489=>"000111111",
        7490=>"111000111",
        7491=>"111111110",
        7492=>"110011000",
        7493=>"010011001",
        7494=>"111010010",
        7495=>"010000111",
        7496=>"111011000",
        7497=>"000010111",
        7498=>"111010000",
        7499=>"000100000",
        7500=>"010001000",
        7501=>"000010111",
        7502=>"110111110",
        7503=>"111010000",
        7504=>"100010010",
        7505=>"110100111",
        7506=>"111000010",
        7507=>"011001111",
        7508=>"000110110",
        7509=>"000000000",
        7510=>"111011111",
        7511=>"010111001",
        7512=>"101000001",
        7513=>"000100100",
        7514=>"000111011",
        7515=>"000000000",
        7516=>"111111010",
        7517=>"110100110",
        7518=>"000101111",
        7519=>"101111111",
        7520=>"111111000",
        7521=>"011000000",
        7522=>"000010111",
        7523=>"010000000",
        7524=>"000000000",
        7525=>"100000000",
        7526=>"110001000",
        7527=>"010000000",
        7528=>"001011111",
        7529=>"011101100",
        7530=>"110111001",
        7531=>"000000010",
        7532=>"000101000",
        7533=>"111001001",
        7534=>"111011110",
        7535=>"000001110",
        7536=>"111000000",
        7537=>"000000000",
        7538=>"000111111",
        7539=>"111000000",
        7540=>"001111110",
        7541=>"101000100",
        7542=>"000000001",
        7543=>"001001001",
        7544=>"111100111",
        7545=>"010000000",
        7546=>"110110101",
        7547=>"111000000",
        7548=>"000111111",
        7549=>"000000110",
        7550=>"111111010",
        7551=>"111010000",
        7552=>"000001111",
        7553=>"111111000",
        7554=>"111010000",
        7555=>"000001111",
        7556=>"001000000",
        7557=>"000111010",
        7558=>"000000111",
        7559=>"111000000",
        7560=>"000111000",
        7561=>"000001111",
        7562=>"011010000",
        7563=>"011100100",
        7564=>"111000000",
        7565=>"110110110",
        7566=>"100001011",
        7567=>"100000001",
        7568=>"111101101",
        7569=>"000100110",
        7570=>"000000100",
        7571=>"110000001",
        7572=>"000000111",
        7573=>"000000000",
        7574=>"000100000",
        7575=>"000000001",
        7576=>"000000001",
        7577=>"110101010",
        7578=>"111101110",
        7579=>"000111101",
        7580=>"000101010",
        7581=>"000000001",
        7582=>"100111111",
        7583=>"000001011",
        7584=>"111111111",
        7585=>"111001000",
        7586=>"011000000",
        7587=>"000000011",
        7588=>"001111111",
        7589=>"011111111",
        7590=>"111111000",
        7591=>"001000101",
        7592=>"110000010",
        7593=>"001010011",
        7594=>"111111011",
        7595=>"110000001",
        7596=>"001000111",
        7597=>"000000011",
        7598=>"000000001",
        7599=>"111000101",
        7600=>"111010011",
        7601=>"110000000",
        7602=>"011100110",
        7603=>"000001111",
        7604=>"100100100",
        7605=>"000111111",
        7606=>"011011000",
        7607=>"000110010",
        7608=>"010000101",
        7609=>"000000111",
        7610=>"100100111",
        7611=>"011011001",
        7612=>"000000111",
        7613=>"001111111",
        7614=>"001100110",
        7615=>"100101111",
        7616=>"100010100",
        7617=>"011000101",
        7618=>"101010111",
        7619=>"000000111",
        7620=>"100101111",
        7621=>"000110011",
        7622=>"101101110",
        7623=>"000000000",
        7624=>"110001000",
        7625=>"000000111",
        7626=>"010010111",
        7627=>"000000010",
        7628=>"111111010",
        7629=>"000000000",
        7630=>"001011010",
        7631=>"111010000",
        7632=>"111000100",
        7633=>"111011000",
        7634=>"111010000",
        7635=>"110101001",
        7636=>"000111110",
        7637=>"111110000",
        7638=>"000111101",
        7639=>"100110110",
        7640=>"110110111",
        7641=>"000111110",
        7642=>"111111011",
        7643=>"000000111",
        7644=>"011010000",
        7645=>"011000101",
        7646=>"111001001",
        7647=>"000001111",
        7648=>"100100110",
        7649=>"011011100",
        7650=>"010000010",
        7651=>"111000010",
        7652=>"111111110",
        7653=>"111000000",
        7654=>"111000000",
        7655=>"010000000",
        7656=>"110011111",
        7657=>"111000000",
        7658=>"001001110",
        7659=>"111111111",
        7660=>"000010000",
        7661=>"010000000",
        7662=>"000001100",
        7663=>"001101110",
        7664=>"000000010",
        7665=>"000000000",
        7666=>"111111000",
        7667=>"111011000",
        7668=>"000111111",
        7669=>"110100000",
        7670=>"000000000",
        7671=>"110010011",
        7672=>"110010110",
        7673=>"111000001",
        7674=>"111110100",
        7675=>"111011000",
        7676=>"111111111",
        7677=>"001010111",
        7678=>"010000101",
        7679=>"100111111",
        7680=>"010110110",
        7681=>"110010000",
        7682=>"101100000",
        7683=>"100101110",
        7684=>"101101000",
        7685=>"010001111",
        7686=>"110011010",
        7687=>"101001010",
        7688=>"000100101",
        7689=>"000111111",
        7690=>"010110101",
        7691=>"000011011",
        7692=>"000001000",
        7693=>"010010010",
        7694=>"011001111",
        7695=>"001000110",
        7696=>"100000001",
        7697=>"011001000",
        7698=>"110001111",
        7699=>"101100100",
        7700=>"010000010",
        7701=>"110001111",
        7702=>"101100000",
        7703=>"000000110",
        7704=>"111111100",
        7705=>"001100111",
        7706=>"101100001",
        7707=>"111110001",
        7708=>"100110110",
        7709=>"101101100",
        7710=>"011110100",
        7711=>"001000101",
        7712=>"000110111",
        7713=>"011110000",
        7714=>"000111101",
        7715=>"111001100",
        7716=>"000000011",
        7717=>"110010000",
        7718=>"101100000",
        7719=>"101101001",
        7720=>"001010101",
        7721=>"000000000",
        7722=>"101000000",
        7723=>"101101101",
        7724=>"000011000",
        7725=>"111001111",
        7726=>"000011010",
        7727=>"111101111",
        7728=>"010010111",
        7729=>"101101000",
        7730=>"101001101",
        7731=>"001000000",
        7732=>"100111001",
        7733=>"000001100",
        7734=>"010100000",
        7735=>"101001010",
        7736=>"000000000",
        7737=>"010001001",
        7738=>"100110111",
        7739=>"000110010",
        7740=>"111101101",
        7741=>"101100101",
        7742=>"111011100",
        7743=>"011000000",
        7744=>"011111001",
        7745=>"111101101",
        7746=>"010000000",
        7747=>"000010111",
        7748=>"000101101",
        7749=>"111000100",
        7750=>"010010000",
        7751=>"110010010",
        7752=>"000000100",
        7753=>"010011000",
        7754=>"000011000",
        7755=>"101101100",
        7756=>"101111010",
        7757=>"010100000",
        7758=>"000111111",
        7759=>"000000111",
        7760=>"000000010",
        7761=>"001001000",
        7762=>"010011010",
        7763=>"100100000",
        7764=>"010010001",
        7765=>"101111111",
        7766=>"010010011",
        7767=>"000000111",
        7768=>"011100000",
        7769=>"000111111",
        7770=>"011001000",
        7771=>"010100101",
        7772=>"101101101",
        7773=>"100001011",
        7774=>"001001100",
        7775=>"111111101",
        7776=>"000000100",
        7777=>"001010000",
        7778=>"000110110",
        7779=>"000000000",
        7780=>"111111000",
        7781=>"000000000",
        7782=>"100100000",
        7783=>"101111000",
        7784=>"011000000",
        7785=>"100100101",
        7786=>"111101101",
        7787=>"000000010",
        7788=>"111000000",
        7789=>"001001001",
        7790=>"100110000",
        7791=>"111001101",
        7792=>"000101111",
        7793=>"111100001",
        7794=>"100000101",
        7795=>"101101000",
        7796=>"100111111",
        7797=>"000000000",
        7798=>"111011000",
        7799=>"101100100",
        7800=>"000000011",
        7801=>"010111010",
        7802=>"111001100",
        7803=>"001000000",
        7804=>"100000101",
        7805=>"111111110",
        7806=>"010100110",
        7807=>"001111101",
        7808=>"111111110",
        7809=>"111000000",
        7810=>"000110010",
        7811=>"010110010",
        7812=>"010110110",
        7813=>"011101110",
        7814=>"111111011",
        7815=>"000001001",
        7816=>"010110110",
        7817=>"000111111",
        7818=>"001000001",
        7819=>"011000000",
        7820=>"000000000",
        7821=>"110111010",
        7822=>"000000000",
        7823=>"000011001",
        7824=>"000110110",
        7825=>"011110010",
        7826=>"000000000",
        7827=>"110111111",
        7828=>"000011111",
        7829=>"000001000",
        7830=>"000000000",
        7831=>"000000110",
        7832=>"000110111",
        7833=>"100000011",
        7834=>"000100110",
        7835=>"111111111",
        7836=>"110111001",
        7837=>"100110110",
        7838=>"101111111",
        7839=>"111111111",
        7840=>"000000001",
        7841=>"000000001",
        7842=>"001100000",
        7843=>"000000000",
        7844=>"000100000",
        7845=>"000100101",
        7846=>"111000111",
        7847=>"010111111",
        7848=>"000000110",
        7849=>"010000110",
        7850=>"000000001",
        7851=>"011110110",
        7852=>"011001110",
        7853=>"010010110",
        7854=>"100111000",
        7855=>"011011010",
        7856=>"010110111",
        7857=>"000000000",
        7858=>"000000100",
        7859=>"000001011",
        7860=>"000010010",
        7861=>"000000111",
        7862=>"000000010",
        7863=>"000010010",
        7864=>"011000100",
        7865=>"100000101",
        7866=>"000100111",
        7867=>"000000111",
        7868=>"111011001",
        7869=>"101111111",
        7870=>"101101111",
        7871=>"011110001",
        7872=>"000111111",
        7873=>"000000000",
        7874=>"000000000",
        7875=>"000000000",
        7876=>"110111111",
        7877=>"001111111",
        7878=>"010011001",
        7879=>"110010000",
        7880=>"000101011",
        7881=>"000110000",
        7882=>"011011010",
        7883=>"000000000",
        7884=>"111110110",
        7885=>"000110000",
        7886=>"010011111",
        7887=>"000111111",
        7888=>"010110111",
        7889=>"000000001",
        7890=>"000000000",
        7891=>"001011111",
        7892=>"100111111",
        7893=>"000111011",
        7894=>"010011110",
        7895=>"010101010",
        7896=>"000000000",
        7897=>"000010010",
        7898=>"001001011",
        7899=>"010110010",
        7900=>"110111010",
        7901=>"001011100",
        7902=>"000000001",
        7903=>"000000000",
        7904=>"011111111",
        7905=>"010111110",
        7906=>"000111011",
        7907=>"010111000",
        7908=>"011111111",
        7909=>"111000000",
        7910=>"000000100",
        7911=>"110000010",
        7912=>"111000111",
        7913=>"000000000",
        7914=>"001111001",
        7915=>"010101111",
        7916=>"010111010",
        7917=>"010000000",
        7918=>"000000000",
        7919=>"000000010",
        7920=>"000111000",
        7921=>"000000000",
        7922=>"111101001",
        7923=>"000000000",
        7924=>"111011011",
        7925=>"001000001",
        7926=>"000000000",
        7927=>"000000000",
        7928=>"011011011",
        7929=>"000000000",
        7930=>"100001111",
        7931=>"010011011",
        7932=>"100100111",
        7933=>"111000000",
        7934=>"000000100",
        7935=>"100000101",
        7936=>"111001011",
        7937=>"001000100",
        7938=>"001000000",
        7939=>"111000011",
        7940=>"011001001",
        7941=>"100100100",
        7942=>"111011001",
        7943=>"101100011",
        7944=>"000000000",
        7945=>"000000100",
        7946=>"001001000",
        7947=>"011001000",
        7948=>"000000010",
        7949=>"111111011",
        7950=>"100011001",
        7951=>"100100111",
        7952=>"000011011",
        7953=>"001000000",
        7954=>"011001001",
        7955=>"100111111",
        7956=>"110111100",
        7957=>"100010100",
        7958=>"000111110",
        7959=>"110000001",
        7960=>"100111111",
        7961=>"000001011",
        7962=>"111001011",
        7963=>"111111010",
        7964=>"001100100",
        7965=>"000101101",
        7966=>"011000000",
        7967=>"110100110",
        7968=>"011000001",
        7969=>"110111111",
        7970=>"001001000",
        7971=>"000000001",
        7972=>"010000100",
        7973=>"110100100",
        7974=>"110110110",
        7975=>"100110111",
        7976=>"011000000",
        7977=>"000011111",
        7978=>"000000011",
        7979=>"000001000",
        7980=>"011000100",
        7981=>"100100000",
        7982=>"000010010",
        7983=>"011001011",
        7984=>"100111111",
        7985=>"001000000",
        7986=>"111100010",
        7987=>"000111111",
        7988=>"001001101",
        7989=>"101100000",
        7990=>"111001110",
        7991=>"111100110",
        7992=>"001000100",
        7993=>"011111111",
        7994=>"011101011",
        7995=>"001001000",
        7996=>"001100000",
        7997=>"100100100",
        7998=>"000100111",
        7999=>"110111111",
        8000=>"100000000",
        8001=>"001100100",
        8002=>"000000011",
        8003=>"000000000",
        8004=>"111001000",
        8005=>"111001001",
        8006=>"110100000",
        8007=>"001000100",
        8008=>"111101100",
        8009=>"101100010",
        8010=>"111000100",
        8011=>"101100100",
        8012=>"110100110",
        8013=>"111111011",
        8014=>"110110110",
        8015=>"110110010",
        8016=>"100110110",
        8017=>"100110000",
        8018=>"110100000",
        8019=>"100000000",
        8020=>"000110110",
        8021=>"110100000",
        8022=>"011110100",
        8023=>"110100100",
        8024=>"101101011",
        8025=>"001001101",
        8026=>"000000000",
        8027=>"100110010",
        8028=>"000011011",
        8029=>"111011101",
        8030=>"100000000",
        8031=>"001101011",
        8032=>"110111111",
        8033=>"111000000",
        8034=>"111011111",
        8035=>"001001001",
        8036=>"111100010",
        8037=>"110010011",
        8038=>"011000100",
        8039=>"000100100",
        8040=>"000100100",
        8041=>"001000000",
        8042=>"000001011",
        8043=>"110100100",
        8044=>"011011001",
        8045=>"111110111",
        8046=>"011100100",
        8047=>"011001001",
        8048=>"111011000",
        8049=>"110100101",
        8050=>"001100000",
        8051=>"000000000",
        8052=>"111110110",
        8053=>"000000000",
        8054=>"110000000",
        8055=>"001011111",
        8056=>"011111100",
        8057=>"100000011",
        8058=>"000001000",
        8059=>"011011011",
        8060=>"101100100",
        8061=>"001000000",
        8062=>"110011001",
        8063=>"110000000",
        8064=>"101000000",
        8065=>"000110110",
        8066=>"000000011",
        8067=>"111101111",
        8068=>"101001000",
        8069=>"000000010",
        8070=>"111010000",
        8071=>"000100111",
        8072=>"011100100",
        8073=>"100001100",
        8074=>"010001111",
        8075=>"100110001",
        8076=>"001011111",
        8077=>"110111110",
        8078=>"011000000",
        8079=>"000011111",
        8080=>"100100000",
        8081=>"110111111",
        8082=>"110101001",
        8083=>"001001010",
        8084=>"000111111",
        8085=>"101111111",
        8086=>"000000011",
        8087=>"111111111",
        8088=>"111111001",
        8089=>"011110100",
        8090=>"000000000",
        8091=>"100000001",
        8092=>"010110111",
        8093=>"111001000",
        8094=>"111111110",
        8095=>"000000000",
        8096=>"111101000",
        8097=>"000000000",
        8098=>"111000101",
        8099=>"111111101",
        8100=>"111000111",
        8101=>"010111000",
        8102=>"000000010",
        8103=>"111010010",
        8104=>"111111101",
        8105=>"110111101",
        8106=>"111001111",
        8107=>"110101000",
        8108=>"100111000",
        8109=>"001101101",
        8110=>"111101010",
        8111=>"111000010",
        8112=>"101100100",
        8113=>"000000010",
        8114=>"001100100",
        8115=>"000001011",
        8116=>"010100000",
        8117=>"101000000",
        8118=>"000011000",
        8119=>"000000000",
        8120=>"111111101",
        8121=>"111111001",
        8122=>"001111000",
        8123=>"000111111",
        8124=>"000000000",
        8125=>"111000000",
        8126=>"000000010",
        8127=>"110100100",
        8128=>"111110100",
        8129=>"011000000",
        8130=>"011001001",
        8131=>"001010111",
        8132=>"111110111",
        8133=>"111011011",
        8134=>"000000010",
        8135=>"010110000",
        8136=>"001011011",
        8137=>"111100000",
        8138=>"001101000",
        8139=>"000000111",
        8140=>"000110110",
        8141=>"010111000",
        8142=>"110111111",
        8143=>"000000111",
        8144=>"000010000",
        8145=>"111000110",
        8146=>"111000000",
        8147=>"000011011",
        8148=>"111100100",
        8149=>"000111111",
        8150=>"100000011",
        8151=>"000000000",
        8152=>"011001101",
        8153=>"010000110",
        8154=>"111001000",
        8155=>"000000111",
        8156=>"111101000",
        8157=>"001110011",
        8158=>"001000000",
        8159=>"011100000",
        8160=>"101000001",
        8161=>"011001100",
        8162=>"000000101",
        8163=>"000000100",
        8164=>"101000001",
        8165=>"000001000",
        8166=>"101100010",
        8167=>"111101101",
        8168=>"000111111",
        8169=>"000000010",
        8170=>"111001000",
        8171=>"111101111",
        8172=>"111000101",
        8173=>"000100010",
        8174=>"111111001",
        8175=>"110111011",
        8176=>"000000111",
        8177=>"010000110",
        8178=>"111000000",
        8179=>"110111110",
        8180=>"000010110",
        8181=>"000010110",
        8182=>"000000111",
        8183=>"100001001",
        8184=>"010011000",
        8185=>"000101001",
        8186=>"001110111",
        8187=>"000111100",
        8188=>"110000110",
        8189=>"110111100",
        8190=>"100110000",
        8191=>"111000000",
        8192=>"000000000",
        8193=>"010000000",
        8194=>"000011010",
        8195=>"111111111",
        8196=>"000001100",
        8197=>"010100101",
        8198=>"000000000",
        8199=>"001000101",
        8200=>"101110111",
        8201=>"111011011",
        8202=>"000001001",
        8203=>"110111100",
        8204=>"101111111",
        8205=>"010111000",
        8206=>"111110111",
        8207=>"110110011",
        8208=>"011011101",
        8209=>"111111111",
        8210=>"011001001",
        8211=>"100000000",
        8212=>"010110000",
        8213=>"000000010",
        8214=>"111100101",
        8215=>"111101010",
        8216=>"100011001",
        8217=>"110111001",
        8218=>"111100111",
        8219=>"111110111",
        8220=>"111101000",
        8221=>"100100100",
        8222=>"000111111",
        8223=>"000000000",
        8224=>"111111111",
        8225=>"000000000",
        8226=>"011011111",
        8227=>"000000000",
        8228=>"000000000",
        8229=>"010111000",
        8230=>"111111111",
        8231=>"111111101",
        8232=>"111001101",
        8233=>"111101011",
        8234=>"111011011",
        8235=>"100000001",
        8236=>"001000000",
        8237=>"000000000",
        8238=>"000000000",
        8239=>"110111111",
        8240=>"111000000",
        8241=>"000111100",
        8242=>"000110101",
        8243=>"100000001",
        8244=>"001001011",
        8245=>"000011110",
        8246=>"010000110",
        8247=>"000100111",
        8248=>"000000000",
        8249=>"010000111",
        8250=>"010101110",
        8251=>"110111000",
        8252=>"000000000",
        8253=>"000000000",
        8254=>"011111011",
        8255=>"110101000",
        8256=>"111110111",
        8257=>"000010111",
        8258=>"111000000",
        8259=>"101101000",
        8260=>"000000000",
        8261=>"000000000",
        8262=>"000000000",
        8263=>"110111111",
        8264=>"111111111",
        8265=>"000111101",
        8266=>"101000100",
        8267=>"111111111",
        8268=>"000000000",
        8269=>"000010000",
        8270=>"000000000",
        8271=>"010111111",
        8272=>"011011111",
        8273=>"111111111",
        8274=>"100000000",
        8275=>"010111011",
        8276=>"000000000",
        8277=>"111111001",
        8278=>"000000110",
        8279=>"001011011",
        8280=>"111111101",
        8281=>"111100110",
        8282=>"001111011",
        8283=>"100011100",
        8284=>"100000001",
        8285=>"011111111",
        8286=>"111111111",
        8287=>"000000000",
        8288=>"100010100",
        8289=>"001001000",
        8290=>"001000000",
        8291=>"000010010",
        8292=>"111101111",
        8293=>"101111110",
        8294=>"101111101",
        8295=>"111101001",
        8296=>"110110011",
        8297=>"000000101",
        8298=>"101000000",
        8299=>"110111111",
        8300=>"111110010",
        8301=>"101000000",
        8302=>"010110111",
        8303=>"111111111",
        8304=>"001111011",
        8305=>"010010011",
        8306=>"110110011",
        8307=>"111111110",
        8308=>"111111111",
        8309=>"110011100",
        8310=>"000000111",
        8311=>"110111111",
        8312=>"011000101",
        8313=>"111111111",
        8314=>"011110111",
        8315=>"011111111",
        8316=>"100110010",
        8317=>"111110001",
        8318=>"111111111",
        8319=>"111110111",
        8320=>"010010110",
        8321=>"110111110",
        8322=>"000000000",
        8323=>"110011111",
        8324=>"000100100",
        8325=>"111111111",
        8326=>"010110111",
        8327=>"111101101",
        8328=>"001100111",
        8329=>"110011111",
        8330=>"111111111",
        8331=>"011110110",
        8332=>"111111111",
        8333=>"010111110",
        8334=>"101111111",
        8335=>"111101001",
        8336=>"110110110",
        8337=>"010001000",
        8338=>"010000000",
        8339=>"010010010",
        8340=>"111111010",
        8341=>"110010000",
        8342=>"000000000",
        8343=>"111010110",
        8344=>"101011001",
        8345=>"111111010",
        8346=>"000100011",
        8347=>"110110001",
        8348=>"111110110",
        8349=>"111111000",
        8350=>"011011000",
        8351=>"000000000",
        8352=>"011000000",
        8353=>"110000000",
        8354=>"110101011",
        8355=>"000000111",
        8356=>"000000100",
        8357=>"111110000",
        8358=>"000111111",
        8359=>"010111111",
        8360=>"000111010",
        8361=>"110110111",
        8362=>"111111110",
        8363=>"110110100",
        8364=>"011000110",
        8365=>"111111110",
        8366=>"100000111",
        8367=>"110111110",
        8368=>"111011111",
        8369=>"000110001",
        8370=>"111111001",
        8371=>"000000000",
        8372=>"001011011",
        8373=>"011111011",
        8374=>"110000000",
        8375=>"101101111",
        8376=>"010010010",
        8377=>"011111010",
        8378=>"111111110",
        8379=>"000000000",
        8380=>"000111111",
        8381=>"000000000",
        8382=>"101010100",
        8383=>"000011000",
        8384=>"000000000",
        8385=>"100000000",
        8386=>"010111111",
        8387=>"111111111",
        8388=>"111011111",
        8389=>"011011111",
        8390=>"010000000",
        8391=>"110111111",
        8392=>"111011011",
        8393=>"000000001",
        8394=>"111001001",
        8395=>"111111111",
        8396=>"000000000",
        8397=>"000000000",
        8398=>"000000000",
        8399=>"110110110",
        8400=>"000000000",
        8401=>"110111111",
        8402=>"010000000",
        8403=>"111111111",
        8404=>"110110110",
        8405=>"101101111",
        8406=>"111111111",
        8407=>"000000010",
        8408=>"001011110",
        8409=>"000111111",
        8410=>"000100110",
        8411=>"000000000",
        8412=>"000001001",
        8413=>"011000100",
        8414=>"100110110",
        8415=>"010000010",
        8416=>"110111110",
        8417=>"000000000",
        8418=>"000000101",
        8419=>"110110110",
        8420=>"000001001",
        8421=>"111101111",
        8422=>"111110111",
        8423=>"000000000",
        8424=>"011111011",
        8425=>"111001001",
        8426=>"110001001",
        8427=>"111011101",
        8428=>"000000000",
        8429=>"110001001",
        8430=>"000000000",
        8431=>"101111111",
        8432=>"000000111",
        8433=>"000011000",
        8434=>"101111111",
        8435=>"111000011",
        8436=>"000011111",
        8437=>"111001101",
        8438=>"110010101",
        8439=>"001011000",
        8440=>"111000100",
        8441=>"111010100",
        8442=>"111111110",
        8443=>"111111000",
        8444=>"000111011",
        8445=>"111111010",
        8446=>"010010000",
        8447=>"100000000",
        8448=>"001111111",
        8449=>"111001001",
        8450=>"000011001",
        8451=>"010111111",
        8452=>"111001111",
        8453=>"000010011",
        8454=>"010111111",
        8455=>"000101001",
        8456=>"000110101",
        8457=>"001011011",
        8458=>"111000100",
        8459=>"001010010",
        8460=>"000000110",
        8461=>"111101010",
        8462=>"100100111",
        8463=>"111111100",
        8464=>"000110111",
        8465=>"010010110",
        8466=>"000000111",
        8467=>"100100111",
        8468=>"010110000",
        8469=>"000001011",
        8470=>"010111001",
        8471=>"111111011",
        8472=>"000100111",
        8473=>"100010110",
        8474=>"000000111",
        8475=>"101101100",
        8476=>"111111010",
        8477=>"000000111",
        8478=>"000001011",
        8479=>"000000111",
        8480=>"000001111",
        8481=>"000100110",
        8482=>"000011111",
        8483=>"000000010",
        8484=>"011111010",
        8485=>"000111100",
        8486=>"010011001",
        8487=>"011111100",
        8488=>"111000010",
        8489=>"100000110",
        8490=>"000111111",
        8491=>"000100111",
        8492=>"000011111",
        8493=>"110011010",
        8494=>"000000000",
        8495=>"111101111",
        8496=>"111111000",
        8497=>"111111000",
        8498=>"000111111",
        8499=>"100110110",
        8500=>"000001111",
        8501=>"000000110",
        8502=>"001001101",
        8503=>"111111001",
        8504=>"110000000",
        8505=>"000000010",
        8506=>"000100110",
        8507=>"111101000",
        8508=>"111010000",
        8509=>"000000111",
        8510=>"111101011",
        8511=>"000000011",
        8512=>"000000111",
        8513=>"010111111",
        8514=>"111111111",
        8515=>"110010000",
        8516=>"000111011",
        8517=>"000100111",
        8518=>"110111001",
        8519=>"000000010",
        8520=>"000001111",
        8521=>"000110110",
        8522=>"011011011",
        8523=>"000000111",
        8524=>"001000110",
        8525=>"001111111",
        8526=>"000111111",
        8527=>"110111000",
        8528=>"111111000",
        8529=>"111101100",
        8530=>"000000011",
        8531=>"011101000",
        8532=>"000101111",
        8533=>"111101000",
        8534=>"000011110",
        8535=>"001000000",
        8536=>"001001111",
        8537=>"000111111",
        8538=>"000000110",
        8539=>"011111000",
        8540=>"000100111",
        8541=>"011111001",
        8542=>"000001110",
        8543=>"000010010",
        8544=>"010101100",
        8545=>"001001001",
        8546=>"111111000",
        8547=>"100000000",
        8548=>"000110111",
        8549=>"000001111",
        8550=>"111001001",
        8551=>"010110110",
        8552=>"111000000",
        8553=>"111000000",
        8554=>"000100111",
        8555=>"111110111",
        8556=>"000000111",
        8557=>"111001000",
        8558=>"000000000",
        8559=>"000000110",
        8560=>"111101000",
        8561=>"000000001",
        8562=>"000010111",
        8563=>"111100000",
        8564=>"111111000",
        8565=>"010110001",
        8566=>"010000010",
        8567=>"001111110",
        8568=>"001011011",
        8569=>"011011010",
        8570=>"111011001",
        8571=>"000000111",
        8572=>"000010011",
        8573=>"000110110",
        8574=>"111100000",
        8575=>"011010110",
        8576=>"100010110",
        8577=>"011001101",
        8578=>"011001001",
        8579=>"010010010",
        8580=>"110111100",
        8581=>"000010001",
        8582=>"100100110",
        8583=>"001001001",
        8584=>"100110010",
        8585=>"110101101",
        8586=>"100100100",
        8587=>"000111011",
        8588=>"010100111",
        8589=>"110010100",
        8590=>"101111011",
        8591=>"001000000",
        8592=>"000111111",
        8593=>"000000000",
        8594=>"100000100",
        8595=>"000000010",
        8596=>"100100100",
        8597=>"100001011",
        8598=>"000000000",
        8599=>"010100101",
        8600=>"001001101",
        8601=>"100101000",
        8602=>"000000000",
        8603=>"010010001",
        8604=>"100000010",
        8605=>"010000000",
        8606=>"111111010",
        8607=>"100100000",
        8608=>"110110100",
        8609=>"111001111",
        8610=>"111101011",
        8611=>"100100111",
        8612=>"000000000",
        8613=>"000100100",
        8614=>"010001101",
        8615=>"100010000",
        8616=>"111011001",
        8617=>"100000110",
        8618=>"000110110",
        8619=>"000000000",
        8620=>"110111011",
        8621=>"001100001",
        8622=>"010011111",
        8623=>"111011111",
        8624=>"100110110",
        8625=>"111011000",
        8626=>"000001100",
        8627=>"000000110",
        8628=>"100110110",
        8629=>"000011011",
        8630=>"000111000",
        8631=>"000001011",
        8632=>"010011001",
        8633=>"110000110",
        8634=>"100011001",
        8635=>"110100000",
        8636=>"000000001",
        8637=>"000010110",
        8638=>"100000010",
        8639=>"000100100",
        8640=>"110110100",
        8641=>"011001001",
        8642=>"000100100",
        8643=>"111100100",
        8644=>"100110111",
        8645=>"101101000",
        8646=>"110010101",
        8647=>"100111100",
        8648=>"010110100",
        8649=>"100010010",
        8650=>"110110010",
        8651=>"000001000",
        8652=>"101111110",
        8653=>"001011001",
        8654=>"000100100",
        8655=>"011011011",
        8656=>"000100110",
        8657=>"011001001",
        8658=>"000100110",
        8659=>"000010010",
        8660=>"100100111",
        8661=>"111101001",
        8662=>"000000000",
        8663=>"100010001",
        8664=>"011011101",
        8665=>"111111011",
        8666=>"010001111",
        8667=>"101111111",
        8668=>"111111111",
        8669=>"101101000",
        8670=>"110011011",
        8671=>"111001011",
        8672=>"001100001",
        8673=>"111101111",
        8674=>"011011011",
        8675=>"011001000",
        8676=>"011111001",
        8677=>"000000100",
        8678=>"011001001",
        8679=>"001011011",
        8680=>"011111110",
        8681=>"011001000",
        8682=>"100111111",
        8683=>"101000010",
        8684=>"101001000",
        8685=>"001001001",
        8686=>"111011111",
        8687=>"001000111",
        8688=>"111110001",
        8689=>"000111011",
        8690=>"111001011",
        8691=>"010011000",
        8692=>"011000000",
        8693=>"010000011",
        8694=>"001100001",
        8695=>"100000110",
        8696=>"000100000",
        8697=>"001001111",
        8698=>"000000100",
        8699=>"001000000",
        8700=>"111001001",
        8701=>"100110101",
        8702=>"101010001",
        8703=>"100001000",
        8704=>"000010011",
        8705=>"110111111",
        8706=>"101000000",
        8707=>"100000100",
        8708=>"111001000",
        8709=>"111111010",
        8710=>"010110010",
        8711=>"101000110",
        8712=>"111001000",
        8713=>"111110110",
        8714=>"110010000",
        8715=>"001001001",
        8716=>"000000101",
        8717=>"000111000",
        8718=>"000101100",
        8719=>"100000011",
        8720=>"001000101",
        8721=>"111111000",
        8722=>"000100100",
        8723=>"001100101",
        8724=>"110110000",
        8725=>"000010000",
        8726=>"000000110",
        8727=>"000000110",
        8728=>"001101100",
        8729=>"100000100",
        8730=>"100101111",
        8731=>"100100111",
        8732=>"110111110",
        8733=>"100111011",
        8734=>"111111111",
        8735=>"000111111",
        8736=>"110000000",
        8737=>"101111101",
        8738=>"111000000",
        8739=>"111101101",
        8740=>"000010010",
        8741=>"110110010",
        8742=>"101000000",
        8743=>"000000000",
        8744=>"000000000",
        8745=>"110100000",
        8746=>"000100101",
        8747=>"100101111",
        8748=>"011101010",
        8749=>"001000000",
        8750=>"001000000",
        8751=>"111111111",
        8752=>"000101111",
        8753=>"001000001",
        8754=>"101101100",
        8755=>"011101001",
        8756=>"011101100",
        8757=>"110111111",
        8758=>"111110010",
        8759=>"010110000",
        8760=>"000010011",
        8761=>"111111111",
        8762=>"101111111",
        8763=>"000000000",
        8764=>"000000111",
        8765=>"001001000",
        8766=>"111111111",
        8767=>"111011010",
        8768=>"011111000",
        8769=>"111111110",
        8770=>"111111000",
        8771=>"110011011",
        8772=>"111111101",
        8773=>"010010011",
        8774=>"000110110",
        8775=>"000010010",
        8776=>"100000000",
        8777=>"011111111",
        8778=>"011000100",
        8779=>"011101101",
        8780=>"000101110",
        8781=>"000111100",
        8782=>"001000000",
        8783=>"000101111",
        8784=>"000000000",
        8785=>"000000000",
        8786=>"111111110",
        8787=>"010100101",
        8788=>"010110000",
        8789=>"000000000",
        8790=>"110011111",
        8791=>"111111111",
        8792=>"011001000",
        8793=>"111000000",
        8794=>"111000001",
        8795=>"000111101",
        8796=>"100101001",
        8797=>"000000000",
        8798=>"101001001",
        8799=>"010001110",
        8800=>"000110100",
        8801=>"000000100",
        8802=>"000010011",
        8803=>"101111111",
        8804=>"100111111",
        8805=>"000000101",
        8806=>"000000000",
        8807=>"111011001",
        8808=>"000000001",
        8809=>"101100101",
        8810=>"000111101",
        8811=>"011111111",
        8812=>"010010000",
        8813=>"001000101",
        8814=>"001111110",
        8815=>"011101101",
        8816=>"000000000",
        8817=>"100000000",
        8818=>"000000111",
        8819=>"111000000",
        8820=>"000000000",
        8821=>"000000110",
        8822=>"000000000",
        8823=>"100100001",
        8824=>"011011000",
        8825=>"000000010",
        8826=>"000000100",
        8827=>"101101111",
        8828=>"011000100",
        8829=>"111100010",
        8830=>"110111101",
        8831=>"111111011",
        8832=>"000110111",
        8833=>"011100100",
        8834=>"001100101",
        8835=>"000011001",
        8836=>"001101111",
        8837=>"001000101",
        8838=>"110011010",
        8839=>"110001000",
        8840=>"000100111",
        8841=>"110110111",
        8842=>"110101101",
        8843=>"011011001",
        8844=>"000011011",
        8845=>"011111110",
        8846=>"000110101",
        8847=>"111001100",
        8848=>"010010010",
        8849=>"010010001",
        8850=>"001100001",
        8851=>"100001101",
        8852=>"000011011",
        8853=>"100110101",
        8854=>"000000000",
        8855=>"011001010",
        8856=>"100111010",
        8857=>"000001110",
        8858=>"000100100",
        8859=>"000110010",
        8860=>"111010011",
        8861=>"100100011",
        8862=>"001100111",
        8863=>"110011111",
        8864=>"001111111",
        8865=>"111111000",
        8866=>"100111100",
        8867=>"011001001",
        8868=>"000111001",
        8869=>"000011011",
        8870=>"001101001",
        8871=>"101100111",
        8872=>"011001000",
        8873=>"111011000",
        8874=>"001101101",
        8875=>"000100110",
        8876=>"000011011",
        8877=>"111101101",
        8878=>"000000001",
        8879=>"111100000",
        8880=>"110111011",
        8881=>"100101001",
        8882=>"010111011",
        8883=>"000000100",
        8884=>"000100110",
        8885=>"000011000",
        8886=>"111011100",
        8887=>"000000011",
        8888=>"011100110",
        8889=>"010001101",
        8890=>"001001000",
        8891=>"010000000",
        8892=>"001100100",
        8893=>"000000001",
        8894=>"100010000",
        8895=>"110001101",
        8896=>"111010000",
        8897=>"001000011",
        8898=>"011011001",
        8899=>"001110011",
        8900=>"111011011",
        8901=>"001000111",
        8902=>"010110000",
        8903=>"011111000",
        8904=>"000000001",
        8905=>"000010111",
        8906=>"011001011",
        8907=>"100010000",
        8908=>"110000100",
        8909=>"100100011",
        8910=>"001001001",
        8911=>"100100000",
        8912=>"001001011",
        8913=>"001000110",
        8914=>"001100100",
        8915=>"100111010",
        8916=>"100010011",
        8917=>"001000000",
        8918=>"110011010",
        8919=>"100000101",
        8920=>"000101011",
        8921=>"100000001",
        8922=>"000001001",
        8923=>"000010000",
        8924=>"100110010",
        8925=>"000011011",
        8926=>"101110001",
        8927=>"000100100",
        8928=>"100010000",
        8929=>"000100101",
        8930=>"101000101",
        8931=>"010001011",
        8932=>"011111000",
        8933=>"001011011",
        8934=>"000110011",
        8935=>"010010100",
        8936=>"011100110",
        8937=>"111100100",
        8938=>"101110110",
        8939=>"111111000",
        8940=>"000100011",
        8941=>"101001001",
        8942=>"000001001",
        8943=>"101110001",
        8944=>"001000011",
        8945=>"000011100",
        8946=>"001110111",
        8947=>"110100011",
        8948=>"101100111",
        8949=>"000000000",
        8950=>"110010100",
        8951=>"110010111",
        8952=>"011011000",
        8953=>"011011001",
        8954=>"000001100",
        8955=>"010001100",
        8956=>"000110111",
        8957=>"011100000",
        8958=>"111000000",
        8959=>"111000000",
        8960=>"110111100",
        8961=>"000000110",
        8962=>"001111111",
        8963=>"011000100",
        8964=>"001111100",
        8965=>"110000000",
        8966=>"011111110",
        8967=>"000001100",
        8968=>"111110101",
        8969=>"100110000",
        8970=>"000000011",
        8971=>"001000000",
        8972=>"110000000",
        8973=>"110100110",
        8974=>"111110100",
        8975=>"001100000",
        8976=>"110000011",
        8977=>"111100000",
        8978=>"111111010",
        8979=>"000000111",
        8980=>"111000000",
        8981=>"011111111",
        8982=>"000110000",
        8983=>"000000011",
        8984=>"101011010",
        8985=>"100000000",
        8986=>"110100000",
        8987=>"000000000",
        8988=>"010111111",
        8989=>"000101111",
        8990=>"100100101",
        8991=>"101100001",
        8992=>"111000010",
        8993=>"110100000",
        8994=>"111000000",
        8995=>"000101111",
        8996=>"000111011",
        8997=>"110000000",
        8998=>"100000000",
        8999=>"101000110",
        9000=>"100110011",
        9001=>"100101111",
        9002=>"011011000",
        9003=>"111101000",
        9004=>"111111100",
        9005=>"000001101",
        9006=>"100111111",
        9007=>"101111110",
        9008=>"000101110",
        9009=>"001111111",
        9010=>"110000100",
        9011=>"110000000",
        9012=>"111010000",
        9013=>"100000000",
        9014=>"110000000",
        9015=>"000010011",
        9016=>"111000110",
        9017=>"100111111",
        9018=>"001001101",
        9019=>"000111111",
        9020=>"110011001",
        9021=>"111000000",
        9022=>"110010000",
        9023=>"111000000",
        9024=>"001000101",
        9025=>"001000001",
        9026=>"001010101",
        9027=>"000110111",
        9028=>"111110110",
        9029=>"000001101",
        9030=>"111101100",
        9031=>"000000010",
        9032=>"110001110",
        9033=>"000111100",
        9034=>"111110111",
        9035=>"111000000",
        9036=>"001000110",
        9037=>"001000111",
        9038=>"001111101",
        9039=>"000111111",
        9040=>"110001110",
        9041=>"000000000",
        9042=>"100100000",
        9043=>"111010100",
        9044=>"110010000",
        9045=>"110011001",
        9046=>"111010010",
        9047=>"000010110",
        9048=>"011001100",
        9049=>"100101011",
        9050=>"001001011",
        9051=>"000001001",
        9052=>"000000000",
        9053=>"000000111",
        9054=>"111000000",
        9055=>"100101111",
        9056=>"111101000",
        9057=>"000100100",
        9058=>"001110110",
        9059=>"000111111",
        9060=>"001000000",
        9061=>"110000000",
        9062=>"000000000",
        9063=>"110111110",
        9064=>"110110110",
        9065=>"000101100",
        9066=>"000100010",
        9067=>"011000010",
        9068=>"110110001",
        9069=>"001000111",
        9070=>"110110000",
        9071=>"100110110",
        9072=>"000110111",
        9073=>"001101111",
        9074=>"110001111",
        9075=>"010000000",
        9076=>"000000011",
        9077=>"110111011",
        9078=>"110110001",
        9079=>"110110111",
        9080=>"000000000",
        9081=>"111000100",
        9082=>"101001000",
        9083=>"000000000",
        9084=>"110110011",
        9085=>"001001100",
        9086=>"100000110",
        9087=>"111001000",
        9088=>"110111111",
        9089=>"000111111",
        9090=>"000010111",
        9091=>"000000000",
        9092=>"111011001",
        9093=>"111111111",
        9094=>"000100101",
        9095=>"100000101",
        9096=>"100000011",
        9097=>"011111100",
        9098=>"111111111",
        9099=>"111001000",
        9100=>"110111010",
        9101=>"010111010",
        9102=>"000001001",
        9103=>"110100111",
        9104=>"100111100",
        9105=>"101000101",
        9106=>"111111011",
        9107=>"100100000",
        9108=>"000110110",
        9109=>"000000010",
        9110=>"000000010",
        9111=>"111111010",
        9112=>"111101100",
        9113=>"100101000",
        9114=>"101101101",
        9115=>"110000000",
        9116=>"000101101",
        9117=>"000111111",
        9118=>"111011101",
        9119=>"010010111",
        9120=>"010111001",
        9121=>"000100100",
        9122=>"011111111",
        9123=>"101000000",
        9124=>"011111111",
        9125=>"000111111",
        9126=>"100111111",
        9127=>"000000111",
        9128=>"100000000",
        9129=>"110000000",
        9130=>"011000000",
        9131=>"110100100",
        9132=>"111101000",
        9133=>"111111110",
        9134=>"110000000",
        9135=>"110100111",
        9136=>"110010000",
        9137=>"110111111",
        9138=>"111000100",
        9139=>"110011101",
        9140=>"000100101",
        9141=>"101101000",
        9142=>"111110110",
        9143=>"000110010",
        9144=>"110110010",
        9145=>"000101111",
        9146=>"110110010",
        9147=>"000000000",
        9148=>"111110000",
        9149=>"001001111",
        9150=>"111000100",
        9151=>"000000000",
        9152=>"000110111",
        9153=>"000000000",
        9154=>"000100000",
        9155=>"000000000",
        9156=>"010000000",
        9157=>"011111110",
        9158=>"110101000",
        9159=>"111111111",
        9160=>"000110001",
        9161=>"000111111",
        9162=>"101011000",
        9163=>"111000000",
        9164=>"000000000",
        9165=>"111000001",
        9166=>"010000001",
        9167=>"000000000",
        9168=>"100010111",
        9169=>"110000000",
        9170=>"000000000",
        9171=>"110111010",
        9172=>"100100110",
        9173=>"010111000",
        9174=>"100000111",
        9175=>"001101111",
        9176=>"011001000",
        9177=>"101111010",
        9178=>"000001001",
        9179=>"001000000",
        9180=>"100111111",
        9181=>"001000000",
        9182=>"001101101",
        9183=>"010111111",
        9184=>"101111101",
        9185=>"011011011",
        9186=>"000111111",
        9187=>"110110000",
        9188=>"000001100",
        9189=>"000000111",
        9190=>"001101001",
        9191=>"111011000",
        9192=>"000000000",
        9193=>"111011010",
        9194=>"110100101",
        9195=>"111111100",
        9196=>"011111111",
        9197=>"000011110",
        9198=>"110000001",
        9199=>"000000100",
        9200=>"000010110",
        9201=>"001000010",
        9202=>"101111001",
        9203=>"000110110",
        9204=>"000010110",
        9205=>"111001111",
        9206=>"000000000",
        9207=>"111111001",
        9208=>"111011100",
        9209=>"111110000",
        9210=>"000100111",
        9211=>"111111111",
        9212=>"001100100",
        9213=>"000110010",
        9214=>"101111111",
        9215=>"100111111",
        9216=>"111111110",
        9217=>"001101011",
        9218=>"000000101",
        9219=>"111010001",
        9220=>"111111111",
        9221=>"010000000",
        9222=>"101000000",
        9223=>"010000000",
        9224=>"111001110",
        9225=>"100000101",
        9226=>"100101111",
        9227=>"011001111",
        9228=>"000000111",
        9229=>"111111010",
        9230=>"010011100",
        9231=>"000000111",
        9232=>"001001001",
        9233=>"100000110",
        9234=>"011001000",
        9235=>"110011001",
        9236=>"101001010",
        9237=>"101000000",
        9238=>"101000000",
        9239=>"000110010",
        9240=>"110000000",
        9241=>"110001111",
        9242=>"111100000",
        9243=>"011011100",
        9244=>"001011111",
        9245=>"010011000",
        9246=>"011011000",
        9247=>"010111111",
        9248=>"000001000",
        9249=>"000000000",
        9250=>"111110111",
        9251=>"010111000",
        9252=>"010000000",
        9253=>"111001001",
        9254=>"000101111",
        9255=>"000000000",
        9256=>"001000010",
        9257=>"110001001",
        9258=>"011111011",
        9259=>"110111000",
        9260=>"010111010",
        9261=>"011011000",
        9262=>"000010000",
        9263=>"111000000",
        9264=>"101000011",
        9265=>"001000001",
        9266=>"000110110",
        9267=>"000001000",
        9268=>"001111110",
        9269=>"111000000",
        9270=>"110111111",
        9271=>"010000000",
        9272=>"011000100",
        9273=>"000111010",
        9274=>"001000000",
        9275=>"000101111",
        9276=>"000000001",
        9277=>"000011110",
        9278=>"110110001",
        9279=>"101011111",
        9280=>"010000000",
        9281=>"000000000",
        9282=>"010000111",
        9283=>"111010010",
        9284=>"100001111",
        9285=>"110110110",
        9286=>"101000000",
        9287=>"010100110",
        9288=>"100000100",
        9289=>"100110010",
        9290=>"011100000",
        9291=>"111101000",
        9292=>"000000010",
        9293=>"000101111",
        9294=>"010110111",
        9295=>"100101110",
        9296=>"000010111",
        9297=>"101001000",
        9298=>"000000000",
        9299=>"000100100",
        9300=>"011011011",
        9301=>"000000110",
        9302=>"011111000",
        9303=>"111110000",
        9304=>"011100100",
        9305=>"100000110",
        9306=>"101011111",
        9307=>"000000111",
        9308=>"001111101",
        9309=>"001100000",
        9310=>"100000111",
        9311=>"001111101",
        9312=>"110000001",
        9313=>"100100100",
        9314=>"111010111",
        9315=>"000101111",
        9316=>"110101100",
        9317=>"010100000",
        9318=>"101100000",
        9319=>"011011111",
        9320=>"100100011",
        9321=>"100000101",
        9322=>"110000001",
        9323=>"000000000",
        9324=>"101001000",
        9325=>"001001101",
        9326=>"111100100",
        9327=>"110110000",
        9328=>"010010000",
        9329=>"010011111",
        9330=>"100000000",
        9331=>"111111111",
        9332=>"100111111",
        9333=>"000000001",
        9334=>"100111111",
        9335=>"100111111",
        9336=>"011010000",
        9337=>"000110111",
        9338=>"010000100",
        9339=>"111101101",
        9340=>"101000110",
        9341=>"111101111",
        9342=>"111110000",
        9343=>"111011111",
        9344=>"111010111",
        9345=>"001001001",
        9346=>"110110010",
        9347=>"011011010",
        9348=>"000000100",
        9349=>"111111000",
        9350=>"111000110",
        9351=>"111111111",
        9352=>"111111111",
        9353=>"000000101",
        9354=>"001101101",
        9355=>"000000000",
        9356=>"010110010",
        9357=>"010111010",
        9358=>"111111111",
        9359=>"100011001",
        9360=>"001110110",
        9361=>"010010110",
        9362=>"000000100",
        9363=>"000100000",
        9364=>"000000000",
        9365=>"010111111",
        9366=>"001100101",
        9367=>"000000000",
        9368=>"000001001",
        9369=>"000000001",
        9370=>"100000001",
        9371=>"010110011",
        9372=>"000000000",
        9373=>"101001101",
        9374=>"111011011",
        9375=>"101111111",
        9376=>"111111111",
        9377=>"111110110",
        9378=>"010111110",
        9379=>"000000000",
        9380=>"110111011",
        9381=>"001111000",
        9382=>"001000000",
        9383=>"101101001",
        9384=>"000000000",
        9385=>"000000000",
        9386=>"010011001",
        9387=>"001001101",
        9388=>"101100101",
        9389=>"001000000",
        9390=>"111111110",
        9391=>"110010011",
        9392=>"110100000",
        9393=>"010111011",
        9394=>"011111110",
        9395=>"110000000",
        9396=>"011111111",
        9397=>"000000010",
        9398=>"111111111",
        9399=>"000100000",
        9400=>"100000000",
        9401=>"000110011",
        9402=>"010000000",
        9403=>"000000001",
        9404=>"000010010",
        9405=>"101101010",
        9406=>"110011110",
        9407=>"111001111",
        9408=>"101000101",
        9409=>"000000000",
        9410=>"101000000",
        9411=>"001000010",
        9412=>"011111111",
        9413=>"001000110",
        9414=>"110111111",
        9415=>"111111111",
        9416=>"110111011",
        9417=>"101101001",
        9418=>"000000100",
        9419=>"001000101",
        9420=>"000000000",
        9421=>"111101000",
        9422=>"111111111",
        9423=>"110110000",
        9424=>"101000000",
        9425=>"000001001",
        9426=>"100000100",
        9427=>"000110100",
        9428=>"110001011",
        9429=>"000000000",
        9430=>"000001111",
        9431=>"111111101",
        9432=>"000000001",
        9433=>"111111111",
        9434=>"001001001",
        9435=>"011111110",
        9436=>"100000011",
        9437=>"001000100",
        9438=>"101111111",
        9439=>"000111010",
        9440=>"111110000",
        9441=>"110000000",
        9442=>"000110111",
        9443=>"000000010",
        9444=>"111111001",
        9445=>"111110110",
        9446=>"001100100",
        9447=>"111101101",
        9448=>"001000000",
        9449=>"001000000",
        9450=>"100101101",
        9451=>"111100110",
        9452=>"011001000",
        9453=>"101000000",
        9454=>"000001000",
        9455=>"111111110",
        9456=>"010110111",
        9457=>"101001111",
        9458=>"111111101",
        9459=>"000000000",
        9460=>"000011010",
        9461=>"000000100",
        9462=>"111111111",
        9463=>"110110010",
        9464=>"000000100",
        9465=>"100100000",
        9466=>"100000000",
        9467=>"110111111",
        9468=>"100111100",
        9469=>"000000000",
        9470=>"000000001",
        9471=>"000100110",
        9472=>"111111110",
        9473=>"000111000",
        9474=>"000100111",
        9475=>"101100111",
        9476=>"011000100",
        9477=>"100110000",
        9478=>"111010000",
        9479=>"111000100",
        9480=>"001001101",
        9481=>"110110000",
        9482=>"111000010",
        9483=>"111011110",
        9484=>"101101001",
        9485=>"111111000",
        9486=>"000000001",
        9487=>"110100011",
        9488=>"001001111",
        9489=>"000101111",
        9490=>"100001000",
        9491=>"100100001",
        9492=>"110101011",
        9493=>"010111010",
        9494=>"111100111",
        9495=>"000000000",
        9496=>"111110100",
        9497=>"111100001",
        9498=>"000110100",
        9499=>"000001010",
        9500=>"000101001",
        9501=>"000011000",
        9502=>"001011010",
        9503=>"111111111",
        9504=>"111000101",
        9505=>"100001011",
        9506=>"111101111",
        9507=>"000000010",
        9508=>"000101101",
        9509=>"101101111",
        9510=>"101100111",
        9511=>"101101100",
        9512=>"000000000",
        9513=>"101000011",
        9514=>"000101110",
        9515=>"010101001",
        9516=>"010001111",
        9517=>"111010000",
        9518=>"010000000",
        9519=>"010000100",
        9520=>"011101110",
        9521=>"000000000",
        9522=>"000001110",
        9523=>"010010000",
        9524=>"000010000",
        9525=>"000000000",
        9526=>"011000001",
        9527=>"001000000",
        9528=>"100010011",
        9529=>"000011010",
        9530=>"011010000",
        9531=>"000111100",
        9532=>"101000100",
        9533=>"000000011",
        9534=>"100110110",
        9535=>"011011011",
        9536=>"000000001",
        9537=>"110100100",
        9538=>"111010100",
        9539=>"101101101",
        9540=>"111101111",
        9541=>"101100100",
        9542=>"000000100",
        9543=>"000000000",
        9544=>"110110101",
        9545=>"000100010",
        9546=>"100000110",
        9547=>"101101000",
        9548=>"111000000",
        9549=>"011111000",
        9550=>"000000011",
        9551=>"000000100",
        9552=>"100000111",
        9553=>"100100001",
        9554=>"000001000",
        9555=>"011001000",
        9556=>"100001001",
        9557=>"101000101",
        9558=>"000011011",
        9559=>"110110010",
        9560=>"001101100",
        9561=>"001010100",
        9562=>"000110000",
        9563=>"110101111",
        9564=>"110111000",
        9565=>"011011000",
        9566=>"000000000",
        9567=>"000001011",
        9568=>"110110101",
        9569=>"000100110",
        9570=>"111100101",
        9571=>"110100100",
        9572=>"011110101",
        9573=>"000010011",
        9574=>"001000100",
        9575=>"000000011",
        9576=>"101100111",
        9577=>"010000000",
        9578=>"000101001",
        9579=>"111110000",
        9580=>"001100001",
        9581=>"100000011",
        9582=>"001000000",
        9583=>"000110100",
        9584=>"011000101",
        9585=>"000000000",
        9586=>"101011000",
        9587=>"100100111",
        9588=>"100000000",
        9589=>"000000100",
        9590=>"111111111",
        9591=>"110100011",
        9592=>"011101100",
        9593=>"000001010",
        9594=>"000000110",
        9595=>"101010111",
        9596=>"000000011",
        9597=>"110000010",
        9598=>"101011010",
        9599=>"100001011",
        9600=>"100011011",
        9601=>"110110000",
        9602=>"000000000",
        9603=>"111111111",
        9604=>"001111111",
        9605=>"111011100",
        9606=>"111111111",
        9607=>"100110111",
        9608=>"001011101",
        9609=>"111010110",
        9610=>"000000000",
        9611=>"001000000",
        9612=>"000111111",
        9613=>"000111010",
        9614=>"000001111",
        9615=>"010110111",
        9616=>"111110000",
        9617=>"010111010",
        9618=>"110111110",
        9619=>"110111011",
        9620=>"000000000",
        9621=>"000000100",
        9622=>"011000000",
        9623=>"110111111",
        9624=>"101110011",
        9625=>"000001001",
        9626=>"000000000",
        9627=>"001001001",
        9628=>"111111111",
        9629=>"000000000",
        9630=>"000101010",
        9631=>"111010101",
        9632=>"001000000",
        9633=>"111101001",
        9634=>"010000010",
        9635=>"000011111",
        9636=>"111111101",
        9637=>"101000000",
        9638=>"011111111",
        9639=>"000000000",
        9640=>"000001000",
        9641=>"000100110",
        9642=>"000000001",
        9643=>"110011011",
        9644=>"000110110",
        9645=>"011111011",
        9646=>"010110101",
        9647=>"010110010",
        9648=>"111000011",
        9649=>"000000000",
        9650=>"001000110",
        9651=>"100000011",
        9652=>"111111010",
        9653=>"011001000",
        9654=>"111111101",
        9655=>"000010011",
        9656=>"110111010",
        9657=>"010000111",
        9658=>"001100100",
        9659=>"111111111",
        9660=>"000000000",
        9661=>"111111011",
        9662=>"110100010",
        9663=>"111111111",
        9664=>"000000000",
        9665=>"111001000",
        9666=>"011011000",
        9667=>"100101111",
        9668=>"111111101",
        9669=>"001111111",
        9670=>"000010110",
        9671=>"011111000",
        9672=>"111111000",
        9673=>"101101101",
        9674=>"001000000",
        9675=>"000000000",
        9676=>"111111011",
        9677=>"010011001",
        9678=>"111111111",
        9679=>"100100111",
        9680=>"010111111",
        9681=>"100000001",
        9682=>"000100000",
        9683=>"101111111",
        9684=>"110111111",
        9685=>"000111111",
        9686=>"111011011",
        9687=>"001111010",
        9688=>"001000011",
        9689=>"101010000",
        9690=>"000000000",
        9691=>"111111111",
        9692=>"111110011",
        9693=>"001111010",
        9694=>"000000000",
        9695=>"000000000",
        9696=>"101110000",
        9697=>"000011110",
        9698=>"000000000",
        9699=>"010111110",
        9700=>"010011111",
        9701=>"100001011",
        9702=>"000000000",
        9703=>"101100000",
        9704=>"110111000",
        9705=>"110000000",
        9706=>"110100000",
        9707=>"000011110",
        9708=>"000101000",
        9709=>"000000000",
        9710=>"101000000",
        9711=>"010110011",
        9712=>"101001111",
        9713=>"000001000",
        9714=>"000001000",
        9715=>"000000111",
        9716=>"000000000",
        9717=>"000111000",
        9718=>"010111111",
        9719=>"100111001",
        9720=>"000000000",
        9721=>"001111111",
        9722=>"111111100",
        9723=>"111111001",
        9724=>"000000100",
        9725=>"011011001",
        9726=>"000010000",
        9727=>"000001001",
        9728=>"111111111",
        9729=>"000000001",
        9730=>"000000001",
        9731=>"111010110",
        9732=>"111011100",
        9733=>"110110110",
        9734=>"110110110",
        9735=>"101111001",
        9736=>"111111000",
        9737=>"011110110",
        9738=>"001001011",
        9739=>"001100100",
        9740=>"100000000",
        9741=>"010110000",
        9742=>"110001001",
        9743=>"000000000",
        9744=>"110111000",
        9745=>"001000000",
        9746=>"011001011",
        9747=>"100000001",
        9748=>"000101111",
        9749=>"000001010",
        9750=>"000000000",
        9751=>"110000000",
        9752=>"011011011",
        9753=>"000000000",
        9754=>"001001100",
        9755=>"010100100",
        9756=>"101001010",
        9757=>"111111011",
        9758=>"000000101",
        9759=>"111111111",
        9760=>"110110111",
        9761=>"111001101",
        9762=>"011101001",
        9763=>"001101111",
        9764=>"000000000",
        9765=>"010000000",
        9766=>"111111111",
        9767=>"000000001",
        9768=>"000000000",
        9769=>"000010111",
        9770=>"011011000",
        9771=>"101001111",
        9772=>"011001100",
        9773=>"111101111",
        9774=>"000000110",
        9775=>"111111111",
        9776=>"111111110",
        9777=>"010110000",
        9778=>"110110000",
        9779=>"110000110",
        9780=>"111110011",
        9781=>"001000000",
        9782=>"010110110",
        9783=>"000000000",
        9784=>"000000001",
        9785=>"000000100",
        9786=>"111000010",
        9787=>"110110100",
        9788=>"000101000",
        9789=>"110110010",
        9790=>"100100001",
        9791=>"100111011",
        9792=>"000001111",
        9793=>"011010010",
        9794=>"110110110",
        9795=>"011001010",
        9796=>"111101110",
        9797=>"111111110",
        9798=>"111111100",
        9799=>"110100000",
        9800=>"011110010",
        9801=>"110111111",
        9802=>"010000110",
        9803=>"001000000",
        9804=>"110100110",
        9805=>"001000000",
        9806=>"111111110",
        9807=>"100110110",
        9808=>"110110000",
        9809=>"110110101",
        9810=>"001111111",
        9811=>"111000000",
        9812=>"111011111",
        9813=>"000000000",
        9814=>"010110100",
        9815=>"001001111",
        9816=>"001001001",
        9817=>"101110000",
        9818=>"001000011",
        9819=>"000010000",
        9820=>"011011011",
        9821=>"000000100",
        9822=>"000011000",
        9823=>"010000000",
        9824=>"111110000",
        9825=>"111111000",
        9826=>"010110000",
        9827=>"111101000",
        9828=>"001110110",
        9829=>"111110000",
        9830=>"111111111",
        9831=>"000000101",
        9832=>"110110010",
        9833=>"000000001",
        9834=>"000011111",
        9835=>"000100110",
        9836=>"000110110",
        9837=>"100111001",
        9838=>"001011011",
        9839=>"011110101",
        9840=>"000000001",
        9841=>"000000100",
        9842=>"110110000",
        9843=>"110111110",
        9844=>"011001111",
        9845=>"000000111",
        9846=>"000000110",
        9847=>"110111000",
        9848=>"111110011",
        9849=>"100110110",
        9850=>"100100100",
        9851=>"111110110",
        9852=>"000001011",
        9853=>"111111111",
        9854=>"000000000",
        9855=>"111111110",
        9856=>"111110000",
        9857=>"111000001",
        9858=>"011100001",
        9859=>"011011110",
        9860=>"010000000",
        9861=>"011011010",
        9862=>"011010000",
        9863=>"000111111",
        9864=>"011110000",
        9865=>"000000001",
        9866=>"000000011",
        9867=>"011000001",
        9868=>"100111010",
        9869=>"011111110",
        9870=>"011111110",
        9871=>"110110110",
        9872=>"000000000",
        9873=>"001001011",
        9874=>"001011011",
        9875=>"011011010",
        9876=>"010000000",
        9877=>"010101010",
        9878=>"000100001",
        9879=>"011000000",
        9880=>"101111110",
        9881=>"100111111",
        9882=>"011100000",
        9883=>"101111111",
        9884=>"111111011",
        9885=>"011011010",
        9886=>"010000000",
        9887=>"000000111",
        9888=>"011111011",
        9889=>"101011111",
        9890=>"100000011",
        9891=>"110010110",
        9892=>"011000100",
        9893=>"111111001",
        9894=>"011111101",
        9895=>"111110000",
        9896=>"110100100",
        9897=>"101011110",
        9898=>"101000010",
        9899=>"101011010",
        9900=>"000000000",
        9901=>"110111010",
        9902=>"100001111",
        9903=>"000111110",
        9904=>"011000010",
        9905=>"110100011",
        9906=>"110100001",
        9907=>"101000100",
        9908=>"001010110",
        9909=>"000000010",
        9910=>"000100110",
        9911=>"011111001",
        9912=>"011100000",
        9913=>"110000100",
        9914=>"011101011",
        9915=>"000100001",
        9916=>"100100001",
        9917=>"000001001",
        9918=>"100100000",
        9919=>"010010000",
        9920=>"001001110",
        9921=>"101000000",
        9922=>"000110110",
        9923=>"010000001",
        9924=>"111011111",
        9925=>"111010000",
        9926=>"010111000",
        9927=>"100100100",
        9928=>"000111110",
        9929=>"011000000",
        9930=>"000000100",
        9931=>"000001001",
        9932=>"000111110",
        9933=>"000111110",
        9934=>"010111100",
        9935=>"100100000",
        9936=>"010010001",
        9937=>"111110000",
        9938=>"100100110",
        9939=>"111111100",
        9940=>"110000001",
        9941=>"110100001",
        9942=>"000011010",
        9943=>"011101001",
        9944=>"111110011",
        9945=>"100000000",
        9946=>"011011000",
        9947=>"001000001",
        9948=>"101011110",
        9949=>"000000101",
        9950=>"001000000",
        9951=>"000010000",
        9952=>"001011010",
        9953=>"110110111",
        9954=>"110100100",
        9955=>"111111100",
        9956=>"000010110",
        9957=>"000010000",
        9958=>"100100001",
        9959=>"101011110",
        9960=>"100100100",
        9961=>"111000001",
        9962=>"001011110",
        9963=>"010001110",
        9964=>"100000000",
        9965=>"110001000",
        9966=>"011111000",
        9967=>"001011011",
        9968=>"100111111",
        9969=>"111001000",
        9970=>"111000000",
        9971=>"000110010",
        9972=>"011001001",
        9973=>"000000000",
        9974=>"111001111",
        9975=>"100111111",
        9976=>"000000111",
        9977=>"101000100",
        9978=>"111111001",
        9979=>"000000111",
        9980=>"000100000",
        9981=>"111100100",
        9982=>"111100001",
        9983=>"111011010",
        9984=>"101100000",
        9985=>"110000000",
        9986=>"101101100",
        9987=>"000111111",
        9988=>"110000111",
        9989=>"101111111",
        9990=>"010011111",
        9991=>"000010000",
        9992=>"110100110",
        9993=>"100000001",
        9994=>"111000100",
        9995=>"001001101",
        9996=>"111110111",
        9997=>"010010111",
        9998=>"011110100",
        9999=>"000001100",
        10000=>"110111011",
        10001=>"010001111",
        10002=>"000001001",
        10003=>"000001101",
        10004=>"000000001",
        10005=>"000100010",
        10006=>"000000100",
        10007=>"000001101",
        10008=>"000100000",
        10009=>"011110100",
        10010=>"000000000",
        10011=>"100000100",
        10012=>"111101111",
        10013=>"011111111",
        10014=>"111100001",
        10015=>"111101101",
        10016=>"101111111",
        10017=>"000000000",
        10018=>"011011101",
        10019=>"100101111",
        10020=>"001101001",
        10021=>"101101111",
        10022=>"010010000",
        10023=>"110110010",
        10024=>"111111101",
        10025=>"100011111",
        10026=>"110011110",
        10027=>"011101110",
        10028=>"010111001",
        10029=>"111001000",
        10030=>"000000000",
        10031=>"111111111",
        10032=>"000000000",
        10033=>"000000000",
        10034=>"001001101",
        10035=>"000011000",
        10036=>"110110110",
        10037=>"110010101",
        10038=>"001000101",
        10039=>"110101111",
        10040=>"100001101",
        10041=>"110100111",
        10042=>"000000100",
        10043=>"100010100",
        10044=>"000001001",
        10045=>"000001101",
        10046=>"001000001",
        10047=>"011001100",
        10048=>"011011000",
        10049=>"000000000",
        10050=>"000111101",
        10051=>"011101111",
        10052=>"111111011",
        10053=>"000000000",
        10054=>"000010010",
        10055=>"000101100",
        10056=>"011111110",
        10057=>"111110100",
        10058=>"000011001",
        10059=>"000000000",
        10060=>"001001111",
        10061=>"010000110",
        10062=>"110011001",
        10063=>"000000111",
        10064=>"010010000",
        10065=>"011010110",
        10066=>"000111110",
        10067=>"010111111",
        10068=>"000001000",
        10069=>"000000000",
        10070=>"111111110",
        10071=>"101101111",
        10072=>"000100100",
        10073=>"000000110",
        10074=>"110110110",
        10075=>"000001000",
        10076=>"001011010",
        10077=>"000110110",
        10078=>"011111011",
        10079=>"101101001",
        10080=>"011011111",
        10081=>"000100000",
        10082=>"111110010",
        10083=>"000101101",
        10084=>"000100101",
        10085=>"000110111",
        10086=>"110110111",
        10087=>"001001100",
        10088=>"110010111",
        10089=>"110101010",
        10090=>"001100101",
        10091=>"000000100",
        10092=>"000000000",
        10093=>"001101111",
        10094=>"100001000",
        10095=>"110010011",
        10096=>"000101111",
        10097=>"111111111",
        10098=>"011011010",
        10099=>"100101111",
        10100=>"010000111",
        10101=>"000010001",
        10102=>"000000000",
        10103=>"000101100",
        10104=>"100110111",
        10105=>"000101001",
        10106=>"011110111",
        10107=>"010010010",
        10108=>"010010110",
        10109=>"000000000",
        10110=>"100000000",
        10111=>"110000001",
        10112=>"111111000",
        10113=>"110010001",
        10114=>"111111100",
        10115=>"000000000",
        10116=>"000000110",
        10117=>"100101000",
        10118=>"001111000",
        10119=>"000000101",
        10120=>"001011110",
        10121=>"100000001",
        10122=>"111000000",
        10123=>"001100100",
        10124=>"000011111",
        10125=>"111110110",
        10126=>"100111111",
        10127=>"010000111",
        10128=>"111111010",
        10129=>"000110111",
        10130=>"011100000",
        10131=>"100000001",
        10132=>"111001001",
        10133=>"000001000",
        10134=>"000101011",
        10135=>"001010111",
        10136=>"110001011",
        10137=>"100001011",
        10138=>"100100111",
        10139=>"010111100",
        10140=>"000010010",
        10141=>"011111111",
        10142=>"100100111",
        10143=>"010111100",
        10144=>"001101111",
        10145=>"010100000",
        10146=>"000100000",
        10147=>"000001001",
        10148=>"011101000",
        10149=>"001001011",
        10150=>"000111111",
        10151=>"111000000",
        10152=>"000000001",
        10153=>"110000001",
        10154=>"101101011",
        10155=>"110011011",
        10156=>"000111111",
        10157=>"001000101",
        10158=>"000000000",
        10159=>"000111111",
        10160=>"010000010",
        10161=>"111010001",
        10162=>"001000110",
        10163=>"000000001",
        10164=>"100011111",
        10165=>"000000000",
        10166=>"111000000",
        10167=>"000101001",
        10168=>"111111101",
        10169=>"111010111",
        10170=>"000000110",
        10171=>"001100100",
        10172=>"000011111",
        10173=>"110111000",
        10174=>"111110101",
        10175=>"111010000",
        10176=>"100000000",
        10177=>"000000011",
        10178=>"111111111",
        10179=>"111000000",
        10180=>"111100011",
        10181=>"110110000",
        10182=>"111010010",
        10183=>"000000000",
        10184=>"011011011",
        10185=>"111111000",
        10186=>"000000111",
        10187=>"000101111",
        10188=>"111111010",
        10189=>"111011000",
        10190=>"101111010",
        10191=>"111111000",
        10192=>"010000000",
        10193=>"000000111",
        10194=>"000000000",
        10195=>"000101111",
        10196=>"011000000",
        10197=>"101000000",
        10198=>"101011000",
        10199=>"000101101",
        10200=>"110001000",
        10201=>"001001001",
        10202=>"011001111",
        10203=>"000111111",
        10204=>"111111000",
        10205=>"101100000",
        10206=>"000000110",
        10207=>"111111010",
        10208=>"111011011",
        10209=>"011001100",
        10210=>"111000000",
        10211=>"000010011",
        10212=>"000011101",
        10213=>"111010111",
        10214=>"001001111",
        10215=>"010000001",
        10216=>"110000101",
        10217=>"100100010",
        10218=>"110001001",
        10219=>"000101011",
        10220=>"110000000",
        10221=>"001000111",
        10222=>"101000001",
        10223=>"000111111",
        10224=>"111000000",
        10225=>"111110111",
        10226=>"011000000",
        10227=>"111000100",
        10228=>"111011000",
        10229=>"000000000",
        10230=>"000000101",
        10231=>"001011011",
        10232=>"111011101",
        10233=>"000000000",
        10234=>"010001011",
        10235=>"000111011",
        10236=>"100100011",
        10237=>"110011111",
        10238=>"111000001",
        10239=>"000000111",
        10240=>"000000000",
        10241=>"111111011",
        10242=>"000000101",
        10243=>"110111111",
        10244=>"000111111",
        10245=>"110000110",
        10246=>"111111111",
        10247=>"001000101",
        10248=>"100110000",
        10249=>"000100000",
        10250=>"111001001",
        10251=>"011011111",
        10252=>"000111011",
        10253=>"010010010",
        10254=>"101100000",
        10255=>"100100000",
        10256=>"011011010",
        10257=>"000000000",
        10258=>"001000000",
        10259=>"000011001",
        10260=>"000000000",
        10261=>"000000000",
        10262=>"001000000",
        10263=>"010000000",
        10264=>"110011010",
        10265=>"000011001",
        10266=>"100001100",
        10267=>"000010001",
        10268=>"111001110",
        10269=>"010010011",
        10270=>"001111011",
        10271=>"000000000",
        10272=>"000010111",
        10273=>"111111011",
        10274=>"000011111",
        10275=>"000000000",
        10276=>"111011101",
        10277=>"000010000",
        10278=>"010111010",
        10279=>"000111010",
        10280=>"011000010",
        10281=>"000000000",
        10282=>"011111010",
        10283=>"100100100",
        10284=>"011000000",
        10285=>"000000000",
        10286=>"000111110",
        10287=>"010010000",
        10288=>"110111000",
        10289=>"000010011",
        10290=>"000111010",
        10291=>"110000010",
        10292=>"110111101",
        10293=>"000000000",
        10294=>"010000100",
        10295=>"000010000",
        10296=>"000000000",
        10297=>"000000000",
        10298=>"011001001",
        10299=>"111111111",
        10300=>"011000000",
        10301=>"100000100",
        10302=>"010000100",
        10303=>"011111011",
        10304=>"000000000",
        10305=>"100101001",
        10306=>"011000000",
        10307=>"010110000",
        10308=>"100100000",
        10309=>"011011000",
        10310=>"101000000",
        10311=>"010110111",
        10312=>"110110010",
        10313=>"000001100",
        10314=>"100110000",
        10315=>"010000000",
        10316=>"100011000",
        10317=>"000000000",
        10318=>"100000000",
        10319=>"110010000",
        10320=>"000000000",
        10321=>"111110000",
        10322=>"011111011",
        10323=>"000000111",
        10324=>"100000000",
        10325=>"000010010",
        10326=>"011010000",
        10327=>"010010110",
        10328=>"100100100",
        10329=>"111011000",
        10330=>"101011111",
        10331=>"000000000",
        10332=>"000001011",
        10333=>"010010010",
        10334=>"110100111",
        10335=>"000010000",
        10336=>"011001011",
        10337=>"110111010",
        10338=>"000010010",
        10339=>"000000000",
        10340=>"000000000",
        10341=>"010010000",
        10342=>"111011110",
        10343=>"110110111",
        10344=>"010011111",
        10345=>"001000101",
        10346=>"001111100",
        10347=>"010110111",
        10348=>"110111111",
        10349=>"001000000",
        10350=>"111000010",
        10351=>"111111100",
        10352=>"000010000",
        10353=>"010010000",
        10354=>"110010010",
        10355=>"110010000",
        10356=>"111111101",
        10357=>"101001101",
        10358=>"111111010",
        10359=>"011110100",
        10360=>"000010111",
        10361=>"110010000",
        10362=>"011000001",
        10363=>"011010110",
        10364=>"101111111",
        10365=>"101110111",
        10366=>"100000001",
        10367=>"011111110",
        10368=>"111011011",
        10369=>"100100100",
        10370=>"011001001",
        10371=>"010011011",
        10372=>"010010100",
        10373=>"100100111",
        10374=>"011000010",
        10375=>"100100110",
        10376=>"101101111",
        10377=>"001011011",
        10378=>"100100100",
        10379=>"101110010",
        10380=>"111100110",
        10381=>"110100110",
        10382=>"011001000",
        10383=>"100100110",
        10384=>"000011011",
        10385=>"100100110",
        10386=>"111001000",
        10387=>"001101000",
        10388=>"100100111",
        10389=>"010000000",
        10390=>"001000000",
        10391=>"000011011",
        10392=>"110000110",
        10393=>"001010001",
        10394=>"111110101",
        10395=>"110110011",
        10396=>"000100110",
        10397=>"011001001",
        10398=>"011011011",
        10399=>"011011011",
        10400=>"011000001",
        10401=>"111110101",
        10402=>"111011011",
        10403=>"001011011",
        10404=>"011001001",
        10405=>"100100110",
        10406=>"001100000",
        10407=>"010010011",
        10408=>"011000110",
        10409=>"001011000",
        10410=>"100110100",
        10411=>"011011001",
        10412=>"011011001",
        10413=>"001001011",
        10414=>"000001011",
        10415=>"010111111",
        10416=>"011011001",
        10417=>"000001110",
        10418=>"011010001",
        10419=>"011001001",
        10420=>"100100111",
        10421=>"011010011",
        10422=>"010110011",
        10423=>"110110100",
        10424=>"011110110",
        10425=>"001011011",
        10426=>"011010000",
        10427=>"110000001",
        10428=>"100100110",
        10429=>"001000100",
        10430=>"110111011",
        10431=>"110010011",
        10432=>"000111011",
        10433=>"011011001",
        10434=>"011000010",
        10435=>"000000011",
        10436=>"011011000",
        10437=>"010001000",
        10438=>"011010000",
        10439=>"100000000",
        10440=>"001001000",
        10441=>"110110000",
        10442=>"011011001",
        10443=>"000100010",
        10444=>"000011000",
        10445=>"011001010",
        10446=>"001011001",
        10447=>"011011001",
        10448=>"001001001",
        10449=>"011100110",
        10450=>"000000100",
        10451=>"100110110",
        10452=>"001001001",
        10453=>"100100100",
        10454=>"111001000",
        10455=>"011011011",
        10456=>"001111011",
        10457=>"011011011",
        10458=>"010100111",
        10459=>"011000000",
        10460=>"111011001",
        10461=>"100110110",
        10462=>"100100100",
        10463=>"111101101",
        10464=>"011000000",
        10465=>"011011001",
        10466=>"011001001",
        10467=>"001011001",
        10468=>"011011011",
        10469=>"011001010",
        10470=>"010000100",
        10471=>"011011000",
        10472=>"100100100",
        10473=>"100010110",
        10474=>"011011001",
        10475=>"100010100",
        10476=>"011011011",
        10477=>"100100110",
        10478=>"000000010",
        10479=>"101001001",
        10480=>"001001001",
        10481=>"001001100",
        10482=>"000000111",
        10483=>"100100110",
        10484=>"100100100",
        10485=>"000100111",
        10486=>"110110110",
        10487=>"001011011",
        10488=>"111011011",
        10489=>"000100000",
        10490=>"000100110",
        10491=>"001000101",
        10492=>"100011000",
        10493=>"110110111",
        10494=>"111111100",
        10495=>"010001111",
        10496=>"111011110",
        10497=>"111000011",
        10498=>"110101101",
        10499=>"000100000",
        10500=>"101100110",
        10501=>"110110001",
        10502=>"111010110",
        10503=>"010010011",
        10504=>"111001001",
        10505=>"000100000",
        10506=>"111011010",
        10507=>"001000000",
        10508=>"111001000",
        10509=>"111110110",
        10510=>"111000001",
        10511=>"000000011",
        10512=>"100100100",
        10513=>"000010000",
        10514=>"000101101",
        10515=>"000111111",
        10516=>"000111000",
        10517=>"001001001",
        10518=>"000000010",
        10519=>"000110010",
        10520=>"001110111",
        10521=>"000010001",
        10522=>"101101011",
        10523=>"111111011",
        10524=>"111100110",
        10525=>"101101101",
        10526=>"100000100",
        10527=>"110111110",
        10528=>"001111111",
        10529=>"111111000",
        10530=>"110110000",
        10531=>"100110011",
        10532=>"001111010",
        10533=>"000001111",
        10534=>"111111111",
        10535=>"101001111",
        10536=>"101010000",
        10537=>"001111111",
        10538=>"111111110",
        10539=>"011010100",
        10540=>"110110000",
        10541=>"101101000",
        10542=>"000000000",
        10543=>"100111111",
        10544=>"011111111",
        10545=>"000011101",
        10546=>"100111100",
        10547=>"001001000",
        10548=>"010000000",
        10549=>"001000000",
        10550=>"000010110",
        10551=>"110000111",
        10552=>"001010110",
        10553=>"000010110",
        10554=>"000001000",
        10555=>"000000000",
        10556=>"000000100",
        10557=>"110010010",
        10558=>"110111110",
        10559=>"010101111",
        10560=>"110001100",
        10561=>"111110000",
        10562=>"110111010",
        10563=>"000000010",
        10564=>"000101000",
        10565=>"010010001",
        10566=>"101111110",
        10567=>"000010010",
        10568=>"000001001",
        10569=>"111101101",
        10570=>"110110110",
        10571=>"000111111",
        10572=>"000101000",
        10573=>"001000000",
        10574=>"100000000",
        10575=>"111000110",
        10576=>"011000011",
        10577=>"011000110",
        10578=>"100110000",
        10579=>"011000111",
        10580=>"010010000",
        10581=>"000000111",
        10582=>"111111110",
        10583=>"010110100",
        10584=>"100101100",
        10585=>"000000001",
        10586=>"001011110",
        10587=>"000000110",
        10588=>"110001001",
        10589=>"000100101",
        10590=>"111001011",
        10591=>"101001111",
        10592=>"111100100",
        10593=>"100001001",
        10594=>"111101111",
        10595=>"000010110",
        10596=>"110010010",
        10597=>"100101000",
        10598=>"100000101",
        10599=>"101110011",
        10600=>"100000011",
        10601=>"100100111",
        10602=>"010001001",
        10603=>"000000001",
        10604=>"000000000",
        10605=>"001000111",
        10606=>"000001101",
        10607=>"111101001",
        10608=>"000000101",
        10609=>"100011111",
        10610=>"000000000",
        10611=>"101101100",
        10612=>"001001111",
        10613=>"100000000",
        10614=>"001001010",
        10615=>"000011011",
        10616=>"010100110",
        10617=>"000010010",
        10618=>"011000100",
        10619=>"000000001",
        10620=>"110100100",
        10621=>"010110010",
        10622=>"000000100",
        10623=>"011111000",
        10624=>"010100000",
        10625=>"000100101",
        10626=>"011101001",
        10627=>"111101111",
        10628=>"100010001",
        10629=>"111110110",
        10630=>"111101010",
        10631=>"101001100",
        10632=>"101111100",
        10633=>"101000100",
        10634=>"000000000",
        10635=>"101000111",
        10636=>"101101111",
        10637=>"111111111",
        10638=>"001011001",
        10639=>"000001000",
        10640=>"100101100",
        10641=>"000000000",
        10642=>"111100100",
        10643=>"101100100",
        10644=>"000010000",
        10645=>"011000001",
        10646=>"101000000",
        10647=>"101000011",
        10648=>"011001110",
        10649=>"111001111",
        10650=>"000000001",
        10651=>"001000010",
        10652=>"110111111",
        10653=>"111001110",
        10654=>"111111011",
        10655=>"011001001",
        10656=>"010000100",
        10657=>"000010001",
        10658=>"011011111",
        10659=>"111100010",
        10660=>"010000111",
        10661=>"101000010",
        10662=>"000000111",
        10663=>"101101101",
        10664=>"101001011",
        10665=>"111101100",
        10666=>"110100010",
        10667=>"000011011",
        10668=>"000100110",
        10669=>"011101000",
        10670=>"111010000",
        10671=>"111101000",
        10672=>"010110111",
        10673=>"111001101",
        10674=>"011101101",
        10675=>"111000100",
        10676=>"111111100",
        10677=>"100000110",
        10678=>"001000000",
        10679=>"010100000",
        10680=>"101000101",
        10681=>"111001000",
        10682=>"111000111",
        10683=>"111001111",
        10684=>"111000101",
        10685=>"010011000",
        10686=>"000000111",
        10687=>"000010000",
        10688=>"111001011",
        10689=>"111001011",
        10690=>"000001001",
        10691=>"110011010",
        10692=>"111000010",
        10693=>"011011111",
        10694=>"111000001",
        10695=>"001010010",
        10696=>"001000000",
        10697=>"000010010",
        10698=>"101001011",
        10699=>"110000000",
        10700=>"010101000",
        10701=>"111111001",
        10702=>"100111001",
        10703=>"111101111",
        10704=>"111000001",
        10705=>"000001001",
        10706=>"000101001",
        10707=>"011100000",
        10708=>"111110111",
        10709=>"001000000",
        10710=>"110101111",
        10711=>"111000000",
        10712=>"011000011",
        10713=>"001000001",
        10714=>"000001101",
        10715=>"000000000",
        10716=>"100100001",
        10717=>"000000001",
        10718=>"000000101",
        10719=>"111100000",
        10720=>"111101001",
        10721=>"001000010",
        10722=>"111001001",
        10723=>"010000000",
        10724=>"001000010",
        10725=>"000000100",
        10726=>"011100100",
        10727=>"001000111",
        10728=>"000000000",
        10729=>"000110101",
        10730=>"111100000",
        10731=>"111010101",
        10732=>"000100000",
        10733=>"100000111",
        10734=>"000110110",
        10735=>"111100100",
        10736=>"110000000",
        10737=>"011011001",
        10738=>"011101101",
        10739=>"001001001",
        10740=>"010111010",
        10741=>"000000000",
        10742=>"011101111",
        10743=>"010001101",
        10744=>"000000001",
        10745=>"000000010",
        10746=>"100000000",
        10747=>"101101001",
        10748=>"010001001",
        10749=>"000000000",
        10750=>"000001000",
        10751=>"111111010",
        10752=>"111111110",
        10753=>"000000000",
        10754=>"000000000",
        10755=>"111001000",
        10756=>"011111111",
        10757=>"111111111",
        10758=>"001000010",
        10759=>"111111111",
        10760=>"011111111",
        10761=>"111111100",
        10762=>"111111110",
        10763=>"100011100",
        10764=>"000000000",
        10765=>"010111110",
        10766=>"101001001",
        10767=>"000000001",
        10768=>"001000000",
        10769=>"001101101",
        10770=>"111011101",
        10771=>"110110100",
        10772=>"000010000",
        10773=>"000111011",
        10774=>"011011101",
        10775=>"111000000",
        10776=>"100101101",
        10777=>"000000000",
        10778=>"000000000",
        10779=>"001010110",
        10780=>"000010000",
        10781=>"000101001",
        10782=>"000101100",
        10783=>"000000000",
        10784=>"010000110",
        10785=>"000000000",
        10786=>"011011100",
        10787=>"000000000",
        10788=>"000000000",
        10789=>"010111111",
        10790=>"010111110",
        10791=>"011111001",
        10792=>"100000101",
        10793=>"000100000",
        10794=>"111000010",
        10795=>"100100101",
        10796=>"111011000",
        10797=>"011001000",
        10798=>"111110010",
        10799=>"001000000",
        10800=>"011111111",
        10801=>"011111111",
        10802=>"011100111",
        10803=>"111100000",
        10804=>"110110110",
        10805=>"000000101",
        10806=>"011111111",
        10807=>"010111111",
        10808=>"000000111",
        10809=>"000000000",
        10810=>"011011011",
        10811=>"111111111",
        10812=>"001111000",
        10813=>"010010000",
        10814=>"111010010",
        10815=>"111011111",
        10816=>"111111000",
        10817=>"000000000",
        10818=>"000010111",
        10819=>"101001000",
        10820=>"000000000",
        10821=>"100000001",
        10822=>"000000000",
        10823=>"111000000",
        10824=>"000000000",
        10825=>"010111111",
        10826=>"111111101",
        10827=>"000001101",
        10828=>"000000000",
        10829=>"000010010",
        10830=>"000000000",
        10831=>"010111011",
        10832=>"001101111",
        10833=>"000000001",
        10834=>"000011111",
        10835=>"000010110",
        10836=>"000000110",
        10837=>"111111111",
        10838=>"101111011",
        10839=>"101111000",
        10840=>"110111011",
        10841=>"110111101",
        10842=>"001001000",
        10843=>"111111111",
        10844=>"100100001",
        10845=>"000000000",
        10846=>"100100000",
        10847=>"111111111",
        10848=>"011101101",
        10849=>"111111111",
        10850=>"101101111",
        10851=>"111011111",
        10852=>"000001110",
        10853=>"111111100",
        10854=>"001101100",
        10855=>"111111111",
        10856=>"000000000",
        10857=>"000000101",
        10858=>"100111001",
        10859=>"111000101",
        10860=>"101001101",
        10861=>"000110000",
        10862=>"110100000",
        10863=>"100101101",
        10864=>"000010111",
        10865=>"001000110",
        10866=>"100000000",
        10867=>"010111111",
        10868=>"010111111",
        10869=>"010100001",
        10870=>"000000000",
        10871=>"100111111",
        10872=>"011000010",
        10873=>"010000000",
        10874=>"000000000",
        10875=>"111000000",
        10876=>"000000000",
        10877=>"000000010",
        10878=>"111010110",
        10879=>"110111010",
        10880=>"011011011",
        10881=>"110110000",
        10882=>"000110100",
        10883=>"100111111",
        10884=>"110110110",
        10885=>"111011010",
        10886=>"011011011",
        10887=>"100100100",
        10888=>"011011111",
        10889=>"000000111",
        10890=>"110100000",
        10891=>"001100110",
        10892=>"110001011",
        10893=>"100100100",
        10894=>"001000010",
        10895=>"100100100",
        10896=>"000001100",
        10897=>"111001111",
        10898=>"000010001",
        10899=>"000001001",
        10900=>"001001001",
        10901=>"010000100",
        10902=>"000001001",
        10903=>"100100101",
        10904=>"000000101",
        10905=>"001111110",
        10906=>"100110110",
        10907=>"000111011",
        10908=>"010111100",
        10909=>"011011010",
        10910=>"111011011",
        10911=>"011110110",
        10912=>"101110100",
        10913=>"101000100",
        10914=>"001000000",
        10915=>"111010111",
        10916=>"001001011",
        10917=>"001001000",
        10918=>"110100000",
        10919=>"001001011",
        10920=>"000110110",
        10921=>"000010111",
        10922=>"011010000",
        10923=>"000000001",
        10924=>"110010100",
        10925=>"110110110",
        10926=>"011001011",
        10927=>"100101100",
        10928=>"000000100",
        10929=>"100100100",
        10930=>"111110101",
        10931=>"100001001",
        10932=>"000000000",
        10933=>"000000000",
        10934=>"110110100",
        10935=>"010000100",
        10936=>"010111110",
        10937=>"111110010",
        10938=>"001011001",
        10939=>"100100100",
        10940=>"110110000",
        10941=>"000001011",
        10942=>"111000000",
        10943=>"000001010",
        10944=>"010011101",
        10945=>"100110001",
        10946=>"100100100",
        10947=>"110011011",
        10948=>"011011111",
        10949=>"000011011",
        10950=>"000001110",
        10951=>"001100100",
        10952=>"100001011",
        10953=>"000000000",
        10954=>"110110100",
        10955=>"000000001",
        10956=>"111111110",
        10957=>"000110111",
        10958=>"010001011",
        10959=>"001100100",
        10960=>"100110100",
        10961=>"001001010",
        10962=>"100110100",
        10963=>"111001001",
        10964=>"011001000",
        10965=>"100000100",
        10966=>"001001011",
        10967=>"011001000",
        10968=>"011010000",
        10969=>"000000001",
        10970=>"000100101",
        10971=>"001001000",
        10972=>"001011111",
        10973=>"110001001",
        10974=>"000110100",
        10975=>"110001101",
        10976=>"000000001",
        10977=>"011000000",
        10978=>"101100110",
        10979=>"001011011",
        10980=>"101110000",
        10981=>"010110100",
        10982=>"010001000",
        10983=>"111110110",
        10984=>"111011101",
        10985=>"000110100",
        10986=>"001011011",
        10987=>"101001100",
        10988=>"001100100",
        10989=>"100000001",
        10990=>"000101010",
        10991=>"001001011",
        10992=>"101100110",
        10993=>"110000000",
        10994=>"101111011",
        10995=>"101111111",
        10996=>"110100100",
        10997=>"110110111",
        10998=>"111111000",
        10999=>"110100101",
        11000=>"110100000",
        11001=>"100110100",
        11002=>"001010110",
        11003=>"110100100",
        11004=>"111111011",
        11005=>"000000110",
        11006=>"100110111",
        11007=>"001010100",
        11008=>"011001000",
        11009=>"111000010",
        11010=>"111111111",
        11011=>"111111111",
        11012=>"000000000",
        11013=>"000000000",
        11014=>"101111111",
        11015=>"000010110",
        11016=>"100100001",
        11017=>"111101100",
        11018=>"001100101",
        11019=>"110101101",
        11020=>"000101001",
        11021=>"100000000",
        11022=>"000000000",
        11023=>"110010000",
        11024=>"110100111",
        11025=>"011111111",
        11026=>"011111111",
        11027=>"100000001",
        11028=>"110111010",
        11029=>"101000000",
        11030=>"000000000",
        11031=>"000000000",
        11032=>"100101111",
        11033=>"110101001",
        11034=>"110101111",
        11035=>"011000110",
        11036=>"000000000",
        11037=>"000100101",
        11038=>"011101101",
        11039=>"000100000",
        11040=>"110001000",
        11041=>"101101101",
        11042=>"011101101",
        11043=>"111111110",
        11044=>"100011011",
        11045=>"011111110",
        11046=>"101101111",
        11047=>"000000000",
        11048=>"111101111",
        11049=>"111101111",
        11050=>"000000010",
        11051=>"000101101",
        11052=>"010001001",
        11053=>"010010111",
        11054=>"000000000",
        11055=>"101100100",
        11056=>"100111010",
        11057=>"111111111",
        11058=>"111101111",
        11059=>"101011101",
        11060=>"000000001",
        11061=>"000000000",
        11062=>"000000100",
        11063=>"000000000",
        11064=>"110000000",
        11065=>"101000000",
        11066=>"011010000",
        11067=>"010010000",
        11068=>"101000000",
        11069=>"100011010",
        11070=>"110111101",
        11071=>"010101000",
        11072=>"111111111",
        11073=>"111111011",
        11074=>"000000000",
        11075=>"000000000",
        11076=>"110001000",
        11077=>"011111111",
        11078=>"100100110",
        11079=>"110111111",
        11080=>"001000110",
        11081=>"000000000",
        11082=>"000000000",
        11083=>"011111111",
        11084=>"011111111",
        11085=>"111111111",
        11086=>"000111111",
        11087=>"111110000",
        11088=>"000011011",
        11089=>"111000000",
        11090=>"000101111",
        11091=>"000000000",
        11092=>"100110111",
        11093=>"000000000",
        11094=>"000111000",
        11095=>"000000000",
        11096=>"010111110",
        11097=>"100111101",
        11098=>"001001011",
        11099=>"101111010",
        11100=>"000101111",
        11101=>"001000000",
        11102=>"001101111",
        11103=>"110100000",
        11104=>"010100100",
        11105=>"001111101",
        11106=>"000110000",
        11107=>"111001000",
        11108=>"111101111",
        11109=>"111110111",
        11110=>"001000100",
        11111=>"111111001",
        11112=>"111100100",
        11113=>"100100101",
        11114=>"110101111",
        11115=>"110101000",
        11116=>"000000000",
        11117=>"111111011",
        11118=>"111010011",
        11119=>"000000000",
        11120=>"000000000",
        11121=>"111110011",
        11122=>"010011111",
        11123=>"000000101",
        11124=>"110100000",
        11125=>"001001000",
        11126=>"000000111",
        11127=>"011111011",
        11128=>"111001100",
        11129=>"000000111",
        11130=>"111100100",
        11131=>"000100101",
        11132=>"010110110",
        11133=>"110000010",
        11134=>"111111111",
        11135=>"110111111",
        11136=>"010010111",
        11137=>"000110110",
        11138=>"110100000",
        11139=>"001001111",
        11140=>"011000110",
        11141=>"000010111",
        11142=>"010110010",
        11143=>"111101000",
        11144=>"101100000",
        11145=>"110000000",
        11146=>"101010011",
        11147=>"101000001",
        11148=>"110000101",
        11149=>"111010111",
        11150=>"000100010",
        11151=>"101100100",
        11152=>"111100110",
        11153=>"000000011",
        11154=>"011000000",
        11155=>"000010110",
        11156=>"000011111",
        11157=>"011000100",
        11158=>"000000100",
        11159=>"110100100",
        11160=>"101001000",
        11161=>"111010100",
        11162=>"000110111",
        11163=>"100011101",
        11164=>"000011000",
        11165=>"000000111",
        11166=>"001110010",
        11167=>"010111101",
        11168=>"001010000",
        11169=>"000000000",
        11170=>"001011111",
        11171=>"111110001",
        11172=>"011100000",
        11173=>"000000011",
        11174=>"111101111",
        11175=>"111100100",
        11176=>"001101000",
        11177=>"111111100",
        11178=>"000010111",
        11179=>"111111111",
        11180=>"000011110",
        11181=>"111101000",
        11182=>"000110101",
        11183=>"110101111",
        11184=>"011001000",
        11185=>"000000001",
        11186=>"100110101",
        11187=>"011111100",
        11188=>"000111111",
        11189=>"000000110",
        11190=>"111000110",
        11191=>"111000110",
        11192=>"111111111",
        11193=>"111101011",
        11194=>"001000100",
        11195=>"000000111",
        11196=>"000000011",
        11197=>"000000000",
        11198=>"110101000",
        11199=>"000111111",
        11200=>"000011011",
        11201=>"100100100",
        11202=>"111100101",
        11203=>"010100010",
        11204=>"111010000",
        11205=>"110001000",
        11206=>"000000011",
        11207=>"111010000",
        11208=>"010010111",
        11209=>"011011011",
        11210=>"011111111",
        11211=>"010000000",
        11212=>"000000010",
        11213=>"111100000",
        11214=>"011000000",
        11215=>"111100000",
        11216=>"000000000",
        11217=>"000001001",
        11218=>"000110111",
        11219=>"000010011",
        11220=>"111010011",
        11221=>"000000001",
        11222=>"100110011",
        11223=>"111001000",
        11224=>"011000001",
        11225=>"000000010",
        11226=>"101101000",
        11227=>"111100000",
        11228=>"100000001",
        11229=>"000100011",
        11230=>"001100110",
        11231=>"011000100",
        11232=>"001011110",
        11233=>"011111000",
        11234=>"110110101",
        11235=>"110000000",
        11236=>"100111000",
        11237=>"000101101",
        11238=>"000000100",
        11239=>"111101000",
        11240=>"000101111",
        11241=>"100000000",
        11242=>"110111111",
        11243=>"100100010",
        11244=>"111111011",
        11245=>"111100001",
        11246=>"010000100",
        11247=>"000010000",
        11248=>"010000001",
        11249=>"111011100",
        11250=>"111100100",
        11251=>"000000111",
        11252=>"000000000",
        11253=>"111101101",
        11254=>"111111100",
        11255=>"011000000",
        11256=>"000001111",
        11257=>"100000111",
        11258=>"000100011",
        11259=>"111100000",
        11260=>"000001001",
        11261=>"000001011",
        11262=>"111100100",
        11263=>"101110110",
        11264=>"010000000",
        11265=>"000000000",
        11266=>"000000000",
        11267=>"000111000",
        11268=>"000001000",
        11269=>"000010111",
        11270=>"100101011",
        11271=>"101000000",
        11272=>"011111111",
        11273=>"001011111",
        11274=>"011100000",
        11275=>"010111111",
        11276=>"111001101",
        11277=>"000111110",
        11278=>"100001101",
        11279=>"001001000",
        11280=>"110100001",
        11281=>"000101011",
        11282=>"101000000",
        11283=>"000000000",
        11284=>"000101001",
        11285=>"111000001",
        11286=>"000000000",
        11287=>"100001010",
        11288=>"011000000",
        11289=>"010100110",
        11290=>"111000010",
        11291=>"111101100",
        11292=>"011111111",
        11293=>"110110010",
        11294=>"101001110",
        11295=>"110001000",
        11296=>"110110111",
        11297=>"111000100",
        11298=>"110110111",
        11299=>"111111110",
        11300=>"001111111",
        11301=>"110111001",
        11302=>"010110110",
        11303=>"100001000",
        11304=>"011100001",
        11305=>"000000000",
        11306=>"111111111",
        11307=>"100101101",
        11308=>"111111101",
        11309=>"000000000",
        11310=>"110110111",
        11311=>"000100000",
        11312=>"000100000",
        11313=>"000000000",
        11314=>"010111110",
        11315=>"000000000",
        11316=>"011111110",
        11317=>"111111111",
        11318=>"110110111",
        11319=>"111110111",
        11320=>"010000000",
        11321=>"000000000",
        11322=>"110110111",
        11323=>"000001111",
        11324=>"010000000",
        11325=>"010100001",
        11326=>"111000001",
        11327=>"000101111",
        11328=>"101101111",
        11329=>"000000000",
        11330=>"000011111",
        11331=>"101101000",
        11332=>"110111011",
        11333=>"110111100",
        11334=>"000101100",
        11335=>"110111101",
        11336=>"011000000",
        11337=>"000110111",
        11338=>"001101110",
        11339=>"111101111",
        11340=>"011100001",
        11341=>"001111101",
        11342=>"001001000",
        11343=>"000000000",
        11344=>"010000000",
        11345=>"100000000",
        11346=>"110111111",
        11347=>"111111111",
        11348=>"011111111",
        11349=>"000010000",
        11350=>"111001000",
        11351=>"001100111",
        11352=>"101110100",
        11353=>"000011111",
        11354=>"101000111",
        11355=>"000000011",
        11356=>"101000110",
        11357=>"100100000",
        11358=>"110100000",
        11359=>"011111111",
        11360=>"110110111",
        11361=>"000001000",
        11362=>"000000000",
        11363=>"000000000",
        11364=>"010000000",
        11365=>"111000000",
        11366=>"000000000",
        11367=>"000010000",
        11368=>"110100001",
        11369=>"110000000",
        11370=>"011001010",
        11371=>"111110111",
        11372=>"000000000",
        11373=>"000000000",
        11374=>"000000001",
        11375=>"111100111",
        11376=>"001000000",
        11377=>"001000000",
        11378=>"000000000",
        11379=>"000110000",
        11380=>"000011011",
        11381=>"000000000",
        11382=>"111011111",
        11383=>"011111111",
        11384=>"000000110",
        11385=>"111000000",
        11386=>"111001100",
        11387=>"111111111",
        11388=>"001001111",
        11389=>"010111100",
        11390=>"010100010",
        11391=>"111111110",
        11392=>"101110010",
        11393=>"101101111",
        11394=>"000000111",
        11395=>"101111111",
        11396=>"001100111",
        11397=>"011000000",
        11398=>"111000000",
        11399=>"001000000",
        11400=>"100000000",
        11401=>"000000000",
        11402=>"100011001",
        11403=>"000001001",
        11404=>"010010100",
        11405=>"111111110",
        11406=>"001011000",
        11407=>"000001001",
        11408=>"111110111",
        11409=>"110000111",
        11410=>"100111100",
        11411=>"100001011",
        11412=>"110000000",
        11413=>"111000000",
        11414=>"100100111",
        11415=>"110110111",
        11416=>"011111011",
        11417=>"100010100",
        11418=>"000100101",
        11419=>"011101111",
        11420=>"000000000",
        11421=>"000000001",
        11422=>"111111111",
        11423=>"111111001",
        11424=>"101110000",
        11425=>"111110110",
        11426=>"000010000",
        11427=>"000000000",
        11428=>"111010011",
        11429=>"110101111",
        11430=>"000000000",
        11431=>"001001101",
        11432=>"110111111",
        11433=>"000000000",
        11434=>"111111111",
        11435=>"101100100",
        11436=>"010001101",
        11437=>"001000000",
        11438=>"000000011",
        11439=>"000000000",
        11440=>"000000000",
        11441=>"111111110",
        11442=>"110011000",
        11443=>"101001111",
        11444=>"000001101",
        11445=>"100000000",
        11446=>"111111100",
        11447=>"011111110",
        11448=>"001000001",
        11449=>"100010110",
        11450=>"000000010",
        11451=>"010000101",
        11452=>"000000000",
        11453=>"000000000",
        11454=>"110101101",
        11455=>"111100110",
        11456=>"111101110",
        11457=>"011110011",
        11458=>"111111001",
        11459=>"010110000",
        11460=>"110110111",
        11461=>"110110110",
        11462=>"011000100",
        11463=>"011111011",
        11464=>"111011001",
        11465=>"111111111",
        11466=>"011010001",
        11467=>"110101101",
        11468=>"110111111",
        11469=>"010000000",
        11470=>"000011010",
        11471=>"111110100",
        11472=>"101000011",
        11473=>"100001111",
        11474=>"111111000",
        11475=>"101101111",
        11476=>"001011011",
        11477=>"111000111",
        11478=>"111111111",
        11479=>"000100001",
        11480=>"001000000",
        11481=>"000101010",
        11482=>"000000011",
        11483=>"010001111",
        11484=>"110001001",
        11485=>"001100000",
        11486=>"001100011",
        11487=>"000000111",
        11488=>"010000000",
        11489=>"101101111",
        11490=>"000000000",
        11491=>"111000000",
        11492=>"011110101",
        11493=>"000000000",
        11494=>"110100100",
        11495=>"000000100",
        11496=>"110100000",
        11497=>"000000101",
        11498=>"101100100",
        11499=>"110001111",
        11500=>"101101111",
        11501=>"101000001",
        11502=>"111011101",
        11503=>"001101101",
        11504=>"010000000",
        11505=>"000000000",
        11506=>"100000110",
        11507=>"000001101",
        11508=>"000100000",
        11509=>"110000011",
        11510=>"010111010",
        11511=>"000111011",
        11512=>"001000100",
        11513=>"000010000",
        11514=>"110000000",
        11515=>"000000000",
        11516=>"000000100",
        11517=>"011111001",
        11518=>"101111110",
        11519=>"001010000",
        11520=>"011011111",
        11521=>"110100111",
        11522=>"100110111",
        11523=>"011111111",
        11524=>"000111011",
        11525=>"001000000",
        11526=>"000010011",
        11527=>"100101001",
        11528=>"011000000",
        11529=>"000000011",
        11530=>"101101011",
        11531=>"011000111",
        11532=>"001101000",
        11533=>"101101100",
        11534=>"001000000",
        11535=>"100100110",
        11536=>"001001000",
        11537=>"100100000",
        11538=>"111111100",
        11539=>"111000011",
        11540=>"110000001",
        11541=>"000000001",
        11542=>"100100110",
        11543=>"001010011",
        11544=>"011100000",
        11545=>"011001000",
        11546=>"001001001",
        11547=>"001111011",
        11548=>"001111010",
        11549=>"001001000",
        11550=>"100001001",
        11551=>"111101110",
        11552=>"011011001",
        11553=>"111111001",
        11554=>"001100100",
        11555=>"000000000",
        11556=>"011011110",
        11557=>"111111110",
        11558=>"100110011",
        11559=>"010100010",
        11560=>"001000000",
        11561=>"011001001",
        11562=>"011000001",
        11563=>"011000001",
        11564=>"101011111",
        11565=>"100100111",
        11566=>"001000011",
        11567=>"110110110",
        11568=>"001011001",
        11569=>"100110110",
        11570=>"001011111",
        11571=>"111011101",
        11572=>"001001001",
        11573=>"011001001",
        11574=>"001001000",
        11575=>"100100110",
        11576=>"100100110",
        11577=>"001011111",
        11578=>"001011001",
        11579=>"110100111",
        11580=>"101110011",
        11581=>"010010010",
        11582=>"000000011",
        11583=>"011101101",
        11584=>"011001110",
        11585=>"011000000",
        11586=>"001001001",
        11587=>"100100000",
        11588=>"010010111",
        11589=>"100011000",
        11590=>"100110010",
        11591=>"011011000",
        11592=>"011001000",
        11593=>"101110000",
        11594=>"100001011",
        11595=>"000110000",
        11596=>"011001001",
        11597=>"101111111",
        11598=>"111011001",
        11599=>"100110110",
        11600=>"000100110",
        11601=>"011100011",
        11602=>"001000001",
        11603=>"011011001",
        11604=>"101100101",
        11605=>"100100110",
        11606=>"100010111",
        11607=>"101100100",
        11608=>"001111101",
        11609=>"011011110",
        11610=>"100000000",
        11611=>"100110100",
        11612=>"010000000",
        11613=>"100110010",
        11614=>"100100100",
        11615=>"100110010",
        11616=>"000010001",
        11617=>"000001010",
        11618=>"100100111",
        11619=>"000111011",
        11620=>"011001011",
        11621=>"000001001",
        11622=>"000000110",
        11623=>"011011001",
        11624=>"100001000",
        11625=>"100100010",
        11626=>"111000001",
        11627=>"011000110",
        11628=>"000100100",
        11629=>"000100010",
        11630=>"110011111",
        11631=>"101111111",
        11632=>"001100111",
        11633=>"000011011",
        11634=>"011100000",
        11635=>"000010010",
        11636=>"110110111",
        11637=>"011000101",
        11638=>"100001001",
        11639=>"011011011",
        11640=>"001000110",
        11641=>"010001001",
        11642=>"111100100",
        11643=>"110011011",
        11644=>"110100101",
        11645=>"011011111",
        11646=>"001101110",
        11647=>"010111001",
        11648=>"111111111",
        11649=>"111111111",
        11650=>"110111010",
        11651=>"000000000",
        11652=>"111001100",
        11653=>"001001111",
        11654=>"010111010",
        11655=>"000000100",
        11656=>"100100100",
        11657=>"000000001",
        11658=>"111111001",
        11659=>"000000100",
        11660=>"111111110",
        11661=>"101101000",
        11662=>"111101100",
        11663=>"101111101",
        11664=>"000000000",
        11665=>"111101111",
        11666=>"111111110",
        11667=>"111111101",
        11668=>"001001000",
        11669=>"000111111",
        11670=>"000000000",
        11671=>"111111110",
        11672=>"111101001",
        11673=>"000000001",
        11674=>"100000000",
        11675=>"000000000",
        11676=>"111111111",
        11677=>"011011110",
        11678=>"000100111",
        11679=>"111111000",
        11680=>"000000000",
        11681=>"111101100",
        11682=>"000000000",
        11683=>"000110100",
        11684=>"010000111",
        11685=>"101111111",
        11686=>"101001001",
        11687=>"111000000",
        11688=>"111100111",
        11689=>"111011101",
        11690=>"001000000",
        11691=>"110110110",
        11692=>"000101100",
        11693=>"000110110",
        11694=>"000000000",
        11695=>"100101111",
        11696=>"000000000",
        11697=>"110100010",
        11698=>"000000000",
        11699=>"100101001",
        11700=>"100000000",
        11701=>"000000101",
        11702=>"101111111",
        11703=>"000000111",
        11704=>"111111111",
        11705=>"111100001",
        11706=>"000000100",
        11707=>"000000000",
        11708=>"111111111",
        11709=>"000000010",
        11710=>"000000000",
        11711=>"101010101",
        11712=>"000101100",
        11713=>"110110000",
        11714=>"111101001",
        11715=>"111101110",
        11716=>"000000000",
        11717=>"100000000",
        11718=>"001101000",
        11719=>"110101111",
        11720=>"000000000",
        11721=>"111000000",
        11722=>"001111111",
        11723=>"000101000",
        11724=>"111000000",
        11725=>"000000001",
        11726=>"110110011",
        11727=>"010000010",
        11728=>"111111010",
        11729=>"001111111",
        11730=>"100100101",
        11731=>"110111101",
        11732=>"000010010",
        11733=>"000000110",
        11734=>"000100000",
        11735=>"000110111",
        11736=>"100111111",
        11737=>"000000101",
        11738=>"000001100",
        11739=>"010110100",
        11740=>"101001101",
        11741=>"100101111",
        11742=>"111111111",
        11743=>"111111111",
        11744=>"011001001",
        11745=>"001000001",
        11746=>"111111110",
        11747=>"111111111",
        11748=>"000000011",
        11749=>"011111010",
        11750=>"000011011",
        11751=>"111000000",
        11752=>"000000000",
        11753=>"000000100",
        11754=>"111011011",
        11755=>"010101101",
        11756=>"000110111",
        11757=>"110100111",
        11758=>"111011111",
        11759=>"111101101",
        11760=>"111111010",
        11761=>"111111111",
        11762=>"111111000",
        11763=>"000010111",
        11764=>"000111010",
        11765=>"000000111",
        11766=>"000000000",
        11767=>"000000000",
        11768=>"110110111",
        11769=>"010111111",
        11770=>"000000000",
        11771=>"001111111",
        11772=>"111111100",
        11773=>"111011111",
        11774=>"100111011",
        11775=>"111101101",
        11776=>"000010000",
        11777=>"111010100",
        11778=>"110010001",
        11779=>"100111110",
        11780=>"111000000",
        11781=>"111110110",
        11782=>"000011110",
        11783=>"111010010",
        11784=>"100101100",
        11785=>"111000000",
        11786=>"011001100",
        11787=>"111011000",
        11788=>"011001011",
        11789=>"111011111",
        11790=>"000000011",
        11791=>"000001111",
        11792=>"011001000",
        11793=>"000110100",
        11794=>"000001000",
        11795=>"000100111",
        11796=>"111111100",
        11797=>"011111010",
        11798=>"010100100",
        11799=>"000001111",
        11800=>"000001001",
        11801=>"000001011",
        11802=>"000100101",
        11803=>"110000000",
        11804=>"110000000",
        11805=>"000001011",
        11806=>"111001100",
        11807=>"101001100",
        11808=>"011110000",
        11809=>"000010000",
        11810=>"000000011",
        11811=>"001000011",
        11812=>"111011000",
        11813=>"101110100",
        11814=>"001010011",
        11815=>"110110100",
        11816=>"001111110",
        11817=>"001001011",
        11818=>"000100111",
        11819=>"000001001",
        11820=>"111001000",
        11821=>"011011010",
        11822=>"111001111",
        11823=>"101010100",
        11824=>"110001001",
        11825=>"111110100",
        11826=>"111011000",
        11827=>"010011011",
        11828=>"100001011",
        11829=>"000001000",
        11830=>"000001100",
        11831=>"011110111",
        11832=>"000100110",
        11833=>"111001000",
        11834=>"000000110",
        11835=>"000100000",
        11836=>"110110001",
        11837=>"011010100",
        11838=>"101001000",
        11839=>"010100101",
        11840=>"100110110",
        11841=>"001000001",
        11842=>"110001011",
        11843=>"110000101",
        11844=>"010001111",
        11845=>"000011111",
        11846=>"101111111",
        11847=>"000000000",
        11848=>"000001011",
        11849=>"100111001",
        11850=>"111001001",
        11851=>"000100000",
        11852=>"001110001",
        11853=>"110000000",
        11854=>"001000111",
        11855=>"100110000",
        11856=>"110010010",
        11857=>"110110001",
        11858=>"100001001",
        11859=>"111110110",
        11860=>"000100000",
        11861=>"010100000",
        11862=>"000001001",
        11863=>"111101110",
        11864=>"111000010",
        11865=>"001000000",
        11866=>"111110000",
        11867=>"111111000",
        11868=>"000000110",
        11869=>"111010000",
        11870=>"101111110",
        11871=>"000010000",
        11872=>"011100000",
        11873=>"000000111",
        11874=>"111111110",
        11875=>"000000100",
        11876=>"000001011",
        11877=>"000111110",
        11878=>"000100100",
        11879=>"011001100",
        11880=>"000011111",
        11881=>"100000000",
        11882=>"000100111",
        11883=>"111101110",
        11884=>"101110100",
        11885=>"001110000",
        11886=>"100111111",
        11887=>"100101000",
        11888=>"000001000",
        11889=>"111000101",
        11890=>"011011100",
        11891=>"001011000",
        11892=>"100110111",
        11893=>"000100110",
        11894=>"001110110",
        11895=>"000011111",
        11896=>"011011101",
        11897=>"000000110",
        11898=>"111100000",
        11899=>"001001111",
        11900=>"100100100",
        11901=>"001001111",
        11902=>"111001100",
        11903=>"111101101",
        11904=>"111001001",
        11905=>"101000110",
        11906=>"110000000",
        11907=>"010111000",
        11908=>"100100100",
        11909=>"001111111",
        11910=>"100000000",
        11911=>"111000001",
        11912=>"100100100",
        11913=>"100001111",
        11914=>"101001111",
        11915=>"011000100",
        11916=>"000000000",
        11917=>"110111110",
        11918=>"100001001",
        11919=>"110000101",
        11920=>"100000000",
        11921=>"111000000",
        11922=>"101011000",
        11923=>"001101001",
        11924=>"000000010",
        11925=>"000100000",
        11926=>"101000000",
        11927=>"010011111",
        11928=>"001101000",
        11929=>"100001011",
        11930=>"001100101",
        11931=>"011100100",
        11932=>"000100111",
        11933=>"100101100",
        11934=>"101001100",
        11935=>"110111111",
        11936=>"000000111",
        11937=>"010000001",
        11938=>"001100001",
        11939=>"000010000",
        11940=>"111010010",
        11941=>"000101110",
        11942=>"000000111",
        11943=>"110110000",
        11944=>"010011101",
        11945=>"111111011",
        11946=>"100001000",
        11947=>"001101000",
        11948=>"100110111",
        11949=>"110110000",
        11950=>"000111111",
        11951=>"011001100",
        11952=>"111111000",
        11953=>"110000111",
        11954=>"001001001",
        11955=>"011010000",
        11956=>"010000000",
        11957=>"000000000",
        11958=>"010000111",
        11959=>"000000111",
        11960=>"110001000",
        11961=>"000001111",
        11962=>"011000101",
        11963=>"100000000",
        11964=>"000000111",
        11965=>"000000000",
        11966=>"111011011",
        11967=>"111101000",
        11968=>"101101110",
        11969=>"111010000",
        11970=>"110001111",
        11971=>"000000100",
        11972=>"011111101",
        11973=>"000101001",
        11974=>"111111000",
        11975=>"000000001",
        11976=>"000000011",
        11977=>"001111110",
        11978=>"100110010",
        11979=>"000000000",
        11980=>"000110010",
        11981=>"010110000",
        11982=>"000010110",
        11983=>"110000000",
        11984=>"110010000",
        11985=>"111000000",
        11986=>"100110000",
        11987=>"100000101",
        11988=>"000110000",
        11989=>"101010010",
        11990=>"110000000",
        11991=>"000001001",
        11992=>"111101100",
        11993=>"101001110",
        11994=>"000011110",
        11995=>"010000001",
        11996=>"011101000",
        11997=>"111110100",
        11998=>"000001011",
        11999=>"101001011",
        12000=>"000011111",
        12001=>"111110000",
        12002=>"111111010",
        12003=>"000001111",
        12004=>"110110100",
        12005=>"110101001",
        12006=>"111000000",
        12007=>"110111000",
        12008=>"100000000",
        12009=>"101001111",
        12010=>"100001000",
        12011=>"111111000",
        12012=>"111101010",
        12013=>"110000000",
        12014=>"111111111",
        12015=>"011000000",
        12016=>"010000000",
        12017=>"000111111",
        12018=>"000100111",
        12019=>"111000001",
        12020=>"000001000",
        12021=>"111000000",
        12022=>"000000000",
        12023=>"100110110",
        12024=>"111110000",
        12025=>"111000000",
        12026=>"001000000",
        12027=>"000000111",
        12028=>"000111011",
        12029=>"100000111",
        12030=>"010110001",
        12031=>"011111111",
        12032=>"100101001",
        12033=>"100000001",
        12034=>"101100111",
        12035=>"111101010",
        12036=>"101111100",
        12037=>"110111011",
        12038=>"111111110",
        12039=>"111000110",
        12040=>"010000000",
        12041=>"010110001",
        12042=>"100000000",
        12043=>"100001000",
        12044=>"101001111",
        12045=>"111111110",
        12046=>"100111011",
        12047=>"000000010",
        12048=>"101101101",
        12049=>"111100001",
        12050=>"001101110",
        12051=>"100110001",
        12052=>"111001111",
        12053=>"101100101",
        12054=>"111000110",
        12055=>"111000110",
        12056=>"111101111",
        12057=>"001100000",
        12058=>"101001001",
        12059=>"000000011",
        12060=>"000010000",
        12061=>"111101001",
        12062=>"101100000",
        12063=>"011101000",
        12064=>"111000000",
        12065=>"000001000",
        12066=>"010001001",
        12067=>"111101111",
        12068=>"111111110",
        12069=>"000000000",
        12070=>"011011000",
        12071=>"101101101",
        12072=>"111110010",
        12073=>"110111111",
        12074=>"001100110",
        12075=>"101111111",
        12076=>"111001101",
        12077=>"111100101",
        12078=>"000000000",
        12079=>"010001000",
        12080=>"001000100",
        12081=>"000101100",
        12082=>"100001001",
        12083=>"000000001",
        12084=>"001101001",
        12085=>"000000000",
        12086=>"110010111",
        12087=>"000000011",
        12088=>"101010010",
        12089=>"001000001",
        12090=>"010000001",
        12091=>"110000000",
        12092=>"010101101",
        12093=>"000010000",
        12094=>"000101110",
        12095=>"101011101",
        12096=>"000011111",
        12097=>"001100001",
        12098=>"010000010",
        12099=>"000110110",
        12100=>"111110001",
        12101=>"010110110",
        12102=>"111010110",
        12103=>"011000001",
        12104=>"110001001",
        12105=>"101001001",
        12106=>"001001111",
        12107=>"111000000",
        12108=>"000101101",
        12109=>"101111111",
        12110=>"000100100",
        12111=>"000100010",
        12112=>"000000101",
        12113=>"100100001",
        12114=>"100101100",
        12115=>"101111111",
        12116=>"010011011",
        12117=>"000000000",
        12118=>"001000010",
        12119=>"000110000",
        12120=>"011111111",
        12121=>"110000111",
        12122=>"001000000",
        12123=>"101100011",
        12124=>"111111111",
        12125=>"000001100",
        12126=>"001001101",
        12127=>"111000101",
        12128=>"100001100",
        12129=>"101000111",
        12130=>"111111111",
        12131=>"001010010",
        12132=>"000110110",
        12133=>"010100000",
        12134=>"000001100",
        12135=>"110110100",
        12136=>"111001000",
        12137=>"000000001",
        12138=>"100101111",
        12139=>"000010100",
        12140=>"000000000",
        12141=>"000000100",
        12142=>"000111110",
        12143=>"001000000",
        12144=>"101000100",
        12145=>"111011110",
        12146=>"111111101",
        12147=>"000110000",
        12148=>"111001111",
        12149=>"100101111",
        12150=>"000000011",
        12151=>"001001011",
        12152=>"111001111",
        12153=>"111010111",
        12154=>"100100111",
        12155=>"010001111",
        12156=>"000000000",
        12157=>"100000011",
        12158=>"011000000",
        12159=>"101100100",
        12160=>"000000000",
        12161=>"111000010",
        12162=>"000111111",
        12163=>"000011111",
        12164=>"110001000",
        12165=>"100000000",
        12166=>"010010111",
        12167=>"111000000",
        12168=>"000001111",
        12169=>"011111011",
        12170=>"111101000",
        12171=>"101111101",
        12172=>"000000100",
        12173=>"010111010",
        12174=>"000100100",
        12175=>"101100011",
        12176=>"000111110",
        12177=>"111100000",
        12178=>"111000100",
        12179=>"011110100",
        12180=>"000000111",
        12181=>"000000100",
        12182=>"011011111",
        12183=>"111110000",
        12184=>"010001001",
        12185=>"011111100",
        12186=>"100000000",
        12187=>"101111000",
        12188=>"010000000",
        12189=>"000001001",
        12190=>"110100110",
        12191=>"111001000",
        12192=>"000111010",
        12193=>"111110000",
        12194=>"111101100",
        12195=>"110101000",
        12196=>"000011111",
        12197=>"000010100",
        12198=>"111000000",
        12199=>"000000111",
        12200=>"111111000",
        12201=>"111111000",
        12202=>"001110101",
        12203=>"011110101",
        12204=>"000000100",
        12205=>"000000001",
        12206=>"111111000",
        12207=>"111000110",
        12208=>"011111000",
        12209=>"111010011",
        12210=>"111011101",
        12211=>"000000100",
        12212=>"110100101",
        12213=>"000110111",
        12214=>"011111011",
        12215=>"000010111",
        12216=>"000110111",
        12217=>"111111101",
        12218=>"100111111",
        12219=>"110000000",
        12220=>"111000000",
        12221=>"111100000",
        12222=>"111111000",
        12223=>"111111011",
        12224=>"010000000",
        12225=>"101101100",
        12226=>"000000000",
        12227=>"101111101",
        12228=>"010101111",
        12229=>"000000000",
        12230=>"000111111",
        12231=>"111000000",
        12232=>"000111011",
        12233=>"010011111",
        12234=>"111011000",
        12235=>"100000000",
        12236=>"111111001",
        12237=>"110000000",
        12238=>"111100000",
        12239=>"000011111",
        12240=>"000011011",
        12241=>"000000110",
        12242=>"011100100",
        12243=>"111000000",
        12244=>"000000000",
        12245=>"000110111",
        12246=>"111100011",
        12247=>"000000101",
        12248=>"110001000",
        12249=>"000101111",
        12250=>"111000000",
        12251=>"000111010",
        12252=>"011001111",
        12253=>"100001011",
        12254=>"100000011",
        12255=>"111000101",
        12256=>"000001110",
        12257=>"001011001",
        12258=>"100111111",
        12259=>"000111111",
        12260=>"101011111",
        12261=>"000000100",
        12262=>"100100011",
        12263=>"010111000",
        12264=>"000000011",
        12265=>"111100100",
        12266=>"011110100",
        12267=>"111101111",
        12268=>"011000000",
        12269=>"111000000",
        12270=>"010111111",
        12271=>"001000101",
        12272=>"010000111",
        12273=>"100001000",
        12274=>"000101111",
        12275=>"111011111",
        12276=>"010111111",
        12277=>"100000111",
        12278=>"000000000",
        12279=>"011110001",
        12280=>"000100011",
        12281=>"100111011",
        12282=>"000000110",
        12283=>"111000000",
        12284=>"010000110",
        12285=>"001010010",
        12286=>"011101100",
        12287=>"011100101",
        12288=>"000000000",
        12289=>"111101111",
        12290=>"111111110",
        12291=>"010001000",
        12292=>"000010000",
        12293=>"010011110",
        12294=>"111111111",
        12295=>"000000100",
        12296=>"110010011",
        12297=>"011010011",
        12298=>"101000111",
        12299=>"010010100",
        12300=>"111111011",
        12301=>"110110010",
        12302=>"110111110",
        12303=>"000001001",
        12304=>"110111111",
        12305=>"111100001",
        12306=>"001000000",
        12307=>"100000000",
        12308=>"111111000",
        12309=>"000010000",
        12310=>"110010110",
        12311=>"111111111",
        12312=>"011011000",
        12313=>"011110001",
        12314=>"010111011",
        12315=>"010111011",
        12316=>"000000000",
        12317=>"010111110",
        12318=>"111111000",
        12319=>"000000000",
        12320=>"000000011",
        12321=>"000011110",
        12322=>"010010000",
        12323=>"000000000",
        12324=>"000000101",
        12325=>"110011111",
        12326=>"111111111",
        12327=>"011000000",
        12328=>"000000000",
        12329=>"000000000",
        12330=>"010000000",
        12331=>"111111001",
        12332=>"001000111",
        12333=>"000000000",
        12334=>"000000000",
        12335=>"000000111",
        12336=>"101011111",
        12337=>"111111010",
        12338=>"000110010",
        12339=>"111111111",
        12340=>"110111111",
        12341=>"000000000",
        12342=>"111000111",
        12343=>"000001000",
        12344=>"000000001",
        12345=>"001111111",
        12346=>"110100110",
        12347=>"000000000",
        12348=>"111101111",
        12349=>"001100100",
        12350=>"010110110",
        12351=>"000000010",
        12352=>"111000101",
        12353=>"111111111",
        12354=>"000000000",
        12355=>"000000000",
        12356=>"000000001",
        12357=>"111101000",
        12358=>"011111110",
        12359=>"111101001",
        12360=>"111111111",
        12361=>"101111011",
        12362=>"001001111",
        12363=>"000000000",
        12364=>"001000000",
        12365=>"111011011",
        12366=>"000000011",
        12367=>"010111110",
        12368=>"111111011",
        12369=>"101000011",
        12370=>"111010011",
        12371=>"111111111",
        12372=>"100100101",
        12373=>"001001111",
        12374=>"010101111",
        12375=>"000010010",
        12376=>"000000000",
        12377=>"010010000",
        12378=>"001000000",
        12379=>"101111110",
        12380=>"111111111",
        12381=>"011000110",
        12382=>"000000000",
        12383=>"111111111",
        12384=>"111101110",
        12385=>"111101111",
        12386=>"000001001",
        12387=>"000001111",
        12388=>"111101111",
        12389=>"100000000",
        12390=>"101100100",
        12391=>"001000000",
        12392=>"111111011",
        12393=>"000111000",
        12394=>"101101010",
        12395=>"111111111",
        12396=>"111111011",
        12397=>"000111111",
        12398=>"101100001",
        12399=>"110111111",
        12400=>"000000000",
        12401=>"111111011",
        12402=>"001001000",
        12403=>"110111010",
        12404=>"111111111",
        12405=>"111010010",
        12406=>"011010000",
        12407=>"110111011",
        12408=>"001000011",
        12409=>"000000001",
        12410=>"011111110",
        12411=>"010000111",
        12412=>"000000000",
        12413=>"111110111",
        12414=>"001000000",
        12415=>"001010010",
        12416=>"000001000",
        12417=>"000000101",
        12418=>"111111000",
        12419=>"100101001",
        12420=>"111011110",
        12421=>"111111111",
        12422=>"000100001",
        12423=>"000000000",
        12424=>"001000000",
        12425=>"000000001",
        12426=>"000000100",
        12427=>"000100111",
        12428=>"000000010",
        12429=>"111111000",
        12430=>"001001011",
        12431=>"010000001",
        12432=>"000000110",
        12433=>"101000101",
        12434=>"111101111",
        12435=>"110111001",
        12436=>"000010000",
        12437=>"000100001",
        12438=>"000000111",
        12439=>"011000111",
        12440=>"111111111",
        12441=>"001001111",
        12442=>"001011101",
        12443=>"000000000",
        12444=>"110011111",
        12445=>"001101001",
        12446=>"011111111",
        12447=>"000000000",
        12448=>"001001000",
        12449=>"000001000",
        12450=>"111101110",
        12451=>"111111101",
        12452=>"000000011",
        12453=>"010111110",
        12454=>"001001011",
        12455=>"101110000",
        12456=>"101111111",
        12457=>"001000111",
        12458=>"111001001",
        12459=>"001001001",
        12460=>"000100111",
        12461=>"000000000",
        12462=>"000000000",
        12463=>"101101000",
        12464=>"000000000",
        12465=>"101110100",
        12466=>"000011000",
        12467=>"000010000",
        12468=>"000000110",
        12469=>"000000000",
        12470=>"000000000",
        12471=>"001001000",
        12472=>"000001111",
        12473=>"000101110",
        12474=>"000000111",
        12475=>"001000101",
        12476=>"000100111",
        12477=>"000001000",
        12478=>"000000000",
        12479=>"111011001",
        12480=>"011111010",
        12481=>"110111111",
        12482=>"111111111",
        12483=>"101101111",
        12484=>"000000111",
        12485=>"001001011",
        12486=>"000000000",
        12487=>"100101101",
        12488=>"000000001",
        12489=>"000111010",
        12490=>"001001110",
        12491=>"000000101",
        12492=>"000000000",
        12493=>"001000000",
        12494=>"000000010",
        12495=>"110110001",
        12496=>"000001011",
        12497=>"000001001",
        12498=>"001011000",
        12499=>"011111111",
        12500=>"111001111",
        12501=>"010010000",
        12502=>"000000000",
        12503=>"000000000",
        12504=>"001101100",
        12505=>"000000101",
        12506=>"000000000",
        12507=>"111111010",
        12508=>"001001111",
        12509=>"110000100",
        12510=>"111111111",
        12511=>"001110010",
        12512=>"000000001",
        12513=>"000000000",
        12514=>"010010000",
        12515=>"110110000",
        12516=>"001101111",
        12517=>"000000001",
        12518=>"000000000",
        12519=>"000000011",
        12520=>"101001101",
        12521=>"000000000",
        12522=>"101101001",
        12523=>"110001101",
        12524=>"010010000",
        12525=>"000000100",
        12526=>"110111110",
        12527=>"001001000",
        12528=>"111111010",
        12529=>"110111111",
        12530=>"001001001",
        12531=>"111111101",
        12532=>"111111010",
        12533=>"000000111",
        12534=>"101000111",
        12535=>"000100101",
        12536=>"000000110",
        12537=>"110111111",
        12538=>"001000111",
        12539=>"000000001",
        12540=>"101011001",
        12541=>"000000111",
        12542=>"111111111",
        12543=>"111111110",
        12544=>"000001000",
        12545=>"111000000",
        12546=>"001000000",
        12547=>"000111001",
        12548=>"011001100",
        12549=>"010111111",
        12550=>"000000000",
        12551=>"101000101",
        12552=>"000000000",
        12553=>"001110011",
        12554=>"101000000",
        12555=>"100101111",
        12556=>"001000000",
        12557=>"111111010",
        12558=>"001001001",
        12559=>"101110100",
        12560=>"100101011",
        12561=>"100100011",
        12562=>"101011010",
        12563=>"100000100",
        12564=>"101000010",
        12565=>"000000000",
        12566=>"101000100",
        12567=>"001000101",
        12568=>"000100000",
        12569=>"101110010",
        12570=>"100000000",
        12571=>"111000111",
        12572=>"111011111",
        12573=>"011001101",
        12574=>"000000000",
        12575=>"101100001",
        12576=>"000010111",
        12577=>"000000000",
        12578=>"111111000",
        12579=>"100000010",
        12580=>"100000111",
        12581=>"010110010",
        12582=>"000000111",
        12583=>"000010101",
        12584=>"111111000",
        12585=>"001011011",
        12586=>"101110100",
        12587=>"000000000",
        12588=>"000001001",
        12589=>"111100000",
        12590=>"000100110",
        12591=>"101100111",
        12592=>"000011011",
        12593=>"101000101",
        12594=>"100110000",
        12595=>"000000110",
        12596=>"100100111",
        12597=>"101100000",
        12598=>"000000000",
        12599=>"110000000",
        12600=>"000101111",
        12601=>"000000000",
        12602=>"100111111",
        12603=>"000000110",
        12604=>"000000100",
        12605=>"010101011",
        12606=>"110001111",
        12607=>"111011011",
        12608=>"101100000",
        12609=>"000000100",
        12610=>"100011111",
        12611=>"011111111",
        12612=>"000000001",
        12613=>"011011101",
        12614=>"111111001",
        12615=>"011000000",
        12616=>"001000100",
        12617=>"010011110",
        12618=>"001000000",
        12619=>"101000111",
        12620=>"100000100",
        12621=>"010000000",
        12622=>"000101101",
        12623=>"001100111",
        12624=>"100101000",
        12625=>"000000000",
        12626=>"011111000",
        12627=>"101100100",
        12628=>"010100100",
        12629=>"000010000",
        12630=>"001000101",
        12631=>"000001111",
        12632=>"001100110",
        12633=>"101100100",
        12634=>"000001111",
        12635=>"000000000",
        12636=>"000001001",
        12637=>"101000001",
        12638=>"100101001",
        12639=>"111111001",
        12640=>"000001011",
        12641=>"000110110",
        12642=>"111111111",
        12643=>"100000001",
        12644=>"001000001",
        12645=>"000000111",
        12646=>"000000000",
        12647=>"000000110",
        12648=>"000000011",
        12649=>"101100100",
        12650=>"110100001",
        12651=>"101001000",
        12652=>"011001101",
        12653=>"111000101",
        12654=>"110010110",
        12655=>"000101100",
        12656=>"000000000",
        12657=>"011111111",
        12658=>"100000000",
        12659=>"000111110",
        12660=>"111111101",
        12661=>"000000001",
        12662=>"000000101",
        12663=>"001011101",
        12664=>"111100110",
        12665=>"100000100",
        12666=>"000000110",
        12667=>"111000001",
        12668=>"000000111",
        12669=>"101101111",
        12670=>"111111010",
        12671=>"110111011",
        12672=>"110110110",
        12673=>"001011001",
        12674=>"000111111",
        12675=>"100100111",
        12676=>"000100100",
        12677=>"110011101",
        12678=>"000100110",
        12679=>"010011011",
        12680=>"101000001",
        12681=>"001010011",
        12682=>"111000111",
        12683=>"011000111",
        12684=>"011001000",
        12685=>"011101001",
        12686=>"100000000",
        12687=>"011011001",
        12688=>"111010010",
        12689=>"000011011",
        12690=>"000100000",
        12691=>"111110110",
        12692=>"000011000",
        12693=>"000100000",
        12694=>"011011100",
        12695=>"111111001",
        12696=>"000100110",
        12697=>"101000100",
        12698=>"110100100",
        12699=>"111100100",
        12700=>"000000000",
        12701=>"100110110",
        12702=>"110110111",
        12703=>"010111110",
        12704=>"110110111",
        12705=>"000000000",
        12706=>"101100010",
        12707=>"000000000",
        12708=>"100100110",
        12709=>"010011111",
        12710=>"111011011",
        12711=>"100100100",
        12712=>"010001111",
        12713=>"010100000",
        12714=>"110100000",
        12715=>"100100100",
        12716=>"100100110",
        12717=>"000110100",
        12718=>"010001100",
        12719=>"101110111",
        12720=>"110001001",
        12721=>"001011001",
        12722=>"111110111",
        12723=>"111100000",
        12724=>"011111011",
        12725=>"001001000",
        12726=>"000001001",
        12727=>"111001000",
        12728=>"110100110",
        12729=>"100110110",
        12730=>"100100111",
        12731=>"010010100",
        12732=>"001010000",
        12733=>"010000000",
        12734=>"100100110",
        12735=>"100100101",
        12736=>"000110000",
        12737=>"011101111",
        12738=>"100011011",
        12739=>"011001001",
        12740=>"110100110",
        12741=>"110110110",
        12742=>"111000000",
        12743=>"001100110",
        12744=>"000000000",
        12745=>"111001001",
        12746=>"100110011",
        12747=>"000100000",
        12748=>"001010100",
        12749=>"011001011",
        12750=>"001000000",
        12751=>"111011001",
        12752=>"011011001",
        12753=>"110010000",
        12754=>"001001001",
        12755=>"111010000",
        12756=>"110110000",
        12757=>"011011000",
        12758=>"110000000",
        12759=>"110110111",
        12760=>"100100000",
        12761=>"000100100",
        12762=>"001000000",
        12763=>"100000001",
        12764=>"100100100",
        12765=>"001000010",
        12766=>"110110000",
        12767=>"001001000",
        12768=>"000001000",
        12769=>"100110111",
        12770=>"000100101",
        12771=>"100100110",
        12772=>"110110010",
        12773=>"110100100",
        12774=>"100100110",
        12775=>"100100100",
        12776=>"001001000",
        12777=>"011000000",
        12778=>"100100100",
        12779=>"011010010",
        12780=>"110100100",
        12781=>"001011001",
        12782=>"111111110",
        12783=>"111100110",
        12784=>"011000001",
        12785=>"001101111",
        12786=>"000000000",
        12787=>"011011001",
        12788=>"001000101",
        12789=>"011000001",
        12790=>"001011011",
        12791=>"010000000",
        12792=>"000000101",
        12793=>"011011010",
        12794=>"010011011",
        12795=>"000001011",
        12796=>"110100111",
        12797=>"111011011",
        12798=>"000110111",
        12799=>"110101011",
        12800=>"001001000",
        12801=>"010111010",
        12802=>"100000100",
        12803=>"001000000",
        12804=>"011011101",
        12805=>"111111111",
        12806=>"000000110",
        12807=>"000110100",
        12808=>"001001010",
        12809=>"100101100",
        12810=>"000000100",
        12811=>"111111111",
        12812=>"111111111",
        12813=>"010010010",
        12814=>"101111011",
        12815=>"010001011",
        12816=>"001100100",
        12817=>"111111111",
        12818=>"000000000",
        12819=>"110110101",
        12820=>"010000000",
        12821=>"111110101",
        12822=>"111111111",
        12823=>"010101111",
        12824=>"000000000",
        12825=>"011011001",
        12826=>"111011111",
        12827=>"000000011",
        12828=>"000000000",
        12829=>"111101111",
        12830=>"001000000",
        12831=>"000000000",
        12832=>"011111111",
        12833=>"000000000",
        12834=>"111011110",
        12835=>"000000000",
        12836=>"001000111",
        12837=>"111000101",
        12838=>"111111111",
        12839=>"000000000",
        12840=>"000000000",
        12841=>"000000000",
        12842=>"011101000",
        12843=>"000000000",
        12844=>"100100110",
        12845=>"000000000",
        12846=>"000101000",
        12847=>"000000000",
        12848=>"010001010",
        12849=>"111111000",
        12850=>"111111110",
        12851=>"100001001",
        12852=>"110100111",
        12853=>"111111111",
        12854=>"010111111",
        12855=>"000111111",
        12856=>"111011000",
        12857=>"000000111",
        12858=>"010101110",
        12859=>"111111111",
        12860=>"011111010",
        12861=>"000000000",
        12862=>"000000100",
        12863=>"110000110",
        12864=>"111101011",
        12865=>"000111000",
        12866=>"000111111",
        12867=>"110111111",
        12868=>"000000000",
        12869=>"000000010",
        12870=>"000111001",
        12871=>"101100101",
        12872=>"100100100",
        12873=>"111111110",
        12874=>"000000100",
        12875=>"111101111",
        12876=>"000000000",
        12877=>"000000000",
        12878=>"000000000",
        12879=>"010011011",
        12880=>"011111111",
        12881=>"111000111",
        12882=>"110110010",
        12883=>"110100100",
        12884=>"000000110",
        12885=>"111111000",
        12886=>"000000000",
        12887=>"000000000",
        12888=>"000000000",
        12889=>"110010110",
        12890=>"001111111",
        12891=>"010111110",
        12892=>"000000000",
        12893=>"001000100",
        12894=>"111111100",
        12895=>"111111001",
        12896=>"100100100",
        12897=>"101100000",
        12898=>"111111111",
        12899=>"001011011",
        12900=>"100011111",
        12901=>"011111111",
        12902=>"101101100",
        12903=>"101101111",
        12904=>"111111111",
        12905=>"100000111",
        12906=>"010000001",
        12907=>"000000110",
        12908=>"000000000",
        12909=>"000110110",
        12910=>"110110011",
        12911=>"100000000",
        12912=>"000000111",
        12913=>"011001110",
        12914=>"111000000",
        12915=>"111111111",
        12916=>"111111111",
        12917=>"000000001",
        12918=>"011011111",
        12919=>"111110011",
        12920=>"000111110",
        12921=>"111111011",
        12922=>"111111111",
        12923=>"000000000",
        12924=>"110111001",
        12925=>"100111111",
        12926=>"110000000",
        12927=>"011110100",
        12928=>"111111011",
        12929=>"111000000",
        12930=>"000000000",
        12931=>"000100000",
        12932=>"100101100",
        12933=>"110101111",
        12934=>"011111101",
        12935=>"001000101",
        12936=>"011111111",
        12937=>"110100110",
        12938=>"111111010",
        12939=>"111011000",
        12940=>"001000001",
        12941=>"010111010",
        12942=>"000000111",
        12943=>"101000000",
        12944=>"111111000",
        12945=>"010011011",
        12946=>"011011011",
        12947=>"001001001",
        12948=>"010111010",
        12949=>"000000000",
        12950=>"000000100",
        12951=>"101101111",
        12952=>"110100100",
        12953=>"111100000",
        12954=>"100100100",
        12955=>"001001110",
        12956=>"110111111",
        12957=>"100100100",
        12958=>"000001111",
        12959=>"011000111",
        12960=>"101101101",
        12961=>"011001001",
        12962=>"010001000",
        12963=>"000000111",
        12964=>"101111000",
        12965=>"010010010",
        12966=>"100000000",
        12967=>"000010110",
        12968=>"111011000",
        12969=>"001010011",
        12970=>"100101000",
        12971=>"001011000",
        12972=>"101111111",
        12973=>"000000000",
        12974=>"110010010",
        12975=>"101111011",
        12976=>"111111101",
        12977=>"111001101",
        12978=>"011111110",
        12979=>"000011011",
        12980=>"101011011",
        12981=>"000000000",
        12982=>"111100101",
        12983=>"100101111",
        12984=>"011101000",
        12985=>"000010001",
        12986=>"011011111",
        12987=>"001101000",
        12988=>"000000000",
        12989=>"010010111",
        12990=>"101001000",
        12991=>"000000100",
        12992=>"111111100",
        12993=>"111101000",
        12994=>"111000000",
        12995=>"100111010",
        12996=>"110111011",
        12997=>"001011001",
        12998=>"000000111",
        12999=>"111000000",
        13000=>"110111101",
        13001=>"111000000",
        13002=>"000100110",
        13003=>"000000000",
        13004=>"000000000",
        13005=>"010010001",
        13006=>"000010010",
        13007=>"101000101",
        13008=>"101000000",
        13009=>"000000000",
        13010=>"000000000",
        13011=>"000000000",
        13012=>"110110000",
        13013=>"000000000",
        13014=>"001000000",
        13015=>"111111111",
        13016=>"110100111",
        13017=>"000000000",
        13018=>"011011011",
        13019=>"000010000",
        13020=>"010100100",
        13021=>"101000001",
        13022=>"001001001",
        13023=>"100100000",
        13024=>"101111110",
        13025=>"101111110",
        13026=>"111111010",
        13027=>"000000000",
        13028=>"011000000",
        13029=>"011010000",
        13030=>"000000011",
        13031=>"101001110",
        13032=>"010000001",
        13033=>"111100100",
        13034=>"110001111",
        13035=>"000100000",
        13036=>"011111010",
        13037=>"010000000",
        13038=>"000100000",
        13039=>"111011011",
        13040=>"111101000",
        13041=>"000000010",
        13042=>"010111100",
        13043=>"000000000",
        13044=>"001000101",
        13045=>"000000001",
        13046=>"000000000",
        13047=>"111101111",
        13048=>"011001000",
        13049=>"000000010",
        13050=>"000100100",
        13051=>"000000000",
        13052=>"110110110",
        13053=>"111111111",
        13054=>"000000000",
        13055=>"110100011",
        13056=>"111111111",
        13057=>"001000000",
        13058=>"000000111",
        13059=>"111100001",
        13060=>"000110000",
        13061=>"111000101",
        13062=>"000000000",
        13063=>"000111111",
        13064=>"000100111",
        13065=>"111100010",
        13066=>"111111010",
        13067=>"001011100",
        13068=>"000000111",
        13069=>"010111010",
        13070=>"100110110",
        13071=>"110111011",
        13072=>"011100100",
        13073=>"111111111",
        13074=>"000011001",
        13075=>"000011011",
        13076=>"110000000",
        13077=>"110111010",
        13078=>"111000101",
        13079=>"111111110",
        13080=>"110110100",
        13081=>"100000000",
        13082=>"100101001",
        13083=>"001101001",
        13084=>"111111100",
        13085=>"111111100",
        13086=>"001001000",
        13087=>"111111111",
        13088=>"100101111",
        13089=>"001011000",
        13090=>"001100110",
        13091=>"000000000",
        13092=>"000010000",
        13093=>"111000001",
        13094=>"010111111",
        13095=>"100001000",
        13096=>"011000000",
        13097=>"010010011",
        13098=>"100001001",
        13099=>"000111001",
        13100=>"010111000",
        13101=>"111111000",
        13102=>"000001010",
        13103=>"001010010",
        13104=>"101101011",
        13105=>"000000000",
        13106=>"110100110",
        13107=>"011001001",
        13108=>"111111011",
        13109=>"111000000",
        13110=>"100000000",
        13111=>"001000101",
        13112=>"000011011",
        13113=>"000000010",
        13114=>"001001001",
        13115=>"010110011",
        13116=>"000000000",
        13117=>"000000110",
        13118=>"100101000",
        13119=>"011000111",
        13120=>"111000000",
        13121=>"000000000",
        13122=>"111010010",
        13123=>"101011000",
        13124=>"101000000",
        13125=>"110110100",
        13126=>"110100110",
        13127=>"000000000",
        13128=>"110100000",
        13129=>"000000000",
        13130=>"010011001",
        13131=>"000111111",
        13132=>"000000111",
        13133=>"000000000",
        13134=>"000001000",
        13135=>"000111011",
        13136=>"000000010",
        13137=>"110010000",
        13138=>"010111010",
        13139=>"111000000",
        13140=>"011011011",
        13141=>"000000101",
        13142=>"000001011",
        13143=>"011001001",
        13144=>"110110100",
        13145=>"110001011",
        13146=>"000001010",
        13147=>"110000000",
        13148=>"000001000",
        13149=>"000111110",
        13150=>"001011011",
        13151=>"000000000",
        13152=>"111100100",
        13153=>"111100100",
        13154=>"111100100",
        13155=>"000000000",
        13156=>"010110110",
        13157=>"011111010",
        13158=>"001011000",
        13159=>"101111111",
        13160=>"010001011",
        13161=>"100000000",
        13162=>"111110011",
        13163=>"000000000",
        13164=>"101000101",
        13165=>"111010110",
        13166=>"111111111",
        13167=>"000001001",
        13168=>"010111010",
        13169=>"100100011",
        13170=>"101001000",
        13171=>"001000101",
        13172=>"101001111",
        13173=>"000010011",
        13174=>"000000000",
        13175=>"010001011",
        13176=>"110010110",
        13177=>"101111111",
        13178=>"100010010",
        13179=>"111111111",
        13180=>"100110110",
        13181=>"111000100",
        13182=>"100010010",
        13183=>"001001111",
        13184=>"010111111",
        13185=>"110010010",
        13186=>"100000100",
        13187=>"111111111",
        13188=>"001001100",
        13189=>"011110000",
        13190=>"110010001",
        13191=>"000100111",
        13192=>"111101101",
        13193=>"100000000",
        13194=>"111010101",
        13195=>"100100100",
        13196=>"001000000",
        13197=>"111010100",
        13198=>"111001100",
        13199=>"100100110",
        13200=>"011011001",
        13201=>"000111101",
        13202=>"001001001",
        13203=>"000100000",
        13204=>"010011001",
        13205=>"000000010",
        13206=>"000000010",
        13207=>"010110110",
        13208=>"001001001",
        13209=>"011011000",
        13210=>"011001001",
        13211=>"111110000",
        13212=>"111111000",
        13213=>"011000001",
        13214=>"000101101",
        13215=>"000100010",
        13216=>"011001000",
        13217=>"001000000",
        13218=>"011001001",
        13219=>"000001000",
        13220=>"111011000",
        13221=>"110001100",
        13222=>"111011000",
        13223=>"111011001",
        13224=>"110110110",
        13225=>"101000100",
        13226=>"000010000",
        13227=>"001001001",
        13228=>"001001111",
        13229=>"000110110",
        13230=>"001000000",
        13231=>"111111111",
        13232=>"011001001",
        13233=>"100110101",
        13234=>"100100100",
        13235=>"000100000",
        13236=>"011001101",
        13237=>"011000000",
        13238=>"111011000",
        13239=>"100111111",
        13240=>"110110110",
        13241=>"111011100",
        13242=>"000000000",
        13243=>"010110110",
        13244=>"110100110",
        13245=>"100110100",
        13246=>"000010000",
        13247=>"001111101",
        13248=>"101000000",
        13249=>"011000101",
        13250=>"010011000",
        13251=>"111111101",
        13252=>"011001000",
        13253=>"011100000",
        13254=>"100000110",
        13255=>"010110011",
        13256=>"100100100",
        13257=>"010101001",
        13258=>"111000000",
        13259=>"100110110",
        13260=>"000110100",
        13261=>"000000001",
        13262=>"100010100",
        13263=>"100010110",
        13264=>"011010000",
        13265=>"100110110",
        13266=>"000000001",
        13267=>"011001111",
        13268=>"001011001",
        13269=>"110110010",
        13270=>"000100111",
        13271=>"011110000",
        13272=>"000001001",
        13273=>"011111011",
        13274=>"000100100",
        13275=>"011000000",
        13276=>"001101001",
        13277=>"011011001",
        13278=>"001111111",
        13279=>"000010111",
        13280=>"101101000",
        13281=>"110111111",
        13282=>"111111111",
        13283=>"111111001",
        13284=>"010000000",
        13285=>"100110010",
        13286=>"111001000",
        13287=>"011011111",
        13288=>"011001001",
        13289=>"100100000",
        13290=>"101101001",
        13291=>"011110001",
        13292=>"111111111",
        13293=>"001000010",
        13294=>"110100100",
        13295=>"101101111",
        13296=>"101110110",
        13297=>"100110111",
        13298=>"100111000",
        13299=>"011001011",
        13300=>"111101100",
        13301=>"001100100",
        13302=>"111000010",
        13303=>"001011001",
        13304=>"011111001",
        13305=>"110110110",
        13306=>"100100110",
        13307=>"000110010",
        13308=>"000011101",
        13309=>"011111100",
        13310=>"010111110",
        13311=>"100100000",
        13312=>"101111110",
        13313=>"111100101",
        13314=>"111111000",
        13315=>"000000111",
        13316=>"111011000",
        13317=>"100110111",
        13318=>"010111010",
        13319=>"111011111",
        13320=>"100111011",
        13321=>"110110111",
        13322=>"111001000",
        13323=>"100101111",
        13324=>"000000111",
        13325=>"110111110",
        13326=>"000001011",
        13327=>"000000111",
        13328=>"010001111",
        13329=>"000000101",
        13330=>"100110011",
        13331=>"110000000",
        13332=>"110000100",
        13333=>"010000000",
        13334=>"111010111",
        13335=>"000111111",
        13336=>"011011110",
        13337=>"000111111",
        13338=>"011100100",
        13339=>"011110011",
        13340=>"000000010",
        13341=>"100011011",
        13342=>"110111001",
        13343=>"000111110",
        13344=>"000010111",
        13345=>"001100000",
        13346=>"000101000",
        13347=>"000000000",
        13348=>"111110010",
        13349=>"100000000",
        13350=>"000000111",
        13351=>"111100110",
        13352=>"000000111",
        13353=>"000000000",
        13354=>"000000001",
        13355=>"000111000",
        13356=>"000111111",
        13357=>"111111111",
        13358=>"000001011",
        13359=>"000000101",
        13360=>"101011101",
        13361=>"010111000",
        13362=>"000000111",
        13363=>"010111100",
        13364=>"010100000",
        13365=>"101111101",
        13366=>"010000110",
        13367=>"000010110",
        13368=>"000000000",
        13369=>"000000010",
        13370=>"011111111",
        13371=>"000000111",
        13372=>"111010000",
        13373=>"010011110",
        13374=>"000111011",
        13375=>"011111110",
        13376=>"101000000",
        13377=>"111011000",
        13378=>"000001111",
        13379=>"101001111",
        13380=>"101001011",
        13381=>"000100100",
        13382=>"111111100",
        13383=>"101110101",
        13384=>"110000011",
        13385=>"101111000",
        13386=>"111111111",
        13387=>"000000000",
        13388=>"110000000",
        13389=>"111111000",
        13390=>"011000000",
        13391=>"001110011",
        13392=>"000000000",
        13393=>"111000100",
        13394=>"000111111",
        13395=>"110000001",
        13396=>"000011010",
        13397=>"111001101",
        13398=>"000110010",
        13399=>"111111001",
        13400=>"001001000",
        13401=>"111101010",
        13402=>"000001010",
        13403=>"111000000",
        13404=>"111111000",
        13405=>"011000100",
        13406=>"101111100",
        13407=>"000111111",
        13408=>"110111100",
        13409=>"110111001",
        13410=>"001101111",
        13411=>"111100000",
        13412=>"000111111",
        13413=>"010111011",
        13414=>"010000011",
        13415=>"011000010",
        13416=>"011001111",
        13417=>"111000000",
        13418=>"111011000",
        13419=>"111111101",
        13420=>"111111110",
        13421=>"111000001",
        13422=>"000110110",
        13423=>"000100110",
        13424=>"111111000",
        13425=>"101001111",
        13426=>"110111100",
        13427=>"100000111",
        13428=>"111111101",
        13429=>"010010000",
        13430=>"101000100",
        13431=>"000101110",
        13432=>"010000000",
        13433=>"011100000",
        13434=>"000000010",
        13435=>"010000000",
        13436=>"100101111",
        13437=>"101111111",
        13438=>"001000000",
        13439=>"001111000",
        13440=>"000100111",
        13441=>"000111111",
        13442=>"111101111",
        13443=>"111101111",
        13444=>"100000000",
        13445=>"011111111",
        13446=>"010000010",
        13447=>"101001001",
        13448=>"111100101",
        13449=>"100111100",
        13450=>"111101000",
        13451=>"011011110",
        13452=>"000010000",
        13453=>"010111110",
        13454=>"000000000",
        13455=>"111000001",
        13456=>"100011001",
        13457=>"000000100",
        13458=>"100100100",
        13459=>"001011011",
        13460=>"011000010",
        13461=>"111110010",
        13462=>"000000000",
        13463=>"001000111",
        13464=>"001001000",
        13465=>"110100001",
        13466=>"110100111",
        13467=>"011111000",
        13468=>"000101111",
        13469=>"000000000",
        13470=>"001000000",
        13471=>"100000000",
        13472=>"101101111",
        13473=>"000000100",
        13474=>"000001010",
        13475=>"011000000",
        13476=>"000110010",
        13477=>"000101111",
        13478=>"100101111",
        13479=>"000000000",
        13480=>"101100000",
        13481=>"111100100",
        13482=>"110111110",
        13483=>"101101101",
        13484=>"111001001",
        13485=>"111111000",
        13486=>"111011000",
        13487=>"101000101",
        13488=>"000001111",
        13489=>"000000000",
        13490=>"100110011",
        13491=>"000000010",
        13492=>"000000000",
        13493=>"000010000",
        13494=>"110111000",
        13495=>"010010010",
        13496=>"111111111",
        13497=>"000000010",
        13498=>"011011010",
        13499=>"000110111",
        13500=>"000000000",
        13501=>"111101111",
        13502=>"010011000",
        13503=>"001001111",
        13504=>"111111010",
        13505=>"111001001",
        13506=>"111001000",
        13507=>"001000000",
        13508=>"111111111",
        13509=>"000000100",
        13510=>"111010100",
        13511=>"000001000",
        13512=>"000110100",
        13513=>"000100101",
        13514=>"101001000",
        13515=>"000000000",
        13516=>"100000000",
        13517=>"111000001",
        13518=>"001000000",
        13519=>"011000001",
        13520=>"111101000",
        13521=>"001010110",
        13522=>"101101000",
        13523=>"111100000",
        13524=>"001000001",
        13525=>"000010001",
        13526=>"111000000",
        13527=>"000111111",
        13528=>"111011011",
        13529=>"000110000",
        13530=>"001011111",
        13531=>"101000000",
        13532=>"101001001",
        13533=>"100010001",
        13534=>"011111111",
        13535=>"111110110",
        13536=>"111011000",
        13537=>"100100111",
        13538=>"000001101",
        13539=>"111000000",
        13540=>"111111000",
        13541=>"000000000",
        13542=>"100010011",
        13543=>"101101010",
        13544=>"000110011",
        13545=>"111000000",
        13546=>"001001100",
        13547=>"000000000",
        13548=>"110101111",
        13549=>"000100000",
        13550=>"000111010",
        13551=>"010000000",
        13552=>"101000001",
        13553=>"000000000",
        13554=>"010010010",
        13555=>"000100111",
        13556=>"010111000",
        13557=>"001111010",
        13558=>"111111011",
        13559=>"101101110",
        13560=>"111001101",
        13561=>"000000000",
        13562=>"010010110",
        13563=>"111101001",
        13564=>"110111110",
        13565=>"111001111",
        13566=>"111111111",
        13567=>"000000000",
        13568=>"110100111",
        13569=>"111111110",
        13570=>"011111110",
        13571=>"000100010",
        13572=>"011011101",
        13573=>"100111110",
        13574=>"100010010",
        13575=>"110001011",
        13576=>"111000000",
        13577=>"110111010",
        13578=>"100000100",
        13579=>"000000000",
        13580=>"000110000",
        13581=>"111111111",
        13582=>"000000001",
        13583=>"110001111",
        13584=>"101101000",
        13585=>"111011111",
        13586=>"011110100",
        13587=>"100000001",
        13588=>"000000000",
        13589=>"111110001",
        13590=>"111000111",
        13591=>"000001111",
        13592=>"100100000",
        13593=>"100010110",
        13594=>"111111111",
        13595=>"101111011",
        13596=>"001101100",
        13597=>"110111011",
        13598=>"011100001",
        13599=>"111001000",
        13600=>"001000000",
        13601=>"110000000",
        13602=>"111111101",
        13603=>"110001000",
        13604=>"000010011",
        13605=>"011100101",
        13606=>"111011111",
        13607=>"000100100",
        13608=>"101110010",
        13609=>"110001010",
        13610=>"011100100",
        13611=>"011001001",
        13612=>"111001100",
        13613=>"011010000",
        13614=>"100100001",
        13615=>"111110111",
        13616=>"100100010",
        13617=>"001000100",
        13618=>"000000000",
        13619=>"100001000",
        13620=>"101101100",
        13621=>"000000000",
        13622=>"010010010",
        13623=>"011111010",
        13624=>"111000010",
        13625=>"110001001",
        13626=>"011100110",
        13627=>"000000000",
        13628=>"101100100",
        13629=>"011100111",
        13630=>"010000000",
        13631=>"110010111",
        13632=>"110011010",
        13633=>"101011000",
        13634=>"110001000",
        13635=>"110010110",
        13636=>"111110110",
        13637=>"110110000",
        13638=>"100101111",
        13639=>"011010011",
        13640=>"000000010",
        13641=>"111111100",
        13642=>"100000010",
        13643=>"000000000",
        13644=>"100000011",
        13645=>"001001001",
        13646=>"011011111",
        13647=>"000110100",
        13648=>"010010000",
        13649=>"000000000",
        13650=>"100001110",
        13651=>"111101010",
        13652=>"110111111",
        13653=>"011011010",
        13654=>"000110010",
        13655=>"001001110",
        13656=>"111111110",
        13657=>"010010111",
        13658=>"000001000",
        13659=>"011011000",
        13660=>"001101110",
        13661=>"011111111",
        13662=>"000100101",
        13663=>"001000011",
        13664=>"101111111",
        13665=>"011111111",
        13666=>"000000010",
        13667=>"110100010",
        13668=>"001011111",
        13669=>"000010010",
        13670=>"101111100",
        13671=>"111000011",
        13672=>"111111111",
        13673=>"000000000",
        13674=>"100001101",
        13675=>"111001000",
        13676=>"000001000",
        13677=>"001000001",
        13678=>"011010000",
        13679=>"110011111",
        13680=>"000000001",
        13681=>"011011001",
        13682=>"000100100",
        13683=>"000011010",
        13684=>"111101111",
        13685=>"010001001",
        13686=>"100111011",
        13687=>"111111111",
        13688=>"000110111",
        13689=>"111100010",
        13690=>"000000000",
        13691=>"110001011",
        13692=>"111111111",
        13693=>"111011111",
        13694=>"111100010",
        13695=>"000000000",
        13696=>"100010011",
        13697=>"111111000",
        13698=>"111111011",
        13699=>"011011010",
        13700=>"001000010",
        13701=>"111111000",
        13702=>"000000000",
        13703=>"000000111",
        13704=>"000000101",
        13705=>"010110100",
        13706=>"000000000",
        13707=>"000000100",
        13708=>"100100111",
        13709=>"111111111",
        13710=>"101001000",
        13711=>"110011011",
        13712=>"000000111",
        13713=>"111110010",
        13714=>"111101111",
        13715=>"110011000",
        13716=>"111011011",
        13717=>"010010000",
        13718=>"000000111",
        13719=>"101011010",
        13720=>"111111000",
        13721=>"110001011",
        13722=>"111111100",
        13723=>"000001111",
        13724=>"000010000",
        13725=>"100101101",
        13726=>"111111110",
        13727=>"010011110",
        13728=>"000000000",
        13729=>"100000000",
        13730=>"100100110",
        13731=>"001000111",
        13732=>"111011000",
        13733=>"000100101",
        13734=>"000000000",
        13735=>"111111000",
        13736=>"111101000",
        13737=>"000001111",
        13738=>"000000000",
        13739=>"100101000",
        13740=>"000110010",
        13741=>"000010111",
        13742=>"000000111",
        13743=>"000000001",
        13744=>"000001101",
        13745=>"111111010",
        13746=>"000100110",
        13747=>"111111011",
        13748=>"001001100",
        13749=>"000000101",
        13750=>"100101000",
        13751=>"101111010",
        13752=>"111111110",
        13753=>"000011001",
        13754=>"101101111",
        13755=>"111111110",
        13756=>"000000000",
        13757=>"101010000",
        13758=>"000110111",
        13759=>"101010110",
        13760=>"111101110",
        13761=>"000000000",
        13762=>"110000101",
        13763=>"000010000",
        13764=>"101000100",
        13765=>"000000000",
        13766=>"000100000",
        13767=>"000000000",
        13768=>"100100100",
        13769=>"100000000",
        13770=>"000100010",
        13771=>"111111011",
        13772=>"000000000",
        13773=>"101111111",
        13774=>"010101010",
        13775=>"100101111",
        13776=>"011111111",
        13777=>"100001001",
        13778=>"000000101",
        13779=>"111111111",
        13780=>"000000001",
        13781=>"000000000",
        13782=>"100000000",
        13783=>"101111111",
        13784=>"001100011",
        13785=>"000000000",
        13786=>"001001001",
        13787=>"111111100",
        13788=>"100100001",
        13789=>"011111110",
        13790=>"000000000",
        13791=>"001000101",
        13792=>"000100100",
        13793=>"111110111",
        13794=>"111111011",
        13795=>"010000000",
        13796=>"010111111",
        13797=>"111111000",
        13798=>"000100110",
        13799=>"010000000",
        13800=>"100100010",
        13801=>"111111000",
        13802=>"110011001",
        13803=>"111111101",
        13804=>"101111000",
        13805=>"111000101",
        13806=>"000000000",
        13807=>"001110000",
        13808=>"111111111",
        13809=>"000000110",
        13810=>"100100111",
        13811=>"000000000",
        13812=>"000010000",
        13813=>"000100111",
        13814=>"010000011",
        13815=>"000000011",
        13816=>"000000101",
        13817=>"000000010",
        13818=>"001011110",
        13819=>"000000101",
        13820=>"000000100",
        13821=>"000000000",
        13822=>"111111010",
        13823=>"100001000",
        13824=>"100000000",
        13825=>"000000000",
        13826=>"110110111",
        13827=>"001000000",
        13828=>"001001100",
        13829=>"001000000",
        13830=>"101110111",
        13831=>"001010001",
        13832=>"100100000",
        13833=>"011110110",
        13834=>"110101011",
        13835=>"011001011",
        13836=>"000011000",
        13837=>"010111110",
        13838=>"000000001",
        13839=>"100000011",
        13840=>"001111100",
        13841=>"111110101",
        13842=>"000000000",
        13843=>"111111000",
        13844=>"111110000",
        13845=>"101010010",
        13846=>"001000000",
        13847=>"010000111",
        13848=>"001001010",
        13849=>"100000010",
        13850=>"000000110",
        13851=>"011011111",
        13852=>"111111111",
        13853=>"100000000",
        13854=>"111111111",
        13855=>"000000110",
        13856=>"110000000",
        13857=>"111000110",
        13858=>"001100000",
        13859=>"111111111",
        13860=>"100101001",
        13861=>"111001111",
        13862=>"000010111",
        13863=>"101111001",
        13864=>"000000000",
        13865=>"000000000",
        13866=>"100100001",
        13867=>"001001001",
        13868=>"101111100",
        13869=>"101010111",
        13870=>"010101111",
        13871=>"000000000",
        13872=>"000011111",
        13873=>"000001111",
        13874=>"110111111",
        13875=>"101010101",
        13876=>"000000000",
        13877=>"000000000",
        13878=>"111111110",
        13879=>"000000100",
        13880=>"000000000",
        13881=>"111101111",
        13882=>"011101011",
        13883=>"000000000",
        13884=>"000000000",
        13885=>"111001111",
        13886=>"110110111",
        13887=>"111110111",
        13888=>"011011111",
        13889=>"111111111",
        13890=>"000000110",
        13891=>"101110111",
        13892=>"111111100",
        13893=>"110111111",
        13894=>"110111111",
        13895=>"101010111",
        13896=>"010001011",
        13897=>"111111111",
        13898=>"000000001",
        13899=>"101000000",
        13900=>"111111001",
        13901=>"011011100",
        13902=>"111110101",
        13903=>"110111111",
        13904=>"111111111",
        13905=>"100011001",
        13906=>"000100010",
        13907=>"000100111",
        13908=>"011111111",
        13909=>"000110100",
        13910=>"101110111",
        13911=>"111010110",
        13912=>"000000000",
        13913=>"101111111",
        13914=>"000000000",
        13915=>"111111111",
        13916=>"000000100",
        13917=>"011001000",
        13918=>"000000000",
        13919=>"011101111",
        13920=>"000010100",
        13921=>"110110111",
        13922=>"000000000",
        13923=>"000000000",
        13924=>"111111111",
        13925=>"000000000",
        13926=>"111110100",
        13927=>"001000000",
        13928=>"000010000",
        13929=>"000000000",
        13930=>"000001000",
        13931=>"101110100",
        13932=>"000000000",
        13933=>"111111111",
        13934=>"000000000",
        13935=>"000000100",
        13936=>"101110100",
        13937=>"010000000",
        13938=>"000000000",
        13939=>"000000000",
        13940=>"000111010",
        13941=>"001000000",
        13942=>"001111111",
        13943=>"000001111",
        13944=>"001001000",
        13945=>"000000000",
        13946=>"000000000",
        13947=>"000010010",
        13948=>"000000000",
        13949=>"001010010",
        13950=>"111001100",
        13951=>"110101111",
        13952=>"111111000",
        13953=>"111101100",
        13954=>"010111111",
        13955=>"000010000",
        13956=>"000001001",
        13957=>"111111111",
        13958=>"100000001",
        13959=>"000000111",
        13960=>"111011111",
        13961=>"110110111",
        13962=>"101001000",
        13963=>"100111101",
        13964=>"000001011",
        13965=>"111111000",
        13966=>"100011001",
        13967=>"000000011",
        13968=>"001100110",
        13969=>"111000100",
        13970=>"001001011",
        13971=>"000110001",
        13972=>"101000101",
        13973=>"111010000",
        13974=>"001000101",
        13975=>"000111111",
        13976=>"100100000",
        13977=>"011111001",
        13978=>"100000000",
        13979=>"010100011",
        13980=>"111111110",
        13981=>"100011000",
        13982=>"101000000",
        13983=>"010111000",
        13984=>"010000010",
        13985=>"000000001",
        13986=>"100110000",
        13987=>"100101011",
        13988=>"010111001",
        13989=>"000000000",
        13990=>"000000000",
        13991=>"100101101",
        13992=>"000001000",
        13993=>"000000010",
        13994=>"001001100",
        13995=>"111110110",
        13996=>"001001010",
        13997=>"010000000",
        13998=>"011010000",
        13999=>"010000000",
        14000=>"010000000",
        14001=>"011000000",
        14002=>"000101000",
        14003=>"111101000",
        14004=>"001100000",
        14005=>"100011100",
        14006=>"001111111",
        14007=>"010110000",
        14008=>"111101011",
        14009=>"000000101",
        14010=>"001010000",
        14011=>"111001000",
        14012=>"000000000",
        14013=>"011100000",
        14014=>"100111111",
        14015=>"101111111",
        14016=>"100000100",
        14017=>"000111101",
        14018=>"000000000",
        14019=>"000111111",
        14020=>"110100000",
        14021=>"110110100",
        14022=>"111101111",
        14023=>"000110010",
        14024=>"110000011",
        14025=>"111111000",
        14026=>"111001000",
        14027=>"000000101",
        14028=>"000010111",
        14029=>"000000000",
        14030=>"110100000",
        14031=>"000111110",
        14032=>"000000111",
        14033=>"100000001",
        14034=>"111111110",
        14035=>"000000100",
        14036=>"000011011",
        14037=>"000000111",
        14038=>"000111101",
        14039=>"111111111",
        14040=>"000100110",
        14041=>"111011000",
        14042=>"001001000",
        14043=>"000000000",
        14044=>"000011011",
        14045=>"011000100",
        14046=>"110111000",
        14047=>"111101001",
        14048=>"110100000",
        14049=>"110100100",
        14050=>"010111110",
        14051=>"000000111",
        14052=>"000101110",
        14053=>"001000000",
        14054=>"001000100",
        14055=>"011111110",
        14056=>"101000010",
        14057=>"000000000",
        14058=>"100110001",
        14059=>"010000010",
        14060=>"101000001",
        14061=>"000000111",
        14062=>"111111010",
        14063=>"100110010",
        14064=>"111000000",
        14065=>"001101011",
        14066=>"111101001",
        14067=>"000000000",
        14068=>"010001000",
        14069=>"000010111",
        14070=>"111111000",
        14071=>"000100100",
        14072=>"000010111",
        14073=>"000000110",
        14074=>"000000111",
        14075=>"010111111",
        14076=>"000110000",
        14077=>"111101010",
        14078=>"101010000",
        14079=>"000000000",
        14080=>"000010110",
        14081=>"010110010",
        14082=>"111110000",
        14083=>"111101000",
        14084=>"011000000",
        14085=>"111111111",
        14086=>"101111111",
        14087=>"001111001",
        14088=>"110000000",
        14089=>"001001011",
        14090=>"010111011",
        14091=>"100100100",
        14092=>"010000000",
        14093=>"111011111",
        14094=>"110000000",
        14095=>"111111000",
        14096=>"100000000",
        14097=>"111000111",
        14098=>"010000010",
        14099=>"010111010",
        14100=>"100100100",
        14101=>"110111010",
        14102=>"111111011",
        14103=>"100100000",
        14104=>"010000011",
        14105=>"001000001",
        14106=>"111000111",
        14107=>"111110110",
        14108=>"111110110",
        14109=>"000010011",
        14110=>"101000101",
        14111=>"100000111",
        14112=>"100000000",
        14113=>"111010001",
        14114=>"010000100",
        14115=>"111111111",
        14116=>"101101111",
        14117=>"100110000",
        14118=>"111011111",
        14119=>"000110010",
        14120=>"000101100",
        14121=>"000000000",
        14122=>"000110110",
        14123=>"000000011",
        14124=>"000101110",
        14125=>"100101100",
        14126=>"000001110",
        14127=>"010010010",
        14128=>"100000000",
        14129=>"010111000",
        14130=>"101100001",
        14131=>"100000100",
        14132=>"000000010",
        14133=>"110110000",
        14134=>"110100100",
        14135=>"111011000",
        14136=>"000110010",
        14137=>"101000000",
        14138=>"110100111",
        14139=>"111111110",
        14140=>"010010000",
        14141=>"010001111",
        14142=>"111001001",
        14143=>"010011010",
        14144=>"110111001",
        14145=>"110111111",
        14146=>"101101000",
        14147=>"010111111",
        14148=>"110110110",
        14149=>"111000111",
        14150=>"010111011",
        14151=>"100100000",
        14152=>"000010100",
        14153=>"000000000",
        14154=>"101111000",
        14155=>"000010000",
        14156=>"111111101",
        14157=>"110000000",
        14158=>"000000000",
        14159=>"010111010",
        14160=>"100111100",
        14161=>"010010110",
        14162=>"110110000",
        14163=>"100110000",
        14164=>"111000111",
        14165=>"010111010",
        14166=>"111100100",
        14167=>"000000110",
        14168=>"010000111",
        14169=>"000000111",
        14170=>"110010111",
        14171=>"111111001",
        14172=>"010000010",
        14173=>"110110000",
        14174=>"111010010",
        14175=>"000011000",
        14176=>"000000000",
        14177=>"000000101",
        14178=>"010010010",
        14179=>"010110000",
        14180=>"111101101",
        14181=>"010010000",
        14182=>"110010111",
        14183=>"100000000",
        14184=>"100111110",
        14185=>"011010010",
        14186=>"010000010",
        14187=>"000000000",
        14188=>"111010010",
        14189=>"010111010",
        14190=>"100010010",
        14191=>"000000000",
        14192=>"100110110",
        14193=>"101100000",
        14194=>"111000110",
        14195=>"100110000",
        14196=>"010111010",
        14197=>"100101100",
        14198=>"111111100",
        14199=>"101000110",
        14200=>"000010000",
        14201=>"101111100",
        14202=>"101111010",
        14203=>"101111000",
        14204=>"111001011",
        14205=>"100000000",
        14206=>"000010000",
        14207=>"010010010",
        14208=>"000000111",
        14209=>"000000010",
        14210=>"000101011",
        14211=>"011010111",
        14212=>"111110110",
        14213=>"111111111",
        14214=>"010000101",
        14215=>"110111101",
        14216=>"101011111",
        14217=>"101011111",
        14218=>"111000011",
        14219=>"101011110",
        14220=>"001000001",
        14221=>"001111000",
        14222=>"011100000",
        14223=>"000010001",
        14224=>"011011000",
        14225=>"111111010",
        14226=>"100110010",
        14227=>"001111110",
        14228=>"000001000",
        14229=>"111111111",
        14230=>"000100000",
        14231=>"011000001",
        14232=>"000001000",
        14233=>"101110000",
        14234=>"111111111",
        14235=>"110110000",
        14236=>"000000000",
        14237=>"011011111",
        14238=>"001100111",
        14239=>"111010111",
        14240=>"001010100",
        14241=>"000000100",
        14242=>"101010100",
        14243=>"000000101",
        14244=>"111011000",
        14245=>"000111000",
        14246=>"000000101",
        14247=>"010000000",
        14248=>"101111110",
        14249=>"111111100",
        14250=>"011000000",
        14251=>"110110110",
        14252=>"000110110",
        14253=>"010111111",
        14254=>"111000000",
        14255=>"000000000",
        14256=>"101101001",
        14257=>"100001111",
        14258=>"011011000",
        14259=>"011011011",
        14260=>"111101001",
        14261=>"110101000",
        14262=>"100101000",
        14263=>"110110111",
        14264=>"110100010",
        14265=>"100001000",
        14266=>"100110111",
        14267=>"010010100",
        14268=>"011011011",
        14269=>"000000010",
        14270=>"011001111",
        14271=>"000100010",
        14272=>"000000000",
        14273=>"100000111",
        14274=>"111111111",
        14275=>"000000000",
        14276=>"001000001",
        14277=>"011001010",
        14278=>"000010000",
        14279=>"000000010",
        14280=>"110110111",
        14281=>"110100000",
        14282=>"000100101",
        14283=>"111111010",
        14284=>"111101000",
        14285=>"111101010",
        14286=>"000000000",
        14287=>"111110111",
        14288=>"000100101",
        14289=>"010000000",
        14290=>"111100111",
        14291=>"110110100",
        14292=>"100100110",
        14293=>"000101100",
        14294=>"000000010",
        14295=>"111001010",
        14296=>"011011000",
        14297=>"000011111",
        14298=>"111100101",
        14299=>"001111111",
        14300=>"001011011",
        14301=>"001011000",
        14302=>"110110010",
        14303=>"111110111",
        14304=>"001000110",
        14305=>"110110111",
        14306=>"101101111",
        14307=>"111111010",
        14308=>"000000000",
        14309=>"110101000",
        14310=>"011000000",
        14311=>"101110111",
        14312=>"000000001",
        14313=>"111010000",
        14314=>"110110000",
        14315=>"101101111",
        14316=>"111111011",
        14317=>"111111111",
        14318=>"111101000",
        14319=>"110001000",
        14320=>"111111100",
        14321=>"001001000",
        14322=>"110000101",
        14323=>"000000000",
        14324=>"000111010",
        14325=>"001111101",
        14326=>"000000000",
        14327=>"110110101",
        14328=>"101111110",
        14329=>"100101000",
        14330=>"000001000",
        14331=>"110110101",
        14332=>"100001010",
        14333=>"110111111",
        14334=>"111011111",
        14335=>"101110111",
        14336=>"000110101",
        14337=>"111100110",
        14338=>"000000000",
        14339=>"000000000",
        14340=>"010001100",
        14341=>"000101011",
        14342=>"011101011",
        14343=>"101001101",
        14344=>"001111111",
        14345=>"011111100",
        14346=>"111001001",
        14347=>"011011001",
        14348=>"000111010",
        14349=>"010111111",
        14350=>"000000001",
        14351=>"001000000",
        14352=>"110111011",
        14353=>"101000000",
        14354=>"000011001",
        14355=>"000100011",
        14356=>"101000101",
        14357=>"011010101",
        14358=>"101000101",
        14359=>"100100111",
        14360=>"001100110",
        14361=>"110100000",
        14362=>"000000001",
        14363=>"011111111",
        14364=>"000001100",
        14365=>"011011001",
        14366=>"010001101",
        14367=>"010010010",
        14368=>"000101100",
        14369=>"110100100",
        14370=>"011001001",
        14371=>"000000000",
        14372=>"110111111",
        14373=>"100001000",
        14374=>"101101000",
        14375=>"000010110",
        14376=>"111111101",
        14377=>"110111111",
        14378=>"000101111",
        14379=>"001100010",
        14380=>"011001101",
        14381=>"001000100",
        14382=>"010010111",
        14383=>"110101100",
        14384=>"111110011",
        14385=>"000000000",
        14386=>"000000111",
        14387=>"000010111",
        14388=>"000100111",
        14389=>"110111101",
        14390=>"111111000",
        14391=>"000000000",
        14392=>"000100101",
        14393=>"000111011",
        14394=>"110111001",
        14395=>"001101111",
        14396=>"111101111",
        14397=>"000101010",
        14398=>"111110111",
        14399=>"101101111",
        14400=>"111111010",
        14401=>"000000000",
        14402=>"011000101",
        14403=>"111111101",
        14404=>"001111110",
        14405=>"000110110",
        14406=>"010111000",
        14407=>"110001000",
        14408=>"010111110",
        14409=>"000111111",
        14410=>"010001000",
        14411=>"101001101",
        14412=>"000011111",
        14413=>"000111011",
        14414=>"011111111",
        14415=>"000010000",
        14416=>"000111111",
        14417=>"011000000",
        14418=>"001111111",
        14419=>"000000000",
        14420=>"000010011",
        14421=>"111000000",
        14422=>"111100111",
        14423=>"000000000",
        14424=>"010110011",
        14425=>"101001110",
        14426=>"010001001",
        14427=>"001000000",
        14428=>"000001111",
        14429=>"100000000",
        14430=>"001000001",
        14431=>"111111111",
        14432=>"100111111",
        14433=>"000111110",
        14434=>"010111111",
        14435=>"000000000",
        14436=>"111001101",
        14437=>"001010010",
        14438=>"111000101",
        14439=>"111111000",
        14440=>"011111011",
        14441=>"101000000",
        14442=>"110100110",
        14443=>"110000000",
        14444=>"000111111",
        14445=>"110001001",
        14446=>"111111110",
        14447=>"000001110",
        14448=>"000111010",
        14449=>"111111111",
        14450=>"011000110",
        14451=>"000000000",
        14452=>"000000000",
        14453=>"000000101",
        14454=>"000000000",
        14455=>"101111111",
        14456=>"000110111",
        14457=>"101000101",
        14458=>"001110110",
        14459=>"111111010",
        14460=>"000100110",
        14461=>"110111111",
        14462=>"000010000",
        14463=>"000100000",
        14464=>"000000111",
        14465=>"100001011",
        14466=>"111011111",
        14467=>"000110011",
        14468=>"000001000",
        14469=>"010010010",
        14470=>"000010110",
        14471=>"111100001",
        14472=>"001011110",
        14473=>"000000000",
        14474=>"110000000",
        14475=>"111000011",
        14476=>"000110110",
        14477=>"110110110",
        14478=>"001101001",
        14479=>"000110100",
        14480=>"110000000",
        14481=>"100111001",
        14482=>"001011000",
        14483=>"000100101",
        14484=>"000110110",
        14485=>"100100111",
        14486=>"000000000",
        14487=>"110100110",
        14488=>"100101110",
        14489=>"110110100",
        14490=>"001001000",
        14491=>"001000000",
        14492=>"010010010",
        14493=>"100101011",
        14494=>"111111000",
        14495=>"001111101",
        14496=>"100101011",
        14497=>"100101001",
        14498=>"100100011",
        14499=>"111010000",
        14500=>"000110110",
        14501=>"010101101",
        14502=>"100001110",
        14503=>"000001011",
        14504=>"110110100",
        14505=>"110100111",
        14506=>"111111011",
        14507=>"000011011",
        14508=>"110000010",
        14509=>"000101101",
        14510=>"001100100",
        14511=>"111000000",
        14512=>"000000010",
        14513=>"111000100",
        14514=>"011100100",
        14515=>"000100100",
        14516=>"000011101",
        14517=>"000000100",
        14518=>"111110000",
        14519=>"100000110",
        14520=>"100001000",
        14521=>"110110101",
        14522=>"011011110",
        14523=>"010010110",
        14524=>"111001000",
        14525=>"001011100",
        14526=>"001111100",
        14527=>"000010011",
        14528=>"110010100",
        14529=>"100100110",
        14530=>"110110110",
        14531=>"001011110",
        14532=>"000111111",
        14533=>"000000111",
        14534=>"010001110",
        14535=>"110110100",
        14536=>"000111010",
        14537=>"000001111",
        14538=>"110100000",
        14539=>"001000000",
        14540=>"110100110",
        14541=>"110011111",
        14542=>"111100100",
        14543=>"001001010",
        14544=>"110110110",
        14545=>"000011110",
        14546=>"110000000",
        14547=>"110110110",
        14548=>"110000111",
        14549=>"100100100",
        14550=>"000110110",
        14551=>"000100101",
        14552=>"101111101",
        14553=>"011000001",
        14554=>"001011111",
        14555=>"000000010",
        14556=>"000001001",
        14557=>"111000100",
        14558=>"010001101",
        14559=>"100000000",
        14560=>"000001011",
        14561=>"000100110",
        14562=>"001011011",
        14563=>"010110110",
        14564=>"110111100",
        14565=>"001011110",
        14566=>"100000001",
        14567=>"010100100",
        14568=>"110110011",
        14569=>"101000001",
        14570=>"100011011",
        14571=>"111110101",
        14572=>"000001011",
        14573=>"001011100",
        14574=>"110100110",
        14575=>"000001001",
        14576=>"000000100",
        14577=>"001010110",
        14578=>"000001011",
        14579=>"001001000",
        14580=>"101001111",
        14581=>"000000001",
        14582=>"000100011",
        14583=>"110110010",
        14584=>"011000100",
        14585=>"111110100",
        14586=>"110100111",
        14587=>"010100000",
        14588=>"100000000",
        14589=>"110000000",
        14590=>"111000100",
        14591=>"001011110",
        14592=>"000111010",
        14593=>"111000000",
        14594=>"100010011",
        14595=>"011111111",
        14596=>"011001001",
        14597=>"100000010",
        14598=>"101111111",
        14599=>"110000101",
        14600=>"000000111",
        14601=>"100100110",
        14602=>"000110000",
        14603=>"110001000",
        14604=>"110000000",
        14605=>"010111111",
        14606=>"000110000",
        14607=>"001011000",
        14608=>"001001100",
        14609=>"110111000",
        14610=>"000001101",
        14611=>"000000010",
        14612=>"001101101",
        14613=>"001011010",
        14614=>"111101100",
        14615=>"111101001",
        14616=>"001100100",
        14617=>"011100000",
        14618=>"010000100",
        14619=>"100100100",
        14620=>"000000000",
        14621=>"011100001",
        14622=>"100100010",
        14623=>"000111111",
        14624=>"111111101",
        14625=>"111111110",
        14626=>"010001100",
        14627=>"111111111",
        14628=>"111111001",
        14629=>"110101000",
        14630=>"111101100",
        14631=>"000110111",
        14632=>"111011000",
        14633=>"111010000",
        14634=>"011100000",
        14635=>"000100000",
        14636=>"111001001",
        14637=>"100011001",
        14638=>"000110111",
        14639=>"011111110",
        14640=>"110011000",
        14641=>"100111111",
        14642=>"111001000",
        14643=>"000110110",
        14644=>"011001101",
        14645=>"000000000",
        14646=>"010001000",
        14647=>"100111111",
        14648=>"111100000",
        14649=>"110000000",
        14650=>"011101110",
        14651=>"100110111",
        14652=>"000011000",
        14653=>"000000000",
        14654=>"000001001",
        14655=>"111100100",
        14656=>"111100011",
        14657=>"000000110",
        14658=>"111101101",
        14659=>"000000000",
        14660=>"000111111",
        14661=>"000011001",
        14662=>"000010101",
        14663=>"111000000",
        14664=>"000100001",
        14665=>"011001111",
        14666=>"111100110",
        14667=>"011001101",
        14668=>"100111000",
        14669=>"000010000",
        14670=>"000010111",
        14671=>"000110111",
        14672=>"001010001",
        14673=>"111001110",
        14674=>"001100100",
        14675=>"000001000",
        14676=>"000100100",
        14677=>"101000000",
        14678=>"111101101",
        14679=>"000000101",
        14680=>"110100100",
        14681=>"111000110",
        14682=>"000000001",
        14683=>"000111111",
        14684=>"001000001",
        14685=>"100000100",
        14686=>"000000100",
        14687=>"000000000",
        14688=>"000100110",
        14689=>"000011001",
        14690=>"000010111",
        14691=>"000100000",
        14692=>"111101000",
        14693=>"000001111",
        14694=>"011100000",
        14695=>"011100101",
        14696=>"000000000",
        14697=>"111000000",
        14698=>"000001001",
        14699=>"101111010",
        14700=>"000000110",
        14701=>"000001000",
        14702=>"111101001",
        14703=>"010000000",
        14704=>"000011111",
        14705=>"000100111",
        14706=>"000101101",
        14707=>"111000000",
        14708=>"000110111",
        14709=>"001000111",
        14710=>"100000000",
        14711=>"111100101",
        14712=>"111100101",
        14713=>"111111000",
        14714=>"000000000",
        14715=>"000000000",
        14716=>"000000110",
        14717=>"111100000",
        14718=>"111111000",
        14719=>"111100111",
        14720=>"000001001",
        14721=>"110110110",
        14722=>"110110100",
        14723=>"111111011",
        14724=>"000000000",
        14725=>"110011111",
        14726=>"011001011",
        14727=>"110100100",
        14728=>"100101001",
        14729=>"001011011",
        14730=>"111110110",
        14731=>"001101010",
        14732=>"010000010",
        14733=>"110001100",
        14734=>"000000000",
        14735=>"110110111",
        14736=>"111010010",
        14737=>"110111011",
        14738=>"001001100",
        14739=>"000100110",
        14740=>"100110111",
        14741=>"010000001",
        14742=>"110010110",
        14743=>"110101001",
        14744=>"111011001",
        14745=>"001111111",
        14746=>"101101101",
        14747=>"001001001",
        14748=>"000001001",
        14749=>"000000000",
        14750=>"000001000",
        14751=>"101111100",
        14752=>"011001000",
        14753=>"001100100",
        14754=>"011000000",
        14755=>"011111011",
        14756=>"111011011",
        14757=>"110110101",
        14758=>"110110010",
        14759=>"010001011",
        14760=>"110110110",
        14761=>"001111111",
        14762=>"000000000",
        14763=>"000000000",
        14764=>"111001000",
        14765=>"001110100",
        14766=>"001001001",
        14767=>"010110000",
        14768=>"110100101",
        14769=>"110100110",
        14770=>"011001000",
        14771=>"001101101",
        14772=>"011111101",
        14773=>"001011001",
        14774=>"001001011",
        14775=>"011001000",
        14776=>"110110111",
        14777=>"011001001",
        14778=>"011001101",
        14779=>"000110110",
        14780=>"110110111",
        14781=>"010011111",
        14782=>"011000001",
        14783=>"001001011",
        14784=>"111010001",
        14785=>"110110100",
        14786=>"001001001",
        14787=>"100100111",
        14788=>"101000010",
        14789=>"000000011",
        14790=>"001001011",
        14791=>"111110011",
        14792=>"000110110",
        14793=>"001001001",
        14794=>"111110101",
        14795=>"110000000",
        14796=>"011110010",
        14797=>"001001001",
        14798=>"011101111",
        14799=>"110110110",
        14800=>"110110110",
        14801=>"100110110",
        14802=>"001001001",
        14803=>"010000001",
        14804=>"111000001",
        14805=>"100100101",
        14806=>"001111001",
        14807=>"110001101",
        14808=>"100000000",
        14809=>"001001010",
        14810=>"100100100",
        14811=>"110110100",
        14812=>"001101001",
        14813=>"111100000",
        14814=>"100000000",
        14815=>"001000000",
        14816=>"110000000",
        14817=>"111001001",
        14818=>"100110110",
        14819=>"100110100",
        14820=>"110110011",
        14821=>"000110110",
        14822=>"010000000",
        14823=>"010110110",
        14824=>"110110100",
        14825=>"001001001",
        14826=>"000001001",
        14827=>"001001100",
        14828=>"001001001",
        14829=>"010000001",
        14830=>"011001001",
        14831=>"001001011",
        14832=>"111010110",
        14833=>"101000000",
        14834=>"110110011",
        14835=>"001001001",
        14836=>"111000000",
        14837=>"110110110",
        14838=>"110010000",
        14839=>"001110010",
        14840=>"001100010",
        14841=>"111110110",
        14842=>"110110010",
        14843=>"011110110",
        14844=>"000000100",
        14845=>"011011111",
        14846=>"001001000",
        14847=>"001001000",
        14848=>"011111111",
        14849=>"000011111",
        14850=>"101110111",
        14851=>"000000100",
        14852=>"000001111",
        14853=>"101010011",
        14854=>"100110111",
        14855=>"001001101",
        14856=>"100101011",
        14857=>"100101101",
        14858=>"100000001",
        14859=>"011000011",
        14860=>"000010001",
        14861=>"111001111",
        14862=>"100100100",
        14863=>"010000011",
        14864=>"001011111",
        14865=>"000110110",
        14866=>"100000000",
        14867=>"100100100",
        14868=>"010100100",
        14869=>"000011000",
        14870=>"010111111",
        14871=>"111010000",
        14872=>"110100000",
        14873=>"110100000",
        14874=>"100000010",
        14875=>"000001100",
        14876=>"000001000",
        14877=>"110100101",
        14878=>"100110110",
        14879=>"101111111",
        14880=>"111100000",
        14881=>"100101101",
        14882=>"001001011",
        14883=>"100000100",
        14884=>"010110100",
        14885=>"000000100",
        14886=>"000011111",
        14887=>"001110100",
        14888=>"110100000",
        14889=>"100000000",
        14890=>"111001000",
        14891=>"110100100",
        14892=>"101001001",
        14893=>"110111100",
        14894=>"000000111",
        14895=>"111000100",
        14896=>"110100110",
        14897=>"001011101",
        14898=>"110111110",
        14899=>"001011000",
        14900=>"100001001",
        14901=>"001000000",
        14902=>"111101010",
        14903=>"010111011",
        14904=>"100011111",
        14905=>"111000001",
        14906=>"100100010",
        14907=>"000011011",
        14908=>"000010000",
        14909=>"001000000",
        14910=>"111111101",
        14911=>"101100001",
        14912=>"110100000",
        14913=>"000000010",
        14914=>"110001000",
        14915=>"000011111",
        14916=>"110000110",
        14917=>"110110110",
        14918=>"100000010",
        14919=>"000000011",
        14920=>"111110000",
        14921=>"000001100",
        14922=>"011000000",
        14923=>"000000000",
        14924=>"011000011",
        14925=>"001000111",
        14926=>"011011011",
        14927=>"001011110",
        14928=>"000011011",
        14929=>"100110010",
        14930=>"000000110",
        14931=>"001011110",
        14932=>"111000101",
        14933=>"011011011",
        14934=>"001000000",
        14935=>"010110101",
        14936=>"100100010",
        14937=>"100110111",
        14938=>"000001011",
        14939=>"011010110",
        14940=>"100100000",
        14941=>"001011111",
        14942=>"000001111",
        14943=>"001001011",
        14944=>"111101101",
        14945=>"011111101",
        14946=>"011111100",
        14947=>"100100000",
        14948=>"100010011",
        14949=>"000111000",
        14950=>"001011011",
        14951=>"100100110",
        14952=>"011011111",
        14953=>"100000000",
        14954=>"110100000",
        14955=>"011111010",
        14956=>"001011110",
        14957=>"000011111",
        14958=>"000000000",
        14959=>"001000001",
        14960=>"111001011",
        14961=>"000011111",
        14962=>"000011001",
        14963=>"110100100",
        14964=>"011011111",
        14965=>"001011110",
        14966=>"011111100",
        14967=>"110000000",
        14968=>"100011111",
        14969=>"110100010",
        14970=>"000010110",
        14971=>"111011011",
        14972=>"100100100",
        14973=>"110101010",
        14974=>"110110000",
        14975=>"100100001",
        14976=>"011111111",
        14977=>"010010000",
        14978=>"111010010",
        14979=>"110010010",
        14980=>"000000100",
        14981=>"101010110",
        14982=>"110010110",
        14983=>"101101101",
        14984=>"000001100",
        14985=>"000000001",
        14986=>"111001111",
        14987=>"110100100",
        14988=>"000000100",
        14989=>"111111000",
        14990=>"110110110",
        14991=>"101101101",
        14992=>"111101111",
        14993=>"000111010",
        14994=>"110100111",
        14995=>"000011001",
        14996=>"000000101",
        14997=>"100100000",
        14998=>"000100001",
        14999=>"001101001",
        15000=>"111110101",
        15001=>"001000001",
        15002=>"110010010",
        15003=>"100000000",
        15004=>"110110000",
        15005=>"011010110",
        15006=>"001101111",
        15007=>"101101101",
        15008=>"000000000",
        15009=>"111000000",
        15010=>"000000000",
        15011=>"001111111",
        15012=>"000000000",
        15013=>"011110111",
        15014=>"101111001",
        15015=>"010110010",
        15016=>"010101101",
        15017=>"001011011",
        15018=>"110111111",
        15019=>"001011001",
        15020=>"001100101",
        15021=>"101101101",
        15022=>"000000000",
        15023=>"000111000",
        15024=>"101111101",
        15025=>"000000000",
        15026=>"001101101",
        15027=>"100001111",
        15028=>"110011110",
        15029=>"000000000",
        15030=>"001101000",
        15031=>"110000010",
        15032=>"111011101",
        15033=>"101000001",
        15034=>"000000110",
        15035=>"000100101",
        15036=>"101101101",
        15037=>"000000011",
        15038=>"001000000",
        15039=>"010110111",
        15040=>"111110111",
        15041=>"100101000",
        15042=>"000100101",
        15043=>"101100000",
        15044=>"000000001",
        15045=>"111101100",
        15046=>"000000100",
        15047=>"111100111",
        15048=>"101000101",
        15049=>"110110010",
        15050=>"101100101",
        15051=>"101101000",
        15052=>"101000001",
        15053=>"010011011",
        15054=>"101101001",
        15055=>"111111100",
        15056=>"000101101",
        15057=>"000010000",
        15058=>"000100101",
        15059=>"111011011",
        15060=>"100110111",
        15061=>"001000001",
        15062=>"010010010",
        15063=>"000000010",
        15064=>"000100110",
        15065=>"000101111",
        15066=>"001011000",
        15067=>"100001011",
        15068=>"000100110",
        15069=>"100110000",
        15070=>"111111011",
        15071=>"000000101",
        15072=>"001000000",
        15073=>"111111111",
        15074=>"011011111",
        15075=>"010010000",
        15076=>"001001000",
        15077=>"001101001",
        15078=>"000000000",
        15079=>"101100101",
        15080=>"001010010",
        15081=>"000100000",
        15082=>"011011011",
        15083=>"000101101",
        15084=>"010000110",
        15085=>"001101000",
        15086=>"010100010",
        15087=>"111010011",
        15088=>"100000101",
        15089=>"101110100",
        15090=>"000110010",
        15091=>"111001000",
        15092=>"000001101",
        15093=>"000000100",
        15094=>"011110000",
        15095=>"101110111",
        15096=>"100001101",
        15097=>"101001101",
        15098=>"000000000",
        15099=>"001000000",
        15100=>"111111110",
        15101=>"111001100",
        15102=>"101011111",
        15103=>"000010000",
        15104=>"111101111",
        15105=>"010010010",
        15106=>"111000000",
        15107=>"101111000",
        15108=>"100110111",
        15109=>"111111101",
        15110=>"000010101",
        15111=>"111111010",
        15112=>"111110111",
        15113=>"111111111",
        15114=>"101110000",
        15115=>"100111011",
        15116=>"110110101",
        15117=>"110000000",
        15118=>"010110110",
        15119=>"111101000",
        15120=>"000001001",
        15121=>"111110010",
        15122=>"100111110",
        15123=>"011011110",
        15124=>"000000101",
        15125=>"000000011",
        15126=>"100010000",
        15127=>"000010000",
        15128=>"011111111",
        15129=>"000110100",
        15130=>"010010111",
        15131=>"100000100",
        15132=>"100010000",
        15133=>"000010110",
        15134=>"110111111",
        15135=>"010000100",
        15136=>"000000010",
        15137=>"000000000",
        15138=>"000110011",
        15139=>"001111111",
        15140=>"111101111",
        15141=>"001111101",
        15142=>"111000100",
        15143=>"100111011",
        15144=>"000101010",
        15145=>"001111110",
        15146=>"111000010",
        15147=>"001110110",
        15148=>"100111011",
        15149=>"000101111",
        15150=>"101111111",
        15151=>"111111110",
        15152=>"011010010",
        15153=>"110010000",
        15154=>"000000000",
        15155=>"001010111",
        15156=>"000010011",
        15157=>"000000111",
        15158=>"101101000",
        15159=>"000000000",
        15160=>"111000010",
        15161=>"000000000",
        15162=>"101111111",
        15163=>"110100000",
        15164=>"111001010",
        15165=>"000001000",
        15166=>"001001011",
        15167=>"001101111",
        15168=>"000001111",
        15169=>"010000000",
        15170=>"001000000",
        15171=>"110110000",
        15172=>"101111001",
        15173=>"001011101",
        15174=>"010001110",
        15175=>"101000000",
        15176=>"100110111",
        15177=>"000000111",
        15178=>"101111111",
        15179=>"010010000",
        15180=>"101100000",
        15181=>"000100111",
        15182=>"000010000",
        15183=>"111011000",
        15184=>"000100011",
        15185=>"111110110",
        15186=>"000001111",
        15187=>"100000110",
        15188=>"000100101",
        15189=>"110010011",
        15190=>"000000000",
        15191=>"111101111",
        15192=>"000110011",
        15193=>"111111111",
        15194=>"000100110",
        15195=>"111000000",
        15196=>"000111110",
        15197=>"111111111",
        15198=>"010110010",
        15199=>"010000000",
        15200=>"010010111",
        15201=>"100100000",
        15202=>"111001000",
        15203=>"110111010",
        15204=>"100101000",
        15205=>"000101000",
        15206=>"101111111",
        15207=>"101111101",
        15208=>"101101111",
        15209=>"111111101",
        15210=>"000111110",
        15211=>"111111111",
        15212=>"010001000",
        15213=>"010110111",
        15214=>"000001101",
        15215=>"111110011",
        15216=>"100100000",
        15217=>"000100000",
        15218=>"000010111",
        15219=>"000000100",
        15220=>"111010000",
        15221=>"001101011",
        15222=>"111111100",
        15223=>"000000000",
        15224=>"100101011",
        15225=>"101101000",
        15226=>"101111110",
        15227=>"101000000",
        15228=>"011011010",
        15229=>"110000001",
        15230=>"111111111",
        15231=>"001000010",
        15232=>"010010010",
        15233=>"010000010",
        15234=>"001000101",
        15235=>"111101110",
        15236=>"111011010",
        15237=>"010110110",
        15238=>"000111111",
        15239=>"001001001",
        15240=>"111101011",
        15241=>"100100000",
        15242=>"000000000",
        15243=>"001001100",
        15244=>"001001001",
        15245=>"010111000",
        15246=>"011011111",
        15247=>"101100100",
        15248=>"001101100",
        15249=>"001001111",
        15250=>"001001011",
        15251=>"110100000",
        15252=>"001001011",
        15253=>"110101010",
        15254=>"000001010",
        15255=>"000101110",
        15256=>"000101101",
        15257=>"100001011",
        15258=>"000001101",
        15259=>"011111101",
        15260=>"110110111",
        15261=>"001001010",
        15262=>"110111011",
        15263=>"000011111",
        15264=>"001101111",
        15265=>"000000011",
        15266=>"001010100",
        15267=>"101000111",
        15268=>"000000110",
        15269=>"000000111",
        15270=>"001001111",
        15271=>"111100000",
        15272=>"000001101",
        15273=>"000001000",
        15274=>"101101100",
        15275=>"110100100",
        15276=>"111001001",
        15277=>"111000111",
        15278=>"001000000",
        15279=>"101101111",
        15280=>"001001001",
        15281=>"001001001",
        15282=>"000101100",
        15283=>"111000101",
        15284=>"110110110",
        15285=>"000000110",
        15286=>"110110110",
        15287=>"000000000",
        15288=>"000000111",
        15289=>"111000000",
        15290=>"001001110",
        15291=>"110110000",
        15292=>"101001001",
        15293=>"001001010",
        15294=>"010110101",
        15295=>"101111111",
        15296=>"011110100",
        15297=>"000001010",
        15298=>"101111110",
        15299=>"110111011",
        15300=>"110100111",
        15301=>"000000000",
        15302=>"000001101",
        15303=>"110001000",
        15304=>"001001101",
        15305=>"111110000",
        15306=>"000000000",
        15307=>"000001001",
        15308=>"100111000",
        15309=>"111110000",
        15310=>"101110001",
        15311=>"001001111",
        15312=>"000000000",
        15313=>"000000101",
        15314=>"000000110",
        15315=>"110111111",
        15316=>"001001001",
        15317=>"001001001",
        15318=>"011111111",
        15319=>"111111111",
        15320=>"000000001",
        15321=>"000111111",
        15322=>"001011111",
        15323=>"001111111",
        15324=>"011000110",
        15325=>"001000001",
        15326=>"011011001",
        15327=>"111111110",
        15328=>"011011000",
        15329=>"101100001",
        15330=>"011110000",
        15331=>"110111111",
        15332=>"101000100",
        15333=>"000000101",
        15334=>"100000011",
        15335=>"000001111",
        15336=>"101000100",
        15337=>"111101001",
        15338=>"000011001",
        15339=>"111101000",
        15340=>"001000001",
        15341=>"010010000",
        15342=>"000111000",
        15343=>"000100000",
        15344=>"001000101",
        15345=>"000101101",
        15346=>"111100000",
        15347=>"010110000",
        15348=>"010001010",
        15349=>"101001001",
        15350=>"100001111",
        15351=>"001011110",
        15352=>"001000001",
        15353=>"010000110",
        15354=>"111010000",
        15355=>"101001111",
        15356=>"000000100",
        15357=>"111111110",
        15358=>"000000111",
        15359=>"110011010",
        15360=>"000000000",
        15361=>"000000011",
        15362=>"000011001",
        15363=>"000111101",
        15364=>"111101111",
        15365=>"111010010",
        15366=>"000000000",
        15367=>"000101100",
        15368=>"110001001",
        15369=>"000001111",
        15370=>"000110111",
        15371=>"000101101",
        15372=>"110000000",
        15373=>"110110100",
        15374=>"110111011",
        15375=>"100111111",
        15376=>"111000000",
        15377=>"000000111",
        15378=>"011001000",
        15379=>"011001001",
        15380=>"000001101",
        15381=>"111000000",
        15382=>"000000000",
        15383=>"111110101",
        15384=>"111000001",
        15385=>"110111110",
        15386=>"010000000",
        15387=>"111100100",
        15388=>"111111111",
        15389=>"011001000",
        15390=>"000100100",
        15391=>"101111111",
        15392=>"111110101",
        15393=>"001100000",
        15394=>"111100110",
        15395=>"110000100",
        15396=>"000000000",
        15397=>"110111111",
        15398=>"111111111",
        15399=>"000000000",
        15400=>"000111110",
        15401=>"000100111",
        15402=>"000000100",
        15403=>"001000000",
        15404=>"111110110",
        15405=>"000000100",
        15406=>"111001101",
        15407=>"000111101",
        15408=>"000000100",
        15409=>"000111100",
        15410=>"111111011",
        15411=>"000000000",
        15412=>"111000000",
        15413=>"111111101",
        15414=>"111111111",
        15415=>"110111000",
        15416=>"000000000",
        15417=>"111111101",
        15418=>"000100110",
        15419=>"111000000",
        15420=>"001000100",
        15421=>"110000000",
        15422=>"111011001",
        15423=>"111111000",
        15424=>"011111111",
        15425=>"011001000",
        15426=>"111111111",
        15427=>"100000101",
        15428=>"111100000",
        15429=>"111010000",
        15430=>"111100100",
        15431=>"111000001",
        15432=>"111000000",
        15433=>"000000000",
        15434=>"111100111",
        15435=>"000000100",
        15436=>"100111111",
        15437=>"111111111",
        15438=>"011101000",
        15439=>"000111010",
        15440=>"101101111",
        15441=>"011000001",
        15442=>"111111000",
        15443=>"100111010",
        15444=>"111000000",
        15445=>"111111111",
        15446=>"111111011",
        15447=>"111010000",
        15448=>"000010001",
        15449=>"011100111",
        15450=>"110000100",
        15451=>"000000000",
        15452=>"000000100",
        15453=>"110110110",
        15454=>"000000000",
        15455=>"001001000",
        15456=>"011000010",
        15457=>"000000000",
        15458=>"000100101",
        15459=>"000110111",
        15460=>"111010111",
        15461=>"000000111",
        15462=>"011000000",
        15463=>"000101100",
        15464=>"000000000",
        15465=>"000001011",
        15466=>"000000000",
        15467=>"111111101",
        15468=>"000000000",
        15469=>"000101101",
        15470=>"111111110",
        15471=>"010111100",
        15472=>"000010000",
        15473=>"001000111",
        15474=>"000000000",
        15475=>"011111101",
        15476=>"111111111",
        15477=>"000000100",
        15478=>"101100100",
        15479=>"111111111",
        15480=>"100110111",
        15481=>"100000000",
        15482=>"000000000",
        15483=>"100111010",
        15484=>"000000001",
        15485=>"111111000",
        15486=>"001101111",
        15487=>"011000101",
        15488=>"111111011",
        15489=>"011010011",
        15490=>"000000010",
        15491=>"010110100",
        15492=>"110011011",
        15493=>"100111010",
        15494=>"000000110",
        15495=>"101100000",
        15496=>"110000000",
        15497=>"100000000",
        15498=>"000000110",
        15499=>"011001000",
        15500=>"101111001",
        15501=>"111010010",
        15502=>"110001000",
        15503=>"000101011",
        15504=>"111001000",
        15505=>"111111101",
        15506=>"001000111",
        15507=>"011000100",
        15508=>"000001110",
        15509=>"111111000",
        15510=>"011000000",
        15511=>"000000010",
        15512=>"000000111",
        15513=>"101001000",
        15514=>"111000100",
        15515=>"011111000",
        15516=>"000010111",
        15517=>"010100011",
        15518=>"000101111",
        15519=>"000000011",
        15520=>"011111100",
        15521=>"000000000",
        15522=>"101111100",
        15523=>"000111110",
        15524=>"000110000",
        15525=>"000100011",
        15526=>"111111000",
        15527=>"111100000",
        15528=>"001000010",
        15529=>"001000111",
        15530=>"111110100",
        15531=>"000000110",
        15532=>"000010011",
        15533=>"000001111",
        15534=>"000010100",
        15535=>"111111000",
        15536=>"111001000",
        15537=>"110100111",
        15538=>"101111000",
        15539=>"101111111",
        15540=>"000010110",
        15541=>"000111111",
        15542=>"000000011",
        15543=>"000000111",
        15544=>"100000010",
        15545=>"000000010",
        15546=>"001100100",
        15547=>"111100000",
        15548=>"111000000",
        15549=>"110101000",
        15550=>"010110101",
        15551=>"000001111",
        15552=>"010010011",
        15553=>"111101100",
        15554=>"000000011",
        15555=>"011000000",
        15556=>"101100111",
        15557=>"111110000",
        15558=>"000000111",
        15559=>"010011111",
        15560=>"011100000",
        15561=>"000000111",
        15562=>"000010111",
        15563=>"011101000",
        15564=>"111100101",
        15565=>"000010111",
        15566=>"010111100",
        15567=>"111111001",
        15568=>"011110110",
        15569=>"111000000",
        15570=>"000000111",
        15571=>"000000010",
        15572=>"011011000",
        15573=>"101000000",
        15574=>"110000001",
        15575=>"100011100",
        15576=>"111100011",
        15577=>"011000000",
        15578=>"111011000",
        15579=>"111111000",
        15580=>"111001011",
        15581=>"110000110",
        15582=>"011111100",
        15583=>"000010011",
        15584=>"011001100",
        15585=>"100100011",
        15586=>"101100010",
        15587=>"111000000",
        15588=>"111111111",
        15589=>"111101000",
        15590=>"111100000",
        15591=>"110010111",
        15592=>"111011000",
        15593=>"101100000",
        15594=>"000000000",
        15595=>"110111111",
        15596=>"011001110",
        15597=>"000000000",
        15598=>"000000111",
        15599=>"001000010",
        15600=>"000000111",
        15601=>"001101111",
        15602=>"111100100",
        15603=>"000111111",
        15604=>"011111101",
        15605=>"111101000",
        15606=>"111011000",
        15607=>"110100100",
        15608=>"000001011",
        15609=>"000100000",
        15610=>"111101000",
        15611=>"111000000",
        15612=>"111010001",
        15613=>"110011111",
        15614=>"000000011",
        15615=>"101011111",
        15616=>"000000010",
        15617=>"111111110",
        15618=>"010011000",
        15619=>"111110111",
        15620=>"011000000",
        15621=>"000001010",
        15622=>"110001000",
        15623=>"000111000",
        15624=>"011101001",
        15625=>"111110100",
        15626=>"101111110",
        15627=>"111110000",
        15628=>"000100001",
        15629=>"101100101",
        15630=>"111111110",
        15631=>"011011000",
        15632=>"000000000",
        15633=>"000110000",
        15634=>"111111101",
        15635=>"000000000",
        15636=>"000110111",
        15637=>"000000000",
        15638=>"000110000",
        15639=>"110111100",
        15640=>"110110000",
        15641=>"101000000",
        15642=>"110111000",
        15643=>"111110110",
        15644=>"111101000",
        15645=>"101100000",
        15646=>"111111111",
        15647=>"000000001",
        15648=>"111111110",
        15649=>"000000000",
        15650=>"011000000",
        15651=>"001000000",
        15652=>"111000000",
        15653=>"110000110",
        15654=>"101111111",
        15655=>"111111111",
        15656=>"111110100",
        15657=>"111111110",
        15658=>"000010100",
        15659=>"011111110",
        15660=>"110110011",
        15661=>"111001001",
        15662=>"010000000",
        15663=>"111111111",
        15664=>"111101110",
        15665=>"100111000",
        15666=>"011111011",
        15667=>"010010000",
        15668=>"110000000",
        15669=>"111111001",
        15670=>"000000000",
        15671=>"001001001",
        15672=>"101110111",
        15673=>"111101111",
        15674=>"011010011",
        15675=>"000111111",
        15676=>"001001111",
        15677=>"011111000",
        15678=>"111111011",
        15679=>"000011100",
        15680=>"000000000",
        15681=>"011110100",
        15682=>"000111111",
        15683=>"111111101",
        15684=>"110011000",
        15685=>"111100100",
        15686=>"111111110",
        15687=>"111111000",
        15688=>"100110000",
        15689=>"000000000",
        15690=>"000110010",
        15691=>"000000000",
        15692=>"110000000",
        15693=>"111111100",
        15694=>"000010000",
        15695=>"111000000",
        15696=>"000101001",
        15697=>"000001111",
        15698=>"111111000",
        15699=>"010000000",
        15700=>"101001011",
        15701=>"000101101",
        15702=>"000100000",
        15703=>"111111111",
        15704=>"111111111",
        15705=>"111001000",
        15706=>"111110110",
        15707=>"011000000",
        15708=>"110111011",
        15709=>"011100000",
        15710=>"100111110",
        15711=>"000000000",
        15712=>"101001001",
        15713=>"000000000",
        15714=>"011111010",
        15715=>"111101110",
        15716=>"010000000",
        15717=>"000000000",
        15718=>"100110111",
        15719=>"111110110",
        15720=>"111011010",
        15721=>"110110010",
        15722=>"011011011",
        15723=>"110100011",
        15724=>"000000000",
        15725=>"101101111",
        15726=>"000010001",
        15727=>"110111000",
        15728=>"000001001",
        15729=>"111111000",
        15730=>"111111111",
        15731=>"000000000",
        15732=>"111110100",
        15733=>"011111000",
        15734=>"110100000",
        15735=>"111111110",
        15736=>"111111100",
        15737=>"110000000",
        15738=>"110100110",
        15739=>"111111010",
        15740=>"011111011",
        15741=>"111110000",
        15742=>"111110000",
        15743=>"101100000",
        15744=>"110110001",
        15745=>"111101000",
        15746=>"101101111",
        15747=>"111110101",
        15748=>"001011001",
        15749=>"110100000",
        15750=>"000111011",
        15751=>"001101101",
        15752=>"100100100",
        15753=>"000000000",
        15754=>"001101000",
        15755=>"001001001",
        15756=>"100111111",
        15757=>"100111111",
        15758=>"011000110",
        15759=>"100100100",
        15760=>"001001001",
        15761=>"001100101",
        15762=>"110000011",
        15763=>"001000100",
        15764=>"010010000",
        15765=>"010110111",
        15766=>"111001100",
        15767=>"001001000",
        15768=>"010110110",
        15769=>"100100100",
        15770=>"010000000",
        15771=>"011010110",
        15772=>"000000010",
        15773=>"000000001",
        15774=>"000011011",
        15775=>"111001101",
        15776=>"010111111",
        15777=>"011100001",
        15778=>"010010111",
        15779=>"000001000",
        15780=>"100010100",
        15781=>"001111001",
        15782=>"101101001",
        15783=>"010010010",
        15784=>"111011000",
        15785=>"100111110",
        15786=>"110111111",
        15787=>"000000010",
        15788=>"001001011",
        15789=>"101011001",
        15790=>"000000000",
        15791=>"010000111",
        15792=>"011011000",
        15793=>"100000001",
        15794=>"001011011",
        15795=>"101110110",
        15796=>"000010010",
        15797=>"010010000",
        15798=>"100100000",
        15799=>"111101010",
        15800=>"101101100",
        15801=>"011111101",
        15802=>"100100100",
        15803=>"000000110",
        15804=>"011101101",
        15805=>"000000101",
        15806=>"010001011",
        15807=>"111110000",
        15808=>"100000010",
        15809=>"000010101",
        15810=>"111101101",
        15811=>"100100100",
        15812=>"000011101",
        15813=>"001000110",
        15814=>"111111111",
        15815=>"001100000",
        15816=>"000100100",
        15817=>"010010010",
        15818=>"011001001",
        15819=>"001000000",
        15820=>"110010110",
        15821=>"010111000",
        15822=>"110100101",
        15823=>"000000001",
        15824=>"100100000",
        15825=>"100100100",
        15826=>"011011111",
        15827=>"100011100",
        15828=>"001001000",
        15829=>"101000000",
        15830=>"111110111",
        15831=>"111111000",
        15832=>"011001010",
        15833=>"000010010",
        15834=>"001100100",
        15835=>"100001010",
        15836=>"100100100",
        15837=>"000001001",
        15838=>"011110111",
        15839=>"000111010",
        15840=>"011001001",
        15841=>"010010000",
        15842=>"011001000",
        15843=>"000010001",
        15844=>"001101101",
        15845=>"101000110",
        15846=>"001001001",
        15847=>"101111100",
        15848=>"100100100",
        15849=>"010100001",
        15850=>"000000000",
        15851=>"001010111",
        15852=>"011001000",
        15853=>"101100000",
        15854=>"101010000",
        15855=>"011000001",
        15856=>"101001101",
        15857=>"100001100",
        15858=>"000100100",
        15859=>"100110100",
        15860=>"101000000",
        15861=>"000100000",
        15862=>"111101101",
        15863=>"100100110",
        15864=>"011011001",
        15865=>"101101100",
        15866=>"001001001",
        15867=>"101101101",
        15868=>"000001100",
        15869=>"000100000",
        15870=>"000000000",
        15871=>"010010000",
        15872=>"000111111",
        15873=>"001000010",
        15874=>"101000000",
        15875=>"000011011",
        15876=>"110110010",
        15877=>"000010011",
        15878=>"000001011",
        15879=>"110101101",
        15880=>"000010001",
        15881=>"110110000",
        15882=>"101000001",
        15883=>"000111011",
        15884=>"010010111",
        15885=>"010111010",
        15886=>"001011001",
        15887=>"000000001",
        15888=>"011111110",
        15889=>"000000000",
        15890=>"110110110",
        15891=>"110011011",
        15892=>"001001101",
        15893=>"000001100",
        15894=>"101000001",
        15895=>"001111111",
        15896=>"001111111",
        15897=>"110111111",
        15898=>"101100100",
        15899=>"000011110",
        15900=>"000000000",
        15901=>"110111011",
        15902=>"101110111",
        15903=>"100110110",
        15904=>"000111011",
        15905=>"110111100",
        15906=>"001111111",
        15907=>"111111110",
        15908=>"111010000",
        15909=>"111111111",
        15910=>"100111010",
        15911=>"010000011",
        15912=>"000000000",
        15913=>"111010110",
        15914=>"000011000",
        15915=>"110100100",
        15916=>"111011001",
        15917=>"010011010",
        15918=>"000110110",
        15919=>"110111111",
        15920=>"110110110",
        15921=>"000110010",
        15922=>"000111110",
        15923=>"100111111",
        15924=>"111011100",
        15925=>"101101111",
        15926=>"110111011",
        15927=>"010000000",
        15928=>"110111000",
        15929=>"011111101",
        15930=>"001011010",
        15931=>"010000000",
        15932=>"100100100",
        15933=>"000000000",
        15934=>"000101111",
        15935=>"100101111",
        15936=>"000000000",
        15937=>"101111111",
        15938=>"110111011",
        15939=>"000010111",
        15940=>"111111110",
        15941=>"010110111",
        15942=>"010000000",
        15943=>"001010111",
        15944=>"010111111",
        15945=>"111101001",
        15946=>"001001000",
        15947=>"111111100",
        15948=>"111111100",
        15949=>"000000000",
        15950=>"010000100",
        15951=>"010111111",
        15952=>"000010000",
        15953=>"000000001",
        15954=>"000000000",
        15955=>"000000000",
        15956=>"010111110",
        15957=>"000000000",
        15958=>"000010001",
        15959=>"001011111",
        15960=>"011110011",
        15961=>"000001000",
        15962=>"001001011",
        15963=>"000000000",
        15964=>"000010011",
        15965=>"010001110",
        15966=>"101111101",
        15967=>"000111000",
        15968=>"100111100",
        15969=>"110010111",
        15970=>"100000000",
        15971=>"111111111",
        15972=>"101000000",
        15973=>"111011110",
        15974=>"000000100",
        15975=>"110111111",
        15976=>"010010011",
        15977=>"111000100",
        15978=>"100000010",
        15979=>"110011011",
        15980=>"111000000",
        15981=>"111000000",
        15982=>"101001000",
        15983=>"001100000",
        15984=>"010000000",
        15985=>"000111000",
        15986=>"000111010",
        15987=>"010000000",
        15988=>"111101111",
        15989=>"000000000",
        15990=>"111111111",
        15991=>"000011011",
        15992=>"000000000",
        15993=>"000010001",
        15994=>"000111110",
        15995=>"000111000",
        15996=>"001100111",
        15997=>"010111011",
        15998=>"101111001",
        15999=>"101011111",
        16000=>"110111111",
        16001=>"000110111",
        16002=>"000110101",
        16003=>"110110000",
        16004=>"001011001",
        16005=>"111111111",
        16006=>"111101101",
        16007=>"000010000",
        16008=>"110001101",
        16009=>"111100001",
        16010=>"001001001",
        16011=>"001010000",
        16012=>"001001111",
        16013=>"110111110",
        16014=>"000000001",
        16015=>"000010110",
        16016=>"011100110",
        16017=>"110111000",
        16018=>"110111101",
        16019=>"100010111",
        16020=>"000010000",
        16021=>"000000000",
        16022=>"110000101",
        16023=>"000000000",
        16024=>"000111011",
        16025=>"001001000",
        16026=>"000101101",
        16027=>"111011000",
        16028=>"111111000",
        16029=>"001100001",
        16030=>"000001000",
        16031=>"111111111",
        16032=>"100000101",
        16033=>"111111111",
        16034=>"000000000",
        16035=>"001000110",
        16036=>"111111100",
        16037=>"000000000",
        16038=>"001111111",
        16039=>"000000000",
        16040=>"111111100",
        16041=>"110110111",
        16042=>"100011011",
        16043=>"011011100",
        16044=>"101110111",
        16045=>"111111000",
        16046=>"111001000",
        16047=>"000000100",
        16048=>"110000101",
        16049=>"000000001",
        16050=>"001000110",
        16051=>"100000001",
        16052=>"100101100",
        16053=>"010000000",
        16054=>"111111010",
        16055=>"000010111",
        16056=>"010010101",
        16057=>"001101111",
        16058=>"111011001",
        16059=>"000000000",
        16060=>"111111111",
        16061=>"000000001",
        16062=>"100100000",
        16063=>"101101010",
        16064=>"111111010",
        16065=>"000000000",
        16066=>"111010000",
        16067=>"111000000",
        16068=>"011001010",
        16069=>"001110111",
        16070=>"000000000",
        16071=>"000000000",
        16072=>"110000111",
        16073=>"000111011",
        16074=>"000100111",
        16075=>"001000000",
        16076=>"110001101",
        16077=>"111111000",
        16078=>"111010110",
        16079=>"000000111",
        16080=>"010010110",
        16081=>"100110000",
        16082=>"101001011",
        16083=>"000100100",
        16084=>"100100110",
        16085=>"110110010",
        16086=>"000110100",
        16087=>"110000011",
        16088=>"111110110",
        16089=>"110100000",
        16090=>"001011111",
        16091=>"110110110",
        16092=>"100100010",
        16093=>"111000010",
        16094=>"001001001",
        16095=>"110111111",
        16096=>"001101011",
        16097=>"011000000",
        16098=>"111111101",
        16099=>"000000000",
        16100=>"111111001",
        16101=>"000000100",
        16102=>"001110111",
        16103=>"000000000",
        16104=>"001010111",
        16105=>"110000100",
        16106=>"100011011",
        16107=>"111001111",
        16108=>"010111111",
        16109=>"000010010",
        16110=>"111011000",
        16111=>"001000000",
        16112=>"110110000",
        16113=>"100110001",
        16114=>"000101111",
        16115=>"110010000",
        16116=>"000111011",
        16117=>"000000010",
        16118=>"000000000",
        16119=>"000000011",
        16120=>"111000000",
        16121=>"111100010",
        16122=>"100100111",
        16123=>"000000000",
        16124=>"000101111",
        16125=>"100010011",
        16126=>"111111001",
        16127=>"111101001",
        16128=>"000110100",
        16129=>"101100100",
        16130=>"001011111",
        16131=>"011011011",
        16132=>"001001011",
        16133=>"011001100",
        16134=>"100100000",
        16135=>"000000110",
        16136=>"110001110",
        16137=>"110010001",
        16138=>"011011000",
        16139=>"101001000",
        16140=>"000110000",
        16141=>"000111110",
        16142=>"111111111",
        16143=>"000001001",
        16144=>"010111011",
        16145=>"001101100",
        16146=>"000000000",
        16147=>"001111100",
        16148=>"011011011",
        16149=>"100100000",
        16150=>"011000000",
        16151=>"001110101",
        16152=>"111111011",
        16153=>"001001011",
        16154=>"000000010",
        16155=>"010010100",
        16156=>"101100000",
        16157=>"101001101",
        16158=>"001011111",
        16159=>"011111000",
        16160=>"000111101",
        16161=>"111111100",
        16162=>"001001000",
        16163=>"000000000",
        16164=>"100110000",
        16165=>"100001000",
        16166=>"011001011",
        16167=>"000001011",
        16168=>"011100100",
        16169=>"100100000",
        16170=>"011000000",
        16171=>"011100000",
        16172=>"100100000",
        16173=>"000100100",
        16174=>"110110100",
        16175=>"011011011",
        16176=>"010010110",
        16177=>"011001011",
        16178=>"011001101",
        16179=>"100110110",
        16180=>"101101001",
        16181=>"100100100",
        16182=>"110110100",
        16183=>"001101001",
        16184=>"100100000",
        16185=>"001011001",
        16186=>"100111111",
        16187=>"100011011",
        16188=>"000110110",
        16189=>"111010011",
        16190=>"101101000",
        16191=>"011110100",
        16192=>"011011010",
        16193=>"100011111",
        16194=>"110100110",
        16195=>"100100000",
        16196=>"111111111",
        16197=>"110111111",
        16198=>"010100000",
        16199=>"100001000",
        16200=>"111111111",
        16201=>"100010000",
        16202=>"110110110",
        16203=>"100100000",
        16204=>"100110000",
        16205=>"001011001",
        16206=>"100100110",
        16207=>"001001011",
        16208=>"010111101",
        16209=>"100000100",
        16210=>"001001111",
        16211=>"111001011",
        16212=>"000000001",
        16213=>"000001011",
        16214=>"000010000",
        16215=>"011001000",
        16216=>"111110100",
        16217=>"100010110",
        16218=>"000000000",
        16219=>"100100000",
        16220=>"110110110",
        16221=>"010001110",
        16222=>"011011001",
        16223=>"000101101",
        16224=>"011011111",
        16225=>"001000100",
        16226=>"001011011",
        16227=>"110100100",
        16228=>"001011000",
        16229=>"000010100",
        16230=>"000000010",
        16231=>"010000110",
        16232=>"100100000",
        16233=>"110011110",
        16234=>"000110100",
        16235=>"110001001",
        16236=>"000011011",
        16237=>"100000001",
        16238=>"000100100",
        16239=>"110000000",
        16240=>"011011010",
        16241=>"000101101",
        16242=>"111110011",
        16243=>"001011001",
        16244=>"011001011",
        16245=>"001000000",
        16246=>"111100100",
        16247=>"001011010",
        16248=>"001100100",
        16249=>"110100110",
        16250=>"100110000",
        16251=>"110100110",
        16252=>"001111011",
        16253=>"000111101",
        16254=>"000100101",
        16255=>"001111111",
        16256=>"110111111",
        16257=>"000000111",
        16258=>"111101101",
        16259=>"010010010",
        16260=>"000110010",
        16261=>"000000000",
        16262=>"111111111",
        16263=>"111111111",
        16264=>"111100011",
        16265=>"010011111",
        16266=>"001000000",
        16267=>"011100111",
        16268=>"000001000",
        16269=>"010111010",
        16270=>"111110000",
        16271=>"100000001",
        16272=>"000000000",
        16273=>"010111010",
        16274=>"000010000",
        16275=>"010011011",
        16276=>"000000100",
        16277=>"010000001",
        16278=>"000000000",
        16279=>"100000110",
        16280=>"000011101",
        16281=>"100001011",
        16282=>"111111111",
        16283=>"000000000",
        16284=>"000010110",
        16285=>"101111001",
        16286=>"101111111",
        16287=>"101111110",
        16288=>"111111111",
        16289=>"000000000",
        16290=>"111111110",
        16291=>"000010110",
        16292=>"010010111",
        16293=>"110110100",
        16294=>"111111110",
        16295=>"000111001",
        16296=>"000000001",
        16297=>"100000101",
        16298=>"111111000",
        16299=>"010111001",
        16300=>"110111111",
        16301=>"111111111",
        16302=>"100111110",
        16303=>"111111111",
        16304=>"111000000",
        16305=>"000000000",
        16306=>"000101100",
        16307=>"000001011",
        16308=>"111011010",
        16309=>"000000001",
        16310=>"100000010",
        16311=>"111100110",
        16312=>"011000000",
        16313=>"111111111",
        16314=>"011110110",
        16315=>"000011000",
        16316=>"110111010",
        16317=>"000111000",
        16318=>"000110000",
        16319=>"111000111",
        16320=>"010010111",
        16321=>"000101111",
        16322=>"111111000",
        16323=>"000010000",
        16324=>"001011010",
        16325=>"111111111",
        16326=>"011111001",
        16327=>"111111111",
        16328=>"100000000",
        16329=>"000000000",
        16330=>"000000111",
        16331=>"111111010",
        16332=>"111111111",
        16333=>"001000001",
        16334=>"110111011",
        16335=>"101000000",
        16336=>"000000100",
        16337=>"111111011",
        16338=>"000000101",
        16339=>"110111111",
        16340=>"111111111",
        16341=>"111101100",
        16342=>"000011000",
        16343=>"111111111",
        16344=>"101101100",
        16345=>"000111111",
        16346=>"001001010",
        16347=>"001000000",
        16348=>"100111000",
        16349=>"011110000",
        16350=>"111011010",
        16351=>"000011000",
        16352=>"100000010",
        16353=>"000000000",
        16354=>"000000000",
        16355=>"111110000",
        16356=>"000110010",
        16357=>"000011010",
        16358=>"111110110",
        16359=>"100111111",
        16360=>"010010110",
        16361=>"101000000",
        16362=>"100111100",
        16363=>"110111110",
        16364=>"001000000",
        16365=>"111000000",
        16366=>"000000000",
        16367=>"111111100",
        16368=>"000010110",
        16369=>"000101001",
        16370=>"000000001",
        16371=>"010111000",
        16372=>"000000101",
        16373=>"000000000",
        16374=>"111111111",
        16375=>"000111011",
        16376=>"111100110",
        16377=>"111010010",
        16378=>"010010000",
        16379=>"000000110",
        16380=>"110111011",
        16381=>"111110111",
        16382=>"000000011",
        16383=>"100111010");
        BEGIN
        weight <= ROM_content(to_integer(address));
    END RTL;