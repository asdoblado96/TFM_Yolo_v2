LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L8_14_BNROM IS
  PORT (
    coefs : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    address : IN unsigned(5 DOWNTO 0));
END L8_14_BNROM;

ARCHITECTURE RTL OF L8_14_BNROM IS

  TYPE ROM_mem IS ARRAY (0 TO 63) OF STD_LOGIC_VECTOR(31 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem :=

  --Contenido bias || scale
  (0=>"0001101001010001"&"0010010101101101",
  1=>"0001001001001001"&"0010010001111010",
  2=>"0001000001010101"&"0001111110110010",
  3=>"0001101101110110"&"0010011011110110",
  4=>"0001000111100110"&"0010010111101100",
  5=>"0000110000100011"&"0001111010011010",
  6=>"0000110100011111"&"0010010001101010",
  7=>"1111101100101101"&"0010010001000001",
  8=>"0000101101101000"&"0010010101101100",
  9=>"1111110101000010"&"0001101100010100",
  10=>"0001100001011101"&"0010001000000000",
  11=>"0010011010100010"&"0010010100011001",
  12=>"0010010100010100"&"0001101110101011",
  13=>"0010011100111011"&"0010000100101010",
  14=>"0010010111001001"&"0010010101111011",
  15=>"0001010101001010"&"0010010100110111",
  16=>"0010010011111010"&"0010001100000001",
  17=>"0001011001111100"&"0001111001000011",
  18=>"0010100010110001"&"0010010000101101",
  19=>"0000101110110110"&"0010010010110101",
  20=>"0001001111001100"&"0001111010110101",
  21=>"0000111110101111"&"0001110100001111",
  22=>"1111101101101001"&"0001101100101000",
  23=>"0001101100110000"&"0010011101111001",
  24=>"0001001110110110"&"0010011111100001",
  25=>"0001101110101111"&"0010000010011010",
  26=>"0010011010110011"&"0001110111111100",
  27=>"0001100011010111"&"0010010110110011",
  28=>"0001111011110100"&"0001111010001010",
  29=>"0001010101100010"&"0010011010011010",
  30=>"0000110000101101"&"0010010001001111",
  31=>"0000111101110001"&"0010011101011101",
  32=>"0001011001111111"&"0010011010011100",
  33=>"0000011111011110"&"0010010011010101",
  34=>"0000111111001001"&"0010011011101000",
  35=>"0000011011101100"&"0010000000011001",
  36=>"0010010100111011"&"0010000001110100",
  37=>"0000101100101011"&"0001110010000110",
  38=>"0000111000111100"&"0010001110011101",
  39=>"0001101011110101"&"0010001100110001",
  40=>"0000111000011110"&"0010010000111001",
  41=>"0010001001111101"&"0010010101011000",
  42=>"0010000111000010"&"0001111100010110",
  43=>"0000100111011010"&"0010010010110110",
  44=>"0010000000001010"&"0001110100110000",
  45=>"0000001111110101"&"0010000000100100",
  46=>"0001011110010011"&"0010010111011011",
  47=>"1111100110010101"&"0010010100001011",
  48=>"0000111011111110"&"0010001000100010",
  49=>"0001001100111100"&"0010011000110000",
  50=>"0001100100111110"&"0001110000110101",
  51=>"0000010011101011"&"0010011011110011",
  52=>"0001110110101010"&"0001111001000110",
  53=>"0000100100100101"&"0010011101100100",
  54=>"0001101101001100"&"0010010001011010",
  55=>"0001101111010110"&"0010000110100010",
  56=>"1110111101101101"&"0010000110100010",
  57=>"0010011010100011"&"0010001111010000",
  58=>"0001111111101010"&"0010001111101100",
  59=>"0001011100110100"&"0001111111001000",
  60=>"0000110110100001"&"0010011011010111",
  61=>"0001101001101100"&"0010001111000111",
  62=>"0000110000010111"&"0010100100001001",
  63=>"0000100101000011"&"0010000101101011");

BEGIN
  coefs <= ROM_content(to_integer(address));
END RTL;