LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L8_9_WROM IS
  PORT (
    weight : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
    address : IN unsigned(weightsbitsAddress(8)-1 DOWNTO 0));
END L8_9_WROM;

ARCHITECTURE RTL OF L8_9_WROM IS

  TYPE ROM_mem IS ARRAY (0 TO 65535) OF STD_LOGIC_VECTOR(8 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem := (0=>"101100100",
  1=>"001001101",
  2=>"101110100",
  3=>"110111010",
  4=>"010110011",
  5=>"010100111",
  6=>"110000100",
  7=>"010011000",
  8=>"110100101",
  9=>"010010001",
  10=>"111001011",
  11=>"100011010",
  12=>"010010011",
  13=>"100100010",
  14=>"011110111",
  15=>"101110111",
  16=>"101100111",
  17=>"100001010",
  18=>"000010111",
  19=>"101101110",
  20=>"001100010",
  21=>"100001110",
  22=>"111110000",
  23=>"001101100",
  24=>"100000111",
  25=>"100011000",
  26=>"000100101",
  27=>"011101101",
  28=>"110110110",
  29=>"011101100",
  30=>"011000011",
  31=>"001001011",
  32=>"111101010",
  33=>"000110010",
  34=>"010111110",
  35=>"000011010",
  36=>"101110000",
  37=>"100011011",
  38=>"011011101",
  39=>"000100001",
  40=>"001100100",
  41=>"010011101",
  42=>"111000111",
  43=>"101110101",
  44=>"101010000",
  45=>"110000010",
  46=>"101011011",
  47=>"100011101",
  48=>"001110101",
  49=>"110100111",
  50=>"111110110",
  51=>"010110000",
  52=>"101010011",
  53=>"011010101",
  54=>"010001111",
  55=>"001111011",
  56=>"011000100",
  57=>"000100010",
  58=>"000000001",
  59=>"001100100",
  60=>"010000100",
  61=>"001011010",
  62=>"001001111",
  63=>"000110100",
  64=>"110011101",
  65=>"111001101",
  66=>"111010101",
  67=>"100000001",
  68=>"010101001",
  69=>"100011101",
  70=>"011111011",
  71=>"001001010",
  72=>"011010001",
  73=>"001001000",
  74=>"000100100",
  75=>"111111101",
  76=>"101100000",
  77=>"011001100",
  78=>"111110110",
  79=>"001001110",
  80=>"001001111",
  81=>"101101110",
  82=>"100011111",
  83=>"110111000",
  84=>"000111011",
  85=>"000001111",
  86=>"111101000",
  87=>"001011101",
  88=>"011111000",
  89=>"011110001",
  90=>"111010101",
  91=>"101000000",
  92=>"110110101",
  93=>"011100011",
  94=>"010100111",
  95=>"011011110",
  96=>"001101000",
  97=>"001000100",
  98=>"100100111",
  99=>"000000011",
  100=>"010000111",
  101=>"000100110",
  102=>"000111000",
  103=>"110011010",
  104=>"111010100",
  105=>"110011000",
  106=>"000110101",
  107=>"101111100",
  108=>"100011000",
  109=>"110011101",
  110=>"111101000",
  111=>"111011011",
  112=>"111011100",
  113=>"011011100",
  114=>"000001000",
  115=>"011101101",
  116=>"011101010",
  117=>"100111001",
  118=>"101000001",
  119=>"010110111",
  120=>"010111111",
  121=>"111010001",
  122=>"101001101",
  123=>"110000111",
  124=>"111001011",
  125=>"001010001",
  126=>"011110001",
  127=>"011001011",
  128=>"111001001",
  129=>"011011100",
  130=>"110010101",
  131=>"000001001",
  132=>"010101000",
  133=>"001110110",
  134=>"110001010",
  135=>"001001010",
  136=>"100001100",
  137=>"100100011",
  138=>"011001001",
  139=>"000000001",
  140=>"110010001",
  141=>"111011101",
  142=>"010110011",
  143=>"001110101",
  144=>"010100100",
  145=>"111110011",
  146=>"111001111",
  147=>"010000110",
  148=>"100111011",
  149=>"000010100",
  150=>"010101000",
  151=>"011011011",
  152=>"011001101",
  153=>"111111101",
  154=>"100101001",
  155=>"110011111",
  156=>"000011011",
  157=>"110110100",
  158=>"101010010",
  159=>"010011100",
  160=>"000001001",
  161=>"111011100",
  162=>"110101100",
  163=>"010001100",
  164=>"110100101",
  165=>"100011100",
  166=>"000000111",
  167=>"100111111",
  168=>"110110111",
  169=>"110010101",
  170=>"100011111",
  171=>"001000001",
  172=>"011011110",
  173=>"100000110",
  174=>"100111010",
  175=>"110000000",
  176=>"111110001",
  177=>"100011110",
  178=>"011101111",
  179=>"000010010",
  180=>"000001000",
  181=>"000011000",
  182=>"101100101",
  183=>"101010010",
  184=>"001111111",
  185=>"100110111",
  186=>"101100100",
  187=>"110110011",
  188=>"011011011",
  189=>"001101100",
  190=>"111001001",
  191=>"010000011",
  192=>"010000111",
  193=>"101000101",
  194=>"110001100",
  195=>"111011101",
  196=>"000110011",
  197=>"110001110",
  198=>"101101111",
  199=>"001101000",
  200=>"000000011",
  201=>"000011110",
  202=>"001100001",
  203=>"111011000",
  204=>"101011101",
  205=>"100101101",
  206=>"100101001",
  207=>"001000101",
  208=>"110010001",
  209=>"111111001",
  210=>"100001001",
  211=>"000011010",
  212=>"101001100",
  213=>"101101110",
  214=>"111010001",
  215=>"011110001",
  216=>"101010110",
  217=>"011101100",
  218=>"111010010",
  219=>"000010100",
  220=>"010111000",
  221=>"001110000",
  222=>"111101101",
  223=>"100001010",
  224=>"001001100",
  225=>"001010000",
  226=>"010010001",
  227=>"011101011",
  228=>"110010110",
  229=>"000100110",
  230=>"010011110",
  231=>"011010011",
  232=>"011111111",
  233=>"100011010",
  234=>"100101111",
  235=>"111101011",
  236=>"101100101",
  237=>"011110111",
  238=>"001000111",
  239=>"010111100",
  240=>"111101110",
  241=>"101111011",
  242=>"010000111",
  243=>"110110110",
  244=>"000100001",
  245=>"101110000",
  246=>"110101100",
  247=>"110000010",
  248=>"101001110",
  249=>"000110101",
  250=>"110010000",
  251=>"100010100",
  252=>"100100011",
  253=>"010010010",
  254=>"000010100",
  255=>"010100001",
  256=>"101101100",
  257=>"110111111",
  258=>"000110011",
  259=>"111001010",
  260=>"111011111",
  261=>"001110011",
  262=>"111000111",
  263=>"110010101",
  264=>"110001011",
  265=>"010011111",
  266=>"110000111",
  267=>"101101101",
  268=>"101010011",
  269=>"001000011",
  270=>"010011001",
  271=>"001110001",
  272=>"111100101",
  273=>"110100111",
  274=>"010010010",
  275=>"001001111",
  276=>"000101010",
  277=>"011000100",
  278=>"000100000",
  279=>"000001101",
  280=>"001011001",
  281=>"111000011",
  282=>"100000111",
  283=>"000011001",
  284=>"111101111",
  285=>"101001110",
  286=>"110110100",
  287=>"000101110",
  288=>"000001100",
  289=>"110011011",
  290=>"001010111",
  291=>"100011100",
  292=>"101011010",
  293=>"011100111",
  294=>"100001101",
  295=>"101110011",
  296=>"111001111",
  297=>"011010100",
  298=>"111011000",
  299=>"011011010",
  300=>"100101010",
  301=>"001100000",
  302=>"111000001",
  303=>"000001010",
  304=>"101010101",
  305=>"010111001",
  306=>"000001001",
  307=>"011010011",
  308=>"111010010",
  309=>"010110001",
  310=>"100101110",
  311=>"101111000",
  312=>"000101101",
  313=>"111110001",
  314=>"000010010",
  315=>"110000011",
  316=>"110111000",
  317=>"011111101",
  318=>"010000010",
  319=>"100011100",
  320=>"001100100",
  321=>"011000000",
  322=>"000110001",
  323=>"110001100",
  324=>"000110010",
  325=>"001110100",
  326=>"100100011",
  327=>"111000010",
  328=>"110001110",
  329=>"100010000",
  330=>"100000000",
  331=>"010111111",
  332=>"011011111",
  333=>"000111011",
  334=>"010101110",
  335=>"100101110",
  336=>"101001001",
  337=>"100111101",
  338=>"100111101",
  339=>"000011000",
  340=>"000100011",
  341=>"010010100",
  342=>"010011000",
  343=>"000011001",
  344=>"111110111",
  345=>"011010110",
  346=>"001110011",
  347=>"101100011",
  348=>"111011000",
  349=>"110001110",
  350=>"000000111",
  351=>"100111110",
  352=>"000110110",
  353=>"110110010",
  354=>"111111000",
  355=>"100000010",
  356=>"111110110",
  357=>"000111010",
  358=>"110110011",
  359=>"101011000",
  360=>"001110110",
  361=>"011001100",
  362=>"000010101",
  363=>"000101000",
  364=>"011101111",
  365=>"001110101",
  366=>"111110001",
  367=>"111001011",
  368=>"101100101",
  369=>"110110111",
  370=>"110001010",
  371=>"011110011",
  372=>"001101100",
  373=>"111000010",
  374=>"000000001",
  375=>"011101111",
  376=>"001011000",
  377=>"010110011",
  378=>"011000100",
  379=>"110010000",
  380=>"001010011",
  381=>"110000100",
  382=>"000111101",
  383=>"001100011",
  384=>"000010001",
  385=>"110100010",
  386=>"010111110",
  387=>"111101001",
  388=>"111111101",
  389=>"111110011",
  390=>"100100111",
  391=>"100011000",
  392=>"111110010",
  393=>"011000100",
  394=>"100001010",
  395=>"111111110",
  396=>"111100100",
  397=>"110011001",
  398=>"010010010",
  399=>"101110111",
  400=>"000010101",
  401=>"010011001",
  402=>"000000100",
  403=>"111010010",
  404=>"000011001",
  405=>"011110000",
  406=>"010100101",
  407=>"111100000",
  408=>"010111001",
  409=>"111101010",
  410=>"010000000",
  411=>"111111100",
  412=>"111101001",
  413=>"100110001",
  414=>"110011001",
  415=>"100111000",
  416=>"100001101",
  417=>"111111100",
  418=>"101101111",
  419=>"111111111",
  420=>"000101101",
  421=>"100010100",
  422=>"100010011",
  423=>"100111111",
  424=>"100000000",
  425=>"000100110",
  426=>"001101011",
  427=>"100101101",
  428=>"010011111",
  429=>"001011101",
  430=>"110011101",
  431=>"010011001",
  432=>"110111010",
  433=>"010000011",
  434=>"000010110",
  435=>"010011010",
  436=>"100101000",
  437=>"110001000",
  438=>"111101101",
  439=>"110000010",
  440=>"001111101",
  441=>"010100011",
  442=>"010111101",
  443=>"111001111",
  444=>"011010101",
  445=>"111111100",
  446=>"010000100",
  447=>"111111100",
  448=>"010011001",
  449=>"100100011",
  450=>"110111101",
  451=>"011100110",
  452=>"010010011",
  453=>"010000101",
  454=>"011111000",
  455=>"110100011",
  456=>"100010111",
  457=>"001101011",
  458=>"001001100",
  459=>"000100011",
  460=>"111011001",
  461=>"111100000",
  462=>"001101100",
  463=>"001110001",
  464=>"101101111",
  465=>"101010100",
  466=>"101101001",
  467=>"011010100",
  468=>"000011110",
  469=>"011111010",
  470=>"110000001",
  471=>"000110000",
  472=>"111110000",
  473=>"001001100",
  474=>"010001110",
  475=>"011000001",
  476=>"010110010",
  477=>"101011100",
  478=>"010010001",
  479=>"000010111",
  480=>"110011011",
  481=>"111001011",
  482=>"111100110",
  483=>"101100000",
  484=>"100101101",
  485=>"010100100",
  486=>"101010110",
  487=>"010011001",
  488=>"010011110",
  489=>"110000000",
  490=>"001001111",
  491=>"111101101",
  492=>"100011000",
  493=>"111011001",
  494=>"100010010",
  495=>"101001001",
  496=>"011000110",
  497=>"111001101",
  498=>"100101001",
  499=>"100001010",
  500=>"111000110",
  501=>"101110110",
  502=>"000011000",
  503=>"010011100",
  504=>"101111101",
  505=>"100110100",
  506=>"011111001",
  507=>"011011011",
  508=>"000110000",
  509=>"101011011",
  510=>"111011000",
  511=>"101100101",
  512=>"010101000",
  513=>"101000010",
  514=>"100001011",
  515=>"001100011",
  516=>"100111100",
  517=>"011000110",
  518=>"011010010",
  519=>"100010010",
  520=>"100110101",
  521=>"100010110",
  522=>"111001101",
  523=>"110100011",
  524=>"010100001",
  525=>"001000011",
  526=>"001110000",
  527=>"011000001",
  528=>"100010111",
  529=>"100000000",
  530=>"111000111",
  531=>"111011010",
  532=>"110010100",
  533=>"001010110",
  534=>"010100001",
  535=>"111000010",
  536=>"000101010",
  537=>"000011001",
  538=>"000101101",
  539=>"011011100",
  540=>"011100001",
  541=>"000000001",
  542=>"000001110",
  543=>"101101101",
  544=>"001100010",
  545=>"111100100",
  546=>"011101000",
  547=>"101101000",
  548=>"001111101",
  549=>"111001110",
  550=>"101101011",
  551=>"101000001",
  552=>"100000000",
  553=>"001010110",
  554=>"010110100",
  555=>"101110100",
  556=>"011111010",
  557=>"000111111",
  558=>"101000001",
  559=>"000101110",
  560=>"111100000",
  561=>"101100111",
  562=>"111101110",
  563=>"011001100",
  564=>"001001011",
  565=>"100000010",
  566=>"010011000",
  567=>"000100011",
  568=>"111110011",
  569=>"001110100",
  570=>"110110111",
  571=>"110010111",
  572=>"000111000",
  573=>"100101101",
  574=>"000110111",
  575=>"110010101",
  576=>"000110011",
  577=>"011111001",
  578=>"000000101",
  579=>"100110110",
  580=>"101100000",
  581=>"000111001",
  582=>"000001010",
  583=>"110000101",
  584=>"001010110",
  585=>"011000000",
  586=>"100001000",
  587=>"100110000",
  588=>"011001011",
  589=>"011100111",
  590=>"110111101",
  591=>"111111000",
  592=>"101010000",
  593=>"000111010",
  594=>"000110001",
  595=>"101110010",
  596=>"111111111",
  597=>"110111111",
  598=>"100110100",
  599=>"001000000",
  600=>"001111001",
  601=>"101001000",
  602=>"111100001",
  603=>"110111111",
  604=>"100111100",
  605=>"100010000",
  606=>"111010100",
  607=>"000010000",
  608=>"001001000",
  609=>"001010000",
  610=>"001111111",
  611=>"100101001",
  612=>"111010100",
  613=>"000111000",
  614=>"000010010",
  615=>"100010010",
  616=>"111100110",
  617=>"001001101",
  618=>"110011100",
  619=>"100001101",
  620=>"011001100",
  621=>"101001100",
  622=>"101111100",
  623=>"110110000",
  624=>"011011000",
  625=>"100000100",
  626=>"100110010",
  627=>"110100111",
  628=>"110110101",
  629=>"011010110",
  630=>"001011111",
  631=>"100110010",
  632=>"000110101",
  633=>"111011100",
  634=>"101110111",
  635=>"011000111",
  636=>"111001101",
  637=>"000110111",
  638=>"101111011",
  639=>"001110101",
  640=>"000000000",
  641=>"011000011",
  642=>"111101010",
  643=>"111001100",
  644=>"000111111",
  645=>"001100101",
  646=>"011110000",
  647=>"111001001",
  648=>"010110111",
  649=>"001101000",
  650=>"000100000",
  651=>"010110010",
  652=>"010110101",
  653=>"111110011",
  654=>"010110111",
  655=>"011010010",
  656=>"110110011",
  657=>"111110110",
  658=>"100111101",
  659=>"011010101",
  660=>"111110010",
  661=>"111011011",
  662=>"101111010",
  663=>"011010101",
  664=>"011110010",
  665=>"011110101",
  666=>"011100000",
  667=>"111010101",
  668=>"000000101",
  669=>"100110100",
  670=>"011000100",
  671=>"000001100",
  672=>"100110011",
  673=>"000101000",
  674=>"101101100",
  675=>"110110000",
  676=>"111110100",
  677=>"111011100",
  678=>"101110010",
  679=>"011100101",
  680=>"000000001",
  681=>"010000100",
  682=>"001011010",
  683=>"000001011",
  684=>"101000001",
  685=>"110000010",
  686=>"110010110",
  687=>"000000101",
  688=>"001000000",
  689=>"100101001",
  690=>"001101000",
  691=>"100111011",
  692=>"100001110",
  693=>"001101101",
  694=>"110111000",
  695=>"010010010",
  696=>"000000100",
  697=>"011011100",
  698=>"001000001",
  699=>"111001000",
  700=>"001111110",
  701=>"010011000",
  702=>"001001001",
  703=>"001000101",
  704=>"111110000",
  705=>"000001111",
  706=>"011110100",
  707=>"100110010",
  708=>"111110000",
  709=>"101110010",
  710=>"100000110",
  711=>"101001101",
  712=>"101100101",
  713=>"010001100",
  714=>"110010110",
  715=>"011101000",
  716=>"110100100",
  717=>"111010000",
  718=>"110011111",
  719=>"100110000",
  720=>"000100000",
  721=>"111100100",
  722=>"010010010",
  723=>"101101000",
  724=>"000110010",
  725=>"000110110",
  726=>"001001100",
  727=>"110010000",
  728=>"110100000",
  729=>"100101001",
  730=>"101001000",
  731=>"101011000",
  732=>"101001001",
  733=>"111010011",
  734=>"100100101",
  735=>"011111111",
  736=>"010101111",
  737=>"111001001",
  738=>"110010001",
  739=>"110000011",
  740=>"000111100",
  741=>"010000001",
  742=>"011001001",
  743=>"100011001",
  744=>"011001001",
  745=>"011011100",
  746=>"111100011",
  747=>"110000000",
  748=>"001100000",
  749=>"000111000",
  750=>"001111001",
  751=>"001100010",
  752=>"010000110",
  753=>"110101000",
  754=>"101010011",
  755=>"010100010",
  756=>"110010010",
  757=>"001010001",
  758=>"010100010",
  759=>"000100000",
  760=>"100000110",
  761=>"111010110",
  762=>"010011001",
  763=>"110000000",
  764=>"100101010",
  765=>"010110101",
  766=>"011101000",
  767=>"110001001",
  768=>"101010001",
  769=>"000101101",
  770=>"011101111",
  771=>"110100000",
  772=>"111111110",
  773=>"001010101",
  774=>"000010010",
  775=>"101111001",
  776=>"010101001",
  777=>"101101001",
  778=>"011101010",
  779=>"101000110",
  780=>"011111000",
  781=>"001110101",
  782=>"010001111",
  783=>"111011100",
  784=>"100010111",
  785=>"001100001",
  786=>"111110011",
  787=>"111011110",
  788=>"111010010",
  789=>"011111100",
  790=>"100010011",
  791=>"111000010",
  792=>"011000101",
  793=>"011101101",
  794=>"111000011",
  795=>"010010100",
  796=>"001110111",
  797=>"100000011",
  798=>"000100010",
  799=>"011100111",
  800=>"111101110",
  801=>"110110011",
  802=>"011100000",
  803=>"010011100",
  804=>"111110101",
  805=>"001110001",
  806=>"111101010",
  807=>"000010011",
  808=>"001100001",
  809=>"000010010",
  810=>"100000110",
  811=>"111110111",
  812=>"101010110",
  813=>"101001000",
  814=>"111111101",
  815=>"000110101",
  816=>"101101111",
  817=>"110100101",
  818=>"000001000",
  819=>"101110010",
  820=>"011001000",
  821=>"011011111",
  822=>"111011001",
  823=>"000100110",
  824=>"010010010",
  825=>"000001000",
  826=>"010101000",
  827=>"011010101",
  828=>"101000000",
  829=>"001101101",
  830=>"001100010",
  831=>"011010011",
  832=>"001110001",
  833=>"101111011",
  834=>"111010011",
  835=>"001110001",
  836=>"110011110",
  837=>"100010100",
  838=>"000101000",
  839=>"111111110",
  840=>"011001111",
  841=>"110010001",
  842=>"010010001",
  843=>"010100110",
  844=>"100011010",
  845=>"101101000",
  846=>"001111111",
  847=>"000110001",
  848=>"111000100",
  849=>"101010100",
  850=>"011100000",
  851=>"000001100",
  852=>"001111010",
  853=>"111101110",
  854=>"000011011",
  855=>"001010101",
  856=>"111011100",
  857=>"100001101",
  858=>"011011001",
  859=>"001011111",
  860=>"010100010",
  861=>"111110001",
  862=>"000100001",
  863=>"001011101",
  864=>"100011101",
  865=>"101111100",
  866=>"101110001",
  867=>"010111011",
  868=>"011000111",
  869=>"111001011",
  870=>"110110111",
  871=>"011100100",
  872=>"100001101",
  873=>"111100110",
  874=>"101111011",
  875=>"000101101",
  876=>"100011010",
  877=>"001100010",
  878=>"000000101",
  879=>"011100110",
  880=>"101110110",
  881=>"100011001",
  882=>"111101010",
  883=>"110100000",
  884=>"011110011",
  885=>"100001011",
  886=>"001101100",
  887=>"111010111",
  888=>"001110011",
  889=>"010001110",
  890=>"010111011",
  891=>"011011000",
  892=>"001011110",
  893=>"110111100",
  894=>"000111010",
  895=>"111000111",
  896=>"100111101",
  897=>"110011010",
  898=>"100100100",
  899=>"111111100",
  900=>"100010001",
  901=>"100001001",
  902=>"011111110",
  903=>"011101001",
  904=>"011000000",
  905=>"000111010",
  906=>"011001111",
  907=>"110011000",
  908=>"001000000",
  909=>"011011011",
  910=>"110100111",
  911=>"100101011",
  912=>"000001010",
  913=>"100001110",
  914=>"000100100",
  915=>"000010000",
  916=>"100010001",
  917=>"111010001",
  918=>"011110100",
  919=>"000001101",
  920=>"111011110",
  921=>"011000110",
  922=>"011101010",
  923=>"100010001",
  924=>"000110010",
  925=>"111111111",
  926=>"010000110",
  927=>"001101010",
  928=>"010101001",
  929=>"010101100",
  930=>"011010100",
  931=>"111001011",
  932=>"100000000",
  933=>"001100111",
  934=>"110100100",
  935=>"010010001",
  936=>"010000011",
  937=>"110101100",
  938=>"011011000",
  939=>"110111100",
  940=>"001101111",
  941=>"111111011",
  942=>"001000011",
  943=>"010011001",
  944=>"110100101",
  945=>"101001001",
  946=>"011010101",
  947=>"011011100",
  948=>"101011001",
  949=>"101110010",
  950=>"010111101",
  951=>"011010101",
  952=>"001000011",
  953=>"000000101",
  954=>"110000101",
  955=>"100010001",
  956=>"000100000",
  957=>"000000111",
  958=>"101010100",
  959=>"000010101",
  960=>"010000110",
  961=>"001111100",
  962=>"101101011",
  963=>"000010001",
  964=>"000101100",
  965=>"101011111",
  966=>"101100111",
  967=>"010100011",
  968=>"111001111",
  969=>"001001110",
  970=>"110110110",
  971=>"110001011",
  972=>"100111000",
  973=>"110000001",
  974=>"101101111",
  975=>"010011100",
  976=>"000110111",
  977=>"100110001",
  978=>"100111001",
  979=>"111000000",
  980=>"101101000",
  981=>"111011000",
  982=>"000100000",
  983=>"000010111",
  984=>"110101100",
  985=>"000111000",
  986=>"010001000",
  987=>"000001001",
  988=>"111110111",
  989=>"110100010",
  990=>"100000000",
  991=>"111100010",
  992=>"111101011",
  993=>"010111110",
  994=>"011010111",
  995=>"000010110",
  996=>"010000011",
  997=>"001010000",
  998=>"101001001",
  999=>"100110111",
  1000=>"000111001",
  1001=>"111001101",
  1002=>"110000001",
  1003=>"101101101",
  1004=>"101100000",
  1005=>"001011011",
  1006=>"101101010",
  1007=>"010111100",
  1008=>"101011001",
  1009=>"110001000",
  1010=>"001011010",
  1011=>"001001111",
  1012=>"011000111",
  1013=>"100111110",
  1014=>"001101000",
  1015=>"111101000",
  1016=>"100111110",
  1017=>"001111001",
  1018=>"000101010",
  1019=>"001001101",
  1020=>"000011100",
  1021=>"111110100",
  1022=>"110011000",
  1023=>"010101000",
  1024=>"100001011",
  1025=>"010101011",
  1026=>"110100100",
  1027=>"001000110",
  1028=>"111000111",
  1029=>"110110111",
  1030=>"101001010",
  1031=>"001011001",
  1032=>"100010111",
  1033=>"000100000",
  1034=>"111011111",
  1035=>"000110000",
  1036=>"001100010",
  1037=>"110111111",
  1038=>"010001010",
  1039=>"001101100",
  1040=>"101001001",
  1041=>"011100001",
  1042=>"101000111",
  1043=>"101101100",
  1044=>"111000110",
  1045=>"001101101",
  1046=>"001110110",
  1047=>"101111011",
  1048=>"010011000",
  1049=>"000011011",
  1050=>"000011000",
  1051=>"110000110",
  1052=>"101110011",
  1053=>"101001110",
  1054=>"011111111",
  1055=>"000011100",
  1056=>"100000011",
  1057=>"100010001",
  1058=>"000001001",
  1059=>"100111010",
  1060=>"101000101",
  1061=>"111000101",
  1062=>"010100000",
  1063=>"111110111",
  1064=>"110011011",
  1065=>"010110110",
  1066=>"011011000",
  1067=>"010101101",
  1068=>"110011011",
  1069=>"111011001",
  1070=>"011011010",
  1071=>"011100011",
  1072=>"101100100",
  1073=>"111010000",
  1074=>"100111000",
  1075=>"000000100",
  1076=>"010001001",
  1077=>"101100101",
  1078=>"111111000",
  1079=>"000111000",
  1080=>"101110101",
  1081=>"101010110",
  1082=>"100101100",
  1083=>"100000110",
  1084=>"000010010",
  1085=>"001000101",
  1086=>"011011001",
  1087=>"111101110",
  1088=>"010101111",
  1089=>"001101101",
  1090=>"111001011",
  1091=>"100010001",
  1092=>"001110100",
  1093=>"100001010",
  1094=>"011110010",
  1095=>"101001000",
  1096=>"101111100",
  1097=>"100100001",
  1098=>"011110010",
  1099=>"001111101",
  1100=>"110010000",
  1101=>"100101010",
  1102=>"101111000",
  1103=>"100010101",
  1104=>"010101100",
  1105=>"111010011",
  1106=>"110010000",
  1107=>"100100011",
  1108=>"110101100",
  1109=>"010110110",
  1110=>"000010100",
  1111=>"000111001",
  1112=>"100011001",
  1113=>"100100100",
  1114=>"100000011",
  1115=>"111101001",
  1116=>"101001110",
  1117=>"000001010",
  1118=>"001110110",
  1119=>"111000001",
  1120=>"000001111",
  1121=>"111110110",
  1122=>"010011000",
  1123=>"101101001",
  1124=>"001111011",
  1125=>"100100111",
  1126=>"101000101",
  1127=>"011000011",
  1128=>"101010111",
  1129=>"111001000",
  1130=>"001100110",
  1131=>"010001110",
  1132=>"000111100",
  1133=>"111101001",
  1134=>"101000100",
  1135=>"000101001",
  1136=>"011001110",
  1137=>"000111011",
  1138=>"001111010",
  1139=>"000001011",
  1140=>"111101011",
  1141=>"111100110",
  1142=>"111010110",
  1143=>"011010011",
  1144=>"101000100",
  1145=>"000010000",
  1146=>"011001010",
  1147=>"111111001",
  1148=>"100100001",
  1149=>"110110000",
  1150=>"010110000",
  1151=>"000101000",
  1152=>"011011100",
  1153=>"111000111",
  1154=>"101100001",
  1155=>"100111010",
  1156=>"000000000",
  1157=>"010010010",
  1158=>"010111111",
  1159=>"101000111",
  1160=>"001011111",
  1161=>"001000001",
  1162=>"101111100",
  1163=>"010110101",
  1164=>"111000101",
  1165=>"111110011",
  1166=>"010111001",
  1167=>"010101011",
  1168=>"001100110",
  1169=>"101101110",
  1170=>"101000010",
  1171=>"001000100",
  1172=>"001001000",
  1173=>"110000001",
  1174=>"001111001",
  1175=>"101101110",
  1176=>"010011010",
  1177=>"110001101",
  1178=>"010100110",
  1179=>"001111110",
  1180=>"001111010",
  1181=>"111110100",
  1182=>"000100111",
  1183=>"011010001",
  1184=>"001100111",
  1185=>"110000011",
  1186=>"100101100",
  1187=>"011010000",
  1188=>"000110100",
  1189=>"000100011",
  1190=>"100011001",
  1191=>"000110110",
  1192=>"100001001",
  1193=>"101000000",
  1194=>"001011000",
  1195=>"001011000",
  1196=>"110101101",
  1197=>"111100000",
  1198=>"000000100",
  1199=>"111000101",
  1200=>"011101101",
  1201=>"011011101",
  1202=>"000101111",
  1203=>"101001000",
  1204=>"011110000",
  1205=>"000110001",
  1206=>"000100111",
  1207=>"001000110",
  1208=>"001001101",
  1209=>"000110001",
  1210=>"010100010",
  1211=>"110110100",
  1212=>"011101001",
  1213=>"101001101",
  1214=>"100101111",
  1215=>"101111000",
  1216=>"011001000",
  1217=>"100001100",
  1218=>"111110011",
  1219=>"110101010",
  1220=>"000001111",
  1221=>"110100111",
  1222=>"000110010",
  1223=>"100000110",
  1224=>"011110101",
  1225=>"101001101",
  1226=>"100000101",
  1227=>"110110111",
  1228=>"110000111",
  1229=>"111010110",
  1230=>"001010110",
  1231=>"111000011",
  1232=>"111000011",
  1233=>"011101001",
  1234=>"101010010",
  1235=>"000011100",
  1236=>"101111001",
  1237=>"000110101",
  1238=>"001011000",
  1239=>"111111111",
  1240=>"000000000",
  1241=>"110111011",
  1242=>"001111001",
  1243=>"011101100",
  1244=>"111100010",
  1245=>"101010001",
  1246=>"010010010",
  1247=>"101110011",
  1248=>"111110101",
  1249=>"010101111",
  1250=>"110011011",
  1251=>"000011011",
  1252=>"101001110",
  1253=>"101001011",
  1254=>"010100110",
  1255=>"100010000",
  1256=>"110111110",
  1257=>"110111100",
  1258=>"001110010",
  1259=>"000010011",
  1260=>"010111101",
  1261=>"001101100",
  1262=>"100110000",
  1263=>"000100001",
  1264=>"010000011",
  1265=>"100001110",
  1266=>"010011110",
  1267=>"011000001",
  1268=>"111001011",
  1269=>"000000100",
  1270=>"000000100",
  1271=>"111000111",
  1272=>"001011001",
  1273=>"111010111",
  1274=>"110000101",
  1275=>"100010100",
  1276=>"000010001",
  1277=>"011100110",
  1278=>"111011110",
  1279=>"010001111",
  1280=>"111100111",
  1281=>"100001111",
  1282=>"111010011",
  1283=>"001101010",
  1284=>"100001100",
  1285=>"101001100",
  1286=>"011010100",
  1287=>"110110100",
  1288=>"001110100",
  1289=>"001000001",
  1290=>"010000011",
  1291=>"111001000",
  1292=>"011101000",
  1293=>"000010000",
  1294=>"000001110",
  1295=>"100011000",
  1296=>"110101000",
  1297=>"010100000",
  1298=>"110110101",
  1299=>"100101001",
  1300=>"000111011",
  1301=>"011101001",
  1302=>"001101100",
  1303=>"010111110",
  1304=>"001010010",
  1305=>"110111010",
  1306=>"000010001",
  1307=>"111101100",
  1308=>"000101011",
  1309=>"000001001",
  1310=>"010001100",
  1311=>"100000000",
  1312=>"000000001",
  1313=>"001101101",
  1314=>"110011111",
  1315=>"110000101",
  1316=>"010110110",
  1317=>"010010011",
  1318=>"100000000",
  1319=>"100101111",
  1320=>"000000011",
  1321=>"101110100",
  1322=>"111011010",
  1323=>"011110001",
  1324=>"101101010",
  1325=>"010000011",
  1326=>"010001010",
  1327=>"001000110",
  1328=>"011011100",
  1329=>"011111011",
  1330=>"000101001",
  1331=>"110100101",
  1332=>"100101000",
  1333=>"011010100",
  1334=>"001011111",
  1335=>"111000111",
  1336=>"110101101",
  1337=>"000110111",
  1338=>"101010101",
  1339=>"010010011",
  1340=>"100000100",
  1341=>"101110000",
  1342=>"111101110",
  1343=>"111010101",
  1344=>"001001010",
  1345=>"100100010",
  1346=>"100100001",
  1347=>"111001011",
  1348=>"111111000",
  1349=>"011111101",
  1350=>"011001001",
  1351=>"100000010",
  1352=>"010101010",
  1353=>"100110101",
  1354=>"000001011",
  1355=>"101101011",
  1356=>"000110010",
  1357=>"011000010",
  1358=>"010001111",
  1359=>"111001000",
  1360=>"100011101",
  1361=>"000110000",
  1362=>"100111010",
  1363=>"000001001",
  1364=>"001000100",
  1365=>"001101100",
  1366=>"111000110",
  1367=>"011100101",
  1368=>"010111001",
  1369=>"100010010",
  1370=>"000111111",
  1371=>"110011101",
  1372=>"111111111",
  1373=>"100111101",
  1374=>"000001010",
  1375=>"011101111",
  1376=>"111011110",
  1377=>"111011100",
  1378=>"111101101",
  1379=>"000010101",
  1380=>"001110001",
  1381=>"100110110",
  1382=>"000100001",
  1383=>"100010110",
  1384=>"101111101",
  1385=>"110110110",
  1386=>"001011010",
  1387=>"011111011",
  1388=>"111000010",
  1389=>"111011111",
  1390=>"000000110",
  1391=>"110011000",
  1392=>"001101001",
  1393=>"000010111",
  1394=>"011010110",
  1395=>"000111101",
  1396=>"000000101",
  1397=>"010111000",
  1398=>"111001000",
  1399=>"110110100",
  1400=>"110101111",
  1401=>"100000101",
  1402=>"001100111",
  1403=>"111111011",
  1404=>"111100110",
  1405=>"000001010",
  1406=>"000001000",
  1407=>"000101110",
  1408=>"100010011",
  1409=>"011100111",
  1410=>"011111110",
  1411=>"011100100",
  1412=>"010001111",
  1413=>"100000000",
  1414=>"010001000",
  1415=>"001001011",
  1416=>"011100011",
  1417=>"011001100",
  1418=>"000001010",
  1419=>"101100001",
  1420=>"000000000",
  1421=>"011010001",
  1422=>"001000001",
  1423=>"011000111",
  1424=>"000101111",
  1425=>"010010001",
  1426=>"001110111",
  1427=>"000011001",
  1428=>"110100110",
  1429=>"011001100",
  1430=>"011110000",
  1431=>"101100011",
  1432=>"000110110",
  1433=>"000110010",
  1434=>"000000111",
  1435=>"010001011",
  1436=>"010100011",
  1437=>"001001001",
  1438=>"001111111",
  1439=>"001010110",
  1440=>"101110000",
  1441=>"011100001",
  1442=>"000100010",
  1443=>"101000000",
  1444=>"000111110",
  1445=>"110010111",
  1446=>"001010011",
  1447=>"001000110",
  1448=>"111100110",
  1449=>"001011001",
  1450=>"100011010",
  1451=>"011111001",
  1452=>"101101000",
  1453=>"011111000",
  1454=>"000001011",
  1455=>"000110111",
  1456=>"111101100",
  1457=>"001010001",
  1458=>"010011010",
  1459=>"001011111",
  1460=>"111000100",
  1461=>"101000111",
  1462=>"110000100",
  1463=>"001010110",
  1464=>"111111010",
  1465=>"001000000",
  1466=>"101001000",
  1467=>"000011100",
  1468=>"110111101",
  1469=>"010011110",
  1470=>"001101011",
  1471=>"100011101",
  1472=>"001001110",
  1473=>"000100101",
  1474=>"100101111",
  1475=>"000111110",
  1476=>"001110101",
  1477=>"111111000",
  1478=>"010001001",
  1479=>"100111111",
  1480=>"000010110",
  1481=>"101001101",
  1482=>"101000101",
  1483=>"000001001",
  1484=>"100100100",
  1485=>"011000001",
  1486=>"011101000",
  1487=>"011110100",
  1488=>"011101100",
  1489=>"101001001",
  1490=>"010111000",
  1491=>"010110111",
  1492=>"001110001",
  1493=>"001000011",
  1494=>"101101001",
  1495=>"110000010",
  1496=>"100010011",
  1497=>"111111110",
  1498=>"010110000",
  1499=>"100101111",
  1500=>"010011000",
  1501=>"010011111",
  1502=>"110011100",
  1503=>"000100110",
  1504=>"100001011",
  1505=>"101101100",
  1506=>"110100010",
  1507=>"100100001",
  1508=>"000100001",
  1509=>"011011111",
  1510=>"011010111",
  1511=>"011010010",
  1512=>"101001010",
  1513=>"001110100",
  1514=>"011101101",
  1515=>"111010101",
  1516=>"001110011",
  1517=>"101101101",
  1518=>"110011110",
  1519=>"010101010",
  1520=>"110100011",
  1521=>"010110101",
  1522=>"111101000",
  1523=>"010101010",
  1524=>"100001111",
  1525=>"111111111",
  1526=>"011000001",
  1527=>"000010100",
  1528=>"110000011",
  1529=>"100110011",
  1530=>"001110000",
  1531=>"100111101",
  1532=>"101110101",
  1533=>"001110011",
  1534=>"100101000",
  1535=>"110110110",
  1536=>"110011111",
  1537=>"100100111",
  1538=>"001011111",
  1539=>"001000111",
  1540=>"000000011",
  1541=>"110111000",
  1542=>"010010011",
  1543=>"111000101",
  1544=>"111010100",
  1545=>"010101110",
  1546=>"010101000",
  1547=>"010010111",
  1548=>"011001000",
  1549=>"010000110",
  1550=>"101100001",
  1551=>"001110111",
  1552=>"101100001",
  1553=>"001110010",
  1554=>"011110111",
  1555=>"011101101",
  1556=>"000101001",
  1557=>"000101000",
  1558=>"010100011",
  1559=>"001000101",
  1560=>"010000001",
  1561=>"000111110",
  1562=>"001000101",
  1563=>"010011010",
  1564=>"100001000",
  1565=>"010101000",
  1566=>"111001000",
  1567=>"011110000",
  1568=>"011000010",
  1569=>"100110000",
  1570=>"111001000",
  1571=>"000001100",
  1572=>"001110110",
  1573=>"100000001",
  1574=>"100100001",
  1575=>"111101111",
  1576=>"100101001",
  1577=>"100101100",
  1578=>"000000000",
  1579=>"011110010",
  1580=>"000001010",
  1581=>"110101111",
  1582=>"001010100",
  1583=>"100010110",
  1584=>"000000100",
  1585=>"101101000",
  1586=>"100001000",
  1587=>"011100110",
  1588=>"100000010",
  1589=>"011010010",
  1590=>"011000011",
  1591=>"000000101",
  1592=>"000100101",
  1593=>"111111101",
  1594=>"100000011",
  1595=>"111000000",
  1596=>"011100000",
  1597=>"110110111",
  1598=>"001110111",
  1599=>"111101111",
  1600=>"110110001",
  1601=>"001000101",
  1602=>"001110010",
  1603=>"101111111",
  1604=>"011011110",
  1605=>"001111100",
  1606=>"000000001",
  1607=>"000100001",
  1608=>"101100101",
  1609=>"010101000",
  1610=>"000000101",
  1611=>"001000000",
  1612=>"111100010",
  1613=>"011000101",
  1614=>"010111100",
  1615=>"100000000",
  1616=>"100000010",
  1617=>"001010010",
  1618=>"000101110",
  1619=>"000001000",
  1620=>"101100010",
  1621=>"100010001",
  1622=>"000000110",
  1623=>"101110111",
  1624=>"001000100",
  1625=>"000011100",
  1626=>"000010010",
  1627=>"000010001",
  1628=>"001000100",
  1629=>"010110000",
  1630=>"111100001",
  1631=>"000010101",
  1632=>"010001001",
  1633=>"000010110",
  1634=>"010001001",
  1635=>"101000011",
  1636=>"010011111",
  1637=>"111110001",
  1638=>"001101010",
  1639=>"100111001",
  1640=>"000011110",
  1641=>"000100111",
  1642=>"110111011",
  1643=>"010110100",
  1644=>"000110101",
  1645=>"111001101",
  1646=>"100111101",
  1647=>"111001000",
  1648=>"010000110",
  1649=>"000001111",
  1650=>"001000000",
  1651=>"111010100",
  1652=>"101000110",
  1653=>"111000110",
  1654=>"111110110",
  1655=>"011111111",
  1656=>"111011111",
  1657=>"010100011",
  1658=>"000000101",
  1659=>"011111110",
  1660=>"010010000",
  1661=>"101001110",
  1662=>"111110010",
  1663=>"011110110",
  1664=>"000110001",
  1665=>"111010000",
  1666=>"110111001",
  1667=>"001110110",
  1668=>"100100001",
  1669=>"110011101",
  1670=>"100001110",
  1671=>"101000010",
  1672=>"001100110",
  1673=>"111101101",
  1674=>"100001100",
  1675=>"101010111",
  1676=>"000001001",
  1677=>"000110010",
  1678=>"111110101",
  1679=>"001110011",
  1680=>"101101111",
  1681=>"110010010",
  1682=>"010010101",
  1683=>"111001111",
  1684=>"000100000",
  1685=>"111110111",
  1686=>"000100001",
  1687=>"010000101",
  1688=>"000001100",
  1689=>"000100100",
  1690=>"011101100",
  1691=>"000101001",
  1692=>"111001000",
  1693=>"111011010",
  1694=>"100111011",
  1695=>"010011110",
  1696=>"110110001",
  1697=>"100001101",
  1698=>"000110111",
  1699=>"111011110",
  1700=>"101101001",
  1701=>"101010001",
  1702=>"000001111",
  1703=>"101000110",
  1704=>"011010110",
  1705=>"000111001",
  1706=>"111100010",
  1707=>"010101011",
  1708=>"000001001",
  1709=>"101001011",
  1710=>"111110101",
  1711=>"100011110",
  1712=>"110001011",
  1713=>"011000110",
  1714=>"001100010",
  1715=>"101011101",
  1716=>"000010010",
  1717=>"010111110",
  1718=>"111110100",
  1719=>"010001011",
  1720=>"100000101",
  1721=>"111101100",
  1722=>"101110011",
  1723=>"001011101",
  1724=>"100111010",
  1725=>"111000101",
  1726=>"000000100",
  1727=>"011001011",
  1728=>"101000001",
  1729=>"000111011",
  1730=>"000101001",
  1731=>"011101001",
  1732=>"000011010",
  1733=>"101101111",
  1734=>"100101011",
  1735=>"000011010",
  1736=>"001010011",
  1737=>"011011001",
  1738=>"111011101",
  1739=>"000110110",
  1740=>"000101001",
  1741=>"110101000",
  1742=>"011100001",
  1743=>"111011111",
  1744=>"100000011",
  1745=>"101000101",
  1746=>"111100110",
  1747=>"010011001",
  1748=>"001000001",
  1749=>"001100111",
  1750=>"011100000",
  1751=>"000101001",
  1752=>"000011110",
  1753=>"001011101",
  1754=>"111101111",
  1755=>"011101000",
  1756=>"100101110",
  1757=>"000011000",
  1758=>"100001011",
  1759=>"100010001",
  1760=>"000010010",
  1761=>"111111111",
  1762=>"101011100",
  1763=>"111110111",
  1764=>"001010110",
  1765=>"010000111",
  1766=>"001001010",
  1767=>"010111000",
  1768=>"000001010",
  1769=>"000001001",
  1770=>"101001001",
  1771=>"111001000",
  1772=>"011010000",
  1773=>"101111100",
  1774=>"001111101",
  1775=>"000101111",
  1776=>"001110010",
  1777=>"000110000",
  1778=>"110101101",
  1779=>"001001011",
  1780=>"011011000",
  1781=>"101100001",
  1782=>"010100000",
  1783=>"100001010",
  1784=>"101010111",
  1785=>"010000010",
  1786=>"001100111",
  1787=>"010110010",
  1788=>"011101100",
  1789=>"111010000",
  1790=>"000101111",
  1791=>"000100001",
  1792=>"001011000",
  1793=>"000111111",
  1794=>"011010111",
  1795=>"101001001",
  1796=>"100111001",
  1797=>"100111111",
  1798=>"000110101",
  1799=>"100110100",
  1800=>"111101010",
  1801=>"001111011",
  1802=>"100101110",
  1803=>"111010111",
  1804=>"010111010",
  1805=>"011010001",
  1806=>"110010110",
  1807=>"011100011",
  1808=>"110010000",
  1809=>"111000100",
  1810=>"111011101",
  1811=>"000100000",
  1812=>"111100001",
  1813=>"010010110",
  1814=>"010011110",
  1815=>"111110010",
  1816=>"001111001",
  1817=>"010010101",
  1818=>"100100010",
  1819=>"110001100",
  1820=>"000110000",
  1821=>"000111011",
  1822=>"000010011",
  1823=>"111011111",
  1824=>"101100100",
  1825=>"111011101",
  1826=>"000101011",
  1827=>"010100001",
  1828=>"100111101",
  1829=>"000111001",
  1830=>"110011110",
  1831=>"000011111",
  1832=>"000100000",
  1833=>"110100001",
  1834=>"000000110",
  1835=>"001100101",
  1836=>"100100011",
  1837=>"011001111",
  1838=>"000000001",
  1839=>"010100001",
  1840=>"001111110",
  1841=>"101101111",
  1842=>"011110011",
  1843=>"111110111",
  1844=>"001111000",
  1845=>"001111011",
  1846=>"010011011",
  1847=>"000010100",
  1848=>"111010111",
  1849=>"110101011",
  1850=>"010100001",
  1851=>"100110111",
  1852=>"110000101",
  1853=>"101000001",
  1854=>"111100100",
  1855=>"010111000",
  1856=>"100001100",
  1857=>"010110101",
  1858=>"111111101",
  1859=>"110110000",
  1860=>"101111010",
  1861=>"000000001",
  1862=>"000101111",
  1863=>"010000100",
  1864=>"011100111",
  1865=>"001010010",
  1866=>"000000001",
  1867=>"100011100",
  1868=>"000100101",
  1869=>"110011010",
  1870=>"101100100",
  1871=>"100100011",
  1872=>"011101000",
  1873=>"110001011",
  1874=>"000100010",
  1875=>"111000010",
  1876=>"101000101",
  1877=>"000011001",
  1878=>"000110000",
  1879=>"100100110",
  1880=>"101100011",
  1881=>"110100010",
  1882=>"111010000",
  1883=>"111011100",
  1884=>"001101000",
  1885=>"111101100",
  1886=>"100101000",
  1887=>"001010000",
  1888=>"110100100",
  1889=>"010001100",
  1890=>"110001010",
  1891=>"011110011",
  1892=>"001011100",
  1893=>"100000101",
  1894=>"100010111",
  1895=>"011101111",
  1896=>"001010100",
  1897=>"101101101",
  1898=>"001011001",
  1899=>"000110110",
  1900=>"011110000",
  1901=>"101001000",
  1902=>"000010101",
  1903=>"001100110",
  1904=>"100000111",
  1905=>"110100101",
  1906=>"011000111",
  1907=>"000001101",
  1908=>"010100100",
  1909=>"000100100",
  1910=>"100011101",
  1911=>"010000010",
  1912=>"010011111",
  1913=>"100010000",
  1914=>"011001001",
  1915=>"111100010",
  1916=>"101010100",
  1917=>"001110011",
  1918=>"101000000",
  1919=>"111111111",
  1920=>"111011100",
  1921=>"001000110",
  1922=>"010101010",
  1923=>"000100100",
  1924=>"100011010",
  1925=>"011000101",
  1926=>"100101001",
  1927=>"010000101",
  1928=>"111110101",
  1929=>"111010010",
  1930=>"111110001",
  1931=>"000001100",
  1932=>"000100111",
  1933=>"111010010",
  1934=>"111001010",
  1935=>"100011111",
  1936=>"111010001",
  1937=>"101000100",
  1938=>"010101000",
  1939=>"011011110",
  1940=>"101110010",
  1941=>"110010111",
  1942=>"101010111",
  1943=>"011101001",
  1944=>"100100000",
  1945=>"101011111",
  1946=>"110001110",
  1947=>"110011101",
  1948=>"110100110",
  1949=>"000011001",
  1950=>"011101110",
  1951=>"001000001",
  1952=>"110101110",
  1953=>"101110111",
  1954=>"010101101",
  1955=>"000100010",
  1956=>"000100101",
  1957=>"111010010",
  1958=>"001100000",
  1959=>"010100001",
  1960=>"011110000",
  1961=>"110111111",
  1962=>"110011011",
  1963=>"111001110",
  1964=>"000110101",
  1965=>"000011111",
  1966=>"001101111",
  1967=>"100111100",
  1968=>"000010101",
  1969=>"111011010",
  1970=>"101110010",
  1971=>"101000001",
  1972=>"110000100",
  1973=>"111101111",
  1974=>"111010100",
  1975=>"111101101",
  1976=>"010000110",
  1977=>"100100100",
  1978=>"001100110",
  1979=>"011011101",
  1980=>"110010111",
  1981=>"100010000",
  1982=>"110110010",
  1983=>"100000010",
  1984=>"111000011",
  1985=>"101111011",
  1986=>"110100001",
  1987=>"100111000",
  1988=>"101011010",
  1989=>"110001100",
  1990=>"111000110",
  1991=>"100000100",
  1992=>"000001010",
  1993=>"001100000",
  1994=>"100111101",
  1995=>"100111100",
  1996=>"110100111",
  1997=>"010000000",
  1998=>"100110100",
  1999=>"111101101",
  2000=>"011110111",
  2001=>"011100001",
  2002=>"010110101",
  2003=>"011111011",
  2004=>"111011100",
  2005=>"101111010",
  2006=>"101000001",
  2007=>"001110011",
  2008=>"010111101",
  2009=>"100001110",
  2010=>"010010110",
  2011=>"101101000",
  2012=>"100101010",
  2013=>"111111110",
  2014=>"000000001",
  2015=>"100001100",
  2016=>"101111010",
  2017=>"110011001",
  2018=>"100101101",
  2019=>"101101111",
  2020=>"001100101",
  2021=>"001000110",
  2022=>"011100100",
  2023=>"110100010",
  2024=>"001000000",
  2025=>"011111011",
  2026=>"111101011",
  2027=>"010000000",
  2028=>"001011101",
  2029=>"010101100",
  2030=>"001111101",
  2031=>"100011111",
  2032=>"001001000",
  2033=>"010000000",
  2034=>"000100001",
  2035=>"101110111",
  2036=>"001011001",
  2037=>"100111000",
  2038=>"111011001",
  2039=>"001100111",
  2040=>"101111110",
  2041=>"111100010",
  2042=>"000001101",
  2043=>"100000000",
  2044=>"100110100",
  2045=>"100110011",
  2046=>"010111001",
  2047=>"101001111",
  2048=>"111110011",
  2049=>"110111111",
  2050=>"011111100",
  2051=>"001011111",
  2052=>"000110110",
  2053=>"101001101",
  2054=>"111000001",
  2055=>"101111101",
  2056=>"110110010",
  2057=>"010110010",
  2058=>"000001110",
  2059=>"110000010",
  2060=>"001101000",
  2061=>"011101000",
  2062=>"001001101",
  2063=>"011000000",
  2064=>"000011101",
  2065=>"000100010",
  2066=>"111101010",
  2067=>"100001000",
  2068=>"001111100",
  2069=>"000110101",
  2070=>"010000110",
  2071=>"100100000",
  2072=>"000101100",
  2073=>"000000001",
  2074=>"101101000",
  2075=>"110101011",
  2076=>"111011110",
  2077=>"001101110",
  2078=>"011110011",
  2079=>"110011000",
  2080=>"111010111",
  2081=>"100100000",
  2082=>"101111101",
  2083=>"100000001",
  2084=>"000111010",
  2085=>"001101011",
  2086=>"101000100",
  2087=>"000110110",
  2088=>"010101000",
  2089=>"111001111",
  2090=>"110110011",
  2091=>"100010001",
  2092=>"001000101",
  2093=>"100010011",
  2094=>"111111010",
  2095=>"001000000",
  2096=>"111011101",
  2097=>"000000111",
  2098=>"010101011",
  2099=>"110001110",
  2100=>"010010100",
  2101=>"010100100",
  2102=>"011001010",
  2103=>"011101000",
  2104=>"000000000",
  2105=>"011101100",
  2106=>"100111001",
  2107=>"110000100",
  2108=>"010011011",
  2109=>"010110100",
  2110=>"010010000",
  2111=>"001100110",
  2112=>"100101110",
  2113=>"010011011",
  2114=>"101001000",
  2115=>"001101010",
  2116=>"110011001",
  2117=>"000111100",
  2118=>"001100001",
  2119=>"000011101",
  2120=>"010010110",
  2121=>"100010100",
  2122=>"100010000",
  2123=>"000100110",
  2124=>"011000111",
  2125=>"111110010",
  2126=>"110111010",
  2127=>"111111111",
  2128=>"110101100",
  2129=>"001011011",
  2130=>"001010011",
  2131=>"111110111",
  2132=>"001100111",
  2133=>"101101011",
  2134=>"001000011",
  2135=>"000110111",
  2136=>"100111001",
  2137=>"011100111",
  2138=>"111110110",
  2139=>"011101011",
  2140=>"010011010",
  2141=>"000110000",
  2142=>"000000000",
  2143=>"000011101",
  2144=>"000010100",
  2145=>"001010101",
  2146=>"011100100",
  2147=>"111011011",
  2148=>"110001011",
  2149=>"000101111",
  2150=>"001000101",
  2151=>"011010101",
  2152=>"000100101",
  2153=>"100011011",
  2154=>"111111011",
  2155=>"001100101",
  2156=>"000100001",
  2157=>"011010001",
  2158=>"011010101",
  2159=>"001110101",
  2160=>"110001110",
  2161=>"001000000",
  2162=>"000001110",
  2163=>"011000010",
  2164=>"011101010",
  2165=>"111111010",
  2166=>"110001000",
  2167=>"110010000",
  2168=>"011100000",
  2169=>"001101111",
  2170=>"110110100",
  2171=>"110000111",
  2172=>"001001000",
  2173=>"111100100",
  2174=>"001100101",
  2175=>"101001100",
  2176=>"110001110",
  2177=>"010101111",
  2178=>"011011100",
  2179=>"010010011",
  2180=>"011101000",
  2181=>"110001001",
  2182=>"011011111",
  2183=>"010010000",
  2184=>"110000010",
  2185=>"110101000",
  2186=>"100011011",
  2187=>"110011011",
  2188=>"010010101",
  2189=>"000101110",
  2190=>"100110101",
  2191=>"101111001",
  2192=>"100110001",
  2193=>"110010000",
  2194=>"000001110",
  2195=>"101011100",
  2196=>"010000000",
  2197=>"101110010",
  2198=>"110010110",
  2199=>"011110000",
  2200=>"011000100",
  2201=>"011000100",
  2202=>"110111001",
  2203=>"000110101",
  2204=>"100000111",
  2205=>"111101001",
  2206=>"001010011",
  2207=>"100001011",
  2208=>"100110000",
  2209=>"111011101",
  2210=>"010011010",
  2211=>"101000011",
  2212=>"110001111",
  2213=>"111011110",
  2214=>"000111101",
  2215=>"100101101",
  2216=>"010010011",
  2217=>"101011000",
  2218=>"101010000",
  2219=>"001100011",
  2220=>"111001011",
  2221=>"100110111",
  2222=>"000010111",
  2223=>"111100010",
  2224=>"110111100",
  2225=>"000000001",
  2226=>"000001110",
  2227=>"001000000",
  2228=>"010000000",
  2229=>"111000100",
  2230=>"011000011",
  2231=>"100001010",
  2232=>"000110000",
  2233=>"100101111",
  2234=>"000000000",
  2235=>"011010001",
  2236=>"011110100",
  2237=>"100011011",
  2238=>"010111101",
  2239=>"111101010",
  2240=>"101001000",
  2241=>"110001011",
  2242=>"001111100",
  2243=>"010101001",
  2244=>"010111101",
  2245=>"001000010",
  2246=>"110010101",
  2247=>"001000000",
  2248=>"011011110",
  2249=>"110111110",
  2250=>"000011110",
  2251=>"000100001",
  2252=>"101110111",
  2253=>"001110011",
  2254=>"001101010",
  2255=>"110010010",
  2256=>"011101010",
  2257=>"100001001",
  2258=>"001110101",
  2259=>"000000101",
  2260=>"111110111",
  2261=>"001010101",
  2262=>"011101110",
  2263=>"000000000",
  2264=>"000111110",
  2265=>"110110010",
  2266=>"001110011",
  2267=>"111001110",
  2268=>"101111111",
  2269=>"100011000",
  2270=>"110000000",
  2271=>"100000110",
  2272=>"111111011",
  2273=>"010001010",
  2274=>"011111100",
  2275=>"000011111",
  2276=>"100000101",
  2277=>"110100001",
  2278=>"010100101",
  2279=>"100010000",
  2280=>"101110011",
  2281=>"010100110",
  2282=>"011101100",
  2283=>"000101000",
  2284=>"100101000",
  2285=>"101101010",
  2286=>"110001000",
  2287=>"100000100",
  2288=>"000011110",
  2289=>"110110011",
  2290=>"011010000",
  2291=>"001110011",
  2292=>"110010011",
  2293=>"101001101",
  2294=>"011110011",
  2295=>"011000001",
  2296=>"110100011",
  2297=>"011111010",
  2298=>"000001100",
  2299=>"011100011",
  2300=>"101000010",
  2301=>"101011011",
  2302=>"000011100",
  2303=>"010010110",
  2304=>"110001110",
  2305=>"111010100",
  2306=>"011101000",
  2307=>"100000111",
  2308=>"010100000",
  2309=>"100001110",
  2310=>"000101100",
  2311=>"101100110",
  2312=>"011000001",
  2313=>"000111010",
  2314=>"111110101",
  2315=>"101010011",
  2316=>"010100010",
  2317=>"011011100",
  2318=>"000010100",
  2319=>"011111110",
  2320=>"001101110",
  2321=>"011101101",
  2322=>"001111110",
  2323=>"010010001",
  2324=>"110100010",
  2325=>"001100010",
  2326=>"000011101",
  2327=>"101001101",
  2328=>"010011010",
  2329=>"001000010",
  2330=>"100010100",
  2331=>"111001110",
  2332=>"110101101",
  2333=>"101001101",
  2334=>"101011001",
  2335=>"000010100",
  2336=>"011010000",
  2337=>"011111101",
  2338=>"001111101",
  2339=>"001111001",
  2340=>"100110101",
  2341=>"110010001",
  2342=>"000101101",
  2343=>"110101100",
  2344=>"100010110",
  2345=>"110100110",
  2346=>"010100011",
  2347=>"110000010",
  2348=>"111100111",
  2349=>"010110111",
  2350=>"011111110",
  2351=>"100100000",
  2352=>"010101001",
  2353=>"000101101",
  2354=>"100000010",
  2355=>"010100000",
  2356=>"101011101",
  2357=>"000001000",
  2358=>"101111111",
  2359=>"001000001",
  2360=>"000010010",
  2361=>"010101010",
  2362=>"111100010",
  2363=>"011001000",
  2364=>"011101011",
  2365=>"111101111",
  2366=>"101101111",
  2367=>"010100010",
  2368=>"011010011",
  2369=>"100110101",
  2370=>"111000110",
  2371=>"111111000",
  2372=>"101001000",
  2373=>"101101001",
  2374=>"011100001",
  2375=>"010010000",
  2376=>"111101111",
  2377=>"011100000",
  2378=>"100110100",
  2379=>"000010111",
  2380=>"100100101",
  2381=>"011101000",
  2382=>"111111000",
  2383=>"111100010",
  2384=>"110010111",
  2385=>"111001101",
  2386=>"010011001",
  2387=>"111101101",
  2388=>"101011001",
  2389=>"010010001",
  2390=>"110100100",
  2391=>"011101111",
  2392=>"001011010",
  2393=>"001010111",
  2394=>"100011100",
  2395=>"010000000",
  2396=>"010000010",
  2397=>"110101110",
  2398=>"001110011",
  2399=>"110001100",
  2400=>"011010101",
  2401=>"000010010",
  2402=>"001001011",
  2403=>"000100010",
  2404=>"101011011",
  2405=>"111001101",
  2406=>"010001110",
  2407=>"011110010",
  2408=>"001000100",
  2409=>"110101011",
  2410=>"100110101",
  2411=>"011111010",
  2412=>"010000001",
  2413=>"111110110",
  2414=>"000101010",
  2415=>"010001100",
  2416=>"000101000",
  2417=>"000001100",
  2418=>"001101010",
  2419=>"100000001",
  2420=>"001011000",
  2421=>"110001101",
  2422=>"111100001",
  2423=>"001110101",
  2424=>"111101101",
  2425=>"101010010",
  2426=>"001110001",
  2427=>"000011011",
  2428=>"110000010",
  2429=>"111010111",
  2430=>"110100111",
  2431=>"011000011",
  2432=>"000100000",
  2433=>"001000001",
  2434=>"010001100",
  2435=>"011100010",
  2436=>"000011110",
  2437=>"000000010",
  2438=>"001011001",
  2439=>"011011111",
  2440=>"110110110",
  2441=>"101000011",
  2442=>"010101000",
  2443=>"011000110",
  2444=>"011001010",
  2445=>"000010000",
  2446=>"110100100",
  2447=>"010000010",
  2448=>"011100101",
  2449=>"001011000",
  2450=>"100101101",
  2451=>"000010001",
  2452=>"000101100",
  2453=>"011111010",
  2454=>"111111111",
  2455=>"011110000",
  2456=>"100001000",
  2457=>"000100111",
  2458=>"011110110",
  2459=>"000011100",
  2460=>"111110110",
  2461=>"010011101",
  2462=>"101111101",
  2463=>"000011000",
  2464=>"000101111",
  2465=>"100100011",
  2466=>"110010001",
  2467=>"000000011",
  2468=>"010000011",
  2469=>"101011110",
  2470=>"001100010",
  2471=>"000011010",
  2472=>"100110100",
  2473=>"111011110",
  2474=>"001010111",
  2475=>"101010101",
  2476=>"000111000",
  2477=>"011101010",
  2478=>"000110010",
  2479=>"101111111",
  2480=>"001111011",
  2481=>"101001101",
  2482=>"011111001",
  2483=>"011111100",
  2484=>"010101011",
  2485=>"010110000",
  2486=>"010011110",
  2487=>"110101011",
  2488=>"101100100",
  2489=>"001111110",
  2490=>"110001000",
  2491=>"001000101",
  2492=>"001110101",
  2493=>"001110110",
  2494=>"110111110",
  2495=>"000111111",
  2496=>"000010110",
  2497=>"000000110",
  2498=>"111010110",
  2499=>"011110011",
  2500=>"110110100",
  2501=>"000001001",
  2502=>"000010000",
  2503=>"011101110",
  2504=>"011111100",
  2505=>"101011111",
  2506=>"110001111",
  2507=>"111010000",
  2508=>"000011100",
  2509=>"100110000",
  2510=>"111101010",
  2511=>"111111001",
  2512=>"000000011",
  2513=>"011111111",
  2514=>"010111001",
  2515=>"011101111",
  2516=>"101111000",
  2517=>"011101011",
  2518=>"011111110",
  2519=>"000000100",
  2520=>"000100001",
  2521=>"010011011",
  2522=>"111010001",
  2523=>"101110100",
  2524=>"011100110",
  2525=>"100010100",
  2526=>"101001000",
  2527=>"111111101",
  2528=>"101010010",
  2529=>"111110000",
  2530=>"000100101",
  2531=>"010000101",
  2532=>"011001101",
  2533=>"001000101",
  2534=>"101111110",
  2535=>"101100010",
  2536=>"011110011",
  2537=>"111110101",
  2538=>"000000111",
  2539=>"111010101",
  2540=>"111101110",
  2541=>"001101100",
  2542=>"001010100",
  2543=>"011110100",
  2544=>"010110011",
  2545=>"000011000",
  2546=>"010010010",
  2547=>"011000000",
  2548=>"010111110",
  2549=>"010100010",
  2550=>"010111110",
  2551=>"101000011",
  2552=>"110010111",
  2553=>"000111111",
  2554=>"000111001",
  2555=>"001100010",
  2556=>"100010001",
  2557=>"010000010",
  2558=>"111111010",
  2559=>"101010011",
  2560=>"000000110",
  2561=>"111011000",
  2562=>"110000000",
  2563=>"111010010",
  2564=>"000100111",
  2565=>"010000111",
  2566=>"111000011",
  2567=>"001010100",
  2568=>"011011001",
  2569=>"111011011",
  2570=>"011111100",
  2571=>"100000111",
  2572=>"011111010",
  2573=>"110101001",
  2574=>"111101011",
  2575=>"000101111",
  2576=>"110110010",
  2577=>"111110101",
  2578=>"111011001",
  2579=>"001110000",
  2580=>"001000100",
  2581=>"011110011",
  2582=>"110010111",
  2583=>"010001010",
  2584=>"000100001",
  2585=>"011101011",
  2586=>"010110111",
  2587=>"000111000",
  2588=>"111101001",
  2589=>"101010010",
  2590=>"000101011",
  2591=>"100001001",
  2592=>"000000101",
  2593=>"001000001",
  2594=>"100100100",
  2595=>"110000101",
  2596=>"101101101",
  2597=>"011100010",
  2598=>"110100100",
  2599=>"001001000",
  2600=>"001101111",
  2601=>"110000010",
  2602=>"000000100",
  2603=>"110011111",
  2604=>"001100001",
  2605=>"100001101",
  2606=>"010010111",
  2607=>"001111011",
  2608=>"101011011",
  2609=>"011101100",
  2610=>"010001010",
  2611=>"101111111",
  2612=>"100000000",
  2613=>"111000011",
  2614=>"100011100",
  2615=>"111011100",
  2616=>"001100000",
  2617=>"001100001",
  2618=>"001010011",
  2619=>"001110010",
  2620=>"010001101",
  2621=>"110110000",
  2622=>"001101110",
  2623=>"100100000",
  2624=>"101101111",
  2625=>"110111010",
  2626=>"010000100",
  2627=>"111101100",
  2628=>"011110000",
  2629=>"010001000",
  2630=>"000001010",
  2631=>"000000001",
  2632=>"010110110",
  2633=>"011101110",
  2634=>"101000011",
  2635=>"111100011",
  2636=>"001010101",
  2637=>"100001100",
  2638=>"010110111",
  2639=>"100110110",
  2640=>"111100011",
  2641=>"001111100",
  2642=>"011010111",
  2643=>"000000011",
  2644=>"100001011",
  2645=>"110011101",
  2646=>"000110001",
  2647=>"001011100",
  2648=>"000101101",
  2649=>"001001100",
  2650=>"000101111",
  2651=>"001110111",
  2652=>"100010001",
  2653=>"101001000",
  2654=>"000111100",
  2655=>"000101011",
  2656=>"000001100",
  2657=>"111001111",
  2658=>"110010011",
  2659=>"110101011",
  2660=>"001101011",
  2661=>"010010000",
  2662=>"111011100",
  2663=>"001100110",
  2664=>"001111101",
  2665=>"101110111",
  2666=>"100110111",
  2667=>"111111111",
  2668=>"001111011",
  2669=>"111100100",
  2670=>"010101001",
  2671=>"110011011",
  2672=>"101100010",
  2673=>"011110111",
  2674=>"001011011",
  2675=>"010110000",
  2676=>"110000110",
  2677=>"011100100",
  2678=>"110101011",
  2679=>"100010101",
  2680=>"100001000",
  2681=>"100100110",
  2682=>"110110010",
  2683=>"001001111",
  2684=>"000100101",
  2685=>"001000011",
  2686=>"100001011",
  2687=>"101111101",
  2688=>"100001010",
  2689=>"100000111",
  2690=>"000000110",
  2691=>"010001101",
  2692=>"011101110",
  2693=>"001110000",
  2694=>"000110010",
  2695=>"100100101",
  2696=>"000100000",
  2697=>"101111011",
  2698=>"010010101",
  2699=>"011101110",
  2700=>"010101010",
  2701=>"011001100",
  2702=>"100101100",
  2703=>"011001101",
  2704=>"011111101",
  2705=>"001110111",
  2706=>"111001111",
  2707=>"000010110",
  2708=>"011001011",
  2709=>"010110110",
  2710=>"001000000",
  2711=>"100011000",
  2712=>"000000001",
  2713=>"110100100",
  2714=>"000101101",
  2715=>"101100011",
  2716=>"011001011",
  2717=>"100111000",
  2718=>"010111110",
  2719=>"111001000",
  2720=>"111100111",
  2721=>"111011111",
  2722=>"101001101",
  2723=>"101101111",
  2724=>"110110100",
  2725=>"001110111",
  2726=>"011001001",
  2727=>"111000000",
  2728=>"010001000",
  2729=>"100001010",
  2730=>"100010001",
  2731=>"000011100",
  2732=>"110110001",
  2733=>"000000110",
  2734=>"101001101",
  2735=>"110101101",
  2736=>"000101110",
  2737=>"001010101",
  2738=>"111001011",
  2739=>"111100110",
  2740=>"001111011",
  2741=>"101011000",
  2742=>"110001000",
  2743=>"011100011",
  2744=>"000000110",
  2745=>"111100100",
  2746=>"110100100",
  2747=>"110000100",
  2748=>"001000010",
  2749=>"011011111",
  2750=>"111000011",
  2751=>"101010000",
  2752=>"000100111",
  2753=>"111010001",
  2754=>"100001001",
  2755=>"101111010",
  2756=>"010000111",
  2757=>"000100000",
  2758=>"011100011",
  2759=>"011000101",
  2760=>"111110111",
  2761=>"010110000",
  2762=>"010100010",
  2763=>"110010100",
  2764=>"001111011",
  2765=>"010011100",
  2766=>"001100110",
  2767=>"001010001",
  2768=>"111111111",
  2769=>"000011001",
  2770=>"100111010",
  2771=>"000010001",
  2772=>"111101111",
  2773=>"110010110",
  2774=>"001011101",
  2775=>"100101011",
  2776=>"110000010",
  2777=>"100010000",
  2778=>"000111110",
  2779=>"110000111",
  2780=>"000001001",
  2781=>"001000000",
  2782=>"000011000",
  2783=>"110001101",
  2784=>"111010000",
  2785=>"001100111",
  2786=>"101111011",
  2787=>"000000000",
  2788=>"000001100",
  2789=>"001110001",
  2790=>"011000100",
  2791=>"101111100",
  2792=>"110111111",
  2793=>"101011011",
  2794=>"001011101",
  2795=>"000111010",
  2796=>"101011001",
  2797=>"110111000",
  2798=>"010100100",
  2799=>"001000100",
  2800=>"111000111",
  2801=>"001001100",
  2802=>"010010011",
  2803=>"000101000",
  2804=>"100110010",
  2805=>"000010000",
  2806=>"000101110",
  2807=>"111010000",
  2808=>"000101011",
  2809=>"101101001",
  2810=>"010011011",
  2811=>"011101010",
  2812=>"000100010",
  2813=>"101001100",
  2814=>"100011110",
  2815=>"100001111",
  2816=>"100000011",
  2817=>"111000111",
  2818=>"011001101",
  2819=>"011010101",
  2820=>"000100111",
  2821=>"110100011",
  2822=>"011010001",
  2823=>"010010011",
  2824=>"100000011",
  2825=>"001010111",
  2826=>"010001001",
  2827=>"111111101",
  2828=>"001001110",
  2829=>"010010010",
  2830=>"001110000",
  2831=>"000101000",
  2832=>"000110011",
  2833=>"000010110",
  2834=>"001001110",
  2835=>"001010101",
  2836=>"100010110",
  2837=>"011101101",
  2838=>"011010011",
  2839=>"100011100",
  2840=>"001011011",
  2841=>"100100110",
  2842=>"111100010",
  2843=>"110011100",
  2844=>"000110010",
  2845=>"101101000",
  2846=>"100001111",
  2847=>"011111111",
  2848=>"111010001",
  2849=>"011010110",
  2850=>"110111011",
  2851=>"011111010",
  2852=>"010010000",
  2853=>"000011001",
  2854=>"000001100",
  2855=>"110101011",
  2856=>"110010011",
  2857=>"111000101",
  2858=>"001100010",
  2859=>"101011011",
  2860=>"000010001",
  2861=>"111001000",
  2862=>"100110101",
  2863=>"011001000",
  2864=>"010100000",
  2865=>"011000000",
  2866=>"100000000",
  2867=>"111010001",
  2868=>"001010001",
  2869=>"000100000",
  2870=>"111110111",
  2871=>"010100110",
  2872=>"000011111",
  2873=>"110101000",
  2874=>"011110111",
  2875=>"001001011",
  2876=>"010111010",
  2877=>"010000011",
  2878=>"100110011",
  2879=>"100000001",
  2880=>"001001111",
  2881=>"111110111",
  2882=>"111000100",
  2883=>"110101100",
  2884=>"010101010",
  2885=>"010101000",
  2886=>"000101001",
  2887=>"110010011",
  2888=>"011110101",
  2889=>"010000010",
  2890=>"001010001",
  2891=>"000000101",
  2892=>"011101001",
  2893=>"011111001",
  2894=>"000010011",
  2895=>"000010011",
  2896=>"000000000",
  2897=>"110100110",
  2898=>"110001001",
  2899=>"100001110",
  2900=>"100010000",
  2901=>"101001010",
  2902=>"011111011",
  2903=>"000000001",
  2904=>"111111110",
  2905=>"111111010",
  2906=>"111110011",
  2907=>"110001010",
  2908=>"111110000",
  2909=>"110111111",
  2910=>"111111111",
  2911=>"101001100",
  2912=>"010111101",
  2913=>"110011000",
  2914=>"000000100",
  2915=>"101000001",
  2916=>"000110011",
  2917=>"000001011",
  2918=>"101110000",
  2919=>"001001100",
  2920=>"100100111",
  2921=>"110100011",
  2922=>"111101001",
  2923=>"011100100",
  2924=>"111111101",
  2925=>"000111011",
  2926=>"100110001",
  2927=>"111111101",
  2928=>"110100000",
  2929=>"101100001",
  2930=>"001000010",
  2931=>"000100011",
  2932=>"101111010",
  2933=>"110000011",
  2934=>"101110000",
  2935=>"000110000",
  2936=>"100000011",
  2937=>"110101001",
  2938=>"001110100",
  2939=>"010000100",
  2940=>"111000111",
  2941=>"001001010",
  2942=>"011011110",
  2943=>"000000011",
  2944=>"101011110",
  2945=>"110011001",
  2946=>"110100111",
  2947=>"110001010",
  2948=>"001000010",
  2949=>"011111110",
  2950=>"000010111",
  2951=>"010011011",
  2952=>"001000100",
  2953=>"101010110",
  2954=>"110010100",
  2955=>"100110011",
  2956=>"110100110",
  2957=>"000011011",
  2958=>"111110111",
  2959=>"100100101",
  2960=>"000100011",
  2961=>"010101010",
  2962=>"000000111",
  2963=>"111010001",
  2964=>"110001110",
  2965=>"000010010",
  2966=>"000011101",
  2967=>"101011011",
  2968=>"011011101",
  2969=>"111001101",
  2970=>"011000101",
  2971=>"111000000",
  2972=>"000001001",
  2973=>"100100000",
  2974=>"001001111",
  2975=>"010000011",
  2976=>"010110001",
  2977=>"010001000",
  2978=>"001001010",
  2979=>"001001100",
  2980=>"000100011",
  2981=>"100001100",
  2982=>"101101111",
  2983=>"001100000",
  2984=>"001101000",
  2985=>"000111110",
  2986=>"001001010",
  2987=>"000001001",
  2988=>"100000000",
  2989=>"011011110",
  2990=>"100001110",
  2991=>"000001000",
  2992=>"010110101",
  2993=>"010111011",
  2994=>"100101010",
  2995=>"110110000",
  2996=>"100000101",
  2997=>"001000000",
  2998=>"000000001",
  2999=>"100110000",
  3000=>"000011010",
  3001=>"000100100",
  3002=>"111111101",
  3003=>"000010001",
  3004=>"001101100",
  3005=>"100000101",
  3006=>"111101101",
  3007=>"111101010",
  3008=>"000000111",
  3009=>"111001011",
  3010=>"111011101",
  3011=>"011010100",
  3012=>"010111000",
  3013=>"011100111",
  3014=>"000101110",
  3015=>"110010000",
  3016=>"110110100",
  3017=>"100000001",
  3018=>"010000001",
  3019=>"100101001",
  3020=>"000010001",
  3021=>"111010000",
  3022=>"100111101",
  3023=>"110111110",
  3024=>"001110100",
  3025=>"010101011",
  3026=>"011000110",
  3027=>"010000010",
  3028=>"010011100",
  3029=>"110001110",
  3030=>"010010010",
  3031=>"111101110",
  3032=>"011111101",
  3033=>"100100011",
  3034=>"000010010",
  3035=>"111010011",
  3036=>"100001100",
  3037=>"101110010",
  3038=>"001110000",
  3039=>"101010010",
  3040=>"011011010",
  3041=>"010100000",
  3042=>"000000001",
  3043=>"001101001",
  3044=>"110011100",
  3045=>"000111001",
  3046=>"100010000",
  3047=>"001100101",
  3048=>"110101000",
  3049=>"101111000",
  3050=>"111111011",
  3051=>"101110111",
  3052=>"010010000",
  3053=>"100010000",
  3054=>"000111111",
  3055=>"110011011",
  3056=>"110111111",
  3057=>"100000100",
  3058=>"001100100",
  3059=>"111000001",
  3060=>"011111101",
  3061=>"110001110",
  3062=>"011011100",
  3063=>"011010100",
  3064=>"001111011",
  3065=>"111001000",
  3066=>"100100001",
  3067=>"011101111",
  3068=>"100000000",
  3069=>"100111011",
  3070=>"001001111",
  3071=>"001001111",
  3072=>"110100110",
  3073=>"101100110",
  3074=>"010010010",
  3075=>"110101101",
  3076=>"011010101",
  3077=>"010001100",
  3078=>"110001000",
  3079=>"100101100",
  3080=>"100010100",
  3081=>"101110011",
  3082=>"101110011",
  3083=>"010011111",
  3084=>"011000101",
  3085=>"101001111",
  3086=>"001000111",
  3087=>"000000110",
  3088=>"100111101",
  3089=>"101001101",
  3090=>"100001111",
  3091=>"100011111",
  3092=>"101111111",
  3093=>"010010111",
  3094=>"011001101",
  3095=>"000000100",
  3096=>"110001001",
  3097=>"101100010",
  3098=>"011101001",
  3099=>"011101101",
  3100=>"111000101",
  3101=>"000000000",
  3102=>"000010001",
  3103=>"000001000",
  3104=>"000101010",
  3105=>"000110011",
  3106=>"010100111",
  3107=>"110110010",
  3108=>"110100010",
  3109=>"001001000",
  3110=>"101111111",
  3111=>"110010010",
  3112=>"010001001",
  3113=>"000110000",
  3114=>"001101001",
  3115=>"010100110",
  3116=>"010000001",
  3117=>"100101111",
  3118=>"000001111",
  3119=>"010110101",
  3120=>"110110000",
  3121=>"100110111",
  3122=>"110011001",
  3123=>"100100111",
  3124=>"010010100",
  3125=>"101011000",
  3126=>"001011011",
  3127=>"011011000",
  3128=>"010001110",
  3129=>"011000001",
  3130=>"000110111",
  3131=>"001011101",
  3132=>"100100111",
  3133=>"101101000",
  3134=>"110110101",
  3135=>"110100001",
  3136=>"111011111",
  3137=>"101000100",
  3138=>"110100000",
  3139=>"111110000",
  3140=>"011011011",
  3141=>"101100011",
  3142=>"010100001",
  3143=>"100011110",
  3144=>"110111000",
  3145=>"000010001",
  3146=>"110111110",
  3147=>"011101110",
  3148=>"000101011",
  3149=>"000000011",
  3150=>"100010001",
  3151=>"101001000",
  3152=>"001110100",
  3153=>"011110010",
  3154=>"111011000",
  3155=>"111011101",
  3156=>"010010111",
  3157=>"111111011",
  3158=>"000111011",
  3159=>"010011001",
  3160=>"010011100",
  3161=>"010000010",
  3162=>"000100001",
  3163=>"000111111",
  3164=>"111011111",
  3165=>"101101000",
  3166=>"000011011",
  3167=>"001101111",
  3168=>"001011011",
  3169=>"111101001",
  3170=>"110011010",
  3171=>"011001001",
  3172=>"000100011",
  3173=>"001000110",
  3174=>"011100010",
  3175=>"001110110",
  3176=>"000100010",
  3177=>"110000011",
  3178=>"000111101",
  3179=>"111100010",
  3180=>"000100111",
  3181=>"110001100",
  3182=>"110000000",
  3183=>"101101101",
  3184=>"011101011",
  3185=>"111101111",
  3186=>"001011100",
  3187=>"001110100",
  3188=>"001001101",
  3189=>"000000110",
  3190=>"100010101",
  3191=>"000001000",
  3192=>"000011101",
  3193=>"011011001",
  3194=>"111100100",
  3195=>"101100010",
  3196=>"100100110",
  3197=>"000111110",
  3198=>"100000001",
  3199=>"100101010",
  3200=>"001001000",
  3201=>"100101111",
  3202=>"011100000",
  3203=>"000110001",
  3204=>"000101111",
  3205=>"001000001",
  3206=>"001000010",
  3207=>"000001101",
  3208=>"011001100",
  3209=>"000001010",
  3210=>"001010101",
  3211=>"011000011",
  3212=>"010011100",
  3213=>"100110101",
  3214=>"111101100",
  3215=>"111001000",
  3216=>"100001111",
  3217=>"111010011",
  3218=>"011101000",
  3219=>"011110000",
  3220=>"000111000",
  3221=>"010101110",
  3222=>"001101010",
  3223=>"011001001",
  3224=>"110000010",
  3225=>"101011100",
  3226=>"111110010",
  3227=>"000001101",
  3228=>"100001001",
  3229=>"000011100",
  3230=>"000101101",
  3231=>"100001101",
  3232=>"100111101",
  3233=>"110100011",
  3234=>"100001100",
  3235=>"001011000",
  3236=>"000010100",
  3237=>"111001100",
  3238=>"001100001",
  3239=>"010010110",
  3240=>"101100110",
  3241=>"000110111",
  3242=>"010100001",
  3243=>"110101000",
  3244=>"011000100",
  3245=>"001101101",
  3246=>"101100010",
  3247=>"011011011",
  3248=>"000100001",
  3249=>"001000000",
  3250=>"110011000",
  3251=>"000001011",
  3252=>"111011100",
  3253=>"000001111",
  3254=>"000001001",
  3255=>"001110001",
  3256=>"001000100",
  3257=>"100100110",
  3258=>"010001101",
  3259=>"011111001",
  3260=>"110110101",
  3261=>"010000000",
  3262=>"100011001",
  3263=>"011100101",
  3264=>"101101101",
  3265=>"111111001",
  3266=>"011110001",
  3267=>"100101110",
  3268=>"011011100",
  3269=>"100010100",
  3270=>"111010001",
  3271=>"011000010",
  3272=>"100001100",
  3273=>"110001001",
  3274=>"011011101",
  3275=>"001100100",
  3276=>"101101001",
  3277=>"001111010",
  3278=>"111101011",
  3279=>"000000010",
  3280=>"100001000",
  3281=>"000101011",
  3282=>"010001000",
  3283=>"110010101",
  3284=>"011110100",
  3285=>"001001101",
  3286=>"111101100",
  3287=>"010101010",
  3288=>"100111101",
  3289=>"110011000",
  3290=>"101101011",
  3291=>"111001011",
  3292=>"011001010",
  3293=>"011111001",
  3294=>"111100010",
  3295=>"001100101",
  3296=>"010110001",
  3297=>"010101100",
  3298=>"010000111",
  3299=>"010001110",
  3300=>"111011110",
  3301=>"010100011",
  3302=>"101000010",
  3303=>"001111001",
  3304=>"111001100",
  3305=>"000110101",
  3306=>"010011001",
  3307=>"111100111",
  3308=>"001001111",
  3309=>"011010100",
  3310=>"000001100",
  3311=>"000000011",
  3312=>"010010000",
  3313=>"110101001",
  3314=>"001110100",
  3315=>"110101011",
  3316=>"100011110",
  3317=>"010011000",
  3318=>"111111011",
  3319=>"010011000",
  3320=>"100001111",
  3321=>"011001001",
  3322=>"100100001",
  3323=>"000101000",
  3324=>"110110110",
  3325=>"100000110",
  3326=>"011001100",
  3327=>"100100110",
  3328=>"010001001",
  3329=>"101000001",
  3330=>"100011101",
  3331=>"101001111",
  3332=>"010110001",
  3333=>"100100100",
  3334=>"110011101",
  3335=>"010110110",
  3336=>"000100010",
  3337=>"110111011",
  3338=>"110110011",
  3339=>"000000100",
  3340=>"100110010",
  3341=>"110011101",
  3342=>"101011101",
  3343=>"111000101",
  3344=>"011110100",
  3345=>"100101011",
  3346=>"001101100",
  3347=>"111111010",
  3348=>"001001001",
  3349=>"100010011",
  3350=>"101111001",
  3351=>"100011100",
  3352=>"100011100",
  3353=>"000100011",
  3354=>"001101001",
  3355=>"101111011",
  3356=>"110011001",
  3357=>"111000010",
  3358=>"010110010",
  3359=>"110000100",
  3360=>"010101100",
  3361=>"110110000",
  3362=>"001100110",
  3363=>"010111010",
  3364=>"101101100",
  3365=>"010001010",
  3366=>"000110000",
  3367=>"111110100",
  3368=>"000011101",
  3369=>"100101110",
  3370=>"011101001",
  3371=>"010000110",
  3372=>"000100001",
  3373=>"011000010",
  3374=>"011110100",
  3375=>"011000000",
  3376=>"100010100",
  3377=>"000000001",
  3378=>"000100110",
  3379=>"101011100",
  3380=>"111010001",
  3381=>"001010110",
  3382=>"110000011",
  3383=>"001111101",
  3384=>"000011001",
  3385=>"011110110",
  3386=>"100110110",
  3387=>"110111110",
  3388=>"001011110",
  3389=>"000100111",
  3390=>"000010101",
  3391=>"010011110",
  3392=>"111110100",
  3393=>"001100000",
  3394=>"101000111",
  3395=>"011100101",
  3396=>"110100100",
  3397=>"101100001",
  3398=>"100101000",
  3399=>"100010010",
  3400=>"100101101",
  3401=>"100100000",
  3402=>"011111011",
  3403=>"000001101",
  3404=>"011010011",
  3405=>"111000101",
  3406=>"110000100",
  3407=>"000000110",
  3408=>"011111100",
  3409=>"110100010",
  3410=>"001010111",
  3411=>"100010010",
  3412=>"000001010",
  3413=>"111001011",
  3414=>"000101101",
  3415=>"000110110",
  3416=>"000100100",
  3417=>"101000000",
  3418=>"101000001",
  3419=>"101000000",
  3420=>"010111010",
  3421=>"010110001",
  3422=>"110100001",
  3423=>"000110101",
  3424=>"011001110",
  3425=>"100111100",
  3426=>"010011001",
  3427=>"010101111",
  3428=>"010110110",
  3429=>"110101001",
  3430=>"001111100",
  3431=>"011000111",
  3432=>"111110010",
  3433=>"011101110",
  3434=>"011101111",
  3435=>"101000000",
  3436=>"001111001",
  3437=>"001111011",
  3438=>"100101000",
  3439=>"100101111",
  3440=>"100000100",
  3441=>"110001000",
  3442=>"001000100",
  3443=>"110000010",
  3444=>"010001110",
  3445=>"010111001",
  3446=>"011001110",
  3447=>"101110010",
  3448=>"001110010",
  3449=>"100101010",
  3450=>"110100000",
  3451=>"111000110",
  3452=>"010000011",
  3453=>"101101000",
  3454=>"111110010",
  3455=>"101101100",
  3456=>"110000001",
  3457=>"001101000",
  3458=>"110000000",
  3459=>"100010010",
  3460=>"110011000",
  3461=>"110011100",
  3462=>"100001100",
  3463=>"111111000",
  3464=>"101101010",
  3465=>"000011101",
  3466=>"011000000",
  3467=>"100001100",
  3468=>"000100011",
  3469=>"001110100",
  3470=>"101000100",
  3471=>"011000001",
  3472=>"101100001",
  3473=>"111110000",
  3474=>"110000100",
  3475=>"111010000",
  3476=>"001011000",
  3477=>"010101000",
  3478=>"001111100",
  3479=>"101011110",
  3480=>"111101011",
  3481=>"100110010",
  3482=>"011000111",
  3483=>"111010000",
  3484=>"101101001",
  3485=>"111010100",
  3486=>"101100000",
  3487=>"011111000",
  3488=>"101101100",
  3489=>"101001011",
  3490=>"110101110",
  3491=>"101000101",
  3492=>"001101000",
  3493=>"001011111",
  3494=>"010001111",
  3495=>"000111101",
  3496=>"111110101",
  3497=>"011101000",
  3498=>"001000101",
  3499=>"001010010",
  3500=>"001100100",
  3501=>"010110111",
  3502=>"111011011",
  3503=>"110001101",
  3504=>"010101010",
  3505=>"100011100",
  3506=>"100000100",
  3507=>"010001000",
  3508=>"011101111",
  3509=>"111100010",
  3510=>"011001010",
  3511=>"001001011",
  3512=>"011000101",
  3513=>"000100010",
  3514=>"001001110",
  3515=>"001001101",
  3516=>"000111100",
  3517=>"111010101",
  3518=>"111111101",
  3519=>"001000111",
  3520=>"000111000",
  3521=>"101001000",
  3522=>"110000010",
  3523=>"011110001",
  3524=>"111111111",
  3525=>"010011100",
  3526=>"100001000",
  3527=>"101100111",
  3528=>"101111111",
  3529=>"101101010",
  3530=>"100010111",
  3531=>"000011100",
  3532=>"000110111",
  3533=>"010000110",
  3534=>"001101011",
  3535=>"101001101",
  3536=>"010100010",
  3537=>"100010101",
  3538=>"111010010",
  3539=>"010111001",
  3540=>"001101001",
  3541=>"011010011",
  3542=>"101110111",
  3543=>"110101101",
  3544=>"001001010",
  3545=>"110001010",
  3546=>"111011111",
  3547=>"001001010",
  3548=>"100000101",
  3549=>"101000100",
  3550=>"100000011",
  3551=>"011110100",
  3552=>"010010111",
  3553=>"010100011",
  3554=>"110000010",
  3555=>"111101000",
  3556=>"111101101",
  3557=>"001111001",
  3558=>"011110010",
  3559=>"011000101",
  3560=>"011101110",
  3561=>"000100101",
  3562=>"111010101",
  3563=>"010010110",
  3564=>"101000000",
  3565=>"111010111",
  3566=>"111001000",
  3567=>"000100101",
  3568=>"011101010",
  3569=>"010011100",
  3570=>"100111101",
  3571=>"000111111",
  3572=>"110100100",
  3573=>"110110011",
  3574=>"001110100",
  3575=>"101111010",
  3576=>"010000000",
  3577=>"111100110",
  3578=>"011010010",
  3579=>"001000011",
  3580=>"100110110",
  3581=>"000000111",
  3582=>"111001100",
  3583=>"011011111",
  3584=>"000101000",
  3585=>"001101001",
  3586=>"000011111",
  3587=>"101110010",
  3588=>"010011111",
  3589=>"101001100",
  3590=>"100101111",
  3591=>"100000100",
  3592=>"001010100",
  3593=>"100011111",
  3594=>"011010110",
  3595=>"001010011",
  3596=>"010111001",
  3597=>"000110100",
  3598=>"010101011",
  3599=>"001001000",
  3600=>"101110100",
  3601=>"000101110",
  3602=>"101110010",
  3603=>"101000111",
  3604=>"110011000",
  3605=>"000001010",
  3606=>"001111100",
  3607=>"000100001",
  3608=>"001000110",
  3609=>"010000100",
  3610=>"010111011",
  3611=>"001001010",
  3612=>"010110100",
  3613=>"100000100",
  3614=>"010100001",
  3615=>"001100101",
  3616=>"110110011",
  3617=>"001100111",
  3618=>"001100000",
  3619=>"101110110",
  3620=>"001110100",
  3621=>"000100110",
  3622=>"111000110",
  3623=>"010010001",
  3624=>"000100100",
  3625=>"100011000",
  3626=>"001100000",
  3627=>"100111001",
  3628=>"010110000",
  3629=>"111111111",
  3630=>"000111010",
  3631=>"110010110",
  3632=>"110111001",
  3633=>"110110110",
  3634=>"011000100",
  3635=>"010011110",
  3636=>"011110100",
  3637=>"110000010",
  3638=>"011000001",
  3639=>"010000010",
  3640=>"010110011",
  3641=>"011011101",
  3642=>"010100010",
  3643=>"110101011",
  3644=>"100110011",
  3645=>"100001001",
  3646=>"110111001",
  3647=>"001101000",
  3648=>"011000010",
  3649=>"001010111",
  3650=>"001100110",
  3651=>"111111101",
  3652=>"111101001",
  3653=>"010110011",
  3654=>"100111111",
  3655=>"010111011",
  3656=>"010101011",
  3657=>"111011111",
  3658=>"111110110",
  3659=>"100101101",
  3660=>"101100011",
  3661=>"001100000",
  3662=>"000101010",
  3663=>"100001010",
  3664=>"001000010",
  3665=>"100000100",
  3666=>"000101010",
  3667=>"010000000",
  3668=>"100100100",
  3669=>"010101100",
  3670=>"101100011",
  3671=>"011000101",
  3672=>"111101011",
  3673=>"010010011",
  3674=>"100010101",
  3675=>"111011101",
  3676=>"011001100",
  3677=>"111101010",
  3678=>"101101001",
  3679=>"100011001",
  3680=>"110011000",
  3681=>"100000011",
  3682=>"111000010",
  3683=>"000000001",
  3684=>"010011101",
  3685=>"000100110",
  3686=>"011001001",
  3687=>"100010010",
  3688=>"000001001",
  3689=>"101001101",
  3690=>"111100000",
  3691=>"010011110",
  3692=>"000100011",
  3693=>"101010101",
  3694=>"100110000",
  3695=>"010011001",
  3696=>"101001101",
  3697=>"000001000",
  3698=>"111111010",
  3699=>"000011100",
  3700=>"001011110",
  3701=>"111010011",
  3702=>"000110000",
  3703=>"100110101",
  3704=>"101110011",
  3705=>"000001011",
  3706=>"100010010",
  3707=>"000000001",
  3708=>"111110010",
  3709=>"100000000",
  3710=>"100100010",
  3711=>"000001111",
  3712=>"011111000",
  3713=>"110011010",
  3714=>"010000011",
  3715=>"010010011",
  3716=>"000000010",
  3717=>"110111000",
  3718=>"100001100",
  3719=>"010001010",
  3720=>"011001111",
  3721=>"001100101",
  3722=>"000110010",
  3723=>"100101001",
  3724=>"110111111",
  3725=>"110111111",
  3726=>"111010111",
  3727=>"000100001",
  3728=>"100000100",
  3729=>"101010101",
  3730=>"011111111",
  3731=>"011100011",
  3732=>"010100010",
  3733=>"110111011",
  3734=>"110011010",
  3735=>"110100110",
  3736=>"000111111",
  3737=>"110101101",
  3738=>"110000010",
  3739=>"011101011",
  3740=>"100101111",
  3741=>"110101110",
  3742=>"010101001",
  3743=>"001111010",
  3744=>"101111111",
  3745=>"100100100",
  3746=>"000001101",
  3747=>"100110100",
  3748=>"101011100",
  3749=>"110001011",
  3750=>"011111111",
  3751=>"000000011",
  3752=>"110000101",
  3753=>"010010111",
  3754=>"110010000",
  3755=>"101001010",
  3756=>"100101001",
  3757=>"001000000",
  3758=>"011101010",
  3759=>"101011110",
  3760=>"111010000",
  3761=>"101101010",
  3762=>"001010101",
  3763=>"110101011",
  3764=>"011100001",
  3765=>"010010101",
  3766=>"011101111",
  3767=>"100110100",
  3768=>"011110111",
  3769=>"011011000",
  3770=>"101100001",
  3771=>"010111010",
  3772=>"110100100",
  3773=>"011010000",
  3774=>"001000000",
  3775=>"100011001",
  3776=>"110000101",
  3777=>"010111111",
  3778=>"001110100",
  3779=>"100000100",
  3780=>"100111101",
  3781=>"101111001",
  3782=>"101110101",
  3783=>"000101011",
  3784=>"111111000",
  3785=>"010101010",
  3786=>"001010010",
  3787=>"001110001",
  3788=>"110001111",
  3789=>"010101001",
  3790=>"001101001",
  3791=>"100000110",
  3792=>"001101000",
  3793=>"001011110",
  3794=>"100110001",
  3795=>"010101010",
  3796=>"100101011",
  3797=>"010001100",
  3798=>"111011001",
  3799=>"111001001",
  3800=>"000111010",
  3801=>"101000111",
  3802=>"010010011",
  3803=>"001100111",
  3804=>"011100101",
  3805=>"110001011",
  3806=>"111011110",
  3807=>"000000101",
  3808=>"000010000",
  3809=>"000000100",
  3810=>"110011010",
  3811=>"010100111",
  3812=>"110011110",
  3813=>"011001100",
  3814=>"010110111",
  3815=>"101101111",
  3816=>"001100101",
  3817=>"000111101",
  3818=>"101001010",
  3819=>"010101000",
  3820=>"000011101",
  3821=>"111011101",
  3822=>"000000001",
  3823=>"110001001",
  3824=>"011101000",
  3825=>"011000101",
  3826=>"000111000",
  3827=>"110000010",
  3828=>"011101000",
  3829=>"110110010",
  3830=>"000111101",
  3831=>"010011000",
  3832=>"100100111",
  3833=>"110011000",
  3834=>"001000111",
  3835=>"100110100",
  3836=>"000100000",
  3837=>"011111000",
  3838=>"110000110",
  3839=>"011011111",
  3840=>"100000110",
  3841=>"100111000",
  3842=>"111111001",
  3843=>"110110010",
  3844=>"110100100",
  3845=>"100100111",
  3846=>"000101101",
  3847=>"001111101",
  3848=>"001100011",
  3849=>"001011010",
  3850=>"110010100",
  3851=>"001010010",
  3852=>"110000010",
  3853=>"110111100",
  3854=>"011100100",
  3855=>"101001000",
  3856=>"101000000",
  3857=>"100110000",
  3858=>"100111111",
  3859=>"011110011",
  3860=>"011100101",
  3861=>"010110110",
  3862=>"001111000",
  3863=>"100111000",
  3864=>"101001100",
  3865=>"111111111",
  3866=>"000101011",
  3867=>"101011110",
  3868=>"000011111",
  3869=>"101111110",
  3870=>"010110101",
  3871=>"111111001",
  3872=>"001111011",
  3873=>"100110110",
  3874=>"000100100",
  3875=>"000000100",
  3876=>"001011111",
  3877=>"101000001",
  3878=>"110101110",
  3879=>"001011100",
  3880=>"110011011",
  3881=>"000010011",
  3882=>"100101100",
  3883=>"101010000",
  3884=>"111110000",
  3885=>"000010010",
  3886=>"111001101",
  3887=>"000011011",
  3888=>"011001111",
  3889=>"011100011",
  3890=>"000010010",
  3891=>"111001011",
  3892=>"111010000",
  3893=>"110001100",
  3894=>"001011000",
  3895=>"001000110",
  3896=>"101110100",
  3897=>"000001010",
  3898=>"010001001",
  3899=>"110100000",
  3900=>"110000011",
  3901=>"100000110",
  3902=>"000110011",
  3903=>"101111010",
  3904=>"101100001",
  3905=>"011011011",
  3906=>"101011111",
  3907=>"101100100",
  3908=>"100101011",
  3909=>"100101001",
  3910=>"011100100",
  3911=>"010110001",
  3912=>"111101010",
  3913=>"101100001",
  3914=>"010100101",
  3915=>"000000111",
  3916=>"011111000",
  3917=>"110011110",
  3918=>"100111111",
  3919=>"011101110",
  3920=>"111000110",
  3921=>"011001101",
  3922=>"010011111",
  3923=>"011000010",
  3924=>"101100001",
  3925=>"001000110",
  3926=>"101001010",
  3927=>"101111000",
  3928=>"001001011",
  3929=>"010101111",
  3930=>"111101111",
  3931=>"010100111",
  3932=>"000100010",
  3933=>"000011011",
  3934=>"111100111",
  3935=>"000001011",
  3936=>"111100110",
  3937=>"110101101",
  3938=>"100101011",
  3939=>"110101110",
  3940=>"111110111",
  3941=>"000110001",
  3942=>"000000110",
  3943=>"100100100",
  3944=>"101101111",
  3945=>"000001000",
  3946=>"000011011",
  3947=>"001101100",
  3948=>"011100000",
  3949=>"101001001",
  3950=>"111000000",
  3951=>"011010010",
  3952=>"010110011",
  3953=>"011000011",
  3954=>"111010000",
  3955=>"101011100",
  3956=>"000001000",
  3957=>"000011010",
  3958=>"101110100",
  3959=>"011101101",
  3960=>"000100111",
  3961=>"111111001",
  3962=>"101100011",
  3963=>"100000101",
  3964=>"000010110",
  3965=>"000011110",
  3966=>"010101101",
  3967=>"110010110",
  3968=>"111111001",
  3969=>"001101110",
  3970=>"011000001",
  3971=>"111111011",
  3972=>"000100010",
  3973=>"000001101",
  3974=>"110100011",
  3975=>"001101010",
  3976=>"001000100",
  3977=>"101100111",
  3978=>"110100001",
  3979=>"000000001",
  3980=>"000111101",
  3981=>"101001101",
  3982=>"011111010",
  3983=>"111100100",
  3984=>"101010101",
  3985=>"011111100",
  3986=>"100111100",
  3987=>"001111001",
  3988=>"011111010",
  3989=>"000001101",
  3990=>"010110100",
  3991=>"110011110",
  3992=>"101100010",
  3993=>"000110110",
  3994=>"000001111",
  3995=>"111001111",
  3996=>"001000111",
  3997=>"011101001",
  3998=>"000000110",
  3999=>"010011001",
  4000=>"011001101",
  4001=>"101011110",
  4002=>"111001100",
  4003=>"001000111",
  4004=>"010000000",
  4005=>"101100111",
  4006=>"001110010",
  4007=>"101100101",
  4008=>"000001010",
  4009=>"101000011",
  4010=>"110101111",
  4011=>"100101111",
  4012=>"111111111",
  4013=>"100111111",
  4014=>"111110111",
  4015=>"000100100",
  4016=>"010010000",
  4017=>"100101111",
  4018=>"001001010",
  4019=>"100101111",
  4020=>"110110010",
  4021=>"110010101",
  4022=>"110100101",
  4023=>"111111110",
  4024=>"000100100",
  4025=>"000001110",
  4026=>"011011011",
  4027=>"101101100",
  4028=>"101101101",
  4029=>"000100001",
  4030=>"010000010",
  4031=>"100000110",
  4032=>"000010111",
  4033=>"111111011",
  4034=>"101111011",
  4035=>"111111000",
  4036=>"011111110",
  4037=>"010011010",
  4038=>"110011110",
  4039=>"111001011",
  4040=>"100010010",
  4041=>"110001011",
  4042=>"011100110",
  4043=>"110001000",
  4044=>"010000010",
  4045=>"000101100",
  4046=>"111111111",
  4047=>"100111011",
  4048=>"000100000",
  4049=>"110010000",
  4050=>"111100001",
  4051=>"100010011",
  4052=>"101101000",
  4053=>"100000110",
  4054=>"010011101",
  4055=>"011101111",
  4056=>"100101001",
  4057=>"011000111",
  4058=>"011010010",
  4059=>"110101110",
  4060=>"101001000",
  4061=>"100011111",
  4062=>"111010110",
  4063=>"110010100",
  4064=>"101101100",
  4065=>"100011001",
  4066=>"000111101",
  4067=>"101010100",
  4068=>"101100011",
  4069=>"110110101",
  4070=>"011011111",
  4071=>"010101001",
  4072=>"100101111",
  4073=>"101101111",
  4074=>"000100011",
  4075=>"100010001",
  4076=>"011111011",
  4077=>"001110000",
  4078=>"110001000",
  4079=>"111111111",
  4080=>"000100101",
  4081=>"110001100",
  4082=>"110010100",
  4083=>"001001000",
  4084=>"111111101",
  4085=>"110100011",
  4086=>"000010100",
  4087=>"110010000",
  4088=>"100001100",
  4089=>"000111010",
  4090=>"010110001",
  4091=>"100101111",
  4092=>"111011000",
  4093=>"100110100",
  4094=>"100010100",
  4095=>"000101110",
  4096=>"011100000",
  4097=>"001000110",
  4098=>"010101011",
  4099=>"100011100",
  4100=>"101111001",
  4101=>"111111011",
  4102=>"000001010",
  4103=>"000101101",
  4104=>"011000110",
  4105=>"101010101",
  4106=>"000000100",
  4107=>"111000000",
  4108=>"110101000",
  4109=>"010001100",
  4110=>"001001101",
  4111=>"011001110",
  4112=>"100100000",
  4113=>"011010000",
  4114=>"100100100",
  4115=>"010111011",
  4116=>"010010000",
  4117=>"111000000",
  4118=>"111101010",
  4119=>"111001101",
  4120=>"011100111",
  4121=>"101111010",
  4122=>"010010001",
  4123=>"111100111",
  4124=>"111111000",
  4125=>"010011110",
  4126=>"100000111",
  4127=>"000010000",
  4128=>"010001110",
  4129=>"011101011",
  4130=>"000011111",
  4131=>"000000110",
  4132=>"000100001",
  4133=>"110101010",
  4134=>"110100101",
  4135=>"111001010",
  4136=>"111010101",
  4137=>"000110000",
  4138=>"011000110",
  4139=>"010100010",
  4140=>"101000000",
  4141=>"111000111",
  4142=>"011110011",
  4143=>"010001110",
  4144=>"001111001",
  4145=>"111101111",
  4146=>"000111010",
  4147=>"111011001",
  4148=>"101101111",
  4149=>"001110110",
  4150=>"101000000",
  4151=>"111100000",
  4152=>"000011011",
  4153=>"000101001",
  4154=>"010111001",
  4155=>"011001100",
  4156=>"001110000",
  4157=>"010001010",
  4158=>"100000100",
  4159=>"011010011",
  4160=>"101110111",
  4161=>"110111001",
  4162=>"010101001",
  4163=>"010000110",
  4164=>"001001010",
  4165=>"001110001",
  4166=>"101011111",
  4167=>"011010100",
  4168=>"100110000",
  4169=>"011101110",
  4170=>"000011110",
  4171=>"011000101",
  4172=>"010011111",
  4173=>"101000011",
  4174=>"011110001",
  4175=>"010111101",
  4176=>"010011010",
  4177=>"001000111",
  4178=>"011101101",
  4179=>"110100010",
  4180=>"101001000",
  4181=>"101101000",
  4182=>"000100011",
  4183=>"110011110",
  4184=>"101111110",
  4185=>"001001010",
  4186=>"101011111",
  4187=>"000000101",
  4188=>"111000100",
  4189=>"110111110",
  4190=>"000100011",
  4191=>"100101100",
  4192=>"101001000",
  4193=>"011101010",
  4194=>"001100100",
  4195=>"010101011",
  4196=>"111001001",
  4197=>"000101000",
  4198=>"010110000",
  4199=>"110011010",
  4200=>"100001011",
  4201=>"101011000",
  4202=>"001110100",
  4203=>"110101011",
  4204=>"111111011",
  4205=>"001000001",
  4206=>"100110011",
  4207=>"111111000",
  4208=>"001110111",
  4209=>"101111010",
  4210=>"010111110",
  4211=>"001010010",
  4212=>"000110111",
  4213=>"011111100",
  4214=>"101000001",
  4215=>"010011011",
  4216=>"100111000",
  4217=>"001101100",
  4218=>"101010100",
  4219=>"000100011",
  4220=>"110000000",
  4221=>"011000111",
  4222=>"010001001",
  4223=>"101101001",
  4224=>"110011110",
  4225=>"010101010",
  4226=>"100001001",
  4227=>"111110101",
  4228=>"111000101",
  4229=>"000100011",
  4230=>"000010111",
  4231=>"101010101",
  4232=>"010011010",
  4233=>"011001001",
  4234=>"000011100",
  4235=>"001101100",
  4236=>"111010010",
  4237=>"101100110",
  4238=>"100100001",
  4239=>"110010110",
  4240=>"000010100",
  4241=>"101010010",
  4242=>"101011110",
  4243=>"111100000",
  4244=>"011011111",
  4245=>"101011110",
  4246=>"000101101",
  4247=>"101101010",
  4248=>"000000111",
  4249=>"001011100",
  4250=>"110100100",
  4251=>"000101100",
  4252=>"001100010",
  4253=>"001010011",
  4254=>"001000001",
  4255=>"000001001",
  4256=>"000001101",
  4257=>"010011110",
  4258=>"010101100",
  4259=>"001010100",
  4260=>"001010010",
  4261=>"011011001",
  4262=>"000101000",
  4263=>"011001000",
  4264=>"110101101",
  4265=>"110000000",
  4266=>"101010011",
  4267=>"011111110",
  4268=>"100010011",
  4269=>"101000100",
  4270=>"011110100",
  4271=>"111111100",
  4272=>"001111110",
  4273=>"101100100",
  4274=>"110100011",
  4275=>"010110110",
  4276=>"101000011",
  4277=>"100101100",
  4278=>"000011011",
  4279=>"000001001",
  4280=>"111110101",
  4281=>"001100101",
  4282=>"111100010",
  4283=>"110110100",
  4284=>"011101011",
  4285=>"000000010",
  4286=>"011001100",
  4287=>"100001100",
  4288=>"001000110",
  4289=>"001000010",
  4290=>"011101110",
  4291=>"111101110",
  4292=>"100100111",
  4293=>"100101110",
  4294=>"001100011",
  4295=>"111101010",
  4296=>"000000001",
  4297=>"011001011",
  4298=>"101110110",
  4299=>"101100100",
  4300=>"000101010",
  4301=>"110100010",
  4302=>"001011110",
  4303=>"110111111",
  4304=>"110100110",
  4305=>"110110100",
  4306=>"100101101",
  4307=>"110101011",
  4308=>"011000100",
  4309=>"000101111",
  4310=>"101001011",
  4311=>"111100011",
  4312=>"100000111",
  4313=>"011111100",
  4314=>"101001011",
  4315=>"100101101",
  4316=>"110101111",
  4317=>"101101101",
  4318=>"001000110",
  4319=>"111000000",
  4320=>"000101010",
  4321=>"010001011",
  4322=>"010000100",
  4323=>"111011111",
  4324=>"011000100",
  4325=>"101111011",
  4326=>"001001100",
  4327=>"100010000",
  4328=>"011110000",
  4329=>"100000010",
  4330=>"101000111",
  4331=>"100001000",
  4332=>"001101101",
  4333=>"010101111",
  4334=>"100100001",
  4335=>"101000001",
  4336=>"110011010",
  4337=>"100000010",
  4338=>"110011001",
  4339=>"101001011",
  4340=>"010010001",
  4341=>"001111000",
  4342=>"101001001",
  4343=>"000010110",
  4344=>"101101000",
  4345=>"101010100",
  4346=>"110011110",
  4347=>"000000111",
  4348=>"101001111",
  4349=>"001011101",
  4350=>"101101100",
  4351=>"010111111",
  4352=>"000010110",
  4353=>"111011111",
  4354=>"111101100",
  4355=>"111100101",
  4356=>"000111011",
  4357=>"111010110",
  4358=>"100110010",
  4359=>"000111101",
  4360=>"011000100",
  4361=>"101010100",
  4362=>"001100001",
  4363=>"011011111",
  4364=>"001010011",
  4365=>"101110101",
  4366=>"011011010",
  4367=>"111111100",
  4368=>"000010010",
  4369=>"001100010",
  4370=>"001000010",
  4371=>"010100000",
  4372=>"100111000",
  4373=>"010000011",
  4374=>"100000010",
  4375=>"110000000",
  4376=>"011001011",
  4377=>"101001001",
  4378=>"001100000",
  4379=>"000001110",
  4380=>"111111011",
  4381=>"100100001",
  4382=>"110100001",
  4383=>"010010101",
  4384=>"111101000",
  4385=>"010111001",
  4386=>"010110011",
  4387=>"011110000",
  4388=>"111001010",
  4389=>"011000010",
  4390=>"000100111",
  4391=>"101101101",
  4392=>"001010011",
  4393=>"101011001",
  4394=>"011011001",
  4395=>"101100110",
  4396=>"001100101",
  4397=>"111011010",
  4398=>"011111110",
  4399=>"101110110",
  4400=>"000101010",
  4401=>"000110000",
  4402=>"001000011",
  4403=>"011111100",
  4404=>"001100111",
  4405=>"000000100",
  4406=>"000010100",
  4407=>"111111111",
  4408=>"110010111",
  4409=>"010001100",
  4410=>"100110000",
  4411=>"101010000",
  4412=>"000101000",
  4413=>"000011110",
  4414=>"100000110",
  4415=>"101111101",
  4416=>"110110100",
  4417=>"011111111",
  4418=>"010101011",
  4419=>"000111100",
  4420=>"000010000",
  4421=>"100110000",
  4422=>"111110010",
  4423=>"011010011",
  4424=>"001110100",
  4425=>"110101101",
  4426=>"001000010",
  4427=>"000100101",
  4428=>"110100101",
  4429=>"110011100",
  4430=>"001000010",
  4431=>"010010101",
  4432=>"010100110",
  4433=>"010011001",
  4434=>"001110001",
  4435=>"000001010",
  4436=>"111000100",
  4437=>"010101010",
  4438=>"101101111",
  4439=>"111110111",
  4440=>"001001111",
  4441=>"000111010",
  4442=>"001000100",
  4443=>"011110100",
  4444=>"010111001",
  4445=>"010001000",
  4446=>"100010111",
  4447=>"001100000",
  4448=>"111100010",
  4449=>"001001101",
  4450=>"100101011",
  4451=>"000110010",
  4452=>"111111111",
  4453=>"000010100",
  4454=>"010100000",
  4455=>"011101010",
  4456=>"110100100",
  4457=>"001000110",
  4458=>"001100110",
  4459=>"100111011",
  4460=>"010110001",
  4461=>"111001111",
  4462=>"111011011",
  4463=>"011000111",
  4464=>"001111000",
  4465=>"111111100",
  4466=>"010010100",
  4467=>"010101111",
  4468=>"111110110",
  4469=>"011101100",
  4470=>"001001101",
  4471=>"010110010",
  4472=>"101010100",
  4473=>"101001100",
  4474=>"100000111",
  4475=>"000110101",
  4476=>"010000010",
  4477=>"111001010",
  4478=>"001110001",
  4479=>"100001010",
  4480=>"110011111",
  4481=>"011000000",
  4482=>"001011001",
  4483=>"000100101",
  4484=>"011110111",
  4485=>"001001101",
  4486=>"011111001",
  4487=>"000001110",
  4488=>"001101010",
  4489=>"001010011",
  4490=>"110110101",
  4491=>"110011110",
  4492=>"010100000",
  4493=>"010000100",
  4494=>"000101001",
  4495=>"100010000",
  4496=>"101110011",
  4497=>"000111001",
  4498=>"010010110",
  4499=>"100001000",
  4500=>"110101011",
  4501=>"110101011",
  4502=>"100101110",
  4503=>"000000100",
  4504=>"100010010",
  4505=>"101001100",
  4506=>"100111001",
  4507=>"110110100",
  4508=>"111010111",
  4509=>"110011000",
  4510=>"111101101",
  4511=>"010001010",
  4512=>"010101000",
  4513=>"100001000",
  4514=>"000000111",
  4515=>"110111111",
  4516=>"111010001",
  4517=>"000111000",
  4518=>"001000100",
  4519=>"001011101",
  4520=>"011010000",
  4521=>"110111010",
  4522=>"101001000",
  4523=>"101110110",
  4524=>"101010110",
  4525=>"001100111",
  4526=>"111000001",
  4527=>"111111010",
  4528=>"100011100",
  4529=>"001110101",
  4530=>"101101000",
  4531=>"000101100",
  4532=>"111001111",
  4533=>"111111011",
  4534=>"110010000",
  4535=>"101101101",
  4536=>"011111100",
  4537=>"010110110",
  4538=>"000100101",
  4539=>"010100101",
  4540=>"100011101",
  4541=>"001001100",
  4542=>"111110010",
  4543=>"111010100",
  4544=>"101000101",
  4545=>"101011000",
  4546=>"110001111",
  4547=>"011001100",
  4548=>"111101100",
  4549=>"010111010",
  4550=>"101011011",
  4551=>"000000001",
  4552=>"111011000",
  4553=>"011110011",
  4554=>"001110110",
  4555=>"110010010",
  4556=>"101000001",
  4557=>"011010111",
  4558=>"100000101",
  4559=>"111110011",
  4560=>"111101101",
  4561=>"110011111",
  4562=>"101111111",
  4563=>"110010000",
  4564=>"101101111",
  4565=>"100110010",
  4566=>"011101000",
  4567=>"001101101",
  4568=>"000110010",
  4569=>"010110011",
  4570=>"111100101",
  4571=>"011000001",
  4572=>"001111101",
  4573=>"010010100",
  4574=>"010010110",
  4575=>"101110111",
  4576=>"000110011",
  4577=>"010001001",
  4578=>"011011010",
  4579=>"100110000",
  4580=>"111010010",
  4581=>"000110110",
  4582=>"110011010",
  4583=>"111000011",
  4584=>"001100000",
  4585=>"010001000",
  4586=>"000011110",
  4587=>"000110111",
  4588=>"000110111",
  4589=>"100011010",
  4590=>"010011011",
  4591=>"100111001",
  4592=>"000101100",
  4593=>"011111100",
  4594=>"011000001",
  4595=>"110011010",
  4596=>"100100101",
  4597=>"000111001",
  4598=>"110111001",
  4599=>"000001110",
  4600=>"101111100",
  4601=>"011011001",
  4602=>"001110010",
  4603=>"111010100",
  4604=>"001010010",
  4605=>"100001000",
  4606=>"000010011",
  4607=>"000000001",
  4608=>"101100010",
  4609=>"010000100",
  4610=>"010101110",
  4611=>"010011100",
  4612=>"100000110",
  4613=>"010010110",
  4614=>"011111011",
  4615=>"100000010",
  4616=>"000110110",
  4617=>"111010000",
  4618=>"111000111",
  4619=>"101000111",
  4620=>"010011011",
  4621=>"010110001",
  4622=>"110110101",
  4623=>"101001000",
  4624=>"010100011",
  4625=>"001001101",
  4626=>"010000110",
  4627=>"111101001",
  4628=>"000011010",
  4629=>"011010011",
  4630=>"010100001",
  4631=>"101011101",
  4632=>"101010010",
  4633=>"110111111",
  4634=>"111000011",
  4635=>"101100001",
  4636=>"110100000",
  4637=>"101010001",
  4638=>"001100110",
  4639=>"100100101",
  4640=>"101011101",
  4641=>"110010011",
  4642=>"001000000",
  4643=>"111011011",
  4644=>"011000010",
  4645=>"111010011",
  4646=>"010101000",
  4647=>"100011010",
  4648=>"001110000",
  4649=>"110011111",
  4650=>"011110010",
  4651=>"001010001",
  4652=>"110001011",
  4653=>"000010101",
  4654=>"101111111",
  4655=>"001010001",
  4656=>"000001000",
  4657=>"101000001",
  4658=>"001001001",
  4659=>"101010111",
  4660=>"000011001",
  4661=>"111101011",
  4662=>"000011000",
  4663=>"010110010",
  4664=>"110100101",
  4665=>"011011010",
  4666=>"110000100",
  4667=>"011111110",
  4668=>"010001111",
  4669=>"111111101",
  4670=>"110110100",
  4671=>"010100000",
  4672=>"011101101",
  4673=>"011100100",
  4674=>"001000100",
  4675=>"011110111",
  4676=>"000101000",
  4677=>"101011000",
  4678=>"101110000",
  4679=>"110010001",
  4680=>"000111101",
  4681=>"101000010",
  4682=>"110000001",
  4683=>"001001100",
  4684=>"010110010",
  4685=>"001010011",
  4686=>"110000010",
  4687=>"001001011",
  4688=>"101101111",
  4689=>"010100011",
  4690=>"001101110",
  4691=>"000001100",
  4692=>"000111001",
  4693=>"101111010",
  4694=>"000000010",
  4695=>"000000011",
  4696=>"100101010",
  4697=>"010010000",
  4698=>"011100000",
  4699=>"100101001",
  4700=>"101010100",
  4701=>"101100111",
  4702=>"011010101",
  4703=>"100101110",
  4704=>"001001111",
  4705=>"011111110",
  4706=>"010000000",
  4707=>"010000000",
  4708=>"000010010",
  4709=>"010101000",
  4710=>"011111111",
  4711=>"010111000",
  4712=>"110110000",
  4713=>"111011100",
  4714=>"101010111",
  4715=>"101100000",
  4716=>"101001100",
  4717=>"001100110",
  4718=>"110111111",
  4719=>"001101101",
  4720=>"000110101",
  4721=>"001101110",
  4722=>"111010000",
  4723=>"001101010",
  4724=>"010011001",
  4725=>"111110101",
  4726=>"000010101",
  4727=>"001010100",
  4728=>"100000001",
  4729=>"010011101",
  4730=>"010111000",
  4731=>"010101011",
  4732=>"011001011",
  4733=>"101101101",
  4734=>"101110011",
  4735=>"110110000",
  4736=>"000100111",
  4737=>"111101001",
  4738=>"100001111",
  4739=>"101000000",
  4740=>"001101101",
  4741=>"000010101",
  4742=>"001000001",
  4743=>"011010011",
  4744=>"000011011",
  4745=>"010110100",
  4746=>"100111000",
  4747=>"111010111",
  4748=>"011000001",
  4749=>"010010101",
  4750=>"001100100",
  4751=>"111111000",
  4752=>"111010001",
  4753=>"110101000",
  4754=>"111101101",
  4755=>"101110000",
  4756=>"010000001",
  4757=>"111111010",
  4758=>"100111111",
  4759=>"011000111",
  4760=>"001100001",
  4761=>"110111001",
  4762=>"110000011",
  4763=>"000011101",
  4764=>"010010101",
  4765=>"010100110",
  4766=>"011101000",
  4767=>"100000101",
  4768=>"110101010",
  4769=>"010001011",
  4770=>"000010010",
  4771=>"001001101",
  4772=>"111011001",
  4773=>"111111101",
  4774=>"100010100",
  4775=>"110111011",
  4776=>"010011101",
  4777=>"100011101",
  4778=>"000110101",
  4779=>"111010011",
  4780=>"010000110",
  4781=>"000010000",
  4782=>"010000111",
  4783=>"111100001",
  4784=>"101000110",
  4785=>"010000100",
  4786=>"101101000",
  4787=>"001001100",
  4788=>"001001000",
  4789=>"111001000",
  4790=>"010010111",
  4791=>"010110010",
  4792=>"001000001",
  4793=>"111011010",
  4794=>"110001110",
  4795=>"101100110",
  4796=>"001110100",
  4797=>"001111101",
  4798=>"111001100",
  4799=>"100000100",
  4800=>"000001000",
  4801=>"101111000",
  4802=>"011111110",
  4803=>"011011010",
  4804=>"000110100",
  4805=>"010010100",
  4806=>"110101010",
  4807=>"110110010",
  4808=>"101100011",
  4809=>"011001100",
  4810=>"111001010",
  4811=>"111100001",
  4812=>"111010101",
  4813=>"000100111",
  4814=>"000111110",
  4815=>"101010111",
  4816=>"000000110",
  4817=>"101011101",
  4818=>"111111000",
  4819=>"001000110",
  4820=>"001000111",
  4821=>"101111011",
  4822=>"110001110",
  4823=>"001100111",
  4824=>"010011000",
  4825=>"100000100",
  4826=>"101001100",
  4827=>"011111010",
  4828=>"111011010",
  4829=>"101111100",
  4830=>"010110111",
  4831=>"111110000",
  4832=>"110010110",
  4833=>"100101001",
  4834=>"000010101",
  4835=>"010100011",
  4836=>"110111010",
  4837=>"110100101",
  4838=>"101100101",
  4839=>"100111010",
  4840=>"011011001",
  4841=>"100101001",
  4842=>"011110001",
  4843=>"011011010",
  4844=>"001010010",
  4845=>"100110111",
  4846=>"100101010",
  4847=>"000001010",
  4848=>"011110010",
  4849=>"000110011",
  4850=>"100001010",
  4851=>"011001010",
  4852=>"011100101",
  4853=>"100001100",
  4854=>"001001000",
  4855=>"100010111",
  4856=>"101101110",
  4857=>"001111101",
  4858=>"110101000",
  4859=>"001000010",
  4860=>"000010111",
  4861=>"000011011",
  4862=>"110010010",
  4863=>"010010010",
  4864=>"000010100",
  4865=>"001000010",
  4866=>"001010011",
  4867=>"010001111",
  4868=>"001001011",
  4869=>"001111101",
  4870=>"111010100",
  4871=>"101001100",
  4872=>"101110111",
  4873=>"100011101",
  4874=>"110010110",
  4875=>"100011111",
  4876=>"110110001",
  4877=>"010110110",
  4878=>"111100011",
  4879=>"101001000",
  4880=>"100100100",
  4881=>"111010001",
  4882=>"011011010",
  4883=>"100001111",
  4884=>"100101101",
  4885=>"010001100",
  4886=>"110101000",
  4887=>"111110110",
  4888=>"100111101",
  4889=>"000000000",
  4890=>"101001111",
  4891=>"100000101",
  4892=>"010111111",
  4893=>"110011101",
  4894=>"101000011",
  4895=>"101011110",
  4896=>"011110111",
  4897=>"010010111",
  4898=>"010100111",
  4899=>"111111100",
  4900=>"100100111",
  4901=>"000100101",
  4902=>"111011100",
  4903=>"011011000",
  4904=>"111100000",
  4905=>"000101010",
  4906=>"001111010",
  4907=>"001001000",
  4908=>"111111010",
  4909=>"000001111",
  4910=>"101001111",
  4911=>"101010110",
  4912=>"100100001",
  4913=>"011010111",
  4914=>"110010010",
  4915=>"011101101",
  4916=>"010101000",
  4917=>"101110101",
  4918=>"000000110",
  4919=>"111101101",
  4920=>"011011111",
  4921=>"100100011",
  4922=>"000100110",
  4923=>"100011010",
  4924=>"010111100",
  4925=>"001110011",
  4926=>"111101011",
  4927=>"111010011",
  4928=>"111100000",
  4929=>"100011000",
  4930=>"101001110",
  4931=>"010100100",
  4932=>"101001001",
  4933=>"011010010",
  4934=>"111011101",
  4935=>"111010101",
  4936=>"101011010",
  4937=>"100111110",
  4938=>"011000000",
  4939=>"100001110",
  4940=>"110000011",
  4941=>"001010110",
  4942=>"010101111",
  4943=>"001101111",
  4944=>"010010101",
  4945=>"001100101",
  4946=>"111101110",
  4947=>"011001101",
  4948=>"101100111",
  4949=>"111111011",
  4950=>"011001001",
  4951=>"111101000",
  4952=>"111001000",
  4953=>"111001011",
  4954=>"101000011",
  4955=>"101001001",
  4956=>"100000110",
  4957=>"000000100",
  4958=>"010110110",
  4959=>"001110011",
  4960=>"100010100",
  4961=>"010010000",
  4962=>"000101000",
  4963=>"011100100",
  4964=>"010100001",
  4965=>"000011100",
  4966=>"010101100",
  4967=>"010100000",
  4968=>"001010111",
  4969=>"100111100",
  4970=>"100101000",
  4971=>"010111100",
  4972=>"101101100",
  4973=>"101110011",
  4974=>"110001011",
  4975=>"011001100",
  4976=>"101001011",
  4977=>"010110000",
  4978=>"110011110",
  4979=>"110101001",
  4980=>"000111011",
  4981=>"011010010",
  4982=>"011000101",
  4983=>"111010111",
  4984=>"011100001",
  4985=>"101100110",
  4986=>"000000101",
  4987=>"111111111",
  4988=>"100000110",
  4989=>"010001011",
  4990=>"010001101",
  4991=>"000001001",
  4992=>"001111001",
  4993=>"000000001",
  4994=>"001100011",
  4995=>"000100010",
  4996=>"000100111",
  4997=>"111011010",
  4998=>"101101101",
  4999=>"100110001",
  5000=>"000010001",
  5001=>"101001011",
  5002=>"101010111",
  5003=>"011101000",
  5004=>"111001110",
  5005=>"111011011",
  5006=>"100100101",
  5007=>"110110001",
  5008=>"011011000",
  5009=>"111010100",
  5010=>"100111101",
  5011=>"011101110",
  5012=>"000101111",
  5013=>"111111010",
  5014=>"111101111",
  5015=>"101001110",
  5016=>"101010011",
  5017=>"110010001",
  5018=>"000000011",
  5019=>"000011110",
  5020=>"010111001",
  5021=>"111010111",
  5022=>"100000110",
  5023=>"111011010",
  5024=>"000000011",
  5025=>"001100011",
  5026=>"110001011",
  5027=>"100000110",
  5028=>"111000000",
  5029=>"100110001",
  5030=>"110110011",
  5031=>"110100000",
  5032=>"100011110",
  5033=>"111011110",
  5034=>"010111000",
  5035=>"011001011",
  5036=>"011101000",
  5037=>"001101000",
  5038=>"000010111",
  5039=>"100010101",
  5040=>"010101011",
  5041=>"011110001",
  5042=>"101011100",
  5043=>"011001011",
  5044=>"100110110",
  5045=>"110000110",
  5046=>"110010000",
  5047=>"110111011",
  5048=>"110100010",
  5049=>"110111001",
  5050=>"001111111",
  5051=>"011101101",
  5052=>"110100101",
  5053=>"101000001",
  5054=>"111000010",
  5055=>"010010101",
  5056=>"001010001",
  5057=>"000000000",
  5058=>"111100000",
  5059=>"100100100",
  5060=>"101101011",
  5061=>"110001100",
  5062=>"011001101",
  5063=>"011010101",
  5064=>"001011101",
  5065=>"001101001",
  5066=>"100101100",
  5067=>"101001011",
  5068=>"000100110",
  5069=>"111111001",
  5070=>"000101010",
  5071=>"010110000",
  5072=>"010111111",
  5073=>"010000110",
  5074=>"110111111",
  5075=>"101001111",
  5076=>"000100010",
  5077=>"001111111",
  5078=>"101001000",
  5079=>"100010101",
  5080=>"110001000",
  5081=>"101111010",
  5082=>"100011001",
  5083=>"000011101",
  5084=>"001001000",
  5085=>"011011111",
  5086=>"100000010",
  5087=>"000100110",
  5088=>"011001101",
  5089=>"101011101",
  5090=>"010010111",
  5091=>"001101001",
  5092=>"000010000",
  5093=>"010101011",
  5094=>"100001011",
  5095=>"101000110",
  5096=>"100000000",
  5097=>"011100011",
  5098=>"010001010",
  5099=>"101110001",
  5100=>"011110110",
  5101=>"110001010",
  5102=>"111101101",
  5103=>"100000110",
  5104=>"101000001",
  5105=>"010010011",
  5106=>"001000010",
  5107=>"110111011",
  5108=>"100100011",
  5109=>"010000100",
  5110=>"110100111",
  5111=>"101101110",
  5112=>"011101101",
  5113=>"010110101",
  5114=>"111011001",
  5115=>"110000010",
  5116=>"100111111",
  5117=>"001011100",
  5118=>"011101010",
  5119=>"010011000",
  5120=>"001110111",
  5121=>"100101001",
  5122=>"101001000",
  5123=>"100011110",
  5124=>"101100000",
  5125=>"010101101",
  5126=>"001101100",
  5127=>"001101101",
  5128=>"001110000",
  5129=>"111110000",
  5130=>"100011111",
  5131=>"001010111",
  5132=>"100101011",
  5133=>"000000101",
  5134=>"011010101",
  5135=>"001000011",
  5136=>"110110110",
  5137=>"110000101",
  5138=>"100100101",
  5139=>"100001010",
  5140=>"111000110",
  5141=>"100100101",
  5142=>"010111000",
  5143=>"000101001",
  5144=>"010110101",
  5145=>"111111110",
  5146=>"111110100",
  5147=>"101000111",
  5148=>"110100111",
  5149=>"010000100",
  5150=>"000111010",
  5151=>"110011100",
  5152=>"110100001",
  5153=>"111110011",
  5154=>"111011110",
  5155=>"011111111",
  5156=>"010101100",
  5157=>"101011000",
  5158=>"001111000",
  5159=>"010010111",
  5160=>"011010001",
  5161=>"000111100",
  5162=>"100001111",
  5163=>"011011000",
  5164=>"011010011",
  5165=>"001011100",
  5166=>"010000001",
  5167=>"100011110",
  5168=>"110101000",
  5169=>"010110110",
  5170=>"011111111",
  5171=>"111100010",
  5172=>"101011111",
  5173=>"111011010",
  5174=>"111001101",
  5175=>"101101000",
  5176=>"010111111",
  5177=>"011111011",
  5178=>"111011010",
  5179=>"001000001",
  5180=>"111010101",
  5181=>"100110100",
  5182=>"001101110",
  5183=>"111110011",
  5184=>"101110101",
  5185=>"111111111",
  5186=>"101001110",
  5187=>"101011001",
  5188=>"011101101",
  5189=>"100000000",
  5190=>"011000001",
  5191=>"111111111",
  5192=>"111000010",
  5193=>"010000000",
  5194=>"011010111",
  5195=>"111010010",
  5196=>"010010101",
  5197=>"100100110",
  5198=>"100011001",
  5199=>"000101011",
  5200=>"111101100",
  5201=>"011110000",
  5202=>"100011010",
  5203=>"101110111",
  5204=>"011000111",
  5205=>"001100100",
  5206=>"100100001",
  5207=>"111010100",
  5208=>"000000011",
  5209=>"011000000",
  5210=>"110110110",
  5211=>"011111101",
  5212=>"011110111",
  5213=>"111011100",
  5214=>"000101111",
  5215=>"101101000",
  5216=>"111110110",
  5217=>"001101111",
  5218=>"100000000",
  5219=>"101111101",
  5220=>"111011110",
  5221=>"011110010",
  5222=>"011111010",
  5223=>"111111101",
  5224=>"101110111",
  5225=>"110100101",
  5226=>"111110111",
  5227=>"010001101",
  5228=>"011010111",
  5229=>"111000111",
  5230=>"011100011",
  5231=>"001111010",
  5232=>"111111111",
  5233=>"101000101",
  5234=>"000010101",
  5235=>"000000001",
  5236=>"100110011",
  5237=>"111000101",
  5238=>"000101011",
  5239=>"000000011",
  5240=>"000110100",
  5241=>"110100001",
  5242=>"111000110",
  5243=>"100100100",
  5244=>"111011111",
  5245=>"110100101",
  5246=>"111011000",
  5247=>"100000101",
  5248=>"010111110",
  5249=>"100110001",
  5250=>"011101100",
  5251=>"111110100",
  5252=>"111011011",
  5253=>"011011001",
  5254=>"010000000",
  5255=>"101110000",
  5256=>"001111101",
  5257=>"101001101",
  5258=>"111001111",
  5259=>"111000110",
  5260=>"110000001",
  5261=>"011100011",
  5262=>"010110110",
  5263=>"010011100",
  5264=>"000100110",
  5265=>"000110100",
  5266=>"110100011",
  5267=>"101100001",
  5268=>"001001010",
  5269=>"011100100",
  5270=>"101001010",
  5271=>"101111011",
  5272=>"111101110",
  5273=>"000001010",
  5274=>"000001010",
  5275=>"101100011",
  5276=>"111010000",
  5277=>"011110101",
  5278=>"100010011",
  5279=>"110010010",
  5280=>"100001011",
  5281=>"011111101",
  5282=>"010101011",
  5283=>"000000100",
  5284=>"100010101",
  5285=>"100000011",
  5286=>"000101101",
  5287=>"001011110",
  5288=>"111111110",
  5289=>"000010101",
  5290=>"001100111",
  5291=>"100011001",
  5292=>"001001111",
  5293=>"101001110",
  5294=>"111111011",
  5295=>"111101000",
  5296=>"011111100",
  5297=>"111100010",
  5298=>"011111101",
  5299=>"111001111",
  5300=>"100011000",
  5301=>"010010001",
  5302=>"001000000",
  5303=>"001110000",
  5304=>"011110111",
  5305=>"111111111",
  5306=>"000000010",
  5307=>"100101010",
  5308=>"000011101",
  5309=>"101101100",
  5310=>"010010001",
  5311=>"010101100",
  5312=>"101001000",
  5313=>"001001100",
  5314=>"011101110",
  5315=>"010101010",
  5316=>"010100111",
  5317=>"001101001",
  5318=>"111010100",
  5319=>"010100110",
  5320=>"000101111",
  5321=>"000011001",
  5322=>"010110101",
  5323=>"100110010",
  5324=>"101111101",
  5325=>"101010100",
  5326=>"101100111",
  5327=>"000001011",
  5328=>"011111000",
  5329=>"101011101",
  5330=>"111101010",
  5331=>"010110111",
  5332=>"000010110",
  5333=>"110110011",
  5334=>"010011101",
  5335=>"000001101",
  5336=>"111111111",
  5337=>"000110110",
  5338=>"111011111",
  5339=>"000111011",
  5340=>"111010000",
  5341=>"100111001",
  5342=>"111111011",
  5343=>"100010111",
  5344=>"101100111",
  5345=>"001101111",
  5346=>"000001000",
  5347=>"111111010",
  5348=>"000010000",
  5349=>"110000100",
  5350=>"011101111",
  5351=>"110010000",
  5352=>"101100000",
  5353=>"010111101",
  5354=>"000001001",
  5355=>"111111111",
  5356=>"111001101",
  5357=>"110001101",
  5358=>"110111101",
  5359=>"110111110",
  5360=>"100011101",
  5361=>"110001001",
  5362=>"111011000",
  5363=>"000011101",
  5364=>"001000001",
  5365=>"101001100",
  5366=>"111111011",
  5367=>"111011110",
  5368=>"111010100",
  5369=>"111100011",
  5370=>"001110111",
  5371=>"110100101",
  5372=>"101111111",
  5373=>"101110011",
  5374=>"010111001",
  5375=>"011111101",
  5376=>"100110101",
  5377=>"001000001",
  5378=>"001101110",
  5379=>"111000101",
  5380=>"111101000",
  5381=>"111010011",
  5382=>"100111010",
  5383=>"000001101",
  5384=>"110101000",
  5385=>"111011101",
  5386=>"001110010",
  5387=>"001000000",
  5388=>"011100010",
  5389=>"000011110",
  5390=>"111000100",
  5391=>"111010101",
  5392=>"010010110",
  5393=>"011001001",
  5394=>"100001001",
  5395=>"001000010",
  5396=>"100011010",
  5397=>"110101001",
  5398=>"100010001",
  5399=>"110110011",
  5400=>"110000100",
  5401=>"110100110",
  5402=>"110101110",
  5403=>"010011111",
  5404=>"111100010",
  5405=>"100101111",
  5406=>"101001001",
  5407=>"111111011",
  5408=>"111011011",
  5409=>"110110111",
  5410=>"111011101",
  5411=>"100110010",
  5412=>"110110111",
  5413=>"111100000",
  5414=>"000010010",
  5415=>"000100011",
  5416=>"111001100",
  5417=>"011100100",
  5418=>"000100111",
  5419=>"100111100",
  5420=>"010101011",
  5421=>"101110000",
  5422=>"111001100",
  5423=>"000010001",
  5424=>"010001011",
  5425=>"100111010",
  5426=>"101001010",
  5427=>"111111111",
  5428=>"001011111",
  5429=>"110111010",
  5430=>"000000000",
  5431=>"110000011",
  5432=>"101111110",
  5433=>"100101101",
  5434=>"001000001",
  5435=>"110111110",
  5436=>"010011011",
  5437=>"101001011",
  5438=>"010111000",
  5439=>"100001011",
  5440=>"100000011",
  5441=>"001101001",
  5442=>"101000000",
  5443=>"010000000",
  5444=>"000000100",
  5445=>"100001010",
  5446=>"100110110",
  5447=>"010111110",
  5448=>"100000010",
  5449=>"110110001",
  5450=>"001001000",
  5451=>"111011111",
  5452=>"100011010",
  5453=>"111010101",
  5454=>"011111111",
  5455=>"100011001",
  5456=>"100010100",
  5457=>"101110001",
  5458=>"011111001",
  5459=>"101100100",
  5460=>"011111011",
  5461=>"011001100",
  5462=>"111101101",
  5463=>"100000001",
  5464=>"101111111",
  5465=>"111111111",
  5466=>"001010001",
  5467=>"011010111",
  5468=>"101000001",
  5469=>"111000000",
  5470=>"110001000",
  5471=>"011111000",
  5472=>"101101011",
  5473=>"100100010",
  5474=>"100010000",
  5475=>"101111110",
  5476=>"110110100",
  5477=>"101000111",
  5478=>"111011110",
  5479=>"111001010",
  5480=>"000101111",
  5481=>"101111000",
  5482=>"111111111",
  5483=>"101011000",
  5484=>"101101011",
  5485=>"100001000",
  5486=>"111101011",
  5487=>"110010100",
  5488=>"110101110",
  5489=>"011101001",
  5490=>"000010001",
  5491=>"110011000",
  5492=>"011001111",
  5493=>"101101111",
  5494=>"101111011",
  5495=>"000000010",
  5496=>"110000001",
  5497=>"010010011",
  5498=>"111100101",
  5499=>"011111111",
  5500=>"000110010",
  5501=>"111011001",
  5502=>"000001101",
  5503=>"011011100",
  5504=>"111111101",
  5505=>"010111110",
  5506=>"100110011",
  5507=>"100010000",
  5508=>"110011110",
  5509=>"010001010",
  5510=>"000000000",
  5511=>"001000010",
  5512=>"110111110",
  5513=>"000110000",
  5514=>"011110111",
  5515=>"011100101",
  5516=>"111100110",
  5517=>"001111111",
  5518=>"111000111",
  5519=>"110001001",
  5520=>"001101010",
  5521=>"111111010",
  5522=>"011100111",
  5523=>"010000011",
  5524=>"011001110",
  5525=>"010101010",
  5526=>"111101000",
  5527=>"011001101",
  5528=>"101011111",
  5529=>"101111111",
  5530=>"111111111",
  5531=>"010111110",
  5532=>"001100011",
  5533=>"101000010",
  5534=>"001101000",
  5535=>"011010000",
  5536=>"110001011",
  5537=>"000101000",
  5538=>"011110111",
  5539=>"110011000",
  5540=>"001000110",
  5541=>"111111111",
  5542=>"011101001",
  5543=>"110011111",
  5544=>"111011010",
  5545=>"000100001",
  5546=>"111110110",
  5547=>"010101011",
  5548=>"100011010",
  5549=>"110000010",
  5550=>"111100110",
  5551=>"110110010",
  5552=>"000101001",
  5553=>"011100000",
  5554=>"010010000",
  5555=>"110100010",
  5556=>"101101001",
  5557=>"001101000",
  5558=>"111110111",
  5559=>"111011000",
  5560=>"100111010",
  5561=>"111110011",
  5562=>"111111110",
  5563=>"011011101",
  5564=>"001000011",
  5565=>"001001001",
  5566=>"111110001",
  5567=>"011110001",
  5568=>"101111110",
  5569=>"011101100",
  5570=>"000110111",
  5571=>"111110010",
  5572=>"111110010",
  5573=>"110001000",
  5574=>"100101110",
  5575=>"111111111",
  5576=>"110001000",
  5577=>"101011101",
  5578=>"110110111",
  5579=>"000011000",
  5580=>"010101010",
  5581=>"101101100",
  5582=>"111111111",
  5583=>"111100111",
  5584=>"010111001",
  5585=>"011111011",
  5586=>"110110010",
  5587=>"110110001",
  5588=>"011011000",
  5589=>"110111101",
  5590=>"011000111",
  5591=>"111000010",
  5592=>"111111111",
  5593=>"011010101",
  5594=>"110010011",
  5595=>"101101011",
  5596=>"001110110",
  5597=>"101000110",
  5598=>"110110001",
  5599=>"000110001",
  5600=>"111101010",
  5601=>"101101010",
  5602=>"000101010",
  5603=>"001110011",
  5604=>"010000001",
  5605=>"100000101",
  5606=>"111111111",
  5607=>"101110111",
  5608=>"101101000",
  5609=>"110001100",
  5610=>"111111100",
  5611=>"100000100",
  5612=>"010101010",
  5613=>"010111000",
  5614=>"111111111",
  5615=>"100011110",
  5616=>"111101100",
  5617=>"000100101",
  5618=>"110010000",
  5619=>"111101110",
  5620=>"010101110",
  5621=>"011110000",
  5622=>"000011011",
  5623=>"111111000",
  5624=>"000011111",
  5625=>"111101101",
  5626=>"111010010",
  5627=>"100001111",
  5628=>"100010010",
  5629=>"001001100",
  5630=>"110111011",
  5631=>"001101111",
  5632=>"010100010",
  5633=>"000101010",
  5634=>"001100100",
  5635=>"110101010",
  5636=>"001001100",
  5637=>"101100101",
  5638=>"000100111",
  5639=>"110110001",
  5640=>"111111100",
  5641=>"100100000",
  5642=>"110001100",
  5643=>"111111110",
  5644=>"111011000",
  5645=>"110001010",
  5646=>"111110111",
  5647=>"111101111",
  5648=>"011001101",
  5649=>"111110011",
  5650=>"111000100",
  5651=>"101001010",
  5652=>"111101101",
  5653=>"100100100",
  5654=>"111010000",
  5655=>"110101000",
  5656=>"000111111",
  5657=>"101101000",
  5658=>"111101101",
  5659=>"010010101",
  5660=>"110110000",
  5661=>"111111101",
  5662=>"101111000",
  5663=>"000110100",
  5664=>"000110010",
  5665=>"110111111",
  5666=>"111111000",
  5667=>"110101111",
  5668=>"111111010",
  5669=>"011100110",
  5670=>"000010000",
  5671=>"010110110",
  5672=>"011001111",
  5673=>"101000111",
  5674=>"111111100",
  5675=>"111111001",
  5676=>"010011100",
  5677=>"111111110",
  5678=>"000111101",
  5679=>"111001100",
  5680=>"001000011",
  5681=>"100111100",
  5682=>"101011011",
  5683=>"001110000",
  5684=>"101010110",
  5685=>"010111101",
  5686=>"000111101",
  5687=>"111110110",
  5688=>"111011100",
  5689=>"010001010",
  5690=>"110111111",
  5691=>"101000101",
  5692=>"111110111",
  5693=>"110110001",
  5694=>"110111111",
  5695=>"010100011",
  5696=>"110000101",
  5697=>"101101010",
  5698=>"110110110",
  5699=>"100111000",
  5700=>"110011101",
  5701=>"101000001",
  5702=>"111111110",
  5703=>"101111110",
  5704=>"110100000",
  5705=>"011000110",
  5706=>"011011010",
  5707=>"111100000",
  5708=>"010111001",
  5709=>"111110010",
  5710=>"010001010",
  5711=>"101110110",
  5712=>"110110000",
  5713=>"001110111",
  5714=>"101111000",
  5715=>"001111111",
  5716=>"110011101",
  5717=>"111111111",
  5718=>"011001111",
  5719=>"100001001",
  5720=>"001011111",
  5721=>"110001100",
  5722=>"011110001",
  5723=>"111111010",
  5724=>"010110100",
  5725=>"111110111",
  5726=>"111111000",
  5727=>"000000000",
  5728=>"000001111",
  5729=>"000101100",
  5730=>"010111111",
  5731=>"010000001",
  5732=>"100011101",
  5733=>"110001110",
  5734=>"010111110",
  5735=>"101011000",
  5736=>"110111110",
  5737=>"001111010",
  5738=>"100000001",
  5739=>"110100100",
  5740=>"111110111",
  5741=>"011010010",
  5742=>"010010001",
  5743=>"001101011",
  5744=>"110111011",
  5745=>"101110101",
  5746=>"010100010",
  5747=>"010101111",
  5748=>"110000100",
  5749=>"110101010",
  5750=>"000000001",
  5751=>"100100011",
  5752=>"110110000",
  5753=>"101010100",
  5754=>"111110000",
  5755=>"111001100",
  5756=>"101101111",
  5757=>"111011000",
  5758=>"001010100",
  5759=>"011001111",
  5760=>"110011011",
  5761=>"110110000",
  5762=>"111100010",
  5763=>"110110101",
  5764=>"110001011",
  5765=>"111111010",
  5766=>"101111110",
  5767=>"000110011",
  5768=>"110101001",
  5769=>"011001000",
  5770=>"000010110",
  5771=>"010010001",
  5772=>"110111000",
  5773=>"000111001",
  5774=>"001101000",
  5775=>"111011000",
  5776=>"001011011",
  5777=>"010110000",
  5778=>"001011000",
  5779=>"101000101",
  5780=>"111100011",
  5781=>"000101110",
  5782=>"111101100",
  5783=>"101111101",
  5784=>"101110111",
  5785=>"110000100",
  5786=>"111011011",
  5787=>"001100110",
  5788=>"010111011",
  5789=>"010101010",
  5790=>"111111011",
  5791=>"001100101",
  5792=>"100101101",
  5793=>"010000011",
  5794=>"101011111",
  5795=>"001111000",
  5796=>"110101110",
  5797=>"010010001",
  5798=>"001011010",
  5799=>"011011111",
  5800=>"100110111",
  5801=>"110110111",
  5802=>"111110011",
  5803=>"100110111",
  5804=>"111111101",
  5805=>"100110110",
  5806=>"111110010",
  5807=>"000110011",
  5808=>"111101111",
  5809=>"011001011",
  5810=>"000101100",
  5811=>"110011101",
  5812=>"111011000",
  5813=>"000010001",
  5814=>"011001101",
  5815=>"111111011",
  5816=>"011001010",
  5817=>"110011000",
  5818=>"011110010",
  5819=>"111001001",
  5820=>"110100010",
  5821=>"010010100",
  5822=>"111101111",
  5823=>"111111110",
  5824=>"011010110",
  5825=>"001100001",
  5826=>"011110100",
  5827=>"101100000",
  5828=>"101000011",
  5829=>"101001000",
  5830=>"110110011",
  5831=>"110110110",
  5832=>"101101111",
  5833=>"001101110",
  5834=>"101111011",
  5835=>"111001101",
  5836=>"010001110",
  5837=>"111010110",
  5838=>"110001110",
  5839=>"000001010",
  5840=>"001100100",
  5841=>"110000001",
  5842=>"110100011",
  5843=>"000011100",
  5844=>"000111111",
  5845=>"000110111",
  5846=>"011101000",
  5847=>"001001011",
  5848=>"011011001",
  5849=>"001101001",
  5850=>"001101110",
  5851=>"010001111",
  5852=>"110111001",
  5853=>"101111110",
  5854=>"000000010",
  5855=>"011000000",
  5856=>"101001011",
  5857=>"010110101",
  5858=>"010100101",
  5859=>"011010000",
  5860=>"000111100",
  5861=>"111010101",
  5862=>"001101110",
  5863=>"110111010",
  5864=>"111111110",
  5865=>"000001011",
  5866=>"100111111",
  5867=>"101000111",
  5868=>"111111100",
  5869=>"101010111",
  5870=>"001001100",
  5871=>"110111010",
  5872=>"000000010",
  5873=>"011010100",
  5874=>"101111110",
  5875=>"010010001",
  5876=>"100001111",
  5877=>"001101111",
  5878=>"010110101",
  5879=>"010110011",
  5880=>"110001010",
  5881=>"000011000",
  5882=>"011001100",
  5883=>"110101001",
  5884=>"001010000",
  5885=>"110100110",
  5886=>"001001011",
  5887=>"001000001",
  5888=>"000101111",
  5889=>"100001110",
  5890=>"100000110",
  5891=>"111111100",
  5892=>"000001100",
  5893=>"110110011",
  5894=>"000111110",
  5895=>"100000010",
  5896=>"110010010",
  5897=>"010110000",
  5898=>"001101000",
  5899=>"000110111",
  5900=>"001001110",
  5901=>"111011111",
  5902=>"101000100",
  5903=>"100100000",
  5904=>"111111010",
  5905=>"110010011",
  5906=>"000010010",
  5907=>"011111110",
  5908=>"000001000",
  5909=>"111010011",
  5910=>"110000111",
  5911=>"110110001",
  5912=>"011110110",
  5913=>"111111110",
  5914=>"111111100",
  5915=>"111000011",
  5916=>"111110101",
  5917=>"101111011",
  5918=>"111000101",
  5919=>"010111111",
  5920=>"100000000",
  5921=>"101010000",
  5922=>"011100010",
  5923=>"000000000",
  5924=>"111111100",
  5925=>"101101101",
  5926=>"010001000",
  5927=>"110001100",
  5928=>"011111010",
  5929=>"101010111",
  5930=>"001100101",
  5931=>"111001111",
  5932=>"110110000",
  5933=>"111100100",
  5934=>"001111101",
  5935=>"110000001",
  5936=>"110110111",
  5937=>"011100001",
  5938=>"011111110",
  5939=>"010001100",
  5940=>"110001010",
  5941=>"000000001",
  5942=>"000011010",
  5943=>"111110010",
  5944=>"100001111",
  5945=>"111000001",
  5946=>"011110010",
  5947=>"000101100",
  5948=>"011101110",
  5949=>"101110110",
  5950=>"110110100",
  5951=>"010011111",
  5952=>"111111100",
  5953=>"100100011",
  5954=>"000001111",
  5955=>"111011110",
  5956=>"111110010",
  5957=>"000010001",
  5958=>"011100110",
  5959=>"000001000",
  5960=>"111010000",
  5961=>"100100001",
  5962=>"101100000",
  5963=>"101111100",
  5964=>"000101110",
  5965=>"000000101",
  5966=>"001100001",
  5967=>"100011101",
  5968=>"101101010",
  5969=>"100000000",
  5970=>"111111111",
  5971=>"101011110",
  5972=>"111101111",
  5973=>"010100111",
  5974=>"101111101",
  5975=>"001011110",
  5976=>"101111000",
  5977=>"011000000",
  5978=>"110010100",
  5979=>"111111001",
  5980=>"000000010",
  5981=>"011001111",
  5982=>"001101000",
  5983=>"111111111",
  5984=>"110010101",
  5985=>"110001111",
  5986=>"111111101",
  5987=>"010100111",
  5988=>"101011001",
  5989=>"011111101",
  5990=>"101000011",
  5991=>"100000100",
  5992=>"011011110",
  5993=>"110000100",
  5994=>"111010010",
  5995=>"111011111",
  5996=>"111101101",
  5997=>"101010010",
  5998=>"010111011",
  5999=>"011100100",
  6000=>"011111011",
  6001=>"010100111",
  6002=>"001100011",
  6003=>"111111000",
  6004=>"001111111",
  6005=>"111111010",
  6006=>"101110110",
  6007=>"110011010",
  6008=>"000100110",
  6009=>"010000000",
  6010=>"111110000",
  6011=>"111011011",
  6012=>"111111000",
  6013=>"111000001",
  6014=>"000100001",
  6015=>"000111000",
  6016=>"111011011",
  6017=>"111000110",
  6018=>"111111011",
  6019=>"001100001",
  6020=>"111110111",
  6021=>"100101101",
  6022=>"001011010",
  6023=>"101110010",
  6024=>"000110111",
  6025=>"111101111",
  6026=>"000000110",
  6027=>"011000011",
  6028=>"111110110",
  6029=>"100001010",
  6030=>"001111000",
  6031=>"001001001",
  6032=>"001001110",
  6033=>"111100010",
  6034=>"101111000",
  6035=>"100101110",
  6036=>"011101101",
  6037=>"011000100",
  6038=>"110010110",
  6039=>"001111001",
  6040=>"111100110",
  6041=>"001001000",
  6042=>"000111100",
  6043=>"010110010",
  6044=>"101100110",
  6045=>"001001100",
  6046=>"010011110",
  6047=>"111001101",
  6048=>"100000001",
  6049=>"110000101",
  6050=>"001010011",
  6051=>"111111101",
  6052=>"101111111",
  6053=>"000000000",
  6054=>"010011011",
  6055=>"111101011",
  6056=>"101010101",
  6057=>"010011111",
  6058=>"000000110",
  6059=>"100010001",
  6060=>"101101010",
  6061=>"010100000",
  6062=>"000101010",
  6063=>"011001101",
  6064=>"010111111",
  6065=>"000000001",
  6066=>"111001100",
  6067=>"110111101",
  6068=>"001000001",
  6069=>"010000010",
  6070=>"110000100",
  6071=>"100011001",
  6072=>"000110011",
  6073=>"011110000",
  6074=>"010001111",
  6075=>"010100100",
  6076=>"011101111",
  6077=>"101111001",
  6078=>"111101001",
  6079=>"111100110",
  6080=>"101000001",
  6081=>"100100000",
  6082=>"101100000",
  6083=>"000001011",
  6084=>"011010000",
  6085=>"110010111",
  6086=>"111011101",
  6087=>"011110000",
  6088=>"111111001",
  6089=>"101111111",
  6090=>"100101000",
  6091=>"101001100",
  6092=>"100010001",
  6093=>"110101111",
  6094=>"001100001",
  6095=>"001111101",
  6096=>"110000110",
  6097=>"000110101",
  6098=>"000110100",
  6099=>"001011001",
  6100=>"110111010",
  6101=>"100001100",
  6102=>"011111001",
  6103=>"001011111",
  6104=>"101111000",
  6105=>"110011001",
  6106=>"011111110",
  6107=>"000010111",
  6108=>"000101111",
  6109=>"111010000",
  6110=>"101110010",
  6111=>"010111110",
  6112=>"101100001",
  6113=>"001111110",
  6114=>"110010011",
  6115=>"011110011",
  6116=>"111111101",
  6117=>"111111111",
  6118=>"000001100",
  6119=>"011101110",
  6120=>"010111110",
  6121=>"010010001",
  6122=>"010101101",
  6123=>"000001010",
  6124=>"010101101",
  6125=>"011011011",
  6126=>"101011111",
  6127=>"001010100",
  6128=>"100111011",
  6129=>"010100111",
  6130=>"101100111",
  6131=>"000111100",
  6132=>"111010111",
  6133=>"111111001",
  6134=>"000000000",
  6135=>"101100000",
  6136=>"110111000",
  6137=>"101011010",
  6138=>"101010110",
  6139=>"101001101",
  6140=>"101000111",
  6141=>"111011111",
  6142=>"011010010",
  6143=>"101101001",
  6144=>"011010010",
  6145=>"000100010",
  6146=>"010111001",
  6147=>"000110110",
  6148=>"001100111",
  6149=>"100010100",
  6150=>"110101110",
  6151=>"100010000",
  6152=>"101101110",
  6153=>"110101011",
  6154=>"001110000",
  6155=>"101100000",
  6156=>"110011011",
  6157=>"110001011",
  6158=>"111000011",
  6159=>"000001000",
  6160=>"110101010",
  6161=>"101010000",
  6162=>"110000000",
  6163=>"011111101",
  6164=>"100100110",
  6165=>"100111010",
  6166=>"101011100",
  6167=>"000101100",
  6168=>"110100010",
  6169=>"000000111",
  6170=>"110100010",
  6171=>"011111111",
  6172=>"010010000",
  6173=>"110000100",
  6174=>"101101001",
  6175=>"111111000",
  6176=>"011111010",
  6177=>"001101110",
  6178=>"110010000",
  6179=>"100001011",
  6180=>"110000110",
  6181=>"010101010",
  6182=>"010101101",
  6183=>"001001001",
  6184=>"010001110",
  6185=>"111101010",
  6186=>"010001001",
  6187=>"111100011",
  6188=>"111101001",
  6189=>"001000011",
  6190=>"011111101",
  6191=>"000010101",
  6192=>"011010001",
  6193=>"010111110",
  6194=>"000100001",
  6195=>"100111001",
  6196=>"101011110",
  6197=>"111111010",
  6198=>"000001010",
  6199=>"101000011",
  6200=>"000000000",
  6201=>"110101011",
  6202=>"000111001",
  6203=>"011010010",
  6204=>"101100001",
  6205=>"001001101",
  6206=>"100010000",
  6207=>"001111111",
  6208=>"111000011",
  6209=>"000001101",
  6210=>"000110000",
  6211=>"000000011",
  6212=>"101001111",
  6213=>"001000110",
  6214=>"101001111",
  6215=>"001111000",
  6216=>"010001111",
  6217=>"111111101",
  6218=>"001001101",
  6219=>"111011100",
  6220=>"011111110",
  6221=>"001000111",
  6222=>"110111011",
  6223=>"101111101",
  6224=>"010110111",
  6225=>"000000111",
  6226=>"011110100",
  6227=>"101001000",
  6228=>"110110111",
  6229=>"111111111",
  6230=>"101001000",
  6231=>"010110101",
  6232=>"001101001",
  6233=>"011111110",
  6234=>"001101010",
  6235=>"010110011",
  6236=>"011000000",
  6237=>"010100000",
  6238=>"000010010",
  6239=>"000010011",
  6240=>"010100000",
  6241=>"011111010",
  6242=>"010010111",
  6243=>"010010011",
  6244=>"000111110",
  6245=>"110101101",
  6246=>"101100011",
  6247=>"001110100",
  6248=>"101011011",
  6249=>"000111010",
  6250=>"110100011",
  6251=>"110111101",
  6252=>"001010101",
  6253=>"010101001",
  6254=>"001011100",
  6255=>"000111001",
  6256=>"111000011",
  6257=>"110111000",
  6258=>"111001010",
  6259=>"001010010",
  6260=>"101000100",
  6261=>"001101001",
  6262=>"111111111",
  6263=>"100001011",
  6264=>"101010100",
  6265=>"000000111",
  6266=>"001000110",
  6267=>"001000101",
  6268=>"110001101",
  6269=>"111110010",
  6270=>"000010000",
  6271=>"011000001",
  6272=>"010100111",
  6273=>"111001000",
  6274=>"100011010",
  6275=>"000000101",
  6276=>"100110000",
  6277=>"111110001",
  6278=>"001011100",
  6279=>"001101111",
  6280=>"101011111",
  6281=>"100101011",
  6282=>"011010000",
  6283=>"000000000",
  6284=>"001101010",
  6285=>"100000000",
  6286=>"111111000",
  6287=>"011010000",
  6288=>"000100110",
  6289=>"011001101",
  6290=>"100011101",
  6291=>"011010100",
  6292=>"011101000",
  6293=>"001101100",
  6294=>"111011010",
  6295=>"001101110",
  6296=>"001110100",
  6297=>"100110000",
  6298=>"111010100",
  6299=>"100000011",
  6300=>"000000110",
  6301=>"101101101",
  6302=>"000010100",
  6303=>"000001010",
  6304=>"101110110",
  6305=>"000000010",
  6306=>"011101001",
  6307=>"010001011",
  6308=>"001011111",
  6309=>"001111101",
  6310=>"110110010",
  6311=>"110100000",
  6312=>"101101011",
  6313=>"111111000",
  6314=>"000100000",
  6315=>"001001010",
  6316=>"101100000",
  6317=>"001110011",
  6318=>"110001111",
  6319=>"101101010",
  6320=>"100001111",
  6321=>"000110011",
  6322=>"110110011",
  6323=>"000000100",
  6324=>"110010110",
  6325=>"101010111",
  6326=>"100000000",
  6327=>"010110100",
  6328=>"010110000",
  6329=>"101001101",
  6330=>"000010100",
  6331=>"000010111",
  6332=>"000111101",
  6333=>"010011001",
  6334=>"110001011",
  6335=>"110110111",
  6336=>"000010010",
  6337=>"010100100",
  6338=>"011011110",
  6339=>"100011010",
  6340=>"101000010",
  6341=>"011000001",
  6342=>"011000110",
  6343=>"000011111",
  6344=>"111010001",
  6345=>"101010111",
  6346=>"010001000",
  6347=>"100101001",
  6348=>"111011001",
  6349=>"101000100",
  6350=>"101010000",
  6351=>"011110010",
  6352=>"100111011",
  6353=>"110011011",
  6354=>"010111100",
  6355=>"010010100",
  6356=>"000001010",
  6357=>"111111111",
  6358=>"100101000",
  6359=>"101010000",
  6360=>"101110110",
  6361=>"000011001",
  6362=>"010101010",
  6363=>"110000110",
  6364=>"001000111",
  6365=>"011110010",
  6366=>"110000000",
  6367=>"001010011",
  6368=>"010010101",
  6369=>"100000101",
  6370=>"111111100",
  6371=>"000110011",
  6372=>"000000111",
  6373=>"111101000",
  6374=>"010101000",
  6375=>"101101101",
  6376=>"111011010",
  6377=>"001000101",
  6378=>"111111100",
  6379=>"111010000",
  6380=>"101001110",
  6381=>"111000101",
  6382=>"100010001",
  6383=>"000000000",
  6384=>"101110011",
  6385=>"111111111",
  6386=>"100111111",
  6387=>"100110011",
  6388=>"101111100",
  6389=>"010010100",
  6390=>"010001010",
  6391=>"100010001",
  6392=>"000111000",
  6393=>"111111111",
  6394=>"101111011",
  6395=>"010000000",
  6396=>"000110101",
  6397=>"100111110",
  6398=>"011110000",
  6399=>"101101100",
  6400=>"111011110",
  6401=>"111100000",
  6402=>"100011000",
  6403=>"100011100",
  6404=>"111111100",
  6405=>"010100010",
  6406=>"010000111",
  6407=>"011101000",
  6408=>"101101101",
  6409=>"100101010",
  6410=>"110110010",
  6411=>"101011001",
  6412=>"000001100",
  6413=>"110001101",
  6414=>"101001101",
  6415=>"000001011",
  6416=>"001100100",
  6417=>"010000000",
  6418=>"001000000",
  6419=>"111011001",
  6420=>"100000101",
  6421=>"001111100",
  6422=>"110000111",
  6423=>"001001011",
  6424=>"110110001",
  6425=>"001001000",
  6426=>"000100110",
  6427=>"111000010",
  6428=>"001001010",
  6429=>"100110000",
  6430=>"101011110",
  6431=>"010010110",
  6432=>"100110111",
  6433=>"010000010",
  6434=>"010010100",
  6435=>"010110111",
  6436=>"010100011",
  6437=>"101100110",
  6438=>"100011001",
  6439=>"011110011",
  6440=>"010000010",
  6441=>"000001000",
  6442=>"000010110",
  6443=>"010101010",
  6444=>"010100011",
  6445=>"100110011",
  6446=>"110010011",
  6447=>"110100101",
  6448=>"010100111",
  6449=>"001000100",
  6450=>"100010001",
  6451=>"010010110",
  6452=>"000011101",
  6453=>"000000001",
  6454=>"101111101",
  6455=>"110010001",
  6456=>"111001100",
  6457=>"000111111",
  6458=>"111101101",
  6459=>"111111100",
  6460=>"011101100",
  6461=>"001110000",
  6462=>"100100111",
  6463=>"001001100",
  6464=>"010110100",
  6465=>"100101111",
  6466=>"110111110",
  6467=>"010010111",
  6468=>"110100000",
  6469=>"111011000",
  6470=>"010000101",
  6471=>"111110011",
  6472=>"010000011",
  6473=>"111011101",
  6474=>"100100011",
  6475=>"001101110",
  6476=>"111011001",
  6477=>"110100100",
  6478=>"100110001",
  6479=>"111111110",
  6480=>"001000011",
  6481=>"001100001",
  6482=>"000001111",
  6483=>"000111111",
  6484=>"011100111",
  6485=>"111100100",
  6486=>"110010101",
  6487=>"000100000",
  6488=>"110110000",
  6489=>"100110100",
  6490=>"011000010",
  6491=>"100010001",
  6492=>"001001000",
  6493=>"111011111",
  6494=>"111010111",
  6495=>"000010100",
  6496=>"101000001",
  6497=>"001000011",
  6498=>"010111010",
  6499=>"110111001",
  6500=>"010100011",
  6501=>"001000100",
  6502=>"001100110",
  6503=>"100010101",
  6504=>"101011010",
  6505=>"000000010",
  6506=>"101100001",
  6507=>"011010100",
  6508=>"101001110",
  6509=>"100101101",
  6510=>"100100101",
  6511=>"100000100",
  6512=>"010100000",
  6513=>"111010110",
  6514=>"101001111",
  6515=>"111001100",
  6516=>"010110000",
  6517=>"011000000",
  6518=>"111011011",
  6519=>"111010000",
  6520=>"111110100",
  6521=>"101000000",
  6522=>"110111111",
  6523=>"101011110",
  6524=>"011000010",
  6525=>"111111111",
  6526=>"010110110",
  6527=>"101000100",
  6528=>"101001010",
  6529=>"001011100",
  6530=>"100111100",
  6531=>"110111101",
  6532=>"100011110",
  6533=>"101101011",
  6534=>"001101010",
  6535=>"111100111",
  6536=>"111100000",
  6537=>"100111110",
  6538=>"110100111",
  6539=>"111111110",
  6540=>"110110001",
  6541=>"111001110",
  6542=>"111100100",
  6543=>"111111111",
  6544=>"000100010",
  6545=>"010111111",
  6546=>"101111110",
  6547=>"010011110",
  6548=>"011011110",
  6549=>"000001010",
  6550=>"110111101",
  6551=>"011011100",
  6552=>"000111001",
  6553=>"100000001",
  6554=>"010001011",
  6555=>"010111001",
  6556=>"111000100",
  6557=>"111110100",
  6558=>"110101111",
  6559=>"100011010",
  6560=>"100000100",
  6561=>"001100011",
  6562=>"111101010",
  6563=>"110011000",
  6564=>"101111010",
  6565=>"111011100",
  6566=>"001001100",
  6567=>"110111111",
  6568=>"100111110",
  6569=>"011011100",
  6570=>"001001010",
  6571=>"000010111",
  6572=>"011111110",
  6573=>"010100010",
  6574=>"010101111",
  6575=>"100110110",
  6576=>"110101010",
  6577=>"000110110",
  6578=>"000000010",
  6579=>"111101110",
  6580=>"110101111",
  6581=>"100110101",
  6582=>"110110110",
  6583=>"100011000",
  6584=>"111010001",
  6585=>"000010101",
  6586=>"111010000",
  6587=>"011001100",
  6588=>"101101101",
  6589=>"000100101",
  6590=>"100111111",
  6591=>"000001011",
  6592=>"111010010",
  6593=>"000010010",
  6594=>"001000010",
  6595=>"110111111",
  6596=>"010010001",
  6597=>"101111010",
  6598=>"011111110",
  6599=>"100000000",
  6600=>"000111111",
  6601=>"010000000",
  6602=>"111100110",
  6603=>"011101101",
  6604=>"010110010",
  6605=>"110110111",
  6606=>"000001100",
  6607=>"110011010",
  6608=>"001110001",
  6609=>"010001111",
  6610=>"111111010",
  6611=>"110010111",
  6612=>"110100110",
  6613=>"001000111",
  6614=>"000110101",
  6615=>"110100111",
  6616=>"110001110",
  6617=>"110000101",
  6618=>"000001010",
  6619=>"000001110",
  6620=>"100111100",
  6621=>"110100010",
  6622=>"110000011",
  6623=>"010011011",
  6624=>"011000000",
  6625=>"111010001",
  6626=>"111111000",
  6627=>"110001111",
  6628=>"000101110",
  6629=>"111010011",
  6630=>"010101011",
  6631=>"100011111",
  6632=>"100110110",
  6633=>"110111100",
  6634=>"001000100",
  6635=>"111101100",
  6636=>"010000101",
  6637=>"010101000",
  6638=>"000111010",
  6639=>"010011000",
  6640=>"101000101",
  6641=>"010111110",
  6642=>"010000101",
  6643=>"110000101",
  6644=>"011100000",
  6645=>"101010101",
  6646=>"110011100",
  6647=>"111011011",
  6648=>"101100101",
  6649=>"011101011",
  6650=>"111010000",
  6651=>"010010010",
  6652=>"011011111",
  6653=>"110100010",
  6654=>"110001100",
  6655=>"100001010",
  6656=>"111010101",
  6657=>"110100000",
  6658=>"110010001",
  6659=>"001111100",
  6660=>"100111011",
  6661=>"110000001",
  6662=>"000101100",
  6663=>"011011101",
  6664=>"000010000",
  6665=>"100101101",
  6666=>"011111100",
  6667=>"011111000",
  6668=>"010100011",
  6669=>"000011001",
  6670=>"100001101",
  6671=>"101111011",
  6672=>"111000110",
  6673=>"000100111",
  6674=>"000001100",
  6675=>"000010011",
  6676=>"101001000",
  6677=>"011101000",
  6678=>"010101110",
  6679=>"101001000",
  6680=>"010001010",
  6681=>"001001110",
  6682=>"000011011",
  6683=>"011010011",
  6684=>"101111100",
  6685=>"111111001",
  6686=>"110111101",
  6687=>"101000101",
  6688=>"111000001",
  6689=>"001011011",
  6690=>"011101000",
  6691=>"100111111",
  6692=>"011110111",
  6693=>"001101001",
  6694=>"011001001",
  6695=>"010011000",
  6696=>"010000111",
  6697=>"010010101",
  6698=>"101101000",
  6699=>"101001111",
  6700=>"101100100",
  6701=>"010111110",
  6702=>"010110101",
  6703=>"001011101",
  6704=>"000000101",
  6705=>"011100110",
  6706=>"010000100",
  6707=>"100100111",
  6708=>"011001011",
  6709=>"010000000",
  6710=>"100011101",
  6711=>"011001110",
  6712=>"111001111",
  6713=>"000100100",
  6714=>"000000000",
  6715=>"000010101",
  6716=>"100101101",
  6717=>"000010010",
  6718=>"000001000",
  6719=>"101011000",
  6720=>"011111010",
  6721=>"100000001",
  6722=>"101001001",
  6723=>"110010110",
  6724=>"111000010",
  6725=>"101110000",
  6726=>"000000100",
  6727=>"001001000",
  6728=>"110010100",
  6729=>"010111010",
  6730=>"111110101",
  6731=>"011001111",
  6732=>"110110001",
  6733=>"100100100",
  6734=>"110110101",
  6735=>"110011011",
  6736=>"010010110",
  6737=>"000011110",
  6738=>"101011111",
  6739=>"001010010",
  6740=>"111100111",
  6741=>"101000101",
  6742=>"110001110",
  6743=>"000111001",
  6744=>"011111001",
  6745=>"000100011",
  6746=>"000010001",
  6747=>"010011101",
  6748=>"001100101",
  6749=>"111010000",
  6750=>"110100001",
  6751=>"100000001",
  6752=>"000001001",
  6753=>"100110010",
  6754=>"011000110",
  6755=>"101101011",
  6756=>"100110010",
  6757=>"001010101",
  6758=>"110011110",
  6759=>"001000100",
  6760=>"000111000",
  6761=>"110001000",
  6762=>"110101110",
  6763=>"111011000",
  6764=>"111101111",
  6765=>"010011000",
  6766=>"110000000",
  6767=>"111100011",
  6768=>"000011001",
  6769=>"000001110",
  6770=>"000010110",
  6771=>"001000111",
  6772=>"100101111",
  6773=>"101101010",
  6774=>"110110101",
  6775=>"110100111",
  6776=>"011101010",
  6777=>"000010001",
  6778=>"010001010",
  6779=>"101000100",
  6780=>"110001010",
  6781=>"111111010",
  6782=>"100010110",
  6783=>"110011010",
  6784=>"111001110",
  6785=>"000000000",
  6786=>"100000001",
  6787=>"111110000",
  6788=>"101000010",
  6789=>"111010110",
  6790=>"100111010",
  6791=>"101011000",
  6792=>"000101010",
  6793=>"000010000",
  6794=>"111001111",
  6795=>"111110101",
  6796=>"101111111",
  6797=>"001101000",
  6798=>"010100100",
  6799=>"000000101",
  6800=>"101001110",
  6801=>"110110111",
  6802=>"110000101",
  6803=>"001000100",
  6804=>"001011111",
  6805=>"101100111",
  6806=>"110011011",
  6807=>"101010111",
  6808=>"101000110",
  6809=>"010001000",
  6810=>"000100100",
  6811=>"101110101",
  6812=>"101100011",
  6813=>"110010011",
  6814=>"110100110",
  6815=>"000100101",
  6816=>"100110111",
  6817=>"010011011",
  6818=>"000000111",
  6819=>"001001011",
  6820=>"000010110",
  6821=>"101001001",
  6822=>"010101101",
  6823=>"111011101",
  6824=>"001111001",
  6825=>"100000000",
  6826=>"101100010",
  6827=>"000101111",
  6828=>"111000000",
  6829=>"001100110",
  6830=>"000101101",
  6831=>"011111110",
  6832=>"011011111",
  6833=>"011010001",
  6834=>"101011110",
  6835=>"001010110",
  6836=>"001100011",
  6837=>"110111100",
  6838=>"010000010",
  6839=>"010011010",
  6840=>"101000110",
  6841=>"000000001",
  6842=>"000101111",
  6843=>"110100000",
  6844=>"100101010",
  6845=>"111111011",
  6846=>"011110001",
  6847=>"110111001",
  6848=>"110100111",
  6849=>"001010100",
  6850=>"111110100",
  6851=>"000010000",
  6852=>"100000001",
  6853=>"010011100",
  6854=>"101011111",
  6855=>"111111001",
  6856=>"100001100",
  6857=>"000100000",
  6858=>"111010000",
  6859=>"111000000",
  6860=>"100101111",
  6861=>"011001000",
  6862=>"000000110",
  6863=>"000101111",
  6864=>"011100010",
  6865=>"011000101",
  6866=>"100100101",
  6867=>"010100101",
  6868=>"111001001",
  6869=>"000000101",
  6870=>"011101011",
  6871=>"000100000",
  6872=>"111101110",
  6873=>"101100010",
  6874=>"001000010",
  6875=>"111100010",
  6876=>"111111000",
  6877=>"011011011",
  6878=>"101000101",
  6879=>"111000011",
  6880=>"101000110",
  6881=>"010000011",
  6882=>"000100011",
  6883=>"000000111",
  6884=>"011001011",
  6885=>"110101100",
  6886=>"000010011",
  6887=>"000110110",
  6888=>"011011100",
  6889=>"000101101",
  6890=>"001100010",
  6891=>"001011110",
  6892=>"111100001",
  6893=>"000101011",
  6894=>"001100111",
  6895=>"001000000",
  6896=>"011011100",
  6897=>"000100111",
  6898=>"001101110",
  6899=>"000101000",
  6900=>"110010001",
  6901=>"111110000",
  6902=>"100001101",
  6903=>"011110001",
  6904=>"111001011",
  6905=>"100110101",
  6906=>"001010110",
  6907=>"011100010",
  6908=>"110110100",
  6909=>"001111111",
  6910=>"000011110",
  6911=>"110000000",
  6912=>"101100001",
  6913=>"011100101",
  6914=>"101001000",
  6915=>"000100001",
  6916=>"111100010",
  6917=>"011101111",
  6918=>"001110100",
  6919=>"101110111",
  6920=>"010000010",
  6921=>"110100111",
  6922=>"010101110",
  6923=>"100010110",
  6924=>"110010010",
  6925=>"101011111",
  6926=>"000110101",
  6927=>"010000010",
  6928=>"100110110",
  6929=>"011110100",
  6930=>"001001100",
  6931=>"010101100",
  6932=>"010001110",
  6933=>"111000100",
  6934=>"001101000",
  6935=>"100000010",
  6936=>"111011111",
  6937=>"001011010",
  6938=>"000011011",
  6939=>"101111111",
  6940=>"010110100",
  6941=>"010100000",
  6942=>"110100101",
  6943=>"111110010",
  6944=>"100000100",
  6945=>"011111101",
  6946=>"010011111",
  6947=>"011001111",
  6948=>"111110011",
  6949=>"100111010",
  6950=>"111010011",
  6951=>"001100111",
  6952=>"000010000",
  6953=>"100001011",
  6954=>"010001111",
  6955=>"111110001",
  6956=>"100101110",
  6957=>"111001101",
  6958=>"001010011",
  6959=>"111101010",
  6960=>"100001101",
  6961=>"110100010",
  6962=>"101010110",
  6963=>"110011011",
  6964=>"110101111",
  6965=>"101101011",
  6966=>"111110111",
  6967=>"111110111",
  6968=>"100101010",
  6969=>"001000111",
  6970=>"100100110",
  6971=>"111001110",
  6972=>"000111001",
  6973=>"101011110",
  6974=>"000011100",
  6975=>"101010011",
  6976=>"110110010",
  6977=>"011010000",
  6978=>"001001001",
  6979=>"100001011",
  6980=>"011110100",
  6981=>"100100011",
  6982=>"011000000",
  6983=>"110011111",
  6984=>"101010000",
  6985=>"000101100",
  6986=>"100101101",
  6987=>"011110001",
  6988=>"011111011",
  6989=>"100101011",
  6990=>"100000001",
  6991=>"010001101",
  6992=>"000000000",
  6993=>"000011010",
  6994=>"001001001",
  6995=>"011000100",
  6996=>"111001100",
  6997=>"010101111",
  6998=>"111001000",
  6999=>"110110010",
  7000=>"011111111",
  7001=>"100010000",
  7002=>"001011110",
  7003=>"100011011",
  7004=>"100110100",
  7005=>"111101011",
  7006=>"011100110",
  7007=>"010100010",
  7008=>"110110010",
  7009=>"001001010",
  7010=>"111001000",
  7011=>"100111001",
  7012=>"011001000",
  7013=>"011111011",
  7014=>"001100101",
  7015=>"110110100",
  7016=>"110111000",
  7017=>"010011000",
  7018=>"000101001",
  7019=>"001110100",
  7020=>"101110111",
  7021=>"110011011",
  7022=>"010100010",
  7023=>"111100011",
  7024=>"011011010",
  7025=>"101001011",
  7026=>"101110111",
  7027=>"001101000",
  7028=>"110100111",
  7029=>"100100100",
  7030=>"110100011",
  7031=>"101011110",
  7032=>"010111101",
  7033=>"001101111",
  7034=>"010111110",
  7035=>"001000011",
  7036=>"111110011",
  7037=>"110010010",
  7038=>"010110010",
  7039=>"010011001",
  7040=>"110001001",
  7041=>"101111101",
  7042=>"110000011",
  7043=>"000010010",
  7044=>"001101000",
  7045=>"111110101",
  7046=>"010000100",
  7047=>"110001111",
  7048=>"110010001",
  7049=>"010110111",
  7050=>"111000101",
  7051=>"011001000",
  7052=>"010001011",
  7053=>"110110111",
  7054=>"100101101",
  7055=>"001101111",
  7056=>"101110101",
  7057=>"000100100",
  7058=>"001000001",
  7059=>"110110110",
  7060=>"011110110",
  7061=>"010111001",
  7062=>"001000100",
  7063=>"110011000",
  7064=>"001000010",
  7065=>"000110000",
  7066=>"101010000",
  7067=>"101010110",
  7068=>"000010001",
  7069=>"010100110",
  7070=>"000011010",
  7071=>"011010101",
  7072=>"100111110",
  7073=>"100100010",
  7074=>"000011111",
  7075=>"000110011",
  7076=>"100011101",
  7077=>"011010000",
  7078=>"011011110",
  7079=>"100110110",
  7080=>"101001100",
  7081=>"011000001",
  7082=>"101011110",
  7083=>"100000111",
  7084=>"110110000",
  7085=>"001001111",
  7086=>"011011111",
  7087=>"010001011",
  7088=>"100001011",
  7089=>"000100011",
  7090=>"011110101",
  7091=>"110000101",
  7092=>"011101110",
  7093=>"000001111",
  7094=>"011110101",
  7095=>"010001111",
  7096=>"011111101",
  7097=>"011100111",
  7098=>"111011011",
  7099=>"000010100",
  7100=>"000000110",
  7101=>"111011001",
  7102=>"110111011",
  7103=>"111110101",
  7104=>"100001000",
  7105=>"111000000",
  7106=>"000111101",
  7107=>"111010111",
  7108=>"101111010",
  7109=>"000000011",
  7110=>"000001011",
  7111=>"010111100",
  7112=>"010010100",
  7113=>"110111100",
  7114=>"100000001",
  7115=>"100001001",
  7116=>"011000000",
  7117=>"000000011",
  7118=>"101010001",
  7119=>"011100001",
  7120=>"111111000",
  7121=>"011100101",
  7122=>"110111000",
  7123=>"111111000",
  7124=>"101000000",
  7125=>"000000011",
  7126=>"100111010",
  7127=>"111110111",
  7128=>"000100001",
  7129=>"101001111",
  7130=>"000110011",
  7131=>"001100001",
  7132=>"110000010",
  7133=>"101100111",
  7134=>"000011110",
  7135=>"111000000",
  7136=>"100000100",
  7137=>"010111111",
  7138=>"000011111",
  7139=>"100011010",
  7140=>"010111010",
  7141=>"010100110",
  7142=>"101001101",
  7143=>"010100001",
  7144=>"101000100",
  7145=>"011001001",
  7146=>"110000110",
  7147=>"010011100",
  7148=>"010110010",
  7149=>"011110001",
  7150=>"000110111",
  7151=>"100101110",
  7152=>"110010111",
  7153=>"001100110",
  7154=>"011100010",
  7155=>"110011111",
  7156=>"001111100",
  7157=>"101001101",
  7158=>"100001000",
  7159=>"000011100",
  7160=>"110101101",
  7161=>"101100100",
  7162=>"111011011",
  7163=>"111011001",
  7164=>"111100010",
  7165=>"111100001",
  7166=>"011111100",
  7167=>"010001010",
  7168=>"101111111",
  7169=>"010011010",
  7170=>"100110111",
  7171=>"101101010",
  7172=>"111101101",
  7173=>"101111111",
  7174=>"101111000",
  7175=>"100001101",
  7176=>"000010000",
  7177=>"111011001",
  7178=>"100001000",
  7179=>"010000011",
  7180=>"000010001",
  7181=>"101000100",
  7182=>"000010011",
  7183=>"100111000",
  7184=>"011001111",
  7185=>"010011101",
  7186=>"010101000",
  7187=>"100111111",
  7188=>"010011101",
  7189=>"010110111",
  7190=>"011001100",
  7191=>"110001101",
  7192=>"011110000",
  7193=>"100011111",
  7194=>"100001011",
  7195=>"110101101",
  7196=>"010001001",
  7197=>"000001111",
  7198=>"010011011",
  7199=>"101000111",
  7200=>"000010011",
  7201=>"000100010",
  7202=>"000011000",
  7203=>"111000101",
  7204=>"101000010",
  7205=>"111001000",
  7206=>"101100111",
  7207=>"101100111",
  7208=>"110010010",
  7209=>"100000110",
  7210=>"101100100",
  7211=>"111011010",
  7212=>"111111111",
  7213=>"001001010",
  7214=>"000100001",
  7215=>"001010000",
  7216=>"010011101",
  7217=>"000000100",
  7218=>"111011000",
  7219=>"110011001",
  7220=>"111000001",
  7221=>"001000010",
  7222=>"000010011",
  7223=>"000011011",
  7224=>"000111101",
  7225=>"011111110",
  7226=>"100111101",
  7227=>"100001101",
  7228=>"001101010",
  7229=>"110010111",
  7230=>"111101010",
  7231=>"000111101",
  7232=>"111000000",
  7233=>"101010111",
  7234=>"010011100",
  7235=>"000011110",
  7236=>"001111011",
  7237=>"101011100",
  7238=>"000010100",
  7239=>"100110001",
  7240=>"000100110",
  7241=>"000001111",
  7242=>"000011000",
  7243=>"010011111",
  7244=>"000001100",
  7245=>"011000101",
  7246=>"010001000",
  7247=>"001000010",
  7248=>"011101001",
  7249=>"000001001",
  7250=>"010110001",
  7251=>"111101111",
  7252=>"010100110",
  7253=>"111111101",
  7254=>"001010111",
  7255=>"100000000",
  7256=>"110101111",
  7257=>"000101101",
  7258=>"001110011",
  7259=>"010100110",
  7260=>"110110110",
  7261=>"000101101",
  7262=>"000100111",
  7263=>"001110000",
  7264=>"001010100",
  7265=>"101010101",
  7266=>"000000100",
  7267=>"000001110",
  7268=>"000101111",
  7269=>"011111000",
  7270=>"110101101",
  7271=>"000001101",
  7272=>"010111011",
  7273=>"001001101",
  7274=>"011000111",
  7275=>"010000010",
  7276=>"011101111",
  7277=>"000000001",
  7278=>"001100000",
  7279=>"110110110",
  7280=>"001010101",
  7281=>"000110101",
  7282=>"010001111",
  7283=>"111101111",
  7284=>"011100111",
  7285=>"110100110",
  7286=>"100001111",
  7287=>"110010100",
  7288=>"111110101",
  7289=>"101000001",
  7290=>"001011001",
  7291=>"111111111",
  7292=>"110110010",
  7293=>"111010011",
  7294=>"111111111",
  7295=>"101000011",
  7296=>"101000011",
  7297=>"011010010",
  7298=>"010001101",
  7299=>"011000100",
  7300=>"000001011",
  7301=>"000000000",
  7302=>"011011010",
  7303=>"010100000",
  7304=>"001110011",
  7305=>"010111101",
  7306=>"001011111",
  7307=>"101000001",
  7308=>"100010100",
  7309=>"110001111",
  7310=>"110100111",
  7311=>"110011011",
  7312=>"001001111",
  7313=>"000111011",
  7314=>"101101110",
  7315=>"010001001",
  7316=>"110110000",
  7317=>"110111100",
  7318=>"001111111",
  7319=>"100001111",
  7320=>"111100101",
  7321=>"110100100",
  7322=>"111000010",
  7323=>"001101000",
  7324=>"000000011",
  7325=>"111101110",
  7326=>"111100111",
  7327=>"000100010",
  7328=>"110110110",
  7329=>"011101101",
  7330=>"111001010",
  7331=>"001111001",
  7332=>"000011000",
  7333=>"110110100",
  7334=>"000010111",
  7335=>"010110001",
  7336=>"100100011",
  7337=>"000011100",
  7338=>"100100001",
  7339=>"101100100",
  7340=>"101100111",
  7341=>"001000111",
  7342=>"000100100",
  7343=>"111101110",
  7344=>"001110100",
  7345=>"001101110",
  7346=>"000000100",
  7347=>"110100101",
  7348=>"011100110",
  7349=>"011000101",
  7350=>"001001011",
  7351=>"011111101",
  7352=>"101011100",
  7353=>"101000010",
  7354=>"111111110",
  7355=>"010011110",
  7356=>"111100000",
  7357=>"000000000",
  7358=>"000011110",
  7359=>"110010111",
  7360=>"111010001",
  7361=>"101100110",
  7362=>"110011100",
  7363=>"101001100",
  7364=>"000111110",
  7365=>"101000011",
  7366=>"100000101",
  7367=>"101101001",
  7368=>"000111010",
  7369=>"101110100",
  7370=>"010110101",
  7371=>"110010110",
  7372=>"100110110",
  7373=>"101101001",
  7374=>"010001111",
  7375=>"110100110",
  7376=>"001011110",
  7377=>"010000111",
  7378=>"000111110",
  7379=>"010011111",
  7380=>"110101110",
  7381=>"110001110",
  7382=>"110111111",
  7383=>"011100010",
  7384=>"000000100",
  7385=>"100011101",
  7386=>"000100000",
  7387=>"111110010",
  7388=>"111100001",
  7389=>"110010111",
  7390=>"101101011",
  7391=>"010111110",
  7392=>"010100010",
  7393=>"001110100",
  7394=>"111101100",
  7395=>"001000000",
  7396=>"010000010",
  7397=>"000110000",
  7398=>"101110100",
  7399=>"101111011",
  7400=>"010110010",
  7401=>"101000101",
  7402=>"010110001",
  7403=>"001110110",
  7404=>"000010011",
  7405=>"111010010",
  7406=>"100101001",
  7407=>"011110100",
  7408=>"011000100",
  7409=>"011110000",
  7410=>"101101101",
  7411=>"011001001",
  7412=>"100101100",
  7413=>"101011100",
  7414=>"000000110",
  7415=>"101101010",
  7416=>"110010111",
  7417=>"110101001",
  7418=>"001110010",
  7419=>"010001010",
  7420=>"000011101",
  7421=>"010010111",
  7422=>"100001001",
  7423=>"011010101",
  7424=>"000001111",
  7425=>"000000100",
  7426=>"111111101",
  7427=>"111011101",
  7428=>"100000011",
  7429=>"101110010",
  7430=>"010101011",
  7431=>"111110100",
  7432=>"000111111",
  7433=>"000001000",
  7434=>"001110000",
  7435=>"000000000",
  7436=>"100110011",
  7437=>"001000000",
  7438=>"100110100",
  7439=>"000000101",
  7440=>"011110100",
  7441=>"101111111",
  7442=>"011101000",
  7443=>"001011100",
  7444=>"101010110",
  7445=>"101000111",
  7446=>"100100111",
  7447=>"110010000",
  7448=>"110110100",
  7449=>"010101111",
  7450=>"000001111",
  7451=>"111001000",
  7452=>"100001100",
  7453=>"101000011",
  7454=>"000100111",
  7455=>"010000111",
  7456=>"010110101",
  7457=>"011111110",
  7458=>"011111110",
  7459=>"010000000",
  7460=>"101100010",
  7461=>"010111011",
  7462=>"110011010",
  7463=>"000101101",
  7464=>"101010000",
  7465=>"011110011",
  7466=>"101100001",
  7467=>"100010011",
  7468=>"001100011",
  7469=>"010010010",
  7470=>"000001000",
  7471=>"110100101",
  7472=>"000110000",
  7473=>"001010110",
  7474=>"001010100",
  7475=>"000101001",
  7476=>"110111101",
  7477=>"100110001",
  7478=>"010010011",
  7479=>"111000100",
  7480=>"000010010",
  7481=>"110010111",
  7482=>"001100000",
  7483=>"101011101",
  7484=>"001100110",
  7485=>"110110001",
  7486=>"010100110",
  7487=>"111110101",
  7488=>"110111110",
  7489=>"011110111",
  7490=>"000111000",
  7491=>"000110110",
  7492=>"111110010",
  7493=>"111111110",
  7494=>"110101001",
  7495=>"111100000",
  7496=>"110110100",
  7497=>"011101000",
  7498=>"000000010",
  7499=>"011011000",
  7500=>"000110001",
  7501=>"101110111",
  7502=>"011000100",
  7503=>"011111110",
  7504=>"101111010",
  7505=>"110001100",
  7506=>"101111101",
  7507=>"110010101",
  7508=>"110110010",
  7509=>"001001110",
  7510=>"000000001",
  7511=>"000010111",
  7512=>"010101000",
  7513=>"001000101",
  7514=>"000001001",
  7515=>"010000011",
  7516=>"001010100",
  7517=>"000100000",
  7518=>"000010110",
  7519=>"000001100",
  7520=>"000111111",
  7521=>"111010011",
  7522=>"101101010",
  7523=>"001010000",
  7524=>"111111011",
  7525=>"011011111",
  7526=>"100000111",
  7527=>"010010001",
  7528=>"001110100",
  7529=>"100001001",
  7530=>"000000001",
  7531=>"001100010",
  7532=>"010111111",
  7533=>"000110011",
  7534=>"001011000",
  7535=>"010000001",
  7536=>"110101101",
  7537=>"000001100",
  7538=>"111010010",
  7539=>"100000010",
  7540=>"110101001",
  7541=>"000000101",
  7542=>"011000110",
  7543=>"110001100",
  7544=>"010011101",
  7545=>"110111101",
  7546=>"111111100",
  7547=>"100110001",
  7548=>"011111101",
  7549=>"000010011",
  7550=>"000110000",
  7551=>"000001101",
  7552=>"101011111",
  7553=>"010001010",
  7554=>"110101100",
  7555=>"110110110",
  7556=>"101110010",
  7557=>"101101001",
  7558=>"000101110",
  7559=>"000000010",
  7560=>"001010111",
  7561=>"010011001",
  7562=>"011110100",
  7563=>"000010000",
  7564=>"111010110",
  7565=>"110010110",
  7566=>"000000100",
  7567=>"100101000",
  7568=>"110100000",
  7569=>"001001110",
  7570=>"011010111",
  7571=>"001101111",
  7572=>"101111111",
  7573=>"000110101",
  7574=>"101101101",
  7575=>"010011100",
  7576=>"110011110",
  7577=>"111000001",
  7578=>"111101010",
  7579=>"011000000",
  7580=>"010111101",
  7581=>"101011111",
  7582=>"110111000",
  7583=>"110111100",
  7584=>"110100100",
  7585=>"000010110",
  7586=>"000011011",
  7587=>"101001010",
  7588=>"101011111",
  7589=>"010000111",
  7590=>"110011011",
  7591=>"000001001",
  7592=>"100000011",
  7593=>"110001111",
  7594=>"010101011",
  7595=>"111001010",
  7596=>"001011001",
  7597=>"011101001",
  7598=>"100011101",
  7599=>"000011011",
  7600=>"100100000",
  7601=>"101101111",
  7602=>"001010100",
  7603=>"001000110",
  7604=>"101000110",
  7605=>"100011000",
  7606=>"110111001",
  7607=>"111010101",
  7608=>"110011010",
  7609=>"101110000",
  7610=>"111000001",
  7611=>"000111000",
  7612=>"100111110",
  7613=>"001000100",
  7614=>"011000010",
  7615=>"110111111",
  7616=>"111111100",
  7617=>"101001001",
  7618=>"010111101",
  7619=>"110101001",
  7620=>"110111101",
  7621=>"110011100",
  7622=>"001010001",
  7623=>"011100110",
  7624=>"000011001",
  7625=>"010100010",
  7626=>"101101101",
  7627=>"001101101",
  7628=>"011101111",
  7629=>"000001011",
  7630=>"100100000",
  7631=>"011100011",
  7632=>"110101010",
  7633=>"110111110",
  7634=>"100010101",
  7635=>"011011111",
  7636=>"011111001",
  7637=>"110110011",
  7638=>"010001100",
  7639=>"011101000",
  7640=>"000000101",
  7641=>"000011010",
  7642=>"110010001",
  7643=>"101010110",
  7644=>"000011010",
  7645=>"010000111",
  7646=>"111010010",
  7647=>"001110111",
  7648=>"000110111",
  7649=>"011111111",
  7650=>"110101100",
  7651=>"110011110",
  7652=>"100111010",
  7653=>"001111111",
  7654=>"110001001",
  7655=>"000001110",
  7656=>"100000110",
  7657=>"010001000",
  7658=>"010101010",
  7659=>"100000011",
  7660=>"000000011",
  7661=>"010010110",
  7662=>"110011110",
  7663=>"101011011",
  7664=>"110000000",
  7665=>"101111010",
  7666=>"100110100",
  7667=>"001111001",
  7668=>"110000001",
  7669=>"001101100",
  7670=>"011010110",
  7671=>"111100111",
  7672=>"111100011",
  7673=>"000111011",
  7674=>"100000101",
  7675=>"100110000",
  7676=>"001010001",
  7677=>"011010100",
  7678=>"110110011",
  7679=>"000001010",
  7680=>"111111111",
  7681=>"001111011",
  7682=>"111111100",
  7683=>"101011101",
  7684=>"000000111",
  7685=>"100100010",
  7686=>"010010011",
  7687=>"110000001",
  7688=>"010111011",
  7689=>"101101000",
  7690=>"000001101",
  7691=>"111000110",
  7692=>"000110010",
  7693=>"011100110",
  7694=>"100001100",
  7695=>"100110001",
  7696=>"010000110",
  7697=>"101111001",
  7698=>"011001001",
  7699=>"110001111",
  7700=>"110000001",
  7701=>"110111010",
  7702=>"001100111",
  7703=>"111111110",
  7704=>"010010111",
  7705=>"011110101",
  7706=>"101100001",
  7707=>"111101110",
  7708=>"111101000",
  7709=>"011010100",
  7710=>"001101101",
  7711=>"000000111",
  7712=>"000010100",
  7713=>"010011111",
  7714=>"100100011",
  7715=>"010011001",
  7716=>"011011101",
  7717=>"001010101",
  7718=>"001110101",
  7719=>"111101011",
  7720=>"100000111",
  7721=>"010011101",
  7722=>"100101100",
  7723=>"111000011",
  7724=>"110110111",
  7725=>"100101101",
  7726=>"110001101",
  7727=>"100000001",
  7728=>"001000110",
  7729=>"010000000",
  7730=>"001000111",
  7731=>"100110010",
  7732=>"000111000",
  7733=>"111111101",
  7734=>"111011000",
  7735=>"111000000",
  7736=>"111110011",
  7737=>"101111000",
  7738=>"011010000",
  7739=>"100000110",
  7740=>"100110110",
  7741=>"011000001",
  7742=>"110011011",
  7743=>"101011000",
  7744=>"100101010",
  7745=>"010001000",
  7746=>"101001111",
  7747=>"010000000",
  7748=>"110101000",
  7749=>"011110111",
  7750=>"001000010",
  7751=>"011110111",
  7752=>"111011100",
  7753=>"111001001",
  7754=>"101110000",
  7755=>"101001010",
  7756=>"101111001",
  7757=>"001100001",
  7758=>"101000100",
  7759=>"001101011",
  7760=>"001000100",
  7761=>"010101101",
  7762=>"100011011",
  7763=>"000111110",
  7764=>"110011011",
  7765=>"000001011",
  7766=>"010111010",
  7767=>"111010010",
  7768=>"101010111",
  7769=>"100000000",
  7770=>"000011100",
  7771=>"100100110",
  7772=>"100000001",
  7773=>"100001000",
  7774=>"100001010",
  7775=>"101101011",
  7776=>"100000101",
  7777=>"101011001",
  7778=>"111100100",
  7779=>"001110100",
  7780=>"110100010",
  7781=>"100001010",
  7782=>"000001100",
  7783=>"110111110",
  7784=>"000100010",
  7785=>"010010001",
  7786=>"111001101",
  7787=>"011101111",
  7788=>"110010000",
  7789=>"101100101",
  7790=>"111011111",
  7791=>"100011000",
  7792=>"000110000",
  7793=>"011000100",
  7794=>"001111101",
  7795=>"001111111",
  7796=>"110101101",
  7797=>"110100011",
  7798=>"000111101",
  7799=>"011101001",
  7800=>"011001001",
  7801=>"111000101",
  7802=>"010101100",
  7803=>"010001100",
  7804=>"100000110",
  7805=>"000100001",
  7806=>"110000000",
  7807=>"000011101",
  7808=>"000101001",
  7809=>"100101100",
  7810=>"111101111",
  7811=>"001001111",
  7812=>"001010000",
  7813=>"010101110",
  7814=>"110001111",
  7815=>"101111111",
  7816=>"101111011",
  7817=>"010001010",
  7818=>"010011000",
  7819=>"110100101",
  7820=>"010100000",
  7821=>"010001101",
  7822=>"011001000",
  7823=>"111001011",
  7824=>"100100100",
  7825=>"111110011",
  7826=>"100010000",
  7827=>"111101100",
  7828=>"000000000",
  7829=>"010010000",
  7830=>"001000011",
  7831=>"011010100",
  7832=>"101011110",
  7833=>"001101010",
  7834=>"110000111",
  7835=>"100001110",
  7836=>"111001100",
  7837=>"101111110",
  7838=>"101100010",
  7839=>"101110101",
  7840=>"110110101",
  7841=>"101101100",
  7842=>"101111111",
  7843=>"001101010",
  7844=>"111010110",
  7845=>"111001101",
  7846=>"110000000",
  7847=>"111001000",
  7848=>"101011111",
  7849=>"111001010",
  7850=>"100111000",
  7851=>"111001001",
  7852=>"101011010",
  7853=>"110011000",
  7854=>"011110111",
  7855=>"010010010",
  7856=>"110110111",
  7857=>"000100101",
  7858=>"110000111",
  7859=>"111010111",
  7860=>"111100111",
  7861=>"100000011",
  7862=>"111001110",
  7863=>"000111110",
  7864=>"101000111",
  7865=>"011111010",
  7866=>"111101111",
  7867=>"101110100",
  7868=>"101001000",
  7869=>"010011110",
  7870=>"000010010",
  7871=>"000010001",
  7872=>"111011111",
  7873=>"010101101",
  7874=>"000011100",
  7875=>"101100001",
  7876=>"011110001",
  7877=>"000001100",
  7878=>"010010001",
  7879=>"000001101",
  7880=>"011101001",
  7881=>"110010101",
  7882=>"000001000",
  7883=>"101001110",
  7884=>"011000111",
  7885=>"100110011",
  7886=>"110010101",
  7887=>"111000011",
  7888=>"000000101",
  7889=>"100100111",
  7890=>"001011100",
  7891=>"101001011",
  7892=>"011100000",
  7893=>"111010010",
  7894=>"011001010",
  7895=>"111111010",
  7896=>"000111101",
  7897=>"101100011",
  7898=>"110110101",
  7899=>"101101101",
  7900=>"100100011",
  7901=>"101000110",
  7902=>"110110001",
  7903=>"000001000",
  7904=>"100000000",
  7905=>"110101001",
  7906=>"110101101",
  7907=>"011100111",
  7908=>"011011110",
  7909=>"111000011",
  7910=>"101000001",
  7911=>"100000011",
  7912=>"000100001",
  7913=>"110001010",
  7914=>"000000001",
  7915=>"111000111",
  7916=>"101011111",
  7917=>"001011010",
  7918=>"001111101",
  7919=>"011111001",
  7920=>"011010100",
  7921=>"111011110",
  7922=>"000010100",
  7923=>"100111011",
  7924=>"110111011",
  7925=>"000001100",
  7926=>"000011000",
  7927=>"010000001",
  7928=>"011100000",
  7929=>"001101111",
  7930=>"100101010",
  7931=>"001001001",
  7932=>"110101010",
  7933=>"011111010",
  7934=>"111101110",
  7935=>"111001110",
  7936=>"011001011",
  7937=>"000011010",
  7938=>"000000100",
  7939=>"010010000",
  7940=>"100000010",
  7941=>"110101101",
  7942=>"000100110",
  7943=>"000111100",
  7944=>"011111101",
  7945=>"100100101",
  7946=>"100100010",
  7947=>"101000110",
  7948=>"110101111",
  7949=>"010110001",
  7950=>"100000100",
  7951=>"001110111",
  7952=>"000010001",
  7953=>"001000000",
  7954=>"110000000",
  7955=>"001101100",
  7956=>"111100100",
  7957=>"011110000",
  7958=>"101111111",
  7959=>"001111011",
  7960=>"101101001",
  7961=>"100011100",
  7962=>"111010111",
  7963=>"110011111",
  7964=>"010001000",
  7965=>"000100101",
  7966=>"101110101",
  7967=>"100001110",
  7968=>"000101001",
  7969=>"010001110",
  7970=>"010101101",
  7971=>"101111010",
  7972=>"110101000",
  7973=>"111101011",
  7974=>"110100100",
  7975=>"001100000",
  7976=>"001011010",
  7977=>"100111100",
  7978=>"001011010",
  7979=>"110011111",
  7980=>"110110100",
  7981=>"110010101",
  7982=>"100011110",
  7983=>"111000100",
  7984=>"001000000",
  7985=>"100001100",
  7986=>"010001000",
  7987=>"011010100",
  7988=>"011000000",
  7989=>"000100110",
  7990=>"101001111",
  7991=>"011110100",
  7992=>"111011100",
  7993=>"100110010",
  7994=>"010110110",
  7995=>"000001100",
  7996=>"110000001",
  7997=>"110000010",
  7998=>"101001000",
  7999=>"110010010",
  8000=>"111100001",
  8001=>"010110001",
  8002=>"011010111",
  8003=>"110000101",
  8004=>"011101110",
  8005=>"000000111",
  8006=>"111001100",
  8007=>"111011010",
  8008=>"011100101",
  8009=>"010111111",
  8010=>"011011001",
  8011=>"111110100",
  8012=>"100000000",
  8013=>"010111100",
  8014=>"100001000",
  8015=>"011111010",
  8016=>"111001001",
  8017=>"110001000",
  8018=>"000001000",
  8019=>"001001001",
  8020=>"101101000",
  8021=>"001011100",
  8022=>"110110100",
  8023=>"111010010",
  8024=>"000110010",
  8025=>"111000001",
  8026=>"110001111",
  8027=>"010001110",
  8028=>"110011011",
  8029=>"010111010",
  8030=>"011111001",
  8031=>"000010001",
  8032=>"101000000",
  8033=>"110110111",
  8034=>"000000100",
  8035=>"000111010",
  8036=>"001010010",
  8037=>"111011101",
  8038=>"100000100",
  8039=>"011110001",
  8040=>"000000000",
  8041=>"110110101",
  8042=>"011000110",
  8043=>"100101000",
  8044=>"000100100",
  8045=>"011110110",
  8046=>"110101100",
  8047=>"010110110",
  8048=>"010111000",
  8049=>"001101000",
  8050=>"010101101",
  8051=>"000011001",
  8052=>"010011011",
  8053=>"111111001",
  8054=>"101010110",
  8055=>"000000011",
  8056=>"101110011",
  8057=>"101100000",
  8058=>"110000001",
  8059=>"011001111",
  8060=>"111101111",
  8061=>"111000001",
  8062=>"100011010",
  8063=>"111111111",
  8064=>"101000010",
  8065=>"100111111",
  8066=>"010110011",
  8067=>"000010101",
  8068=>"000100110",
  8069=>"001101001",
  8070=>"011101011",
  8071=>"111010100",
  8072=>"110101111",
  8073=>"010000010",
  8074=>"010110100",
  8075=>"110000000",
  8076=>"110100000",
  8077=>"010010011",
  8078=>"000000110",
  8079=>"100000010",
  8080=>"110101011",
  8081=>"011100100",
  8082=>"100010111",
  8083=>"000100100",
  8084=>"000001001",
  8085=>"111111101",
  8086=>"111100110",
  8087=>"100010101",
  8088=>"101110101",
  8089=>"001000000",
  8090=>"000010100",
  8091=>"100001110",
  8092=>"110000001",
  8093=>"001110101",
  8094=>"111011011",
  8095=>"011000101",
  8096=>"111100001",
  8097=>"001001100",
  8098=>"011010111",
  8099=>"101101101",
  8100=>"000011010",
  8101=>"110100101",
  8102=>"001000011",
  8103=>"111111010",
  8104=>"010011100",
  8105=>"011100111",
  8106=>"111110110",
  8107=>"011001000",
  8108=>"000001100",
  8109=>"110110111",
  8110=>"000100010",
  8111=>"001010010",
  8112=>"011101111",
  8113=>"110101010",
  8114=>"001000001",
  8115=>"001110000",
  8116=>"000111111",
  8117=>"110101001",
  8118=>"110110001",
  8119=>"111011101",
  8120=>"000010100",
  8121=>"001111000",
  8122=>"001001000",
  8123=>"111110000",
  8124=>"011011111",
  8125=>"001010010",
  8126=>"110111110",
  8127=>"111111001",
  8128=>"001111111",
  8129=>"110111101",
  8130=>"010011001",
  8131=>"100001000",
  8132=>"110010001",
  8133=>"011001010",
  8134=>"001001000",
  8135=>"110110111",
  8136=>"001001010",
  8137=>"110110111",
  8138=>"011011100",
  8139=>"001110111",
  8140=>"011100100",
  8141=>"011000111",
  8142=>"000011011",
  8143=>"000000001",
  8144=>"000100110",
  8145=>"110110111",
  8146=>"110111010",
  8147=>"101101100",
  8148=>"110101110",
  8149=>"011011000",
  8150=>"100010010",
  8151=>"010111110",
  8152=>"001010010",
  8153=>"100000001",
  8154=>"011000000",
  8155=>"010001100",
  8156=>"010000111",
  8157=>"111111110",
  8158=>"011100101",
  8159=>"001000001",
  8160=>"111001001",
  8161=>"010000000",
  8162=>"001101000",
  8163=>"010110101",
  8164=>"001011111",
  8165=>"001101001",
  8166=>"100011100",
  8167=>"101011001",
  8168=>"000101010",
  8169=>"110011100",
  8170=>"000010100",
  8171=>"111001000",
  8172=>"011011011",
  8173=>"111010011",
  8174=>"110011100",
  8175=>"111111111",
  8176=>"011010011",
  8177=>"001110010",
  8178=>"110101110",
  8179=>"111100101",
  8180=>"111101000",
  8181=>"010101100",
  8182=>"111111011",
  8183=>"001000101",
  8184=>"001010111",
  8185=>"001011001",
  8186=>"000111110",
  8187=>"100001010",
  8188=>"110010001",
  8189=>"110010101",
  8190=>"100010100",
  8191=>"010011101",
  8192=>"101111100",
  8193=>"100000111",
  8194=>"100000011",
  8195=>"101000011",
  8196=>"110110001",
  8197=>"110010010",
  8198=>"001001100",
  8199=>"010011000",
  8200=>"101000001",
  8201=>"001101001",
  8202=>"000001111",
  8203=>"011110000",
  8204=>"101101000",
  8205=>"011010101",
  8206=>"010110011",
  8207=>"000010101",
  8208=>"110100100",
  8209=>"000111001",
  8210=>"110000010",
  8211=>"111000001",
  8212=>"011001111",
  8213=>"000111001",
  8214=>"011000111",
  8215=>"001000010",
  8216=>"110101100",
  8217=>"000011110",
  8218=>"011101100",
  8219=>"101111011",
  8220=>"101111000",
  8221=>"110110111",
  8222=>"000010000",
  8223=>"011000001",
  8224=>"001001111",
  8225=>"000111010",
  8226=>"111101100",
  8227=>"010001011",
  8228=>"011100100",
  8229=>"001010000",
  8230=>"110100010",
  8231=>"100100110",
  8232=>"110001110",
  8233=>"001101111",
  8234=>"001111011",
  8235=>"001000001",
  8236=>"100100010",
  8237=>"111111101",
  8238=>"010011110",
  8239=>"001101100",
  8240=>"110111000",
  8241=>"010101000",
  8242=>"111010111",
  8243=>"100100111",
  8244=>"100000010",
  8245=>"101100000",
  8246=>"111011110",
  8247=>"101111110",
  8248=>"000000100",
  8249=>"011101000",
  8250=>"100110100",
  8251=>"001100111",
  8252=>"111001111",
  8253=>"000001100",
  8254=>"010001100",
  8255=>"011011001",
  8256=>"110101111",
  8257=>"101001110",
  8258=>"010000001",
  8259=>"001001101",
  8260=>"000001000",
  8261=>"011001111",
  8262=>"100101001",
  8263=>"001010000",
  8264=>"001011001",
  8265=>"110011001",
  8266=>"100010010",
  8267=>"101101011",
  8268=>"111110000",
  8269=>"110001110",
  8270=>"000000101",
  8271=>"111110010",
  8272=>"110101010",
  8273=>"111001110",
  8274=>"011001111",
  8275=>"000011110",
  8276=>"010101110",
  8277=>"011101010",
  8278=>"100010010",
  8279=>"011111111",
  8280=>"111110101",
  8281=>"110100101",
  8282=>"111100110",
  8283=>"001000110",
  8284=>"000000010",
  8285=>"000001011",
  8286=>"110101001",
  8287=>"001000011",
  8288=>"111111111",
  8289=>"010100001",
  8290=>"111101010",
  8291=>"111001100",
  8292=>"010000001",
  8293=>"001111011",
  8294=>"110100000",
  8295=>"011100001",
  8296=>"111111111",
  8297=>"011110000",
  8298=>"011011001",
  8299=>"111100000",
  8300=>"011001110",
  8301=>"110110000",
  8302=>"100000100",
  8303=>"111110110",
  8304=>"000110010",
  8305=>"010011111",
  8306=>"111011110",
  8307=>"101011001",
  8308=>"001111011",
  8309=>"101110000",
  8310=>"111000111",
  8311=>"000110110",
  8312=>"011010100",
  8313=>"000001010",
  8314=>"011000010",
  8315=>"101111110",
  8316=>"100111101",
  8317=>"100100100",
  8318=>"110001100",
  8319=>"000001100",
  8320=>"011001100",
  8321=>"110110111",
  8322=>"100110000",
  8323=>"100010111",
  8324=>"001001100",
  8325=>"001101101",
  8326=>"111001000",
  8327=>"110001011",
  8328=>"111111001",
  8329=>"010011111",
  8330=>"100010001",
  8331=>"010100110",
  8332=>"100000001",
  8333=>"101101101",
  8334=>"011100110",
  8335=>"010000010",
  8336=>"111111010",
  8337=>"111111001",
  8338=>"111110111",
  8339=>"010000110",
  8340=>"100001111",
  8341=>"101000111",
  8342=>"001011001",
  8343=>"001101001",
  8344=>"011101110",
  8345=>"111011110",
  8346=>"000101111",
  8347=>"101101000",
  8348=>"001001010",
  8349=>"100100000",
  8350=>"001111000",
  8351=>"010111000",
  8352=>"100011010",
  8353=>"100000010",
  8354=>"011110110",
  8355=>"110010010",
  8356=>"110000010",
  8357=>"110011000",
  8358=>"101111001",
  8359=>"100000001",
  8360=>"010111011",
  8361=>"101010011",
  8362=>"010100100",
  8363=>"111010011",
  8364=>"011111110",
  8365=>"101100110",
  8366=>"110000100",
  8367=>"011111010",
  8368=>"000110011",
  8369=>"000001010",
  8370=>"111110100",
  8371=>"001000100",
  8372=>"011100001",
  8373=>"010001001",
  8374=>"110010000",
  8375=>"001001011",
  8376=>"100001110",
  8377=>"100011001",
  8378=>"100100000",
  8379=>"111001001",
  8380=>"001000000",
  8381=>"110000101",
  8382=>"110000000",
  8383=>"010001011",
  8384=>"001011101",
  8385=>"111111111",
  8386=>"111010010",
  8387=>"110010001",
  8388=>"010011000",
  8389=>"111101010",
  8390=>"111000110",
  8391=>"110101010",
  8392=>"001100001",
  8393=>"110100111",
  8394=>"000010001",
  8395=>"111111111",
  8396=>"101010111",
  8397=>"100110010",
  8398=>"000011011",
  8399=>"000011000",
  8400=>"010001101",
  8401=>"000010000",
  8402=>"011001111",
  8403=>"011101001",
  8404=>"000100010",
  8405=>"011001001",
  8406=>"010101101",
  8407=>"100000001",
  8408=>"110110000",
  8409=>"101110111",
  8410=>"001010111",
  8411=>"101010100",
  8412=>"110011100",
  8413=>"001000100",
  8414=>"100011000",
  8415=>"101001110",
  8416=>"100000001",
  8417=>"001001001",
  8418=>"010110111",
  8419=>"101011001",
  8420=>"100011011",
  8421=>"011111011",
  8422=>"100001101",
  8423=>"011111110",
  8424=>"011110010",
  8425=>"011101000",
  8426=>"101010000",
  8427=>"001111111",
  8428=>"010000010",
  8429=>"001010101",
  8430=>"001001011",
  8431=>"100000110",
  8432=>"001101111",
  8433=>"110111101",
  8434=>"001001100",
  8435=>"111100101",
  8436=>"110110000",
  8437=>"100000110",
  8438=>"101000000",
  8439=>"010111010",
  8440=>"111101111",
  8441=>"110011101",
  8442=>"111011111",
  8443=>"001010011",
  8444=>"100000000",
  8445=>"000011011",
  8446=>"001111001",
  8447=>"100101000",
  8448=>"110111000",
  8449=>"011010111",
  8450=>"101110110",
  8451=>"101000010",
  8452=>"100011110",
  8453=>"100100111",
  8454=>"110111010",
  8455=>"100100001",
  8456=>"101000010",
  8457=>"111111010",
  8458=>"000010011",
  8459=>"111111000",
  8460=>"011011110",
  8461=>"011100110",
  8462=>"011111101",
  8463=>"111010001",
  8464=>"110110100",
  8465=>"101101110",
  8466=>"101010001",
  8467=>"001000110",
  8468=>"010011001",
  8469=>"001010011",
  8470=>"001000010",
  8471=>"110010101",
  8472=>"000001010",
  8473=>"001100110",
  8474=>"110011110",
  8475=>"110001101",
  8476=>"001011110",
  8477=>"101000000",
  8478=>"010011100",
  8479=>"011001010",
  8480=>"100100100",
  8481=>"111011001",
  8482=>"101011110",
  8483=>"111010011",
  8484=>"101000100",
  8485=>"001011100",
  8486=>"010010011",
  8487=>"101110110",
  8488=>"110001000",
  8489=>"001000111",
  8490=>"101101000",
  8491=>"100100011",
  8492=>"100000011",
  8493=>"001000000",
  8494=>"110011010",
  8495=>"110110000",
  8496=>"100011010",
  8497=>"100110000",
  8498=>"101100110",
  8499=>"000010001",
  8500=>"101111001",
  8501=>"101100000",
  8502=>"000000011",
  8503=>"111110011",
  8504=>"000111010",
  8505=>"111111110",
  8506=>"101011000",
  8507=>"110110100",
  8508=>"100011101",
  8509=>"100101110",
  8510=>"001111000",
  8511=>"001101000",
  8512=>"100011111",
  8513=>"101000100",
  8514=>"000011110",
  8515=>"111111001",
  8516=>"001111110",
  8517=>"111110000",
  8518=>"000010101",
  8519=>"110011010",
  8520=>"000001001",
  8521=>"001001011",
  8522=>"110011101",
  8523=>"001001110",
  8524=>"100001000",
  8525=>"110100111",
  8526=>"101010111",
  8527=>"011001101",
  8528=>"000001010",
  8529=>"001100101",
  8530=>"110000100",
  8531=>"101111110",
  8532=>"100101101",
  8533=>"000111110",
  8534=>"100011111",
  8535=>"101011010",
  8536=>"101101101",
  8537=>"110100110",
  8538=>"001101101",
  8539=>"000100011",
  8540=>"011011001",
  8541=>"111001101",
  8542=>"111000010",
  8543=>"001111110",
  8544=>"011000101",
  8545=>"001010000",
  8546=>"000011000",
  8547=>"000101111",
  8548=>"001110111",
  8549=>"000101000",
  8550=>"100001001",
  8551=>"100011110",
  8552=>"101111111",
  8553=>"000101010",
  8554=>"100101001",
  8555=>"001101110",
  8556=>"001000111",
  8557=>"001010010",
  8558=>"000101001",
  8559=>"010101101",
  8560=>"011001111",
  8561=>"010000111",
  8562=>"011101001",
  8563=>"111100001",
  8564=>"101001101",
  8565=>"011011111",
  8566=>"100011111",
  8567=>"110010101",
  8568=>"101010010",
  8569=>"110000100",
  8570=>"101111111",
  8571=>"111000011",
  8572=>"011100110",
  8573=>"110101110",
  8574=>"010101110",
  8575=>"111101010",
  8576=>"001001111",
  8577=>"011110100",
  8578=>"111111101",
  8579=>"101110000",
  8580=>"011001101",
  8581=>"111011000",
  8582=>"101100111",
  8583=>"101011110",
  8584=>"110011010",
  8585=>"011110110",
  8586=>"101100111",
  8587=>"111110001",
  8588=>"000111010",
  8589=>"000010001",
  8590=>"001011110",
  8591=>"010000110",
  8592=>"001111111",
  8593=>"010001000",
  8594=>"101101000",
  8595=>"011000011",
  8596=>"011101011",
  8597=>"110100111",
  8598=>"001001001",
  8599=>"001001011",
  8600=>"101001100",
  8601=>"101001011",
  8602=>"101111101",
  8603=>"001011111",
  8604=>"101101000",
  8605=>"111011100",
  8606=>"000011111",
  8607=>"110000010",
  8608=>"101101100",
  8609=>"011011010",
  8610=>"111000010",
  8611=>"000111110",
  8612=>"011110001",
  8613=>"101100111",
  8614=>"110001000",
  8615=>"111110100",
  8616=>"001100111",
  8617=>"000110011",
  8618=>"000010111",
  8619=>"000010010",
  8620=>"100100100",
  8621=>"000101111",
  8622=>"111101100",
  8623=>"000011011",
  8624=>"100100101",
  8625=>"011111111",
  8626=>"000001101",
  8627=>"010001000",
  8628=>"100100000",
  8629=>"001000101",
  8630=>"101000011",
  8631=>"101111111",
  8632=>"001011111",
  8633=>"000100101",
  8634=>"001011000",
  8635=>"000100001",
  8636=>"001000101",
  8637=>"111101011",
  8638=>"110010100",
  8639=>"010100100",
  8640=>"011101001",
  8641=>"000000010",
  8642=>"111011010",
  8643=>"101000101",
  8644=>"010000011",
  8645=>"101110100",
  8646=>"111001011",
  8647=>"101001000",
  8648=>"000010110",
  8649=>"000000100",
  8650=>"101010001",
  8651=>"010111111",
  8652=>"011011101",
  8653=>"100001010",
  8654=>"001010001",
  8655=>"001110010",
  8656=>"010101100",
  8657=>"001110011",
  8658=>"000010101",
  8659=>"111000110",
  8660=>"111100001",
  8661=>"101010011",
  8662=>"010010110",
  8663=>"000100010",
  8664=>"100111010",
  8665=>"010001000",
  8666=>"001101010",
  8667=>"000100000",
  8668=>"111000001",
  8669=>"011000011",
  8670=>"010001111",
  8671=>"011010011",
  8672=>"100101111",
  8673=>"111010101",
  8674=>"100110001",
  8675=>"111110000",
  8676=>"111111010",
  8677=>"011110100",
  8678=>"101100010",
  8679=>"111110101",
  8680=>"101001011",
  8681=>"110110000",
  8682=>"100100001",
  8683=>"110100001",
  8684=>"101111100",
  8685=>"011111100",
  8686=>"110100000",
  8687=>"111100100",
  8688=>"001001011",
  8689=>"010111100",
  8690=>"100100001",
  8691=>"111001000",
  8692=>"111101100",
  8693=>"110011100",
  8694=>"110010010",
  8695=>"010010000",
  8696=>"111111010",
  8697=>"101110001",
  8698=>"001001000",
  8699=>"110000110",
  8700=>"111111111",
  8701=>"111110111",
  8702=>"001100101",
  8703=>"100110111",
  8704=>"011000101",
  8705=>"111010000",
  8706=>"001010100",
  8707=>"111000001",
  8708=>"011111100",
  8709=>"101011001",
  8710=>"010001011",
  8711=>"111001011",
  8712=>"011010111",
  8713=>"110000001",
  8714=>"011101101",
  8715=>"001000100",
  8716=>"100110100",
  8717=>"110011011",
  8718=>"000011111",
  8719=>"010110100",
  8720=>"100010101",
  8721=>"111110110",
  8722=>"010001100",
  8723=>"010110011",
  8724=>"000011001",
  8725=>"000010101",
  8726=>"001010000",
  8727=>"011000101",
  8728=>"000110110",
  8729=>"100010011",
  8730=>"101001011",
  8731=>"000011110",
  8732=>"000011111",
  8733=>"111111000",
  8734=>"001110011",
  8735=>"100010110",
  8736=>"001001000",
  8737=>"001001000",
  8738=>"010001010",
  8739=>"101111010",
  8740=>"110001111",
  8741=>"010101100",
  8742=>"001010000",
  8743=>"000011011",
  8744=>"100111110",
  8745=>"000101010",
  8746=>"101101101",
  8747=>"011010001",
  8748=>"000010100",
  8749=>"010100000",
  8750=>"111101100",
  8751=>"110011100",
  8752=>"101000110",
  8753=>"111001101",
  8754=>"011000111",
  8755=>"011110010",
  8756=>"101011010",
  8757=>"010000011",
  8758=>"101010010",
  8759=>"000111101",
  8760=>"000010011",
  8761=>"110111010",
  8762=>"111101111",
  8763=>"101110111",
  8764=>"111111100",
  8765=>"110000100",
  8766=>"101011001",
  8767=>"010011001",
  8768=>"010111100",
  8769=>"110011110",
  8770=>"100000001",
  8771=>"110110000",
  8772=>"100100001",
  8773=>"111001010",
  8774=>"101111110",
  8775=>"000000100",
  8776=>"100110010",
  8777=>"011001110",
  8778=>"001010111",
  8779=>"101000011",
  8780=>"001000100",
  8781=>"100001000",
  8782=>"100011101",
  8783=>"011011111",
  8784=>"010101110",
  8785=>"011101101",
  8786=>"001000111",
  8787=>"001110001",
  8788=>"010100000",
  8789=>"000101110",
  8790=>"100100001",
  8791=>"001011010",
  8792=>"010100010",
  8793=>"001001000",
  8794=>"011101101",
  8795=>"110100001",
  8796=>"100101010",
  8797=>"000100011",
  8798=>"011111011",
  8799=>"001110011",
  8800=>"001111011",
  8801=>"001000100",
  8802=>"101111101",
  8803=>"000010100",
  8804=>"101111010",
  8805=>"110010001",
  8806=>"010001101",
  8807=>"011011101",
  8808=>"100010000",
  8809=>"111011000",
  8810=>"001101000",
  8811=>"011111010",
  8812=>"011100111",
  8813=>"000100100",
  8814=>"110110011",
  8815=>"001101010",
  8816=>"011000001",
  8817=>"011000001",
  8818=>"110001010",
  8819=>"100010001",
  8820=>"011101110",
  8821=>"000010111",
  8822=>"011011011",
  8823=>"110011010",
  8824=>"001011001",
  8825=>"010010101",
  8826=>"101110100",
  8827=>"010111001",
  8828=>"001010010",
  8829=>"010001110",
  8830=>"011100110",
  8831=>"100000001",
  8832=>"011110001",
  8833=>"111011111",
  8834=>"001011001",
  8835=>"000001011",
  8836=>"111111111",
  8837=>"011000110",
  8838=>"010000100",
  8839=>"110011110",
  8840=>"101110100",
  8841=>"000000111",
  8842=>"010011110",
  8843=>"111001010",
  8844=>"000111000",
  8845=>"110101111",
  8846=>"000110010",
  8847=>"000011011",
  8848=>"101011111",
  8849=>"010101110",
  8850=>"111000000",
  8851=>"011110111",
  8852=>"000101011",
  8853=>"111110111",
  8854=>"100001000",
  8855=>"010100111",
  8856=>"100110001",
  8857=>"011011010",
  8858=>"101000001",
  8859=>"101011010",
  8860=>"011011011",
  8861=>"111011001",
  8862=>"110100000",
  8863=>"111001010",
  8864=>"011111101",
  8865=>"001011001",
  8866=>"100101010",
  8867=>"101101100",
  8868=>"001111011",
  8869=>"001011000",
  8870=>"111011010",
  8871=>"100001010",
  8872=>"101100000",
  8873=>"001000001",
  8874=>"100001111",
  8875=>"011001001",
  8876=>"010000010",
  8877=>"101110000",
  8878=>"110001101",
  8879=>"000010011",
  8880=>"001011111",
  8881=>"010111110",
  8882=>"110001111",
  8883=>"110101100",
  8884=>"100000000",
  8885=>"111011100",
  8886=>"011011011",
  8887=>"100011000",
  8888=>"010101111",
  8889=>"001011011",
  8890=>"100111000",
  8891=>"001101101",
  8892=>"010011111",
  8893=>"011010000",
  8894=>"100000111",
  8895=>"011001000",
  8896=>"001010010",
  8897=>"011000010",
  8898=>"101011011",
  8899=>"110000111",
  8900=>"011010011",
  8901=>"001010110",
  8902=>"010011010",
  8903=>"001010111",
  8904=>"011000001",
  8905=>"111101100",
  8906=>"011100101",
  8907=>"001001101",
  8908=>"101110010",
  8909=>"100000100",
  8910=>"001001100",
  8911=>"011001011",
  8912=>"000000001",
  8913=>"101101110",
  8914=>"001110011",
  8915=>"001111100",
  8916=>"000010101",
  8917=>"000101100",
  8918=>"110110001",
  8919=>"000001001",
  8920=>"111001111",
  8921=>"110111010",
  8922=>"111001100",
  8923=>"001001011",
  8924=>"101101111",
  8925=>"000101010",
  8926=>"111100111",
  8927=>"010111101",
  8928=>"111101110",
  8929=>"100110010",
  8930=>"100000101",
  8931=>"001001001",
  8932=>"111000001",
  8933=>"101100000",
  8934=>"010001111",
  8935=>"010011100",
  8936=>"100100001",
  8937=>"001111010",
  8938=>"011111101",
  8939=>"011110000",
  8940=>"010100100",
  8941=>"001110111",
  8942=>"011100010",
  8943=>"011000001",
  8944=>"010011001",
  8945=>"111110100",
  8946=>"000000110",
  8947=>"100101111",
  8948=>"111100100",
  8949=>"010011100",
  8950=>"010010000",
  8951=>"110011001",
  8952=>"100101111",
  8953=>"010010110",
  8954=>"110110100",
  8955=>"011000001",
  8956=>"110001110",
  8957=>"100100010",
  8958=>"001110101",
  8959=>"011010010",
  8960=>"000000111",
  8961=>"111100000",
  8962=>"110110001",
  8963=>"011100010",
  8964=>"101001111",
  8965=>"001011001",
  8966=>"100110010",
  8967=>"001000010",
  8968=>"000000101",
  8969=>"100111111",
  8970=>"011000011",
  8971=>"000000001",
  8972=>"101101010",
  8973=>"110010010",
  8974=>"110000011",
  8975=>"101100010",
  8976=>"010011101",
  8977=>"101101101",
  8978=>"110111001",
  8979=>"111110100",
  8980=>"100101001",
  8981=>"100111010",
  8982=>"110000101",
  8983=>"000100111",
  8984=>"001011011",
  8985=>"110000111",
  8986=>"110110001",
  8987=>"100101101",
  8988=>"010111011",
  8989=>"010011001",
  8990=>"010000111",
  8991=>"000000001",
  8992=>"011100101",
  8993=>"100111100",
  8994=>"111100101",
  8995=>"010111011",
  8996=>"110101110",
  8997=>"100100110",
  8998=>"100010100",
  8999=>"001111111",
  9000=>"001001111",
  9001=>"010101010",
  9002=>"001100111",
  9003=>"010111011",
  9004=>"101110011",
  9005=>"111010010",
  9006=>"001011111",
  9007=>"010011111",
  9008=>"110010111",
  9009=>"000101110",
  9010=>"111011000",
  9011=>"001100111",
  9012=>"011111001",
  9013=>"100000100",
  9014=>"100101101",
  9015=>"000110100",
  9016=>"100001100",
  9017=>"101001011",
  9018=>"100101001",
  9019=>"100100010",
  9020=>"011010010",
  9021=>"000101111",
  9022=>"000001100",
  9023=>"010011001",
  9024=>"110010000",
  9025=>"100001001",
  9026=>"011000101",
  9027=>"010001001",
  9028=>"101000110",
  9029=>"100010010",
  9030=>"111101111",
  9031=>"100011000",
  9032=>"111110111",
  9033=>"011100001",
  9034=>"010110011",
  9035=>"110000100",
  9036=>"001101010",
  9037=>"010110111",
  9038=>"110000111",
  9039=>"111011000",
  9040=>"000111010",
  9041=>"101000011",
  9042=>"001001110",
  9043=>"011010010",
  9044=>"110001001",
  9045=>"000011110",
  9046=>"000100000",
  9047=>"010110011",
  9048=>"100100001",
  9049=>"001100101",
  9050=>"100111000",
  9051=>"101000111",
  9052=>"010000110",
  9053=>"110000000",
  9054=>"000111001",
  9055=>"101011111",
  9056=>"001001010",
  9057=>"001101011",
  9058=>"101010101",
  9059=>"011110010",
  9060=>"001111011",
  9061=>"100011001",
  9062=>"011000100",
  9063=>"100010101",
  9064=>"100000011",
  9065=>"111000000",
  9066=>"111111111",
  9067=>"000101111",
  9068=>"011101001",
  9069=>"001001111",
  9070=>"111010110",
  9071=>"011111100",
  9072=>"010101001",
  9073=>"011011000",
  9074=>"011111111",
  9075=>"001001100",
  9076=>"001010101",
  9077=>"011010000",
  9078=>"010011001",
  9079=>"010011110",
  9080=>"010000000",
  9081=>"110100100",
  9082=>"010111011",
  9083=>"101101011",
  9084=>"011000000",
  9085=>"011000000",
  9086=>"001000101",
  9087=>"110010111",
  9088=>"010111100",
  9089=>"100011100",
  9090=>"010101011",
  9091=>"001011011",
  9092=>"101000000",
  9093=>"011011101",
  9094=>"000011010",
  9095=>"010011001",
  9096=>"100001110",
  9097=>"100110100",
  9098=>"111000001",
  9099=>"111101001",
  9100=>"011000100",
  9101=>"110010010",
  9102=>"011011001",
  9103=>"110011100",
  9104=>"000010111",
  9105=>"110101011",
  9106=>"000000011",
  9107=>"100110011",
  9108=>"011101111",
  9109=>"000100000",
  9110=>"001000001",
  9111=>"100000010",
  9112=>"100010110",
  9113=>"111100101",
  9114=>"110011110",
  9115=>"010100100",
  9116=>"000110010",
  9117=>"000100010",
  9118=>"000101111",
  9119=>"110011000",
  9120=>"011101010",
  9121=>"001001100",
  9122=>"101000100",
  9123=>"000000110",
  9124=>"100001111",
  9125=>"101101001",
  9126=>"001011101",
  9127=>"010110011",
  9128=>"010000100",
  9129=>"101001000",
  9130=>"100000110",
  9131=>"011011110",
  9132=>"010001100",
  9133=>"111011000",
  9134=>"111111100",
  9135=>"010110000",
  9136=>"100011010",
  9137=>"001000010",
  9138=>"011100110",
  9139=>"101111001",
  9140=>"001000100",
  9141=>"011111001",
  9142=>"101001111",
  9143=>"101001011",
  9144=>"001100001",
  9145=>"100110010",
  9146=>"011101110",
  9147=>"011100010",
  9148=>"111111111",
  9149=>"110001110",
  9150=>"000111111",
  9151=>"110000010",
  9152=>"001101101",
  9153=>"100111110",
  9154=>"111001100",
  9155=>"010001111",
  9156=>"010111011",
  9157=>"101010100",
  9158=>"011001001",
  9159=>"111101000",
  9160=>"100111010",
  9161=>"001001001",
  9162=>"100001010",
  9163=>"101101111",
  9164=>"001110111",
  9165=>"011010000",
  9166=>"000100100",
  9167=>"010100000",
  9168=>"111000101",
  9169=>"011000010",
  9170=>"110010001",
  9171=>"011110010",
  9172=>"111001000",
  9173=>"011110011",
  9174=>"010001101",
  9175=>"011101011",
  9176=>"111001100",
  9177=>"111101000",
  9178=>"101100000",
  9179=>"100001001",
  9180=>"000001011",
  9181=>"010110011",
  9182=>"110010001",
  9183=>"000100010",
  9184=>"110010000",
  9185=>"111101110",
  9186=>"100001000",
  9187=>"110011100",
  9188=>"111111101",
  9189=>"000011010",
  9190=>"111000010",
  9191=>"000100101",
  9192=>"001101011",
  9193=>"110111010",
  9194=>"000000111",
  9195=>"101010011",
  9196=>"010101000",
  9197=>"000000010",
  9198=>"110001110",
  9199=>"011100011",
  9200=>"011001111",
  9201=>"000001100",
  9202=>"000110110",
  9203=>"011111101",
  9204=>"101001111",
  9205=>"100111001",
  9206=>"000001000",
  9207=>"111111011",
  9208=>"011001100",
  9209=>"101101111",
  9210=>"110101001",
  9211=>"111010111",
  9212=>"011111011",
  9213=>"000111111",
  9214=>"111110000",
  9215=>"111010001",
  9216=>"010010110",
  9217=>"010010010",
  9218=>"111111111",
  9219=>"110110000",
  9220=>"001111001",
  9221=>"000000011",
  9222=>"000101100",
  9223=>"100101100",
  9224=>"100001101",
  9225=>"011110000",
  9226=>"001001000",
  9227=>"101001111",
  9228=>"011000001",
  9229=>"010110001",
  9230=>"001100010",
  9231=>"001100111",
  9232=>"110101111",
  9233=>"000101101",
  9234=>"101000100",
  9235=>"011100000",
  9236=>"111101111",
  9237=>"011011111",
  9238=>"000001100",
  9239=>"011111001",
  9240=>"101100111",
  9241=>"110111110",
  9242=>"111000101",
  9243=>"000000111",
  9244=>"000001111",
  9245=>"010000011",
  9246=>"111010001",
  9247=>"010100001",
  9248=>"010100011",
  9249=>"110100001",
  9250=>"010000000",
  9251=>"100101000",
  9252=>"011010001",
  9253=>"010111111",
  9254=>"101100001",
  9255=>"001001100",
  9256=>"001101000",
  9257=>"111100101",
  9258=>"101101100",
  9259=>"111111101",
  9260=>"111000101",
  9261=>"111111011",
  9262=>"100011000",
  9263=>"000100010",
  9264=>"111100110",
  9265=>"101000101",
  9266=>"000011111",
  9267=>"000111000",
  9268=>"000010100",
  9269=>"011100110",
  9270=>"111011101",
  9271=>"100010110",
  9272=>"010010110",
  9273=>"011000110",
  9274=>"010000010",
  9275=>"110111111",
  9276=>"000000011",
  9277=>"100110111",
  9278=>"001110100",
  9279=>"110111100",
  9280=>"111110100",
  9281=>"001100001",
  9282=>"111010000",
  9283=>"111111000",
  9284=>"100101100",
  9285=>"111001001",
  9286=>"101010110",
  9287=>"100110010",
  9288=>"000101001",
  9289=>"010000000",
  9290=>"000111110",
  9291=>"011110100",
  9292=>"111110101",
  9293=>"110101000",
  9294=>"001001010",
  9295=>"110000101",
  9296=>"010011010",
  9297=>"000000010",
  9298=>"000101000",
  9299=>"000110011",
  9300=>"001110100",
  9301=>"010101011",
  9302=>"010100111",
  9303=>"001011100",
  9304=>"101010110",
  9305=>"110110100",
  9306=>"100101100",
  9307=>"000011100",
  9308=>"100101110",
  9309=>"101001010",
  9310=>"100011011",
  9311=>"001000011",
  9312=>"000101101",
  9313=>"100101110",
  9314=>"000101110",
  9315=>"000001100",
  9316=>"011100001",
  9317=>"110001101",
  9318=>"000011011",
  9319=>"001111001",
  9320=>"001000011",
  9321=>"101010011",
  9322=>"000001010",
  9323=>"010001001",
  9324=>"110000000",
  9325=>"011010111",
  9326=>"000100101",
  9327=>"110001110",
  9328=>"001000111",
  9329=>"110010101",
  9330=>"011100000",
  9331=>"100010011",
  9332=>"001000010",
  9333=>"101011011",
  9334=>"010101101",
  9335=>"000001111",
  9336=>"011011101",
  9337=>"000001101",
  9338=>"010001100",
  9339=>"001100000",
  9340=>"010101011",
  9341=>"001111000",
  9342=>"100110010",
  9343=>"101001100",
  9344=>"101100100",
  9345=>"110100101",
  9346=>"001110101",
  9347=>"110111100",
  9348=>"001010011",
  9349=>"000110000",
  9350=>"110101100",
  9351=>"011011101",
  9352=>"001111110",
  9353=>"011110111",
  9354=>"101001011",
  9355=>"110011000",
  9356=>"001011100",
  9357=>"001110101",
  9358=>"000000011",
  9359=>"000111001",
  9360=>"111110000",
  9361=>"010101001",
  9362=>"000010100",
  9363=>"110110110",
  9364=>"110100101",
  9365=>"000010000",
  9366=>"101011010",
  9367=>"000110001",
  9368=>"000011001",
  9369=>"100001001",
  9370=>"010010100",
  9371=>"111101111",
  9372=>"100001101",
  9373=>"110111111",
  9374=>"100001110",
  9375=>"111001111",
  9376=>"000100100",
  9377=>"110011010",
  9378=>"101101111",
  9379=>"100111101",
  9380=>"000011111",
  9381=>"111110010",
  9382=>"100110101",
  9383=>"101100001",
  9384=>"001011110",
  9385=>"000110010",
  9386=>"101000010",
  9387=>"001011111",
  9388=>"010100110",
  9389=>"001010101",
  9390=>"000011010",
  9391=>"000100010",
  9392=>"111100100",
  9393=>"000100011",
  9394=>"111001011",
  9395=>"100110100",
  9396=>"001011001",
  9397=>"011010010",
  9398=>"110110010",
  9399=>"111111111",
  9400=>"011100010",
  9401=>"100000111",
  9402=>"100100001",
  9403=>"010010011",
  9404=>"001001000",
  9405=>"000100111",
  9406=>"001000110",
  9407=>"100000000",
  9408=>"111110110",
  9409=>"100111010",
  9410=>"111000101",
  9411=>"010111001",
  9412=>"010010101",
  9413=>"001010001",
  9414=>"001010111",
  9415=>"010100011",
  9416=>"110111000",
  9417=>"111100100",
  9418=>"110100100",
  9419=>"101111100",
  9420=>"011110111",
  9421=>"100000010",
  9422=>"000001000",
  9423=>"100001101",
  9424=>"011010010",
  9425=>"001110000",
  9426=>"110011100",
  9427=>"100010010",
  9428=>"010000011",
  9429=>"010110010",
  9430=>"000010100",
  9431=>"011101111",
  9432=>"101111000",
  9433=>"000001111",
  9434=>"000011100",
  9435=>"010000001",
  9436=>"100000001",
  9437=>"001100111",
  9438=>"100111110",
  9439=>"010000010",
  9440=>"000000000",
  9441=>"111011000",
  9442=>"000001000",
  9443=>"000001001",
  9444=>"101011100",
  9445=>"111111001",
  9446=>"110011110",
  9447=>"100101100",
  9448=>"101110010",
  9449=>"111010110",
  9450=>"001100100",
  9451=>"000001000",
  9452=>"000100011",
  9453=>"001011100",
  9454=>"111100010",
  9455=>"111001010",
  9456=>"110111000",
  9457=>"011111011",
  9458=>"101100010",
  9459=>"001001011",
  9460=>"011001010",
  9461=>"110010001",
  9462=>"100100010",
  9463=>"000111110",
  9464=>"011111001",
  9465=>"110000011",
  9466=>"000101100",
  9467=>"111101100",
  9468=>"001010011",
  9469=>"011001100",
  9470=>"111011011",
  9471=>"011000101",
  9472=>"111110011",
  9473=>"001111000",
  9474=>"110111111",
  9475=>"110110011",
  9476=>"000001110",
  9477=>"101111100",
  9478=>"000011111",
  9479=>"110000100",
  9480=>"000010100",
  9481=>"001010001",
  9482=>"000000111",
  9483=>"001100111",
  9484=>"001000001",
  9485=>"001011101",
  9486=>"100001011",
  9487=>"000001011",
  9488=>"010101100",
  9489=>"011011101",
  9490=>"000111110",
  9491=>"101111111",
  9492=>"011011100",
  9493=>"111111100",
  9494=>"000001011",
  9495=>"101111111",
  9496=>"111000100",
  9497=>"110001011",
  9498=>"010111111",
  9499=>"001010010",
  9500=>"111101010",
  9501=>"111001000",
  9502=>"000010100",
  9503=>"000010110",
  9504=>"000000010",
  9505=>"011110010",
  9506=>"111111111",
  9507=>"100111001",
  9508=>"011110111",
  9509=>"111100101",
  9510=>"000111101",
  9511=>"101110010",
  9512=>"000000111",
  9513=>"111110111",
  9514=>"000111000",
  9515=>"110101101",
  9516=>"110110011",
  9517=>"010010110",
  9518=>"000010100",
  9519=>"011101110",
  9520=>"101110100",
  9521=>"101010010",
  9522=>"111110011",
  9523=>"101001111",
  9524=>"001100001",
  9525=>"110010101",
  9526=>"011111000",
  9527=>"011100011",
  9528=>"000100000",
  9529=>"101101000",
  9530=>"011011001",
  9531=>"101111110",
  9532=>"010000111",
  9533=>"001110010",
  9534=>"100010101",
  9535=>"100100011",
  9536=>"111111010",
  9537=>"110100001",
  9538=>"011010111",
  9539=>"110111111",
  9540=>"100100001",
  9541=>"000110100",
  9542=>"111011000",
  9543=>"010011001",
  9544=>"011011100",
  9545=>"111101110",
  9546=>"100110011",
  9547=>"100111011",
  9548=>"000001110",
  9549=>"000000111",
  9550=>"010111000",
  9551=>"001111011",
  9552=>"111110100",
  9553=>"100000000",
  9554=>"001110010",
  9555=>"000001111",
  9556=>"010010101",
  9557=>"101111001",
  9558=>"110100000",
  9559=>"001100001",
  9560=>"011011000",
  9561=>"101001100",
  9562=>"000101001",
  9563=>"101011110",
  9564=>"101010000",
  9565=>"100100001",
  9566=>"111101011",
  9567=>"011111011",
  9568=>"110110011",
  9569=>"110011001",
  9570=>"011110011",
  9571=>"011111100",
  9572=>"001111100",
  9573=>"110011101",
  9574=>"010000111",
  9575=>"111010000",
  9576=>"100110001",
  9577=>"110011101",
  9578=>"111001011",
  9579=>"110110010",
  9580=>"111001010",
  9581=>"011000011",
  9582=>"100110010",
  9583=>"101010011",
  9584=>"001100100",
  9585=>"101001001",
  9586=>"100100110",
  9587=>"011100100",
  9588=>"111101110",
  9589=>"100001100",
  9590=>"001000001",
  9591=>"010101100",
  9592=>"101010101",
  9593=>"110100000",
  9594=>"111110100",
  9595=>"000110100",
  9596=>"011101111",
  9597=>"100001100",
  9598=>"110011101",
  9599=>"001101110",
  9600=>"110111101",
  9601=>"111001100",
  9602=>"001001101",
  9603=>"101111101",
  9604=>"011010111",
  9605=>"101001110",
  9606=>"111001010",
  9607=>"000010001",
  9608=>"000010010",
  9609=>"011000101",
  9610=>"001000100",
  9611=>"011111010",
  9612=>"100101100",
  9613=>"011110000",
  9614=>"000010101",
  9615=>"000111111",
  9616=>"100100100",
  9617=>"001000101",
  9618=>"100010100",
  9619=>"001110111",
  9620=>"110110000",
  9621=>"101001000",
  9622=>"101011110",
  9623=>"010101110",
  9624=>"100110100",
  9625=>"010101000",
  9626=>"010110001",
  9627=>"010111111",
  9628=>"001111100",
  9629=>"011100111",
  9630=>"001100000",
  9631=>"110010000",
  9632=>"110000110",
  9633=>"010010011",
  9634=>"110111111",
  9635=>"110110110",
  9636=>"111110010",
  9637=>"011010000",
  9638=>"001011111",
  9639=>"101110010",
  9640=>"100010000",
  9641=>"111001101",
  9642=>"110000110",
  9643=>"000000001",
  9644=>"010001111",
  9645=>"110101111",
  9646=>"111010010",
  9647=>"001011000",
  9648=>"001111110",
  9649=>"001000001",
  9650=>"111011001",
  9651=>"111111000",
  9652=>"100111101",
  9653=>"101100100",
  9654=>"101010111",
  9655=>"001000011",
  9656=>"001000011",
  9657=>"101101011",
  9658=>"000010001",
  9659=>"001101111",
  9660=>"111001000",
  9661=>"111101011",
  9662=>"000001000",
  9663=>"010010000",
  9664=>"001000010",
  9665=>"100010110",
  9666=>"111101011",
  9667=>"001000010",
  9668=>"000001000",
  9669=>"101101110",
  9670=>"000111001",
  9671=>"101111011",
  9672=>"100010011",
  9673=>"001001110",
  9674=>"000110010",
  9675=>"001100001",
  9676=>"111111010",
  9677=>"100000000",
  9678=>"110110100",
  9679=>"111100011",
  9680=>"001000000",
  9681=>"100000010",
  9682=>"011100001",
  9683=>"101101111",
  9684=>"110001101",
  9685=>"100000011",
  9686=>"100000001",
  9687=>"111101100",
  9688=>"111000111",
  9689=>"011100010",
  9690=>"010001100",
  9691=>"101000101",
  9692=>"000100001",
  9693=>"000011110",
  9694=>"111011010",
  9695=>"110011111",
  9696=>"011000111",
  9697=>"110010110",
  9698=>"000011101",
  9699=>"101001011",
  9700=>"010110011",
  9701=>"111111101",
  9702=>"100110011",
  9703=>"101000101",
  9704=>"110001010",
  9705=>"110110011",
  9706=>"101001110",
  9707=>"100011001",
  9708=>"101000001",
  9709=>"101111110",
  9710=>"111100110",
  9711=>"010011110",
  9712=>"010100000",
  9713=>"110101110",
  9714=>"110111001",
  9715=>"110110010",
  9716=>"111111111",
  9717=>"101110101",
  9718=>"010001001",
  9719=>"011110100",
  9720=>"000010110",
  9721=>"111110100",
  9722=>"100110111",
  9723=>"110000000",
  9724=>"110111111",
  9725=>"011010100",
  9726=>"110111110",
  9727=>"100010010",
  9728=>"001100111",
  9729=>"101000111",
  9730=>"101111111",
  9731=>"000001100",
  9732=>"011110001",
  9733=>"010101110",
  9734=>"110010010",
  9735=>"111011010",
  9736=>"111010111",
  9737=>"001010100",
  9738=>"100000110",
  9739=>"011100101",
  9740=>"110111001",
  9741=>"111000111",
  9742=>"100001001",
  9743=>"010001101",
  9744=>"101000001",
  9745=>"000001000",
  9746=>"100111000",
  9747=>"101011110",
  9748=>"011001000",
  9749=>"011011101",
  9750=>"110110011",
  9751=>"011001100",
  9752=>"101110001",
  9753=>"110000001",
  9754=>"101000000",
  9755=>"000001101",
  9756=>"011101010",
  9757=>"000011100",
  9758=>"011110000",
  9759=>"010110111",
  9760=>"000100011",
  9761=>"010001001",
  9762=>"111001100",
  9763=>"011111100",
  9764=>"011110011",
  9765=>"011100000",
  9766=>"000100011",
  9767=>"110110010",
  9768=>"111010010",
  9769=>"001101001",
  9770=>"011010100",
  9771=>"111101000",
  9772=>"110010111",
  9773=>"111110101",
  9774=>"111011111",
  9775=>"111010111",
  9776=>"000101101",
  9777=>"110011010",
  9778=>"011001101",
  9779=>"001010110",
  9780=>"111100101",
  9781=>"111000000",
  9782=>"111100010",
  9783=>"000101001",
  9784=>"111111001",
  9785=>"010111100",
  9786=>"111100000",
  9787=>"111000010",
  9788=>"011000001",
  9789=>"010000101",
  9790=>"000111001",
  9791=>"100010011",
  9792=>"101101101",
  9793=>"000001001",
  9794=>"010001100",
  9795=>"000111001",
  9796=>"000000111",
  9797=>"000001001",
  9798=>"010001110",
  9799=>"011001000",
  9800=>"000000110",
  9801=>"000000110",
  9802=>"110001100",
  9803=>"101011010",
  9804=>"011100010",
  9805=>"001100000",
  9806=>"101010110",
  9807=>"100101111",
  9808=>"111001101",
  9809=>"000100101",
  9810=>"001011010",
  9811=>"010100000",
  9812=>"000011001",
  9813=>"000010111",
  9814=>"111010111",
  9815=>"000101011",
  9816=>"011010010",
  9817=>"011010110",
  9818=>"000010000",
  9819=>"111010010",
  9820=>"101011111",
  9821=>"110001100",
  9822=>"011000000",
  9823=>"010000000",
  9824=>"001101001",
  9825=>"010001000",
  9826=>"111011100",
  9827=>"011001011",
  9828=>"100100100",
  9829=>"111100100",
  9830=>"011000000",
  9831=>"100100101",
  9832=>"010111010",
  9833=>"001111001",
  9834=>"101100000",
  9835=>"101001010",
  9836=>"111000111",
  9837=>"000111110",
  9838=>"110000111",
  9839=>"010011111",
  9840=>"001011010",
  9841=>"000000010",
  9842=>"110011011",
  9843=>"010101100",
  9844=>"100011111",
  9845=>"100001001",
  9846=>"011111111",
  9847=>"001100011",
  9848=>"101010100",
  9849=>"111000011",
  9850=>"110001010",
  9851=>"111110010",
  9852=>"000100000",
  9853=>"011001101",
  9854=>"011111001",
  9855=>"011000010",
  9856=>"001011010",
  9857=>"100001110",
  9858=>"110101101",
  9859=>"111001111",
  9860=>"000010101",
  9861=>"111111011",
  9862=>"000000010",
  9863=>"100011111",
  9864=>"011011111",
  9865=>"010001101",
  9866=>"111111011",
  9867=>"100110011",
  9868=>"000111000",
  9869=>"111110011",
  9870=>"111001010",
  9871=>"001000000",
  9872=>"001000110",
  9873=>"011110001",
  9874=>"001101100",
  9875=>"110011100",
  9876=>"000000011",
  9877=>"001110000",
  9878=>"111010000",
  9879=>"010100110",
  9880=>"110111011",
  9881=>"011111000",
  9882=>"111000011",
  9883=>"001100100",
  9884=>"001011100",
  9885=>"101000100",
  9886=>"101111010",
  9887=>"101110110",
  9888=>"011000100",
  9889=>"000011011",
  9890=>"010000100",
  9891=>"011000001",
  9892=>"000100010",
  9893=>"101011110",
  9894=>"100010110",
  9895=>"011001110",
  9896=>"111111101",
  9897=>"000100111",
  9898=>"111011101",
  9899=>"011010011",
  9900=>"001010001",
  9901=>"100000100",
  9902=>"110001010",
  9903=>"100011010",
  9904=>"011011100",
  9905=>"100001010",
  9906=>"001011000",
  9907=>"001010010",
  9908=>"010010011",
  9909=>"010001011",
  9910=>"101101000",
  9911=>"110010001",
  9912=>"111111000",
  9913=>"101000000",
  9914=>"111000110",
  9915=>"110111011",
  9916=>"001010000",
  9917=>"000001110",
  9918=>"001010101",
  9919=>"111001111",
  9920=>"110100101",
  9921=>"100111101",
  9922=>"001011001",
  9923=>"011100100",
  9924=>"101011101",
  9925=>"111001011",
  9926=>"100101011",
  9927=>"010101000",
  9928=>"011010001",
  9929=>"001101101",
  9930=>"101010110",
  9931=>"011111110",
  9932=>"011011101",
  9933=>"101010010",
  9934=>"001110010",
  9935=>"101001000",
  9936=>"000110000",
  9937=>"100111000",
  9938=>"111011101",
  9939=>"010010101",
  9940=>"010100110",
  9941=>"000010001",
  9942=>"000001010",
  9943=>"111100110",
  9944=>"000010100",
  9945=>"100100101",
  9946=>"111111101",
  9947=>"011111101",
  9948=>"011111010",
  9949=>"111101010",
  9950=>"100110000",
  9951=>"100010101",
  9952=>"010101110",
  9953=>"000001100",
  9954=>"111110001",
  9955=>"000000100",
  9956=>"111011011",
  9957=>"100000101",
  9958=>"100110001",
  9959=>"001000000",
  9960=>"100010100",
  9961=>"110111101",
  9962=>"111110100",
  9963=>"000111101",
  9964=>"011111110",
  9965=>"101000111",
  9966=>"101000100",
  9967=>"100000011",
  9968=>"100010101",
  9969=>"010111100",
  9970=>"010001111",
  9971=>"000001101",
  9972=>"001101101",
  9973=>"001100011",
  9974=>"110101010",
  9975=>"011010011",
  9976=>"100110001",
  9977=>"110110101",
  9978=>"001110010",
  9979=>"010111010",
  9980=>"011000111",
  9981=>"011000010",
  9982=>"101111011",
  9983=>"010101010",
  9984=>"111111101",
  9985=>"000010011",
  9986=>"101110101",
  9987=>"011100110",
  9988=>"011110100",
  9989=>"100100011",
  9990=>"110101111",
  9991=>"111011011",
  9992=>"001001011",
  9993=>"000001010",
  9994=>"001001010",
  9995=>"011100000",
  9996=>"000110000",
  9997=>"010011000",
  9998=>"110110100",
  9999=>"001010100",
  10000=>"010111001",
  10001=>"101001000",
  10002=>"000001110",
  10003=>"011010001",
  10004=>"110101101",
  10005=>"010010101",
  10006=>"011110110",
  10007=>"101110101",
  10008=>"010010100",
  10009=>"010100110",
  10010=>"000010100",
  10011=>"011101111",
  10012=>"001110110",
  10013=>"001001100",
  10014=>"001011001",
  10015=>"101110101",
  10016=>"000101010",
  10017=>"111010101",
  10018=>"001000011",
  10019=>"001011100",
  10020=>"000001000",
  10021=>"010010101",
  10022=>"001110011",
  10023=>"001010111",
  10024=>"011101011",
  10025=>"110110000",
  10026=>"011010010",
  10027=>"101011110",
  10028=>"111000101",
  10029=>"101110100",
  10030=>"111010000",
  10031=>"111010101",
  10032=>"000101001",
  10033=>"101001001",
  10034=>"011011110",
  10035=>"000011100",
  10036=>"001011000",
  10037=>"000111000",
  10038=>"011100010",
  10039=>"000000111",
  10040=>"101100011",
  10041=>"011011010",
  10042=>"101000100",
  10043=>"010101101",
  10044=>"000000000",
  10045=>"101001000",
  10046=>"010111110",
  10047=>"000001110",
  10048=>"110111110",
  10049=>"010100110",
  10050=>"111000100",
  10051=>"011111000",
  10052=>"000110100",
  10053=>"011111011",
  10054=>"111101000",
  10055=>"011011010",
  10056=>"110000010",
  10057=>"100111101",
  10058=>"110111001",
  10059=>"001000101",
  10060=>"010011000",
  10061=>"101101100",
  10062=>"111000010",
  10063=>"111010111",
  10064=>"010110111",
  10065=>"101010011",
  10066=>"000011100",
  10067=>"010101001",
  10068=>"010001100",
  10069=>"110001011",
  10070=>"001001101",
  10071=>"101011100",
  10072=>"011110000",
  10073=>"111010100",
  10074=>"111011010",
  10075=>"100100000",
  10076=>"111000101",
  10077=>"101011010",
  10078=>"100011100",
  10079=>"111010100",
  10080=>"000101110",
  10081=>"110110011",
  10082=>"100101000",
  10083=>"010111111",
  10084=>"010000101",
  10085=>"010001001",
  10086=>"001110000",
  10087=>"100100101",
  10088=>"110001001",
  10089=>"111010010",
  10090=>"110001010",
  10091=>"000110110",
  10092=>"100111011",
  10093=>"000010011",
  10094=>"100101000",
  10095=>"000111100",
  10096=>"101111000",
  10097=>"000101000",
  10098=>"000111001",
  10099=>"110101101",
  10100=>"101000000",
  10101=>"100100010",
  10102=>"000010111",
  10103=>"011101000",
  10104=>"101111010",
  10105=>"100100000",
  10106=>"000101100",
  10107=>"111101001",
  10108=>"101000010",
  10109=>"111101010",
  10110=>"100100010",
  10111=>"111110010",
  10112=>"101110011",
  10113=>"010011101",
  10114=>"011000010",
  10115=>"000011101",
  10116=>"010110000",
  10117=>"011010100",
  10118=>"101011100",
  10119=>"001000100",
  10120=>"100010110",
  10121=>"111001101",
  10122=>"000110111",
  10123=>"001000101",
  10124=>"101001110",
  10125=>"101110111",
  10126=>"100000011",
  10127=>"111000000",
  10128=>"001110111",
  10129=>"100000111",
  10130=>"011101100",
  10131=>"110001101",
  10132=>"111000100",
  10133=>"010001100",
  10134=>"101110010",
  10135=>"111100111",
  10136=>"000011100",
  10137=>"101101010",
  10138=>"100011000",
  10139=>"101100100",
  10140=>"111000100",
  10141=>"000100001",
  10142=>"010011010",
  10143=>"111110011",
  10144=>"111111111",
  10145=>"001101001",
  10146=>"111011110",
  10147=>"111110100",
  10148=>"000100100",
  10149=>"111101010",
  10150=>"100100110",
  10151=>"100001000",
  10152=>"110011101",
  10153=>"000000111",
  10154=>"001011110",
  10155=>"101101100",
  10156=>"000111111",
  10157=>"101010111",
  10158=>"110011101",
  10159=>"000010000",
  10160=>"000010101",
  10161=>"101011111",
  10162=>"110010100",
  10163=>"111011111",
  10164=>"111110111",
  10165=>"111101110",
  10166=>"000000100",
  10167=>"000001000",
  10168=>"010001111",
  10169=>"000010110",
  10170=>"001001001",
  10171=>"100011010",
  10172=>"000111000",
  10173=>"100001101",
  10174=>"000001100",
  10175=>"010111010",
  10176=>"001111111",
  10177=>"101100001",
  10178=>"111010010",
  10179=>"111100001",
  10180=>"001000010",
  10181=>"101011000",
  10182=>"001100111",
  10183=>"101000010",
  10184=>"010100010",
  10185=>"110000011",
  10186=>"101001001",
  10187=>"110011010",
  10188=>"000100001",
  10189=>"100100010",
  10190=>"110011001",
  10191=>"010100101",
  10192=>"101010000",
  10193=>"100110110",
  10194=>"000001110",
  10195=>"000000000",
  10196=>"111110001",
  10197=>"111011100",
  10198=>"100101010",
  10199=>"001001100",
  10200=>"100100110",
  10201=>"011100100",
  10202=>"100110001",
  10203=>"101111010",
  10204=>"100011100",
  10205=>"101010111",
  10206=>"010010110",
  10207=>"100010001",
  10208=>"010011000",
  10209=>"011001000",
  10210=>"101111101",
  10211=>"101111101",
  10212=>"001111000",
  10213=>"111100110",
  10214=>"110100110",
  10215=>"110001001",
  10216=>"001010010",
  10217=>"001100101",
  10218=>"101011111",
  10219=>"110010111",
  10220=>"001011001",
  10221=>"100111010",
  10222=>"101011100",
  10223=>"101101001",
  10224=>"101110001",
  10225=>"011001001",
  10226=>"011110000",
  10227=>"100000010",
  10228=>"011100110",
  10229=>"101000010",
  10230=>"110111110",
  10231=>"110100100",
  10232=>"110000110",
  10233=>"100110001",
  10234=>"011001011",
  10235=>"001001101",
  10236=>"101011010",
  10237=>"100001001",
  10238=>"111110110",
  10239=>"001011101",
  10240=>"101101011",
  10241=>"010011100",
  10242=>"111000101",
  10243=>"101010110",
  10244=>"110111100",
  10245=>"011110101",
  10246=>"111100110",
  10247=>"011001111",
  10248=>"001111011",
  10249=>"100000011",
  10250=>"000000110",
  10251=>"110011111",
  10252=>"010101011",
  10253=>"110011000",
  10254=>"000111010",
  10255=>"111101110",
  10256=>"001110010",
  10257=>"001011011",
  10258=>"100000010",
  10259=>"000010001",
  10260=>"111010100",
  10261=>"111110000",
  10262=>"001110111",
  10263=>"000010100",
  10264=>"000001011",
  10265=>"011101000",
  10266=>"100001100",
  10267=>"100100010",
  10268=>"010100010",
  10269=>"111011111",
  10270=>"000000101",
  10271=>"010110100",
  10272=>"101001110",
  10273=>"101100101",
  10274=>"000001110",
  10275=>"101000100",
  10276=>"101100110",
  10277=>"010110101",
  10278=>"100111101",
  10279=>"100011011",
  10280=>"011010110",
  10281=>"010100010",
  10282=>"011001011",
  10283=>"010111101",
  10284=>"110101101",
  10285=>"011110011",
  10286=>"111000000",
  10287=>"011100111",
  10288=>"001011000",
  10289=>"000000001",
  10290=>"011110011",
  10291=>"100001000",
  10292=>"100001111",
  10293=>"010001101",
  10294=>"000001001",
  10295=>"110111111",
  10296=>"000010010",
  10297=>"110101000",
  10298=>"101110111",
  10299=>"101101100",
  10300=>"010011101",
  10301=>"100000110",
  10302=>"110100011",
  10303=>"010110100",
  10304=>"110011111",
  10305=>"000101000",
  10306=>"010011001",
  10307=>"001111001",
  10308=>"100000101",
  10309=>"100111111",
  10310=>"110001000",
  10311=>"000110000",
  10312=>"111011000",
  10313=>"000001000",
  10314=>"110001100",
  10315=>"101101110",
  10316=>"010101101",
  10317=>"110100010",
  10318=>"111001100",
  10319=>"011010100",
  10320=>"101111011",
  10321=>"011100010",
  10322=>"001110010",
  10323=>"011011111",
  10324=>"010001100",
  10325=>"110001101",
  10326=>"011001100",
  10327=>"101001000",
  10328=>"001111101",
  10329=>"011111101",
  10330=>"000110111",
  10331=>"111000111",
  10332=>"011001101",
  10333=>"101011001",
  10334=>"100001101",
  10335=>"011000011",
  10336=>"111101000",
  10337=>"011100000",
  10338=>"001100101",
  10339=>"000011000",
  10340=>"001101000",
  10341=>"110000110",
  10342=>"010110000",
  10343=>"001011100",
  10344=>"111100100",
  10345=>"110011110",
  10346=>"100001110",
  10347=>"101110110",
  10348=>"101101101",
  10349=>"111101001",
  10350=>"100011111",
  10351=>"000111010",
  10352=>"010000110",
  10353=>"011011101",
  10354=>"001101001",
  10355=>"111111011",
  10356=>"011111011",
  10357=>"000000101",
  10358=>"111100100",
  10359=>"010111111",
  10360=>"011100011",
  10361=>"110111100",
  10362=>"010001101",
  10363=>"110100010",
  10364=>"100001010",
  10365=>"001011111",
  10366=>"111010000",
  10367=>"000110011",
  10368=>"100001110",
  10369=>"001111000",
  10370=>"000111010",
  10371=>"010010111",
  10372=>"100111100",
  10373=>"101110111",
  10374=>"101001000",
  10375=>"111000001",
  10376=>"100010110",
  10377=>"101100000",
  10378=>"010000001",
  10379=>"100100100",
  10380=>"100110110",
  10381=>"101100110",
  10382=>"000011001",
  10383=>"010110111",
  10384=>"101011101",
  10385=>"000011110",
  10386=>"010000011",
  10387=>"010000010",
  10388=>"001101110",
  10389=>"000010000",
  10390=>"000011100",
  10391=>"101100111",
  10392=>"000101111",
  10393=>"101010101",
  10394=>"101110100",
  10395=>"010111010",
  10396=>"001101110",
  10397=>"110001100",
  10398=>"100100000",
  10399=>"111110000",
  10400=>"110011100",
  10401=>"000011111",
  10402=>"111100001",
  10403=>"000100001",
  10404=>"101000110",
  10405=>"000111110",
  10406=>"100001101",
  10407=>"100100000",
  10408=>"110110110",
  10409=>"101111011",
  10410=>"001101110",
  10411=>"001110100",
  10412=>"101010010",
  10413=>"101000000",
  10414=>"100101010",
  10415=>"111110111",
  10416=>"011011100",
  10417=>"000000101",
  10418=>"001100001",
  10419=>"011010000",
  10420=>"000000001",
  10421=>"101001110",
  10422=>"100111111",
  10423=>"111000000",
  10424=>"101011101",
  10425=>"111110110",
  10426=>"101100101",
  10427=>"101101111",
  10428=>"011111101",
  10429=>"111101001",
  10430=>"111000001",
  10431=>"010110111",
  10432=>"111001100",
  10433=>"111100011",
  10434=>"110110101",
  10435=>"011100011",
  10436=>"001000111",
  10437=>"000000011",
  10438=>"010011011",
  10439=>"000001010",
  10440=>"011010100",
  10441=>"100110010",
  10442=>"010100001",
  10443=>"010000011",
  10444=>"100000110",
  10445=>"101001000",
  10446=>"101000110",
  10447=>"101111010",
  10448=>"000000000",
  10449=>"000011100",
  10450=>"010000101",
  10451=>"110011000",
  10452=>"001001101",
  10453=>"001111110",
  10454=>"110110010",
  10455=>"110010101",
  10456=>"111001111",
  10457=>"011000001",
  10458=>"100100100",
  10459=>"000100110",
  10460=>"000111000",
  10461=>"110101011",
  10462=>"110110011",
  10463=>"000101100",
  10464=>"110010110",
  10465=>"010001001",
  10466=>"100001111",
  10467=>"010010101",
  10468=>"110110110",
  10469=>"101011010",
  10470=>"110100101",
  10471=>"001011010",
  10472=>"110011110",
  10473=>"010010000",
  10474=>"001001001",
  10475=>"111000101",
  10476=>"010100111",
  10477=>"000011001",
  10478=>"000100111",
  10479=>"101101000",
  10480=>"000001110",
  10481=>"010000010",
  10482=>"101000010",
  10483=>"010001110",
  10484=>"100001110",
  10485=>"101000010",
  10486=>"010010110",
  10487=>"100100101",
  10488=>"100101111",
  10489=>"100011000",
  10490=>"010101101",
  10491=>"000101011",
  10492=>"010110010",
  10493=>"100010001",
  10494=>"110110011",
  10495=>"110100111",
  10496=>"001011111",
  10497=>"100001100",
  10498=>"100100110",
  10499=>"010110011",
  10500=>"001000010",
  10501=>"000100111",
  10502=>"110111001",
  10503=>"011000000",
  10504=>"011001010",
  10505=>"111010111",
  10506=>"110010101",
  10507=>"101000101",
  10508=>"110110110",
  10509=>"111101010",
  10510=>"001101101",
  10511=>"000101001",
  10512=>"010110110",
  10513=>"011000110",
  10514=>"011010000",
  10515=>"111011101",
  10516=>"100000110",
  10517=>"010101101",
  10518=>"101000010",
  10519=>"011111110",
  10520=>"011011111",
  10521=>"100100111",
  10522=>"101100111",
  10523=>"110111111",
  10524=>"010001011",
  10525=>"110000000",
  10526=>"110011111",
  10527=>"001010010",
  10528=>"000100000",
  10529=>"110001001",
  10530=>"010001110",
  10531=>"101000010",
  10532=>"001110100",
  10533=>"111100001",
  10534=>"110110011",
  10535=>"101101101",
  10536=>"101010111",
  10537=>"011001100",
  10538=>"010110111",
  10539=>"101001011",
  10540=>"100011110",
  10541=>"000100100",
  10542=>"001111010",
  10543=>"100111110",
  10544=>"011000101",
  10545=>"110010111",
  10546=>"111111110",
  10547=>"010000000",
  10548=>"001010010",
  10549=>"001001101",
  10550=>"011011110",
  10551=>"101001110",
  10552=>"000011010",
  10553=>"001101110",
  10554=>"100100100",
  10555=>"001000011",
  10556=>"010101111",
  10557=>"111000000",
  10558=>"110111011",
  10559=>"100010111",
  10560=>"010011110",
  10561=>"100010101",
  10562=>"000101000",
  10563=>"111001101",
  10564=>"011011110",
  10565=>"100011111",
  10566=>"010110100",
  10567=>"101011000",
  10568=>"100111000",
  10569=>"101101001",
  10570=>"011111001",
  10571=>"101011111",
  10572=>"010110011",
  10573=>"011111110",
  10574=>"101001011",
  10575=>"000011001",
  10576=>"010111111",
  10577=>"110111111",
  10578=>"010100001",
  10579=>"101010110",
  10580=>"000111010",
  10581=>"110010000",
  10582=>"000011011",
  10583=>"000111010",
  10584=>"000111110",
  10585=>"101010111",
  10586=>"011000000",
  10587=>"101001001",
  10588=>"010001010",
  10589=>"100111010",
  10590=>"010011010",
  10591=>"000111000",
  10592=>"000000001",
  10593=>"010000110",
  10594=>"100101100",
  10595=>"100001011",
  10596=>"100010110",
  10597=>"010000011",
  10598=>"011000111",
  10599=>"011011111",
  10600=>"110010000",
  10601=>"001000111",
  10602=>"000110101",
  10603=>"111011110",
  10604=>"101011100",
  10605=>"001101001",
  10606=>"111000000",
  10607=>"000101000",
  10608=>"101101000",
  10609=>"111000111",
  10610=>"111101010",
  10611=>"110010111",
  10612=>"101111001",
  10613=>"101111111",
  10614=>"011000100",
  10615=>"001110110",
  10616=>"000010111",
  10617=>"000001110",
  10618=>"000001001",
  10619=>"111111111",
  10620=>"010100011",
  10621=>"110001110",
  10622=>"001010100",
  10623=>"000101000",
  10624=>"001001101",
  10625=>"110010100",
  10626=>"011001010",
  10627=>"000000010",
  10628=>"001110000",
  10629=>"110010100",
  10630=>"111100011",
  10631=>"000001100",
  10632=>"111010010",
  10633=>"011000000",
  10634=>"000011010",
  10635=>"000100011",
  10636=>"101110001",
  10637=>"111101100",
  10638=>"110011100",
  10639=>"011001100",
  10640=>"100011110",
  10641=>"000011011",
  10642=>"010011010",
  10643=>"101001111",
  10644=>"110101001",
  10645=>"010101101",
  10646=>"000101111",
  10647=>"111010001",
  10648=>"010110110",
  10649=>"101000001",
  10650=>"111101000",
  10651=>"101000101",
  10652=>"101011111",
  10653=>"101101011",
  10654=>"001010101",
  10655=>"101111010",
  10656=>"001111101",
  10657=>"111010100",
  10658=>"010111010",
  10659=>"010111010",
  10660=>"011010000",
  10661=>"000000111",
  10662=>"100011001",
  10663=>"010011011",
  10664=>"111011100",
  10665=>"110000111",
  10666=>"100001010",
  10667=>"011101101",
  10668=>"001110000",
  10669=>"001011010",
  10670=>"101101101",
  10671=>"111011001",
  10672=>"101111100",
  10673=>"110111100",
  10674=>"000000111",
  10675=>"011110010",
  10676=>"110001100",
  10677=>"011010010",
  10678=>"111011101",
  10679=>"000000110",
  10680=>"101000000",
  10681=>"010111111",
  10682=>"000110001",
  10683=>"000110100",
  10684=>"000001100",
  10685=>"111010010",
  10686=>"010101100",
  10687=>"011111110",
  10688=>"100001001",
  10689=>"110111010",
  10690=>"111110010",
  10691=>"001110100",
  10692=>"100010011",
  10693=>"111100000",
  10694=>"111111101",
  10695=>"110000100",
  10696=>"111111001",
  10697=>"101111010",
  10698=>"001000001",
  10699=>"110110101",
  10700=>"011001101",
  10701=>"001101110",
  10702=>"010010000",
  10703=>"101010111",
  10704=>"111100010",
  10705=>"011011100",
  10706=>"011010111",
  10707=>"010011011",
  10708=>"001000011",
  10709=>"010010001",
  10710=>"001001010",
  10711=>"110100010",
  10712=>"101100111",
  10713=>"000110001",
  10714=>"011110111",
  10715=>"100011111",
  10716=>"110111111",
  10717=>"000100011",
  10718=>"110001110",
  10719=>"010100011",
  10720=>"110110010",
  10721=>"110111100",
  10722=>"010111111",
  10723=>"101111011",
  10724=>"010101011",
  10725=>"111011000",
  10726=>"110000001",
  10727=>"001111001",
  10728=>"011110110",
  10729=>"011110111",
  10730=>"001100111",
  10731=>"001000111",
  10732=>"011110011",
  10733=>"000001101",
  10734=>"011101100",
  10735=>"101111010",
  10736=>"001110011",
  10737=>"111111011",
  10738=>"000011001",
  10739=>"111100111",
  10740=>"100011011",
  10741=>"010000000",
  10742=>"111100100",
  10743=>"100101001",
  10744=>"100000000",
  10745=>"111010111",
  10746=>"011111001",
  10747=>"000100111",
  10748=>"010000000",
  10749=>"001110010",
  10750=>"001101010",
  10751=>"111000101",
  10752=>"111111111",
  10753=>"011001100",
  10754=>"011101011",
  10755=>"000101001",
  10756=>"010100110",
  10757=>"001010000",
  10758=>"000001001",
  10759=>"000010010",
  10760=>"001101001",
  10761=>"010110100",
  10762=>"010011110",
  10763=>"101101100",
  10764=>"101010000",
  10765=>"001110101",
  10766=>"111100000",
  10767=>"011000100",
  10768=>"010111010",
  10769=>"000010000",
  10770=>"011100111",
  10771=>"110111001",
  10772=>"110011111",
  10773=>"111011110",
  10774=>"001100111",
  10775=>"100101110",
  10776=>"000111101",
  10777=>"111011111",
  10778=>"001000010",
  10779=>"011111111",
  10780=>"111111010",
  10781=>"110100001",
  10782=>"000111001",
  10783=>"011000000",
  10784=>"110010000",
  10785=>"110011001",
  10786=>"000101010",
  10787=>"111000111",
  10788=>"111100010",
  10789=>"001101110",
  10790=>"101100001",
  10791=>"011000101",
  10792=>"111111001",
  10793=>"001010111",
  10794=>"001011010",
  10795=>"011100100",
  10796=>"011011111",
  10797=>"011110001",
  10798=>"001010011",
  10799=>"101101100",
  10800=>"100001001",
  10801=>"011010110",
  10802=>"001111110",
  10803=>"010001110",
  10804=>"100011110",
  10805=>"010010100",
  10806=>"100111001",
  10807=>"101110011",
  10808=>"111000011",
  10809=>"100101010",
  10810=>"110110110",
  10811=>"110001110",
  10812=>"110111010",
  10813=>"101001101",
  10814=>"010110111",
  10815=>"110000000",
  10816=>"000111000",
  10817=>"011101000",
  10818=>"000100001",
  10819=>"011111101",
  10820=>"110001110",
  10821=>"101101001",
  10822=>"001100110",
  10823=>"111000000",
  10824=>"001111010",
  10825=>"110000100",
  10826=>"111000001",
  10827=>"011101011",
  10828=>"100110100",
  10829=>"000110000",
  10830=>"110111001",
  10831=>"111001111",
  10832=>"011001101",
  10833=>"011011000",
  10834=>"101100010",
  10835=>"000110100",
  10836=>"111110111",
  10837=>"010010001",
  10838=>"000101101",
  10839=>"101010100",
  10840=>"101001110",
  10841=>"010100001",
  10842=>"001111101",
  10843=>"010000100",
  10844=>"110001111",
  10845=>"100000100",
  10846=>"101001010",
  10847=>"010000000",
  10848=>"011001110",
  10849=>"101010100",
  10850=>"001101111",
  10851=>"000111000",
  10852=>"000110010",
  10853=>"110100111",
  10854=>"111011011",
  10855=>"101001001",
  10856=>"100000111",
  10857=>"010100100",
  10858=>"111000110",
  10859=>"101010000",
  10860=>"110010110",
  10861=>"101110111",
  10862=>"100000010",
  10863=>"010100111",
  10864=>"010111010",
  10865=>"101000010",
  10866=>"111001110",
  10867=>"010010101",
  10868=>"010000010",
  10869=>"010011011",
  10870=>"101000000",
  10871=>"101001111",
  10872=>"010010100",
  10873=>"001000100",
  10874=>"011011000",
  10875=>"111111000",
  10876=>"010010010",
  10877=>"011111100",
  10878=>"000010101",
  10879=>"110101111",
  10880=>"011100100",
  10881=>"010101000",
  10882=>"101111100",
  10883=>"001001100",
  10884=>"001000110",
  10885=>"011100001",
  10886=>"010000011",
  10887=>"110010100",
  10888=>"001101100",
  10889=>"110010101",
  10890=>"100101001",
  10891=>"101111010",
  10892=>"101111000",
  10893=>"011001000",
  10894=>"001101010",
  10895=>"001110000",
  10896=>"010111100",
  10897=>"101110000",
  10898=>"010100100",
  10899=>"011010000",
  10900=>"000110110",
  10901=>"100010010",
  10902=>"101100011",
  10903=>"111101111",
  10904=>"001010111",
  10905=>"111000101",
  10906=>"100001001",
  10907=>"011001111",
  10908=>"111100010",
  10909=>"111000011",
  10910=>"000000101",
  10911=>"110011010",
  10912=>"001110000",
  10913=>"110110010",
  10914=>"110010000",
  10915=>"010011010",
  10916=>"011101111",
  10917=>"101111000",
  10918=>"100011000",
  10919=>"101000111",
  10920=>"101011111",
  10921=>"011010110",
  10922=>"000100101",
  10923=>"000111110",
  10924=>"101011001",
  10925=>"100101100",
  10926=>"000101101",
  10927=>"010111110",
  10928=>"100010111",
  10929=>"000010100",
  10930=>"001011010",
  10931=>"100010000",
  10932=>"111100111",
  10933=>"011111111",
  10934=>"000101001",
  10935=>"011010001",
  10936=>"001110101",
  10937=>"111101010",
  10938=>"110100011",
  10939=>"100100010",
  10940=>"110010000",
  10941=>"110000010",
  10942=>"000100010",
  10943=>"000111101",
  10944=>"101011011",
  10945=>"101010000",
  10946=>"000000001",
  10947=>"101101101",
  10948=>"011101101",
  10949=>"110110000",
  10950=>"000000111",
  10951=>"101101000",
  10952=>"010110100",
  10953=>"000110001",
  10954=>"010011000",
  10955=>"100110001",
  10956=>"100010111",
  10957=>"011111011",
  10958=>"111010000",
  10959=>"111001100",
  10960=>"101100100",
  10961=>"000100101",
  10962=>"010001110",
  10963=>"101111101",
  10964=>"110000001",
  10965=>"000100110",
  10966=>"111000101",
  10967=>"000010010",
  10968=>"111101010",
  10969=>"010111110",
  10970=>"100010100",
  10971=>"010100100",
  10972=>"100101111",
  10973=>"100111111",
  10974=>"111110101",
  10975=>"101110000",
  10976=>"100111101",
  10977=>"100011100",
  10978=>"111111011",
  10979=>"011111101",
  10980=>"100011010",
  10981=>"010010011",
  10982=>"001111100",
  10983=>"100011110",
  10984=>"100101010",
  10985=>"101101000",
  10986=>"110100011",
  10987=>"101001000",
  10988=>"001111000",
  10989=>"111000011",
  10990=>"101111010",
  10991=>"100011101",
  10992=>"110111011",
  10993=>"101111001",
  10994=>"001001001",
  10995=>"100011011",
  10996=>"000110101",
  10997=>"101110010",
  10998=>"010111100",
  10999=>"111011011",
  11000=>"100001010",
  11001=>"011101001",
  11002=>"111010011",
  11003=>"100111101",
  11004=>"110111110",
  11005=>"010000100",
  11006=>"011111001",
  11007=>"101010001",
  11008=>"111000100",
  11009=>"101100011",
  11010=>"000010101",
  11011=>"100100011",
  11012=>"011111111",
  11013=>"001011111",
  11014=>"111110011",
  11015=>"011101011",
  11016=>"011100101",
  11017=>"101001100",
  11018=>"101010000",
  11019=>"011010111",
  11020=>"100100101",
  11021=>"111110101",
  11022=>"110011111",
  11023=>"110001011",
  11024=>"111011111",
  11025=>"010111110",
  11026=>"000111000",
  11027=>"110101101",
  11028=>"100101110",
  11029=>"010100001",
  11030=>"100000001",
  11031=>"101011000",
  11032=>"000101000",
  11033=>"100101100",
  11034=>"001100000",
  11035=>"100100101",
  11036=>"110100000",
  11037=>"011010110",
  11038=>"000001000",
  11039=>"111010101",
  11040=>"111011001",
  11041=>"011001111",
  11042=>"111001110",
  11043=>"001000110",
  11044=>"110000111",
  11045=>"000100100",
  11046=>"100101100",
  11047=>"001011101",
  11048=>"010111011",
  11049=>"011101110",
  11050=>"000001010",
  11051=>"111111011",
  11052=>"110110100",
  11053=>"110101010",
  11054=>"001001111",
  11055=>"000111001",
  11056=>"011001001",
  11057=>"101110110",
  11058=>"000110000",
  11059=>"010110111",
  11060=>"001011010",
  11061=>"000011110",
  11062=>"011000100",
  11063=>"111100000",
  11064=>"101000111",
  11065=>"111000101",
  11066=>"001011001",
  11067=>"111110111",
  11068=>"010000001",
  11069=>"100010000",
  11070=>"111110101",
  11071=>"111001011",
  11072=>"100111001",
  11073=>"101001110",
  11074=>"001010011",
  11075=>"101001110",
  11076=>"001011111",
  11077=>"111111101",
  11078=>"101101100",
  11079=>"010100001",
  11080=>"001010111",
  11081=>"001001101",
  11082=>"101111111",
  11083=>"000101001",
  11084=>"101110011",
  11085=>"011110100",
  11086=>"000000000",
  11087=>"011101000",
  11088=>"110000001",
  11089=>"010111000",
  11090=>"011010010",
  11091=>"011000011",
  11092=>"001000100",
  11093=>"100000111",
  11094=>"001000011",
  11095=>"110000011",
  11096=>"001100011",
  11097=>"001001110",
  11098=>"010101011",
  11099=>"011001110",
  11100=>"001100001",
  11101=>"100010011",
  11102=>"110100000",
  11103=>"010100011",
  11104=>"111000101",
  11105=>"001100000",
  11106=>"000010110",
  11107=>"101111001",
  11108=>"101101111",
  11109=>"001001110",
  11110=>"100100110",
  11111=>"001111101",
  11112=>"011111110",
  11113=>"001100101",
  11114=>"111000100",
  11115=>"101100101",
  11116=>"101101110",
  11117=>"100100010",
  11118=>"000000111",
  11119=>"001111000",
  11120=>"001000110",
  11121=>"100110111",
  11122=>"010110101",
  11123=>"111100010",
  11124=>"100000010",
  11125=>"111001011",
  11126=>"110000011",
  11127=>"110001001",
  11128=>"011001011",
  11129=>"111010101",
  11130=>"010100101",
  11131=>"111011011",
  11132=>"011010100",
  11133=>"010111111",
  11134=>"100011001",
  11135=>"100110001",
  11136=>"100010000",
  11137=>"011111111",
  11138=>"101000010",
  11139=>"100101001",
  11140=>"010011111",
  11141=>"110001011",
  11142=>"100101111",
  11143=>"010001001",
  11144=>"000110000",
  11145=>"100000110",
  11146=>"110011101",
  11147=>"000000011",
  11148=>"000110100",
  11149=>"010001011",
  11150=>"001010111",
  11151=>"101111110",
  11152=>"000000110",
  11153=>"100101010",
  11154=>"100010100",
  11155=>"001100011",
  11156=>"011111000",
  11157=>"111110011",
  11158=>"110101101",
  11159=>"101110010",
  11160=>"110000101",
  11161=>"101111011",
  11162=>"101010101",
  11163=>"000001100",
  11164=>"100101111",
  11165=>"000110111",
  11166=>"110010101",
  11167=>"010111011",
  11168=>"100001100",
  11169=>"110101111",
  11170=>"000000000",
  11171=>"001101110",
  11172=>"000001010",
  11173=>"011111100",
  11174=>"100111111",
  11175=>"001101110",
  11176=>"001000110",
  11177=>"001001100",
  11178=>"000110000",
  11179=>"011001000",
  11180=>"100011101",
  11181=>"111110110",
  11182=>"000000010",
  11183=>"011111111",
  11184=>"000010010",
  11185=>"101010111",
  11186=>"100100000",
  11187=>"000101001",
  11188=>"110101100",
  11189=>"111001101",
  11190=>"111001101",
  11191=>"011100100",
  11192=>"011010001",
  11193=>"000011100",
  11194=>"110111010",
  11195=>"111110000",
  11196=>"111111101",
  11197=>"111000000",
  11198=>"010000110",
  11199=>"001001010",
  11200=>"111011011",
  11201=>"100011001",
  11202=>"111101110",
  11203=>"001101010",
  11204=>"010000010",
  11205=>"000010110",
  11206=>"100100000",
  11207=>"010100101",
  11208=>"010110100",
  11209=>"111011100",
  11210=>"110000110",
  11211=>"111000110",
  11212=>"010110111",
  11213=>"100100011",
  11214=>"000101110",
  11215=>"001010010",
  11216=>"001010011",
  11217=>"110001001",
  11218=>"010011000",
  11219=>"100110100",
  11220=>"000100001",
  11221=>"111101101",
  11222=>"111000001",
  11223=>"010111110",
  11224=>"110000000",
  11225=>"101010001",
  11226=>"011011001",
  11227=>"010000111",
  11228=>"011011000",
  11229=>"001110101",
  11230=>"011100001",
  11231=>"011111000",
  11232=>"001001101",
  11233=>"110000000",
  11234=>"111010110",
  11235=>"001001010",
  11236=>"111111000",
  11237=>"000001101",
  11238=>"001101000",
  11239=>"000101010",
  11240=>"011001111",
  11241=>"000010101",
  11242=>"111010010",
  11243=>"000111110",
  11244=>"100111000",
  11245=>"101000000",
  11246=>"011011100",
  11247=>"100101000",
  11248=>"101011101",
  11249=>"010001010",
  11250=>"001110100",
  11251=>"110101110",
  11252=>"011010000",
  11253=>"101001100",
  11254=>"110000001",
  11255=>"010001100",
  11256=>"001010111",
  11257=>"111010001",
  11258=>"111111101",
  11259=>"101000101",
  11260=>"101001111",
  11261=>"111001010",
  11262=>"111101111",
  11263=>"101101100",
  11264=>"001010110",
  11265=>"101110011",
  11266=>"000100010",
  11267=>"001010011",
  11268=>"011001101",
  11269=>"110110100",
  11270=>"010101101",
  11271=>"111000001",
  11272=>"111111100",
  11273=>"001011111",
  11274=>"000000110",
  11275=>"010110101",
  11276=>"000110010",
  11277=>"011100000",
  11278=>"011101000",
  11279=>"011100011",
  11280=>"100101101",
  11281=>"100010010",
  11282=>"010110110",
  11283=>"110001101",
  11284=>"001000100",
  11285=>"110111011",
  11286=>"000110011",
  11287=>"101101110",
  11288=>"100010011",
  11289=>"010100100",
  11290=>"001100110",
  11291=>"101100000",
  11292=>"011011000",
  11293=>"100100100",
  11294=>"010000000",
  11295=>"101000001",
  11296=>"010000001",
  11297=>"111010001",
  11298=>"000100001",
  11299=>"010001100",
  11300=>"111010000",
  11301=>"110110110",
  11302=>"011101101",
  11303=>"110000101",
  11304=>"011000110",
  11305=>"110011101",
  11306=>"000001110",
  11307=>"001010001",
  11308=>"101000001",
  11309=>"010100011",
  11310=>"110101010",
  11311=>"111111011",
  11312=>"000001000",
  11313=>"111101101",
  11314=>"011110110",
  11315=>"010000001",
  11316=>"010001011",
  11317=>"100110010",
  11318=>"101100000",
  11319=>"001011110",
  11320=>"101100000",
  11321=>"000000001",
  11322=>"000010110",
  11323=>"000100110",
  11324=>"011000000",
  11325=>"111101100",
  11326=>"000111101",
  11327=>"111110001",
  11328=>"010100010",
  11329=>"000001100",
  11330=>"011110000",
  11331=>"000111000",
  11332=>"111010101",
  11333=>"111101001",
  11334=>"101111010",
  11335=>"111000000",
  11336=>"100111001",
  11337=>"011100100",
  11338=>"000000011",
  11339=>"100111100",
  11340=>"011011010",
  11341=>"110111001",
  11342=>"111001110",
  11343=>"111001000",
  11344=>"111000100",
  11345=>"000010100",
  11346=>"100001001",
  11347=>"101100000",
  11348=>"010001101",
  11349=>"100010010",
  11350=>"011010101",
  11351=>"100010000",
  11352=>"111111101",
  11353=>"110010100",
  11354=>"110011101",
  11355=>"001101101",
  11356=>"101010010",
  11357=>"100110010",
  11358=>"001111110",
  11359=>"100010001",
  11360=>"110011010",
  11361=>"011000101",
  11362=>"001001111",
  11363=>"100100101",
  11364=>"110110000",
  11365=>"001011001",
  11366=>"110111001",
  11367=>"001100010",
  11368=>"001101010",
  11369=>"110110110",
  11370=>"110011010",
  11371=>"111001100",
  11372=>"100100001",
  11373=>"101110010",
  11374=>"101001101",
  11375=>"101000001",
  11376=>"011001011",
  11377=>"011111111",
  11378=>"010010111",
  11379=>"010001010",
  11380=>"010101011",
  11381=>"001000001",
  11382=>"100010100",
  11383=>"101111101",
  11384=>"100101001",
  11385=>"000011100",
  11386=>"110101111",
  11387=>"010110100",
  11388=>"001010100",
  11389=>"011110100",
  11390=>"000000001",
  11391=>"100010010",
  11392=>"000100011",
  11393=>"010100111",
  11394=>"100110100",
  11395=>"001010101",
  11396=>"100000000",
  11397=>"101011001",
  11398=>"101101110",
  11399=>"000110000",
  11400=>"011101110",
  11401=>"001010110",
  11402=>"100000100",
  11403=>"011010110",
  11404=>"001010101",
  11405=>"011101111",
  11406=>"110010010",
  11407=>"110000000",
  11408=>"000100010",
  11409=>"010000001",
  11410=>"011111110",
  11411=>"010011110",
  11412=>"000101101",
  11413=>"100110111",
  11414=>"010000110",
  11415=>"010110101",
  11416=>"010000000",
  11417=>"010011110",
  11418=>"110000011",
  11419=>"100011001",
  11420=>"100111110",
  11421=>"000000100",
  11422=>"111100100",
  11423=>"010001000",
  11424=>"110001100",
  11425=>"101100110",
  11426=>"011001000",
  11427=>"111010100",
  11428=>"011011010",
  11429=>"011110010",
  11430=>"101110000",
  11431=>"010000011",
  11432=>"011010101",
  11433=>"011101001",
  11434=>"001010010",
  11435=>"010001101",
  11436=>"000111111",
  11437=>"101000100",
  11438=>"001001001",
  11439=>"100100101",
  11440=>"010100100",
  11441=>"001011011",
  11442=>"111111110",
  11443=>"000100001",
  11444=>"000101100",
  11445=>"110011101",
  11446=>"100000111",
  11447=>"001011010",
  11448=>"000000101",
  11449=>"000100011",
  11450=>"000101100",
  11451=>"100100011",
  11452=>"100110001",
  11453=>"011010011",
  11454=>"011101111",
  11455=>"101101010",
  11456=>"110001100",
  11457=>"100101001",
  11458=>"111100000",
  11459=>"010110100",
  11460=>"100000010",
  11461=>"110110111",
  11462=>"010000110",
  11463=>"111100111",
  11464=>"110100001",
  11465=>"100110100",
  11466=>"000100100",
  11467=>"111100101",
  11468=>"111101111",
  11469=>"110010110",
  11470=>"001101011",
  11471=>"110000101",
  11472=>"101010110",
  11473=>"001010001",
  11474=>"101100001",
  11475=>"000000011",
  11476=>"001000011",
  11477=>"111010001",
  11478=>"110000001",
  11479=>"110011000",
  11480=>"010010101",
  11481=>"001011001",
  11482=>"010001011",
  11483=>"010000000",
  11484=>"101110110",
  11485=>"010101100",
  11486=>"110010101",
  11487=>"111010001",
  11488=>"010100010",
  11489=>"001001110",
  11490=>"100010001",
  11491=>"011101000",
  11492=>"101000101",
  11493=>"000110100",
  11494=>"111110111",
  11495=>"101110110",
  11496=>"011101011",
  11497=>"000101001",
  11498=>"111101101",
  11499=>"101000000",
  11500=>"000111000",
  11501=>"001001111",
  11502=>"000001101",
  11503=>"000000100",
  11504=>"011011111",
  11505=>"001010100",
  11506=>"101001110",
  11507=>"100111100",
  11508=>"101000010",
  11509=>"011111001",
  11510=>"101000001",
  11511=>"010001010",
  11512=>"110101010",
  11513=>"011010110",
  11514=>"101101001",
  11515=>"010100110",
  11516=>"001000000",
  11517=>"000000010",
  11518=>"101000100",
  11519=>"010001110",
  11520=>"011111101",
  11521=>"100101110",
  11522=>"110010110",
  11523=>"011001110",
  11524=>"101000101",
  11525=>"010000111",
  11526=>"100110101",
  11527=>"100110110",
  11528=>"001111111",
  11529=>"101011011",
  11530=>"011101000",
  11531=>"110011100",
  11532=>"001101011",
  11533=>"010100010",
  11534=>"010100101",
  11535=>"000101011",
  11536=>"000110001",
  11537=>"010101111",
  11538=>"110100110",
  11539=>"100001000",
  11540=>"000010100",
  11541=>"000001111",
  11542=>"101001000",
  11543=>"100001111",
  11544=>"110000010",
  11545=>"101110011",
  11546=>"001000101",
  11547=>"111011010",
  11548=>"011101111",
  11549=>"001001101",
  11550=>"010001000",
  11551=>"111000000",
  11552=>"011101101",
  11553=>"001001001",
  11554=>"111010110",
  11555=>"010110010",
  11556=>"000110001",
  11557=>"100101010",
  11558=>"000101011",
  11559=>"111101011",
  11560=>"001000110",
  11561=>"001101100",
  11562=>"100011000",
  11563=>"001111100",
  11564=>"111100101",
  11565=>"000100110",
  11566=>"100100110",
  11567=>"000010111",
  11568=>"100010110",
  11569=>"000100011",
  11570=>"001011111",
  11571=>"100011001",
  11572=>"100011101",
  11573=>"100110010",
  11574=>"101001101",
  11575=>"110011100",
  11576=>"000000011",
  11577=>"011010000",
  11578=>"100111101",
  11579=>"011001110",
  11580=>"001011001",
  11581=>"100000011",
  11582=>"000111110",
  11583=>"011010011",
  11584=>"011100110",
  11585=>"110110001",
  11586=>"100000111",
  11587=>"111101010",
  11588=>"001110100",
  11589=>"011011110",
  11590=>"001111101",
  11591=>"001110101",
  11592=>"100011110",
  11593=>"011110010",
  11594=>"011011110",
  11595=>"101000101",
  11596=>"001101100",
  11597=>"110011111",
  11598=>"100101110",
  11599=>"111101101",
  11600=>"011110000",
  11601=>"111110000",
  11602=>"000011010",
  11603=>"100100101",
  11604=>"011001000",
  11605=>"001111011",
  11606=>"000000001",
  11607=>"000000011",
  11608=>"101010110",
  11609=>"001110011",
  11610=>"001111111",
  11611=>"100100000",
  11612=>"011000000",
  11613=>"001010001",
  11614=>"001001111",
  11615=>"000000110",
  11616=>"101101101",
  11617=>"110110101",
  11618=>"000001100",
  11619=>"000000111",
  11620=>"111111100",
  11621=>"110000111",
  11622=>"011100100",
  11623=>"111110101",
  11624=>"011011100",
  11625=>"000101111",
  11626=>"000010011",
  11627=>"000111100",
  11628=>"111000000",
  11629=>"010010000",
  11630=>"001000000",
  11631=>"000101000",
  11632=>"010001001",
  11633=>"101110111",
  11634=>"101100111",
  11635=>"100111100",
  11636=>"100110110",
  11637=>"001011010",
  11638=>"000000000",
  11639=>"001011001",
  11640=>"010100010",
  11641=>"011101100",
  11642=>"010110010",
  11643=>"101110111",
  11644=>"000010111",
  11645=>"111111000",
  11646=>"010110100",
  11647=>"011011110",
  11648=>"110001001",
  11649=>"000111000",
  11650=>"100110111",
  11651=>"101001010",
  11652=>"010111011",
  11653=>"110101000",
  11654=>"010111111",
  11655=>"011000101",
  11656=>"100101010",
  11657=>"110111111",
  11658=>"010010100",
  11659=>"001100000",
  11660=>"001011001",
  11661=>"111100000",
  11662=>"001100100",
  11663=>"110110100",
  11664=>"111010110",
  11665=>"010000001",
  11666=>"010000110",
  11667=>"110101101",
  11668=>"100000111",
  11669=>"010010001",
  11670=>"100000000",
  11671=>"011111110",
  11672=>"101111010",
  11673=>"000000101",
  11674=>"010010001",
  11675=>"000000010",
  11676=>"011000000",
  11677=>"000110001",
  11678=>"001100110",
  11679=>"101100111",
  11680=>"111110000",
  11681=>"010010010",
  11682=>"011011101",
  11683=>"100000010",
  11684=>"101000100",
  11685=>"001000010",
  11686=>"001100000",
  11687=>"110001111",
  11688=>"010100011",
  11689=>"110110011",
  11690=>"100000000",
  11691=>"100111000",
  11692=>"011100000",
  11693=>"110000111",
  11694=>"000100100",
  11695=>"110010110",
  11696=>"000110000",
  11697=>"001000010",
  11698=>"111010110",
  11699=>"111010111",
  11700=>"010001011",
  11701=>"100001101",
  11702=>"000011011",
  11703=>"000010100",
  11704=>"000110100",
  11705=>"111001101",
  11706=>"100111011",
  11707=>"111010000",
  11708=>"111100000",
  11709=>"000101001",
  11710=>"001100101",
  11711=>"111001001",
  11712=>"011101100",
  11713=>"100001101",
  11714=>"100101001",
  11715=>"111100001",
  11716=>"101000001",
  11717=>"000001011",
  11718=>"100001011",
  11719=>"010000000",
  11720=>"111010110",
  11721=>"000110100",
  11722=>"101011110",
  11723=>"001000000",
  11724=>"000000010",
  11725=>"111111101",
  11726=>"000001011",
  11727=>"010110100",
  11728=>"100010111",
  11729=>"010110001",
  11730=>"101100000",
  11731=>"110110111",
  11732=>"001110011",
  11733=>"010011111",
  11734=>"001110000",
  11735=>"011000110",
  11736=>"101111010",
  11737=>"110001010",
  11738=>"111001001",
  11739=>"101001000",
  11740=>"100001111",
  11741=>"000100001",
  11742=>"110010001",
  11743=>"111111000",
  11744=>"100100001",
  11745=>"111010000",
  11746=>"101010111",
  11747=>"110110101",
  11748=>"101000001",
  11749=>"001001001",
  11750=>"001010001",
  11751=>"011000110",
  11752=>"001001001",
  11753=>"000111000",
  11754=>"110000001",
  11755=>"101001010",
  11756=>"110101010",
  11757=>"100000110",
  11758=>"111111101",
  11759=>"100000110",
  11760=>"000101001",
  11761=>"000000111",
  11762=>"111000010",
  11763=>"000110100",
  11764=>"001001010",
  11765=>"010101100",
  11766=>"111110111",
  11767=>"001110101",
  11768=>"001010010",
  11769=>"011100000",
  11770=>"101100110",
  11771=>"100110011",
  11772=>"000111110",
  11773=>"110000100",
  11774=>"111111000",
  11775=>"010011110",
  11776=>"101101001",
  11777=>"001101001",
  11778=>"101000011",
  11779=>"110011011",
  11780=>"010000000",
  11781=>"100001000",
  11782=>"110001111",
  11783=>"010000000",
  11784=>"000111001",
  11785=>"110111100",
  11786=>"110001111",
  11787=>"111001011",
  11788=>"000011011",
  11789=>"001001110",
  11790=>"000000000",
  11791=>"010011010",
  11792=>"000011011",
  11793=>"110000111",
  11794=>"001000100",
  11795=>"111100001",
  11796=>"101000101",
  11797=>"011101001",
  11798=>"100011010",
  11799=>"100110111",
  11800=>"100100010",
  11801=>"010000010",
  11802=>"000010000",
  11803=>"110010101",
  11804=>"010110110",
  11805=>"000010001",
  11806=>"110100011",
  11807=>"000101101",
  11808=>"111010001",
  11809=>"010001110",
  11810=>"111000101",
  11811=>"000000101",
  11812=>"011111101",
  11813=>"111110101",
  11814=>"111001111",
  11815=>"000111101",
  11816=>"001001001",
  11817=>"011111100",
  11818=>"010011010",
  11819=>"111000000",
  11820=>"010110111",
  11821=>"101011011",
  11822=>"010000010",
  11823=>"110000110",
  11824=>"110101100",
  11825=>"011011100",
  11826=>"101001101",
  11827=>"011010111",
  11828=>"001011010",
  11829=>"000000010",
  11830=>"100100010",
  11831=>"001101111",
  11832=>"100101100",
  11833=>"101101011",
  11834=>"110101101",
  11835=>"100011111",
  11836=>"011100110",
  11837=>"000110010",
  11838=>"101101000",
  11839=>"101011010",
  11840=>"101100101",
  11841=>"011001000",
  11842=>"101011001",
  11843=>"001010010",
  11844=>"011010001",
  11845=>"100100010",
  11846=>"000000010",
  11847=>"010101001",
  11848=>"111111100",
  11849=>"101110001",
  11850=>"111011001",
  11851=>"100010111",
  11852=>"101110011",
  11853=>"000010011",
  11854=>"111110000",
  11855=>"111111011",
  11856=>"011111101",
  11857=>"000100110",
  11858=>"000100011",
  11859=>"000010000",
  11860=>"010011111",
  11861=>"111000010",
  11862=>"000011110",
  11863=>"001011010",
  11864=>"100000001",
  11865=>"100111010",
  11866=>"110011101",
  11867=>"000101011",
  11868=>"101110111",
  11869=>"011100100",
  11870=>"001011110",
  11871=>"011010111",
  11872=>"011000011",
  11873=>"000001000",
  11874=>"101101110",
  11875=>"100101010",
  11876=>"111100011",
  11877=>"100010011",
  11878=>"111100001",
  11879=>"000000101",
  11880=>"100001001",
  11881=>"100001000",
  11882=>"000001010",
  11883=>"100100011",
  11884=>"100100101",
  11885=>"100111000",
  11886=>"111100011",
  11887=>"110011001",
  11888=>"100101011",
  11889=>"111111111",
  11890=>"011101011",
  11891=>"011010000",
  11892=>"010000101",
  11893=>"010010110",
  11894=>"010101101",
  11895=>"000011011",
  11896=>"110000101",
  11897=>"111001001",
  11898=>"001100001",
  11899=>"111100111",
  11900=>"101100111",
  11901=>"001110010",
  11902=>"111001000",
  11903=>"101000111",
  11904=>"000001100",
  11905=>"011000011",
  11906=>"000010000",
  11907=>"100001111",
  11908=>"001100111",
  11909=>"100000100",
  11910=>"010011111",
  11911=>"111101011",
  11912=>"111110001",
  11913=>"010010111",
  11914=>"001001111",
  11915=>"010111111",
  11916=>"011001010",
  11917=>"110010100",
  11918=>"011000110",
  11919=>"111011000",
  11920=>"111000110",
  11921=>"111010001",
  11922=>"110110110",
  11923=>"110111100",
  11924=>"001100000",
  11925=>"100010110",
  11926=>"101111011",
  11927=>"000001001",
  11928=>"110001110",
  11929=>"001000010",
  11930=>"101000111",
  11931=>"111100010",
  11932=>"001110110",
  11933=>"010010001",
  11934=>"000000100",
  11935=>"100010010",
  11936=>"110111001",
  11937=>"100010110",
  11938=>"100001110",
  11939=>"000011111",
  11940=>"001010011",
  11941=>"000111000",
  11942=>"100010100",
  11943=>"000000101",
  11944=>"011100000",
  11945=>"100001011",
  11946=>"101111011",
  11947=>"010111010",
  11948=>"010110111",
  11949=>"101011010",
  11950=>"010110010",
  11951=>"100110110",
  11952=>"110001111",
  11953=>"100000000",
  11954=>"100010010",
  11955=>"111100011",
  11956=>"001111000",
  11957=>"100100110",
  11958=>"010011000",
  11959=>"111110011",
  11960=>"000011111",
  11961=>"100100011",
  11962=>"110001111",
  11963=>"111101101",
  11964=>"010101000",
  11965=>"001000101",
  11966=>"001010100",
  11967=>"101010011",
  11968=>"010001100",
  11969=>"011001101",
  11970=>"100011010",
  11971=>"001001111",
  11972=>"110101110",
  11973=>"001011111",
  11974=>"111010000",
  11975=>"110010010",
  11976=>"111111000",
  11977=>"001001110",
  11978=>"100000110",
  11979=>"101011101",
  11980=>"100101001",
  11981=>"100011110",
  11982=>"011000111",
  11983=>"110100111",
  11984=>"110010101",
  11985=>"011010010",
  11986=>"011100000",
  11987=>"000010101",
  11988=>"110010001",
  11989=>"101101001",
  11990=>"001111101",
  11991=>"101110000",
  11992=>"000000011",
  11993=>"111110110",
  11994=>"010011111",
  11995=>"011100101",
  11996=>"001000110",
  11997=>"001011000",
  11998=>"000100110",
  11999=>"011100111",
  12000=>"101100110",
  12001=>"100000101",
  12002=>"111111011",
  12003=>"010111000",
  12004=>"000101101",
  12005=>"011111101",
  12006=>"010010111",
  12007=>"000111101",
  12008=>"001001000",
  12009=>"101001111",
  12010=>"000110000",
  12011=>"101010111",
  12012=>"000011101",
  12013=>"100010101",
  12014=>"010011110",
  12015=>"100100100",
  12016=>"101110100",
  12017=>"011010000",
  12018=>"101000110",
  12019=>"100000010",
  12020=>"011111110",
  12021=>"001001101",
  12022=>"111111000",
  12023=>"100000111",
  12024=>"011011001",
  12025=>"010111111",
  12026=>"011111011",
  12027=>"011110001",
  12028=>"011011010",
  12029=>"001110000",
  12030=>"001000000",
  12031=>"000001001",
  12032=>"010001010",
  12033=>"001010011",
  12034=>"110000011",
  12035=>"010110000",
  12036=>"100011101",
  12037=>"001100100",
  12038=>"011101111",
  12039=>"101000000",
  12040=>"100011000",
  12041=>"001100110",
  12042=>"111001011",
  12043=>"000001110",
  12044=>"110101001",
  12045=>"101011101",
  12046=>"000000110",
  12047=>"110100001",
  12048=>"000000111",
  12049=>"000000111",
  12050=>"111010100",
  12051=>"111111110",
  12052=>"111111100",
  12053=>"000000010",
  12054=>"101000110",
  12055=>"111101000",
  12056=>"000001010",
  12057=>"001001110",
  12058=>"001000011",
  12059=>"101001010",
  12060=>"001011111",
  12061=>"110111101",
  12062=>"011111000",
  12063=>"101100111",
  12064=>"111010110",
  12065=>"101100101",
  12066=>"010000000",
  12067=>"101000010",
  12068=>"000101000",
  12069=>"110001100",
  12070=>"011000010",
  12071=>"101010101",
  12072=>"111100011",
  12073=>"011001010",
  12074=>"000110011",
  12075=>"011101111",
  12076=>"001101110",
  12077=>"010010001",
  12078=>"000111111",
  12079=>"011011011",
  12080=>"010100000",
  12081=>"111010100",
  12082=>"100111111",
  12083=>"010000100",
  12084=>"001000001",
  12085=>"100011010",
  12086=>"000111000",
  12087=>"011111001",
  12088=>"111010100",
  12089=>"101101000",
  12090=>"000100000",
  12091=>"000010010",
  12092=>"110101001",
  12093=>"000000110",
  12094=>"111001000",
  12095=>"100000010",
  12096=>"001000010",
  12097=>"110111111",
  12098=>"001101000",
  12099=>"011100111",
  12100=>"110000000",
  12101=>"110110010",
  12102=>"010001001",
  12103=>"010000110",
  12104=>"001000000",
  12105=>"111001100",
  12106=>"010000111",
  12107=>"000110011",
  12108=>"000111110",
  12109=>"110100001",
  12110=>"000100001",
  12111=>"001010011",
  12112=>"111100101",
  12113=>"001110111",
  12114=>"110101101",
  12115=>"000101000",
  12116=>"100001001",
  12117=>"010110011",
  12118=>"001100000",
  12119=>"010010111",
  12120=>"000001101",
  12121=>"111111010",
  12122=>"111000011",
  12123=>"101100111",
  12124=>"001000110",
  12125=>"111001111",
  12126=>"110110101",
  12127=>"010000100",
  12128=>"001010011",
  12129=>"110100000",
  12130=>"000110001",
  12131=>"010001000",
  12132=>"110110010",
  12133=>"110000100",
  12134=>"000111010",
  12135=>"111000110",
  12136=>"001010000",
  12137=>"011010011",
  12138=>"010010001",
  12139=>"000111011",
  12140=>"111011011",
  12141=>"000010111",
  12142=>"011101010",
  12143=>"101010010",
  12144=>"110000111",
  12145=>"011011110",
  12146=>"010010000",
  12147=>"100100100",
  12148=>"000111110",
  12149=>"001011101",
  12150=>"101100010",
  12151=>"000000000",
  12152=>"001111100",
  12153=>"111010010",
  12154=>"001010101",
  12155=>"010010111",
  12156=>"001110011",
  12157=>"101111101",
  12158=>"111010010",
  12159=>"111000000",
  12160=>"010110111",
  12161=>"101000000",
  12162=>"000111001",
  12163=>"101111100",
  12164=>"111110100",
  12165=>"000001000",
  12166=>"011101101",
  12167=>"111001100",
  12168=>"101001110",
  12169=>"000111010",
  12170=>"110011011",
  12171=>"100000110",
  12172=>"001010100",
  12173=>"010000001",
  12174=>"000000011",
  12175=>"001011000",
  12176=>"101100110",
  12177=>"001110010",
  12178=>"010000000",
  12179=>"010001100",
  12180=>"001100111",
  12181=>"111001101",
  12182=>"011101101",
  12183=>"101110000",
  12184=>"100010010",
  12185=>"110001011",
  12186=>"110101111",
  12187=>"100110000",
  12188=>"000010000",
  12189=>"101101111",
  12190=>"010001000",
  12191=>"101111110",
  12192=>"110010010",
  12193=>"000010101",
  12194=>"010101010",
  12195=>"110111001",
  12196=>"000011011",
  12197=>"111111101",
  12198=>"000110110",
  12199=>"100101010",
  12200=>"010101110",
  12201=>"010101010",
  12202=>"111111000",
  12203=>"000110011",
  12204=>"101100000",
  12205=>"100100111",
  12206=>"100111010",
  12207=>"001000111",
  12208=>"100011111",
  12209=>"111111001",
  12210=>"101010011",
  12211=>"001001011",
  12212=>"111100001",
  12213=>"001100101",
  12214=>"111110011",
  12215=>"100010011",
  12216=>"011111111",
  12217=>"100111000",
  12218=>"010101110",
  12219=>"011101111",
  12220=>"110000010",
  12221=>"001100001",
  12222=>"110110000",
  12223=>"000110111",
  12224=>"001001110",
  12225=>"010111101",
  12226=>"110001000",
  12227=>"100000111",
  12228=>"100100101",
  12229=>"110010110",
  12230=>"101111101",
  12231=>"000110011",
  12232=>"101101001",
  12233=>"001111000",
  12234=>"011101011",
  12235=>"001000101",
  12236=>"100110011",
  12237=>"000000010",
  12238=>"100011011",
  12239=>"111010001",
  12240=>"100110101",
  12241=>"000011011",
  12242=>"101010011",
  12243=>"100011110",
  12244=>"010111010",
  12245=>"000000110",
  12246=>"110100100",
  12247=>"100111100",
  12248=>"110010000",
  12249=>"111111110",
  12250=>"001011001",
  12251=>"001000000",
  12252=>"110100101",
  12253=>"110111101",
  12254=>"100000101",
  12255=>"011000101",
  12256=>"101111111",
  12257=>"100000000",
  12258=>"111010001",
  12259=>"101110010",
  12260=>"100010000",
  12261=>"001001011",
  12262=>"000110100",
  12263=>"001001001",
  12264=>"100111101",
  12265=>"001101001",
  12266=>"000001011",
  12267=>"010011010",
  12268=>"100000001",
  12269=>"001010111",
  12270=>"000111010",
  12271=>"010100101",
  12272=>"000111110",
  12273=>"001000100",
  12274=>"001111100",
  12275=>"000111000",
  12276=>"101001111",
  12277=>"001001001",
  12278=>"101000101",
  12279=>"001011011",
  12280=>"010011010",
  12281=>"001101100",
  12282=>"110001011",
  12283=>"010011110",
  12284=>"100101111",
  12285=>"101110001",
  12286=>"110011011",
  12287=>"101001101",
  12288=>"011111111",
  12289=>"010111111",
  12290=>"100000000",
  12291=>"100110000",
  12292=>"010100111",
  12293=>"111001111",
  12294=>"111111000",
  12295=>"001100101",
  12296=>"001100111",
  12297=>"000000101",
  12298=>"000011001",
  12299=>"101100010",
  12300=>"101010100",
  12301=>"110110011",
  12302=>"111111011",
  12303=>"001100111",
  12304=>"000000101",
  12305=>"000000111",
  12306=>"111101101",
  12307=>"110111011",
  12308=>"010110101",
  12309=>"001011111",
  12310=>"000011000",
  12311=>"110111001",
  12312=>"111101101",
  12313=>"011010111",
  12314=>"001000011",
  12315=>"001111101",
  12316=>"111000000",
  12317=>"010100101",
  12318=>"010111110",
  12319=>"000110100",
  12320=>"001111111",
  12321=>"000101001",
  12322=>"111011001",
  12323=>"100101010",
  12324=>"011011110",
  12325=>"000001000",
  12326=>"011101101",
  12327=>"111100010",
  12328=>"010100101",
  12329=>"011010010",
  12330=>"110100110",
  12331=>"101011000",
  12332=>"100000000",
  12333=>"111011100",
  12334=>"010110100",
  12335=>"000001100",
  12336=>"000100100",
  12337=>"100101111",
  12338=>"101111111",
  12339=>"100110010",
  12340=>"011110100",
  12341=>"100000001",
  12342=>"010100000",
  12343=>"000000001",
  12344=>"010000001",
  12345=>"111011110",
  12346=>"011111010",
  12347=>"001010011",
  12348=>"000001011",
  12349=>"000111011",
  12350=>"000001010",
  12351=>"110100110",
  12352=>"111110110",
  12353=>"100100111",
  12354=>"001101110",
  12355=>"110101100",
  12356=>"000110101",
  12357=>"000100011",
  12358=>"101010010",
  12359=>"111001011",
  12360=>"111011101",
  12361=>"010000010",
  12362=>"010000110",
  12363=>"011100001",
  12364=>"100100111",
  12365=>"001111010",
  12366=>"001111000",
  12367=>"101101101",
  12368=>"111110111",
  12369=>"111101111",
  12370=>"100110101",
  12371=>"011010111",
  12372=>"100110110",
  12373=>"010010010",
  12374=>"000000101",
  12375=>"001101011",
  12376=>"111111001",
  12377=>"000010000",
  12378=>"101100000",
  12379=>"010010011",
  12380=>"010101111",
  12381=>"101101000",
  12382=>"000111011",
  12383=>"000010001",
  12384=>"110011101",
  12385=>"111111111",
  12386=>"110101111",
  12387=>"111011111",
  12388=>"110000101",
  12389=>"000101001",
  12390=>"010111100",
  12391=>"011000011",
  12392=>"001001000",
  12393=>"010000000",
  12394=>"010101110",
  12395=>"011100101",
  12396=>"100010010",
  12397=>"000001100",
  12398=>"111111101",
  12399=>"000111101",
  12400=>"100110111",
  12401=>"110001100",
  12402=>"011011011",
  12403=>"111000011",
  12404=>"111111111",
  12405=>"001111011",
  12406=>"000111100",
  12407=>"110111110",
  12408=>"001110111",
  12409=>"001101001",
  12410=>"111111010",
  12411=>"011110010",
  12412=>"101111010",
  12413=>"000000010",
  12414=>"000000010",
  12415=>"111110100",
  12416=>"110110000",
  12417=>"010100111",
  12418=>"001011011",
  12419=>"100110101",
  12420=>"010010110",
  12421=>"001100111",
  12422=>"100111111",
  12423=>"111111100",
  12424=>"101000000",
  12425=>"000010000",
  12426=>"001100110",
  12427=>"011111110",
  12428=>"101001001",
  12429=>"010010011",
  12430=>"001100010",
  12431=>"100000100",
  12432=>"101000110",
  12433=>"111001010",
  12434=>"111000000",
  12435=>"000110001",
  12436=>"101001110",
  12437=>"100101110",
  12438=>"000010100",
  12439=>"010001000",
  12440=>"100110110",
  12441=>"111110101",
  12442=>"101000100",
  12443=>"101111001",
  12444=>"000110100",
  12445=>"100000101",
  12446=>"100011010",
  12447=>"111100001",
  12448=>"010000101",
  12449=>"011011101",
  12450=>"011100101",
  12451=>"100010001",
  12452=>"111011000",
  12453=>"011010001",
  12454=>"111000101",
  12455=>"111101111",
  12456=>"001110111",
  12457=>"100011001",
  12458=>"010010101",
  12459=>"111000001",
  12460=>"010001000",
  12461=>"100000110",
  12462=>"010100111",
  12463=>"111001100",
  12464=>"000011000",
  12465=>"100000000",
  12466=>"110010011",
  12467=>"100001111",
  12468=>"100010111",
  12469=>"110101111",
  12470=>"000001101",
  12471=>"000011001",
  12472=>"010011000",
  12473=>"000010001",
  12474=>"100000000",
  12475=>"110000010",
  12476=>"001110011",
  12477=>"100001010",
  12478=>"111111110",
  12479=>"010000010",
  12480=>"101110110",
  12481=>"100011000",
  12482=>"110110101",
  12483=>"110100010",
  12484=>"000000110",
  12485=>"111011111",
  12486=>"001110001",
  12487=>"111101111",
  12488=>"110100011",
  12489=>"000011011",
  12490=>"110001010",
  12491=>"000001001",
  12492=>"110001000",
  12493=>"001011001",
  12494=>"011000101",
  12495=>"100111000",
  12496=>"111100110",
  12497=>"011010100",
  12498=>"010100100",
  12499=>"101111101",
  12500=>"110001000",
  12501=>"101000111",
  12502=>"001001001",
  12503=>"111111111",
  12504=>"000100101",
  12505=>"000111001",
  12506=>"101111000",
  12507=>"000111011",
  12508=>"100101011",
  12509=>"101101110",
  12510=>"101100001",
  12511=>"101011101",
  12512=>"111101110",
  12513=>"011101101",
  12514=>"101010101",
  12515=>"001000101",
  12516=>"111100010",
  12517=>"000011010",
  12518=>"001111110",
  12519=>"001101011",
  12520=>"001111110",
  12521=>"111100101",
  12522=>"010111110",
  12523=>"001000101",
  12524=>"111001001",
  12525=>"011001111",
  12526=>"010101110",
  12527=>"001000000",
  12528=>"011000000",
  12529=>"000010010",
  12530=>"001110000",
  12531=>"000001101",
  12532=>"000101001",
  12533=>"011101110",
  12534=>"111000010",
  12535=>"011010111",
  12536=>"001011000",
  12537=>"111101111",
  12538=>"110011011",
  12539=>"111011011",
  12540=>"000001010",
  12541=>"000100110",
  12542=>"110101011",
  12543=>"011111110",
  12544=>"101100010",
  12545=>"111001110",
  12546=>"100100001",
  12547=>"011010000",
  12548=>"110101111",
  12549=>"111101111",
  12550=>"010010001",
  12551=>"001000001",
  12552=>"010101011",
  12553=>"110111101",
  12554=>"101100010",
  12555=>"111100101",
  12556=>"111000011",
  12557=>"011100100",
  12558=>"010111100",
  12559=>"110101001",
  12560=>"011001100",
  12561=>"010000001",
  12562=>"111011100",
  12563=>"010011010",
  12564=>"110010100",
  12565=>"001111110",
  12566=>"101010010",
  12567=>"001011001",
  12568=>"010101100",
  12569=>"011010011",
  12570=>"111111110",
  12571=>"101000001",
  12572=>"001001001",
  12573=>"010001001",
  12574=>"101011011",
  12575=>"000000010",
  12576=>"001010011",
  12577=>"110010000",
  12578=>"000110101",
  12579=>"101101010",
  12580=>"110100011",
  12581=>"111111100",
  12582=>"001110010",
  12583=>"000011100",
  12584=>"111001010",
  12585=>"011111111",
  12586=>"001101010",
  12587=>"100100100",
  12588=>"010011000",
  12589=>"010000000",
  12590=>"100011111",
  12591=>"110110010",
  12592=>"111000001",
  12593=>"110110011",
  12594=>"100001111",
  12595=>"000000101",
  12596=>"010001000",
  12597=>"111100010",
  12598=>"110110000",
  12599=>"011001010",
  12600=>"010100010",
  12601=>"110110111",
  12602=>"111100111",
  12603=>"000001000",
  12604=>"000110111",
  12605=>"101111110",
  12606=>"000010001",
  12607=>"001010001",
  12608=>"000100000",
  12609=>"111000001",
  12610=>"111001110",
  12611=>"110101011",
  12612=>"010111100",
  12613=>"111101001",
  12614=>"111101101",
  12615=>"001011111",
  12616=>"101100111",
  12617=>"110000010",
  12618=>"010011101",
  12619=>"000010110",
  12620=>"000100111",
  12621=>"101101000",
  12622=>"110000000",
  12623=>"100010101",
  12624=>"000110110",
  12625=>"010010111",
  12626=>"110110111",
  12627=>"010111111",
  12628=>"010011100",
  12629=>"001110111",
  12630=>"000101000",
  12631=>"010011101",
  12632=>"100000110",
  12633=>"111010100",
  12634=>"111011000",
  12635=>"001111010",
  12636=>"111101110",
  12637=>"101111010",
  12638=>"111011011",
  12639=>"000011010",
  12640=>"000000000",
  12641=>"100001011",
  12642=>"011111110",
  12643=>"100111000",
  12644=>"100010001",
  12645=>"000001101",
  12646=>"101111111",
  12647=>"011011011",
  12648=>"100101100",
  12649=>"111111111",
  12650=>"000100110",
  12651=>"000100111",
  12652=>"000000111",
  12653=>"111010010",
  12654=>"111101100",
  12655=>"110000000",
  12656=>"101101010",
  12657=>"000110101",
  12658=>"101101111",
  12659=>"000111010",
  12660=>"111011101",
  12661=>"111000110",
  12662=>"001011101",
  12663=>"000010001",
  12664=>"101011010",
  12665=>"011010001",
  12666=>"111010100",
  12667=>"100100000",
  12668=>"000010000",
  12669=>"110000001",
  12670=>"100100110",
  12671=>"100110001",
  12672=>"000110001",
  12673=>"000001010",
  12674=>"110111100",
  12675=>"111111111",
  12676=>"010011001",
  12677=>"001000001",
  12678=>"111000100",
  12679=>"011000000",
  12680=>"100110001",
  12681=>"011101001",
  12682=>"110100000",
  12683=>"111111000",
  12684=>"100001000",
  12685=>"111101111",
  12686=>"101011110",
  12687=>"010000111",
  12688=>"101110010",
  12689=>"110010010",
  12690=>"011111100",
  12691=>"000100110",
  12692=>"011111111",
  12693=>"000000110",
  12694=>"111110010",
  12695=>"001111100",
  12696=>"001100011",
  12697=>"100001101",
  12698=>"100111100",
  12699=>"001101111",
  12700=>"100001101",
  12701=>"110010011",
  12702=>"000110010",
  12703=>"000110010",
  12704=>"010010000",
  12705=>"001010000",
  12706=>"111100110",
  12707=>"000101111",
  12708=>"011000011",
  12709=>"010011000",
  12710=>"110010111",
  12711=>"000001110",
  12712=>"011101010",
  12713=>"011000100",
  12714=>"110000001",
  12715=>"001001001",
  12716=>"000000001",
  12717=>"110110100",
  12718=>"011001011",
  12719=>"110100011",
  12720=>"011000000",
  12721=>"001000010",
  12722=>"001011011",
  12723=>"010000111",
  12724=>"110100011",
  12725=>"101011011",
  12726=>"111101011",
  12727=>"110000101",
  12728=>"000111110",
  12729=>"110111011",
  12730=>"010010000",
  12731=>"010001100",
  12732=>"111010000",
  12733=>"111000110",
  12734=>"111101001",
  12735=>"011000000",
  12736=>"111110000",
  12737=>"100111110",
  12738=>"010110000",
  12739=>"001111001",
  12740=>"110001101",
  12741=>"010011001",
  12742=>"001100111",
  12743=>"000011010",
  12744=>"100010000",
  12745=>"001110100",
  12746=>"100110000",
  12747=>"000011110",
  12748=>"101000101",
  12749=>"010111100",
  12750=>"000111100",
  12751=>"111111110",
  12752=>"110100110",
  12753=>"100010101",
  12754=>"000011101",
  12755=>"101001011",
  12756=>"010001101",
  12757=>"101110010",
  12758=>"000000101",
  12759=>"110011110",
  12760=>"100011000",
  12761=>"001110100",
  12762=>"011110100",
  12763=>"000110100",
  12764=>"000001001",
  12765=>"001111001",
  12766=>"101011011",
  12767=>"101010111",
  12768=>"110110011",
  12769=>"100100000",
  12770=>"111100101",
  12771=>"011011011",
  12772=>"111000100",
  12773=>"001000011",
  12774=>"001011010",
  12775=>"110111001",
  12776=>"101100101",
  12777=>"111000111",
  12778=>"111101110",
  12779=>"110101011",
  12780=>"000001001",
  12781=>"010000111",
  12782=>"111101101",
  12783=>"001100101",
  12784=>"101011010",
  12785=>"001110000",
  12786=>"000101100",
  12787=>"010111010",
  12788=>"101000100",
  12789=>"100110011",
  12790=>"101111011",
  12791=>"111110011",
  12792=>"111010001",
  12793=>"000101101",
  12794=>"101011100",
  12795=>"000011100",
  12796=>"010000001",
  12797=>"001000010",
  12798=>"101001001",
  12799=>"111010111",
  12800=>"101001110",
  12801=>"001000101",
  12802=>"110011011",
  12803=>"110101100",
  12804=>"100100001",
  12805=>"100011100",
  12806=>"101010100",
  12807=>"001011111",
  12808=>"100110100",
  12809=>"010000000",
  12810=>"110000000",
  12811=>"111110001",
  12812=>"000101100",
  12813=>"010010000",
  12814=>"100111111",
  12815=>"010000011",
  12816=>"000010110",
  12817=>"000111100",
  12818=>"101011101",
  12819=>"011100010",
  12820=>"001101100",
  12821=>"011010000",
  12822=>"110110000",
  12823=>"111101110",
  12824=>"111111100",
  12825=>"111100000",
  12826=>"011100001",
  12827=>"011100100",
  12828=>"011110000",
  12829=>"010001011",
  12830=>"101111010",
  12831=>"011100010",
  12832=>"011100011",
  12833=>"001011000",
  12834=>"100010110",
  12835=>"000010011",
  12836=>"110100010",
  12837=>"110011111",
  12838=>"010010000",
  12839=>"011010000",
  12840=>"100000001",
  12841=>"001100110",
  12842=>"000000001",
  12843=>"101010101",
  12844=>"110111011",
  12845=>"011001110",
  12846=>"001101111",
  12847=>"001001010",
  12848=>"110101001",
  12849=>"001001101",
  12850=>"000001001",
  12851=>"110011000",
  12852=>"011110101",
  12853=>"001110101",
  12854=>"000101011",
  12855=>"000011101",
  12856=>"110111110",
  12857=>"101110111",
  12858=>"010001001",
  12859=>"000101011",
  12860=>"100001111",
  12861=>"100110000",
  12862=>"100101001",
  12863=>"001100000",
  12864=>"111010111",
  12865=>"111110110",
  12866=>"010010111",
  12867=>"111111110",
  12868=>"001011110",
  12869=>"100101011",
  12870=>"100000101",
  12871=>"010101101",
  12872=>"011110011",
  12873=>"111110110",
  12874=>"001111110",
  12875=>"000010101",
  12876=>"111101011",
  12877=>"010111011",
  12878=>"010000000",
  12879=>"011010011",
  12880=>"110001001",
  12881=>"000100100",
  12882=>"111010000",
  12883=>"101011001",
  12884=>"001000000",
  12885=>"100011100",
  12886=>"000000000",
  12887=>"111000011",
  12888=>"001110101",
  12889=>"010001110",
  12890=>"111001000",
  12891=>"010011011",
  12892=>"000000000",
  12893=>"101100110",
  12894=>"011010110",
  12895=>"111100100",
  12896=>"111100000",
  12897=>"001111100",
  12898=>"000010110",
  12899=>"001011010",
  12900=>"000000001",
  12901=>"010010100",
  12902=>"101001101",
  12903=>"001100010",
  12904=>"000000000",
  12905=>"100110010",
  12906=>"011000101",
  12907=>"101001100",
  12908=>"100111001",
  12909=>"101100111",
  12910=>"001001110",
  12911=>"100100100",
  12912=>"000011110",
  12913=>"001011010",
  12914=>"001001011",
  12915=>"000010110",
  12916=>"011100010",
  12917=>"010000101",
  12918=>"101111111",
  12919=>"000010100",
  12920=>"100010110",
  12921=>"010110000",
  12922=>"001101001",
  12923=>"001010001",
  12924=>"001100110",
  12925=>"001001001",
  12926=>"001111111",
  12927=>"100110011",
  12928=>"111011100",
  12929=>"010111110",
  12930=>"100100010",
  12931=>"111110110",
  12932=>"011110110",
  12933=>"011101001",
  12934=>"100100111",
  12935=>"111110101",
  12936=>"110101101",
  12937=>"000110110",
  12938=>"100110010",
  12939=>"100100000",
  12940=>"011101001",
  12941=>"010011000",
  12942=>"101011111",
  12943=>"001001100",
  12944=>"000001011",
  12945=>"100000100",
  12946=>"001010111",
  12947=>"111101100",
  12948=>"000000010",
  12949=>"101010111",
  12950=>"111110100",
  12951=>"011000000",
  12952=>"110010010",
  12953=>"000100100",
  12954=>"011101011",
  12955=>"010110100",
  12956=>"001000111",
  12957=>"111111001",
  12958=>"111011010",
  12959=>"100110100",
  12960=>"000010100",
  12961=>"101010100",
  12962=>"011000011",
  12963=>"101110010",
  12964=>"010001100",
  12965=>"000000001",
  12966=>"101000000",
  12967=>"011010110",
  12968=>"011010000",
  12969=>"000000110",
  12970=>"110100000",
  12971=>"011101110",
  12972=>"111110001",
  12973=>"010110010",
  12974=>"001011001",
  12975=>"111011010",
  12976=>"011010000",
  12977=>"010111010",
  12978=>"110110000",
  12979=>"101110100",
  12980=>"001010101",
  12981=>"111111110",
  12982=>"111000110",
  12983=>"100000100",
  12984=>"001011001",
  12985=>"110010100",
  12986=>"111110111",
  12987=>"011101100",
  12988=>"100000101",
  12989=>"001011010",
  12990=>"111000011",
  12991=>"011100100",
  12992=>"101111101",
  12993=>"011111101",
  12994=>"001000011",
  12995=>"010101010",
  12996=>"010011101",
  12997=>"001100110",
  12998=>"011111000",
  12999=>"110011100",
  13000=>"111100101",
  13001=>"110010001",
  13002=>"001001011",
  13003=>"100011001",
  13004=>"111011111",
  13005=>"000101010",
  13006=>"001101010",
  13007=>"011100110",
  13008=>"101100100",
  13009=>"110100100",
  13010=>"010110000",
  13011=>"001101110",
  13012=>"001010011",
  13013=>"101110101",
  13014=>"100011111",
  13015=>"000111011",
  13016=>"100000100",
  13017=>"111111101",
  13018=>"110001100",
  13019=>"000101100",
  13020=>"010101100",
  13021=>"110100011",
  13022=>"100011001",
  13023=>"100000010",
  13024=>"010110000",
  13025=>"101110111",
  13026=>"000100000",
  13027=>"110111010",
  13028=>"000000110",
  13029=>"110110110",
  13030=>"010000100",
  13031=>"110101101",
  13032=>"011110100",
  13033=>"100001010",
  13034=>"011100100",
  13035=>"000010000",
  13036=>"010111101",
  13037=>"101111100",
  13038=>"101011010",
  13039=>"100100011",
  13040=>"010000011",
  13041=>"110001100",
  13042=>"010010011",
  13043=>"000000110",
  13044=>"110001101",
  13045=>"011010100",
  13046=>"100110111",
  13047=>"011010000",
  13048=>"101101010",
  13049=>"110110101",
  13050=>"001100100",
  13051=>"100100101",
  13052=>"011000110",
  13053=>"000110001",
  13054=>"101110011",
  13055=>"011011101",
  13056=>"000101101",
  13057=>"011110000",
  13058=>"111000000",
  13059=>"000111000",
  13060=>"010111111",
  13061=>"101100010",
  13062=>"111111110",
  13063=>"011110110",
  13064=>"100010011",
  13065=>"110010101",
  13066=>"100001111",
  13067=>"010000100",
  13068=>"011101000",
  13069=>"101001000",
  13070=>"001000011",
  13071=>"000100001",
  13072=>"110110010",
  13073=>"001001000",
  13074=>"110101111",
  13075=>"011001000",
  13076=>"011101111",
  13077=>"011111101",
  13078=>"001000111",
  13079=>"111101101",
  13080=>"010111100",
  13081=>"101000010",
  13082=>"010111110",
  13083=>"000000000",
  13084=>"100101111",
  13085=>"101000001",
  13086=>"010000101",
  13087=>"100001100",
  13088=>"111100000",
  13089=>"010010011",
  13090=>"101000111",
  13091=>"100100111",
  13092=>"111001001",
  13093=>"110010100",
  13094=>"011100001",
  13095=>"110010010",
  13096=>"100111100",
  13097=>"011100110",
  13098=>"100010101",
  13099=>"000100010",
  13100=>"010010010",
  13101=>"010010100",
  13102=>"010100111",
  13103=>"001000010",
  13104=>"011101100",
  13105=>"001010000",
  13106=>"100001001",
  13107=>"101010100",
  13108=>"100000000",
  13109=>"010111101",
  13110=>"110100000",
  13111=>"000111011",
  13112=>"001011101",
  13113=>"001000101",
  13114=>"000010110",
  13115=>"011000111",
  13116=>"110010010",
  13117=>"100101111",
  13118=>"001100110",
  13119=>"010100100",
  13120=>"000011100",
  13121=>"001011010",
  13122=>"111010100",
  13123=>"100001010",
  13124=>"001100011",
  13125=>"010110011",
  13126=>"101010111",
  13127=>"000110101",
  13128=>"010100111",
  13129=>"000010111",
  13130=>"000011100",
  13131=>"001000000",
  13132=>"110000100",
  13133=>"000000110",
  13134=>"111000100",
  13135=>"111000011",
  13136=>"000100110",
  13137=>"000100010",
  13138=>"100001100",
  13139=>"001111111",
  13140=>"011101100",
  13141=>"111000110",
  13142=>"000100010",
  13143=>"110101110",
  13144=>"000001100",
  13145=>"111101011",
  13146=>"001110000",
  13147=>"110110010",
  13148=>"011010110",
  13149=>"111111011",
  13150=>"111000100",
  13151=>"100101001",
  13152=>"111101110",
  13153=>"101010011",
  13154=>"100100100",
  13155=>"111101101",
  13156=>"011111011",
  13157=>"100010110",
  13158=>"010000100",
  13159=>"010010001",
  13160=>"001100011",
  13161=>"000011110",
  13162=>"110001110",
  13163=>"100100111",
  13164=>"110100101",
  13165=>"101101110",
  13166=>"001101000",
  13167=>"001111111",
  13168=>"111001000",
  13169=>"010000001",
  13170=>"000010110",
  13171=>"111100001",
  13172=>"000100110",
  13173=>"001001100",
  13174=>"111001010",
  13175=>"100101111",
  13176=>"110011101",
  13177=>"110100010",
  13178=>"010110101",
  13179=>"111010100",
  13180=>"000100101",
  13181=>"010110000",
  13182=>"001011100",
  13183=>"011011110",
  13184=>"111011010",
  13185=>"011001110",
  13186=>"001001101",
  13187=>"110101101",
  13188=>"101000101",
  13189=>"000110111",
  13190=>"001101101",
  13191=>"000000010",
  13192=>"101111111",
  13193=>"100111100",
  13194=>"010001101",
  13195=>"000011100",
  13196=>"100001110",
  13197=>"110010011",
  13198=>"011010100",
  13199=>"000111111",
  13200=>"001100000",
  13201=>"000111100",
  13202=>"100101010",
  13203=>"011100100",
  13204=>"010101100",
  13205=>"011111110",
  13206=>"001101100",
  13207=>"011100111",
  13208=>"001101010",
  13209=>"010100111",
  13210=>"011010101",
  13211=>"000111100",
  13212=>"011001011",
  13213=>"111010011",
  13214=>"000010111",
  13215=>"001111111",
  13216=>"000010100",
  13217=>"010010000",
  13218=>"001000011",
  13219=>"100111001",
  13220=>"101100000",
  13221=>"011100010",
  13222=>"011010110",
  13223=>"100110110",
  13224=>"010110001",
  13225=>"000010011",
  13226=>"010011101",
  13227=>"100000111",
  13228=>"111010001",
  13229=>"000010101",
  13230=>"010010100",
  13231=>"011101111",
  13232=>"001101010",
  13233=>"000101010",
  13234=>"010110111",
  13235=>"010100011",
  13236=>"101010110",
  13237=>"011011100",
  13238=>"110000000",
  13239=>"110110000",
  13240=>"000110000",
  13241=>"110001000",
  13242=>"010001000",
  13243=>"110001010",
  13244=>"000000101",
  13245=>"111100011",
  13246=>"010101011",
  13247=>"101000110",
  13248=>"010000101",
  13249=>"001101000",
  13250=>"101100001",
  13251=>"000111010",
  13252=>"100000100",
  13253=>"110101101",
  13254=>"110111110",
  13255=>"111100001",
  13256=>"100001111",
  13257=>"010010001",
  13258=>"001010011",
  13259=>"101000100",
  13260=>"010111001",
  13261=>"000000011",
  13262=>"001110100",
  13263=>"110011011",
  13264=>"001010011",
  13265=>"001011001",
  13266=>"011011010",
  13267=>"001110110",
  13268=>"010001100",
  13269=>"100100011",
  13270=>"011110111",
  13271=>"100010010",
  13272=>"111111000",
  13273=>"111001001",
  13274=>"010011010",
  13275=>"110000100",
  13276=>"111010100",
  13277=>"100011011",
  13278=>"000110101",
  13279=>"000011101",
  13280=>"111011010",
  13281=>"010010110",
  13282=>"110110010",
  13283=>"110110011",
  13284=>"000010010",
  13285=>"111100001",
  13286=>"001100111",
  13287=>"111100111",
  13288=>"100100100",
  13289=>"001011101",
  13290=>"010010001",
  13291=>"000101110",
  13292=>"010111100",
  13293=>"101010110",
  13294=>"101001101",
  13295=>"101100010",
  13296=>"110011111",
  13297=>"011100110",
  13298=>"011011011",
  13299=>"011110110",
  13300=>"001010011",
  13301=>"010001001",
  13302=>"101110001",
  13303=>"110111000",
  13304=>"001111001",
  13305=>"001110011",
  13306=>"101010000",
  13307=>"011111110",
  13308=>"110110111",
  13309=>"000010110",
  13310=>"000011000",
  13311=>"000101011",
  13312=>"110010010",
  13313=>"001100000",
  13314=>"111001000",
  13315=>"000111000",
  13316=>"100111111",
  13317=>"011011111",
  13318=>"101001001",
  13319=>"001000001",
  13320=>"111010000",
  13321=>"111010011",
  13322=>"001100111",
  13323=>"101100110",
  13324=>"001001010",
  13325=>"010101100",
  13326=>"111011010",
  13327=>"101000110",
  13328=>"001111011",
  13329=>"101011100",
  13330=>"101010100",
  13331=>"011000000",
  13332=>"101101111",
  13333=>"001100001",
  13334=>"110011110",
  13335=>"011011100",
  13336=>"011100110",
  13337=>"100100101",
  13338=>"101100000",
  13339=>"000010010",
  13340=>"001110100",
  13341=>"000010011",
  13342=>"111000001",
  13343=>"110110110",
  13344=>"100111010",
  13345=>"011101111",
  13346=>"010101011",
  13347=>"000001110",
  13348=>"000100001",
  13349=>"001010000",
  13350=>"000011010",
  13351=>"010000111",
  13352=>"000101010",
  13353=>"010001101",
  13354=>"011110101",
  13355=>"110101111",
  13356=>"101110101",
  13357=>"111001111",
  13358=>"001101101",
  13359=>"000011111",
  13360=>"001111111",
  13361=>"010111000",
  13362=>"000100010",
  13363=>"011010100",
  13364=>"011110110",
  13365=>"101101110",
  13366=>"001011010",
  13367=>"000110110",
  13368=>"001011101",
  13369=>"011011000",
  13370=>"100010100",
  13371=>"111111101",
  13372=>"011001111",
  13373=>"101010011",
  13374=>"100111001",
  13375=>"011110111",
  13376=>"110000000",
  13377=>"000000010",
  13378=>"001110110",
  13379=>"000111101",
  13380=>"000001101",
  13381=>"101001101",
  13382=>"110001011",
  13383=>"010000001",
  13384=>"011110011",
  13385=>"000000000",
  13386=>"111011111",
  13387=>"000000001",
  13388=>"011000001",
  13389=>"010010010",
  13390=>"110101101",
  13391=>"100000011",
  13392=>"100101010",
  13393=>"010110000",
  13394=>"101101111",
  13395=>"000011001",
  13396=>"000010110",
  13397=>"111101101",
  13398=>"111001100",
  13399=>"001110001",
  13400=>"010100011",
  13401=>"001100010",
  13402=>"001001000",
  13403=>"000110000",
  13404=>"111011110",
  13405=>"100100010",
  13406=>"111011011",
  13407=>"001101100",
  13408=>"101000111",
  13409=>"110011111",
  13410=>"001111100",
  13411=>"001001010",
  13412=>"111111111",
  13413=>"100111010",
  13414=>"111011100",
  13415=>"100111110",
  13416=>"011110110",
  13417=>"011110011",
  13418=>"011011111",
  13419=>"000010001",
  13420=>"111110001",
  13421=>"101001000",
  13422=>"100000011",
  13423=>"010001100",
  13424=>"010101000",
  13425=>"011000010",
  13426=>"100110000",
  13427=>"101100100",
  13428=>"010100111",
  13429=>"001001101",
  13430=>"100010111",
  13431=>"101110111",
  13432=>"110110100",
  13433=>"001011011",
  13434=>"011000100",
  13435=>"011111111",
  13436=>"000110011",
  13437=>"001110011",
  13438=>"011111010",
  13439=>"011100111",
  13440=>"101101000",
  13441=>"111010000",
  13442=>"110011011",
  13443=>"001011100",
  13444=>"110001011",
  13445=>"011001001",
  13446=>"010010110",
  13447=>"111110001",
  13448=>"100001000",
  13449=>"011110010",
  13450=>"110001001",
  13451=>"110010000",
  13452=>"000011001",
  13453=>"011111110",
  13454=>"101010000",
  13455=>"110110000",
  13456=>"100010001",
  13457=>"010001000",
  13458=>"111101101",
  13459=>"001010100",
  13460=>"000010001",
  13461=>"010101000",
  13462=>"000000010",
  13463=>"110101001",
  13464=>"110001010",
  13465=>"001001010",
  13466=>"000011110",
  13467=>"100000000",
  13468=>"011010000",
  13469=>"001011101",
  13470=>"111100010",
  13471=>"111100100",
  13472=>"000110000",
  13473=>"101101110",
  13474=>"101100000",
  13475=>"110111101",
  13476=>"000111111",
  13477=>"001011100",
  13478=>"011101110",
  13479=>"111111011",
  13480=>"101110110",
  13481=>"000010010",
  13482=>"011010000",
  13483=>"100111000",
  13484=>"001000110",
  13485=>"000000001",
  13486=>"100000101",
  13487=>"000010100",
  13488=>"001001110",
  13489=>"011011110",
  13490=>"100111110",
  13491=>"010111000",
  13492=>"101001110",
  13493=>"000101010",
  13494=>"110010000",
  13495=>"110000010",
  13496=>"000111011",
  13497=>"011100101",
  13498=>"000001011",
  13499=>"000101111",
  13500=>"110010001",
  13501=>"100000101",
  13502=>"011011001",
  13503=>"001100000",
  13504=>"010001111",
  13505=>"000101100",
  13506=>"100000000",
  13507=>"110101011",
  13508=>"101101100",
  13509=>"101010001",
  13510=>"100001010",
  13511=>"111100001",
  13512=>"001010111",
  13513=>"000011111",
  13514=>"100100111",
  13515=>"101101111",
  13516=>"100111110",
  13517=>"100011111",
  13518=>"010111101",
  13519=>"110001110",
  13520=>"101000110",
  13521=>"000111000",
  13522=>"010101010",
  13523=>"111100000",
  13524=>"111000011",
  13525=>"100000001",
  13526=>"000111110",
  13527=>"101101001",
  13528=>"000100001",
  13529=>"111000110",
  13530=>"001011011",
  13531=>"100000001",
  13532=>"011101011",
  13533=>"100111001",
  13534=>"111001111",
  13535=>"110001000",
  13536=>"111001000",
  13537=>"111100000",
  13538=>"111110100",
  13539=>"100100010",
  13540=>"010110100",
  13541=>"110000100",
  13542=>"000010101",
  13543=>"010010111",
  13544=>"100111000",
  13545=>"111111100",
  13546=>"011000000",
  13547=>"101110010",
  13548=>"000110001",
  13549=>"100101010",
  13550=>"100001001",
  13551=>"011001000",
  13552=>"001011010",
  13553=>"000000101",
  13554=>"101000111",
  13555=>"010101011",
  13556=>"010101111",
  13557=>"001101000",
  13558=>"101100111",
  13559=>"000100000",
  13560=>"101000010",
  13561=>"101011111",
  13562=>"001100001",
  13563=>"000010001",
  13564=>"000101001",
  13565=>"000000001",
  13566=>"001000100",
  13567=>"010101101",
  13568=>"110010011",
  13569=>"111010011",
  13570=>"010011101",
  13571=>"001011010",
  13572=>"111111010",
  13573=>"000101011",
  13574=>"111100101",
  13575=>"001001000",
  13576=>"011101100",
  13577=>"100000010",
  13578=>"010011100",
  13579=>"010010000",
  13580=>"000001101",
  13581=>"111010010",
  13582=>"011111001",
  13583=>"000111001",
  13584=>"110110010",
  13585=>"001111101",
  13586=>"101110100",
  13587=>"000000111",
  13588=>"101100110",
  13589=>"101101110",
  13590=>"001011011",
  13591=>"101000001",
  13592=>"111101001",
  13593=>"110001100",
  13594=>"010001111",
  13595=>"011111001",
  13596=>"001101001",
  13597=>"011000001",
  13598=>"110111000",
  13599=>"110011010",
  13600=>"000100111",
  13601=>"110001011",
  13602=>"101010100",
  13603=>"111110011",
  13604=>"110001101",
  13605=>"001100010",
  13606=>"111010000",
  13607=>"010100011",
  13608=>"101100101",
  13609=>"110100001",
  13610=>"110011011",
  13611=>"111011110",
  13612=>"000111010",
  13613=>"011011000",
  13614=>"100001011",
  13615=>"110010010",
  13616=>"001111100",
  13617=>"001100111",
  13618=>"100010010",
  13619=>"000010000",
  13620=>"100010000",
  13621=>"000110000",
  13622=>"110110111",
  13623=>"010010001",
  13624=>"000100001",
  13625=>"011100000",
  13626=>"011011011",
  13627=>"100111100",
  13628=>"110101010",
  13629=>"110010111",
  13630=>"101011111",
  13631=>"001011101",
  13632=>"111110000",
  13633=>"011001111",
  13634=>"100010010",
  13635=>"111101010",
  13636=>"110100100",
  13637=>"101010101",
  13638=>"001000110",
  13639=>"011110000",
  13640=>"110100110",
  13641=>"001100110",
  13642=>"111111010",
  13643=>"001011010",
  13644=>"111010111",
  13645=>"100010110",
  13646=>"101110110",
  13647=>"011001000",
  13648=>"101100000",
  13649=>"000010010",
  13650=>"011011101",
  13651=>"110101011",
  13652=>"101110011",
  13653=>"001110110",
  13654=>"110000110",
  13655=>"000110101",
  13656=>"010011111",
  13657=>"000000110",
  13658=>"110000111",
  13659=>"010111001",
  13660=>"010101011",
  13661=>"001100111",
  13662=>"100100110",
  13663=>"100000110",
  13664=>"011000110",
  13665=>"000100010",
  13666=>"110100111",
  13667=>"000010010",
  13668=>"010001011",
  13669=>"001100101",
  13670=>"000001100",
  13671=>"110000000",
  13672=>"100111111",
  13673=>"000100000",
  13674=>"111000010",
  13675=>"000101010",
  13676=>"010011010",
  13677=>"001010011",
  13678=>"001101001",
  13679=>"001010001",
  13680=>"001111001",
  13681=>"001011111",
  13682=>"001100011",
  13683=>"101001010",
  13684=>"110101011",
  13685=>"001111100",
  13686=>"100110100",
  13687=>"000000110",
  13688=>"011100010",
  13689=>"000101101",
  13690=>"111011001",
  13691=>"010100111",
  13692=>"101000110",
  13693=>"010000100",
  13694=>"000011110",
  13695=>"000100000",
  13696=>"101110010",
  13697=>"000110110",
  13698=>"111011011",
  13699=>"100110010",
  13700=>"001001001",
  13701=>"000010010",
  13702=>"101000111",
  13703=>"011001110",
  13704=>"110000110",
  13705=>"000000011",
  13706=>"000000100",
  13707=>"011000111",
  13708=>"111001001",
  13709=>"010110010",
  13710=>"010010001",
  13711=>"111011111",
  13712=>"110101100",
  13713=>"100001010",
  13714=>"111010001",
  13715=>"100101111",
  13716=>"110010111",
  13717=>"000110001",
  13718=>"001010001",
  13719=>"011000011",
  13720=>"101111000",
  13721=>"000111110",
  13722=>"101111110",
  13723=>"010100001",
  13724=>"010011110",
  13725=>"001100111",
  13726=>"110010010",
  13727=>"101100111",
  13728=>"011100010",
  13729=>"111000010",
  13730=>"001001110",
  13731=>"011001101",
  13732=>"110000110",
  13733=>"000111111",
  13734=>"011110001",
  13735=>"001010011",
  13736=>"011001000",
  13737=>"110001111",
  13738=>"000010011",
  13739=>"101011110",
  13740=>"000110000",
  13741=>"001001011",
  13742=>"010000011",
  13743=>"011101101",
  13744=>"101000101",
  13745=>"111010001",
  13746=>"100111011",
  13747=>"110010011",
  13748=>"111000111",
  13749=>"110000111",
  13750=>"001011001",
  13751=>"111110011",
  13752=>"010010000",
  13753=>"110100110",
  13754=>"001101010",
  13755=>"100011010",
  13756=>"111010001",
  13757=>"100100100",
  13758=>"011101110",
  13759=>"101011100",
  13760=>"000101100",
  13761=>"011100111",
  13762=>"000101001",
  13763=>"011010110",
  13764=>"011110010",
  13765=>"010001111",
  13766=>"000001001",
  13767=>"001100000",
  13768=>"100000110",
  13769=>"100011111",
  13770=>"100000101",
  13771=>"110110101",
  13772=>"011111001",
  13773=>"111001110",
  13774=>"000110001",
  13775=>"001001100",
  13776=>"101111001",
  13777=>"110010011",
  13778=>"111001001",
  13779=>"101000011",
  13780=>"111011110",
  13781=>"100111001",
  13782=>"100100111",
  13783=>"110010000",
  13784=>"000010100",
  13785=>"111001111",
  13786=>"010100010",
  13787=>"100100110",
  13788=>"001100011",
  13789=>"101100000",
  13790=>"110111011",
  13791=>"110100111",
  13792=>"101010111",
  13793=>"011110100",
  13794=>"000001011",
  13795=>"001100111",
  13796=>"110010111",
  13797=>"100011001",
  13798=>"111110011",
  13799=>"000100110",
  13800=>"101010000",
  13801=>"100100001",
  13802=>"001001100",
  13803=>"000001011",
  13804=>"001000010",
  13805=>"111000101",
  13806=>"101101110",
  13807=>"100000011",
  13808=>"111000000",
  13809=>"101000011",
  13810=>"111001000",
  13811=>"111110101",
  13812=>"100010001",
  13813=>"001000100",
  13814=>"111111101",
  13815=>"001100000",
  13816=>"110000110",
  13817=>"111000001",
  13818=>"010100011",
  13819=>"100111010",
  13820=>"111110111",
  13821=>"101101010",
  13822=>"101101100",
  13823=>"100011110",
  13824=>"011101010",
  13825=>"010101001",
  13826=>"001000001",
  13827=>"000001001",
  13828=>"011011011",
  13829=>"110000001",
  13830=>"011011011",
  13831=>"010101101",
  13832=>"000000010",
  13833=>"111000000",
  13834=>"110110110",
  13835=>"100011111",
  13836=>"101001111",
  13837=>"000000111",
  13838=>"111100111",
  13839=>"111011010",
  13840=>"111010100",
  13841=>"110100111",
  13842=>"111010011",
  13843=>"111100110",
  13844=>"110000000",
  13845=>"110000011",
  13846=>"010010111",
  13847=>"001111011",
  13848=>"000111000",
  13849=>"101000110",
  13850=>"111101000",
  13851=>"010001010",
  13852=>"101011110",
  13853=>"110101001",
  13854=>"111100000",
  13855=>"100000101",
  13856=>"101110011",
  13857=>"100101001",
  13858=>"011010000",
  13859=>"101111011",
  13860=>"110010101",
  13861=>"000010001",
  13862=>"110100011",
  13863=>"101011100",
  13864=>"110000100",
  13865=>"010111011",
  13866=>"001001010",
  13867=>"111110000",
  13868=>"101000000",
  13869=>"000011111",
  13870=>"010001000",
  13871=>"101001101",
  13872=>"011110101",
  13873=>"010010110",
  13874=>"011001101",
  13875=>"000001101",
  13876=>"011111110",
  13877=>"101010110",
  13878=>"010000001",
  13879=>"001100100",
  13880=>"110010010",
  13881=>"110101110",
  13882=>"011000001",
  13883=>"111101110",
  13884=>"010111010",
  13885=>"000110000",
  13886=>"000010000",
  13887=>"100011001",
  13888=>"010001110",
  13889=>"000010110",
  13890=>"111001011",
  13891=>"010101010",
  13892=>"010110000",
  13893=>"100100011",
  13894=>"010000010",
  13895=>"000011110",
  13896=>"111001001",
  13897=>"000111010",
  13898=>"110000011",
  13899=>"000100001",
  13900=>"101110111",
  13901=>"101111001",
  13902=>"001001101",
  13903=>"010101011",
  13904=>"110101000",
  13905=>"010011100",
  13906=>"000001100",
  13907=>"011001100",
  13908=>"011000100",
  13909=>"110001001",
  13910=>"000011010",
  13911=>"101000111",
  13912=>"111001101",
  13913=>"010001010",
  13914=>"110010101",
  13915=>"011110111",
  13916=>"010010111",
  13917=>"100100000",
  13918=>"100100001",
  13919=>"101110010",
  13920=>"110000010",
  13921=>"101111000",
  13922=>"010111110",
  13923=>"100111001",
  13924=>"011000001",
  13925=>"000000101",
  13926=>"011111011",
  13927=>"011011111",
  13928=>"110101011",
  13929=>"000010101",
  13930=>"111111110",
  13931=>"000001000",
  13932=>"101110011",
  13933=>"010011100",
  13934=>"001000001",
  13935=>"110111110",
  13936=>"110011111",
  13937=>"001000010",
  13938=>"101111100",
  13939=>"011101110",
  13940=>"001100111",
  13941=>"111011101",
  13942=>"111100110",
  13943=>"101111100",
  13944=>"101101000",
  13945=>"100010011",
  13946=>"100111000",
  13947=>"100100110",
  13948=>"111111001",
  13949=>"100001001",
  13950=>"110011001",
  13951=>"001110010",
  13952=>"010111000",
  13953=>"000100011",
  13954=>"110100011",
  13955=>"001000100",
  13956=>"010101101",
  13957=>"010101000",
  13958=>"000011101",
  13959=>"000011000",
  13960=>"000100001",
  13961=>"000111001",
  13962=>"000000110",
  13963=>"000000101",
  13964=>"111001111",
  13965=>"011001010",
  13966=>"001111110",
  13967=>"010000100",
  13968=>"110001000",
  13969=>"110101110",
  13970=>"010100001",
  13971=>"001001010",
  13972=>"011110000",
  13973=>"100001000",
  13974=>"001000111",
  13975=>"110100001",
  13976=>"100010101",
  13977=>"111110000",
  13978=>"111111010",
  13979=>"000110000",
  13980=>"110001011",
  13981=>"001111000",
  13982=>"011011011",
  13983=>"110101011",
  13984=>"100110001",
  13985=>"010011001",
  13986=>"000000001",
  13987=>"101000101",
  13988=>"010111111",
  13989=>"000001001",
  13990=>"100000000",
  13991=>"000001000",
  13992=>"011010010",
  13993=>"101110101",
  13994=>"010010110",
  13995=>"001000000",
  13996=>"010100010",
  13997=>"111000010",
  13998=>"100010110",
  13999=>"011000010",
  14000=>"000110100",
  14001=>"100110101",
  14002=>"111011001",
  14003=>"000000110",
  14004=>"100010010",
  14005=>"110100010",
  14006=>"111111100",
  14007=>"001010010",
  14008=>"101010001",
  14009=>"101100000",
  14010=>"011001001",
  14011=>"111101101",
  14012=>"101100100",
  14013=>"010010000",
  14014=>"010101111",
  14015=>"101000101",
  14016=>"011010100",
  14017=>"101111111",
  14018=>"000001010",
  14019=>"000000111",
  14020=>"000110011",
  14021=>"110011111",
  14022=>"110100001",
  14023=>"000010011",
  14024=>"111010100",
  14025=>"001111100",
  14026=>"000000011",
  14027=>"111011100",
  14028=>"011011110",
  14029=>"111100001",
  14030=>"101111000",
  14031=>"100101001",
  14032=>"000010010",
  14033=>"101111011",
  14034=>"111101000",
  14035=>"010010000",
  14036=>"110001011",
  14037=>"110001001",
  14038=>"011011110",
  14039=>"011110100",
  14040=>"011111101",
  14041=>"000010011",
  14042=>"111000111",
  14043=>"110010011",
  14044=>"101100011",
  14045=>"001010001",
  14046=>"010010101",
  14047=>"100111110",
  14048=>"110100001",
  14049=>"001110000",
  14050=>"000011111",
  14051=>"100111111",
  14052=>"110101101",
  14053=>"001110000",
  14054=>"101001000",
  14055=>"000111110",
  14056=>"000101101",
  14057=>"101111001",
  14058=>"011111111",
  14059=>"110100011",
  14060=>"101101011",
  14061=>"000100011",
  14062=>"001100010",
  14063=>"010110101",
  14064=>"111111110",
  14065=>"100001001",
  14066=>"001101100",
  14067=>"101010100",
  14068=>"111010000",
  14069=>"100010001",
  14070=>"100111010",
  14071=>"111010010",
  14072=>"001110011",
  14073=>"110101000",
  14074=>"110111000",
  14075=>"100010000",
  14076=>"001101010",
  14077=>"111111001",
  14078=>"110011111",
  14079=>"110010110",
  14080=>"100110010",
  14081=>"011110001",
  14082=>"011110110",
  14083=>"010100001",
  14084=>"001111100",
  14085=>"111010111",
  14086=>"001110101",
  14087=>"011011110",
  14088=>"011100111",
  14089=>"010011111",
  14090=>"010111111",
  14091=>"101110001",
  14092=>"100001101",
  14093=>"101100101",
  14094=>"110101010",
  14095=>"001011101",
  14096=>"001100110",
  14097=>"000001011",
  14098=>"011100000",
  14099=>"100011011",
  14100=>"000011111",
  14101=>"110111000",
  14102=>"100100000",
  14103=>"111011100",
  14104=>"010001110",
  14105=>"100100110",
  14106=>"010111011",
  14107=>"011010001",
  14108=>"001001111",
  14109=>"011001110",
  14110=>"100001111",
  14111=>"111110010",
  14112=>"010010111",
  14113=>"000001000",
  14114=>"011010001",
  14115=>"110010111",
  14116=>"110100100",
  14117=>"110110101",
  14118=>"010010101",
  14119=>"101101011",
  14120=>"010100001",
  14121=>"101000100",
  14122=>"101011011",
  14123=>"110101111",
  14124=>"100110011",
  14125=>"001011101",
  14126=>"010010000",
  14127=>"000010011",
  14128=>"000111011",
  14129=>"000010011",
  14130=>"000000101",
  14131=>"001101000",
  14132=>"010011110",
  14133=>"100110100",
  14134=>"110111010",
  14135=>"000011101",
  14136=>"011111100",
  14137=>"011010100",
  14138=>"000111100",
  14139=>"110100000",
  14140=>"000100011",
  14141=>"110101110",
  14142=>"110110001",
  14143=>"101111100",
  14144=>"001010011",
  14145=>"110100001",
  14146=>"100001010",
  14147=>"010011011",
  14148=>"100011101",
  14149=>"001010000",
  14150=>"100111001",
  14151=>"011101101",
  14152=>"100100100",
  14153=>"010001110",
  14154=>"011000110",
  14155=>"110011100",
  14156=>"001000001",
  14157=>"110000100",
  14158=>"000000101",
  14159=>"000000000",
  14160=>"000000111",
  14161=>"110010011",
  14162=>"010010001",
  14163=>"001010101",
  14164=>"010111000",
  14165=>"110101101",
  14166=>"000101110",
  14167=>"001101000",
  14168=>"111000100",
  14169=>"110001100",
  14170=>"011111111",
  14171=>"011111001",
  14172=>"010100000",
  14173=>"100100001",
  14174=>"011111111",
  14175=>"010000000",
  14176=>"000000101",
  14177=>"110101001",
  14178=>"010100011",
  14179=>"100011000",
  14180=>"010011010",
  14181=>"000110001",
  14182=>"110000111",
  14183=>"100110110",
  14184=>"111100001",
  14185=>"010100111",
  14186=>"011101001",
  14187=>"100011010",
  14188=>"010000011",
  14189=>"011011011",
  14190=>"111010111",
  14191=>"011000100",
  14192=>"110100001",
  14193=>"010010011",
  14194=>"011011101",
  14195=>"000111111",
  14196=>"100111000",
  14197=>"001010010",
  14198=>"100010010",
  14199=>"011101101",
  14200=>"000100111",
  14201=>"101010111",
  14202=>"001100101",
  14203=>"010100001",
  14204=>"011011011",
  14205=>"010100100",
  14206=>"010000001",
  14207=>"011001100",
  14208=>"100111111",
  14209=>"101011110",
  14210=>"010001010",
  14211=>"100101011",
  14212=>"110101110",
  14213=>"111101001",
  14214=>"000001101",
  14215=>"000010011",
  14216=>"001110011",
  14217=>"011010000",
  14218=>"110000100",
  14219=>"011110110",
  14220=>"111001001",
  14221=>"111100010",
  14222=>"011110110",
  14223=>"111110100",
  14224=>"000111000",
  14225=>"111111110",
  14226=>"101001100",
  14227=>"110001100",
  14228=>"001100000",
  14229=>"000001000",
  14230=>"100110000",
  14231=>"110111001",
  14232=>"111111001",
  14233=>"000010000",
  14234=>"000110001",
  14235=>"000011001",
  14236=>"100101100",
  14237=>"011100010",
  14238=>"100101101",
  14239=>"001110000",
  14240=>"101010100",
  14241=>"010000101",
  14242=>"100000100",
  14243=>"101000100",
  14244=>"001100010",
  14245=>"110000001",
  14246=>"101000100",
  14247=>"001011100",
  14248=>"000011000",
  14249=>"101000101",
  14250=>"110000111",
  14251=>"000100110",
  14252=>"100110000",
  14253=>"100000011",
  14254=>"101110100",
  14255=>"110100100",
  14256=>"110111011",
  14257=>"010100111",
  14258=>"000100111",
  14259=>"011000011",
  14260=>"010100101",
  14261=>"001001001",
  14262=>"011111101",
  14263=>"100110011",
  14264=>"000010101",
  14265=>"011001011",
  14266=>"111110000",
  14267=>"001010010",
  14268=>"101110110",
  14269=>"010011000",
  14270=>"000111011",
  14271=>"000100010",
  14272=>"001011100",
  14273=>"001001110",
  14274=>"000110000",
  14275=>"100100010",
  14276=>"000110001",
  14277=>"101011010",
  14278=>"111010001",
  14279=>"110100010",
  14280=>"111011001",
  14281=>"010100011",
  14282=>"100111111",
  14283=>"101111101",
  14284=>"111010101",
  14285=>"110000110",
  14286=>"001001101",
  14287=>"011100001",
  14288=>"010111101",
  14289=>"001010111",
  14290=>"111000111",
  14291=>"011011000",
  14292=>"011110111",
  14293=>"111000110",
  14294=>"010011111",
  14295=>"100001000",
  14296=>"010000111",
  14297=>"000010010",
  14298=>"010110110",
  14299=>"101110010",
  14300=>"001100110",
  14301=>"111111011",
  14302=>"100110111",
  14303=>"111101100",
  14304=>"000000000",
  14305=>"101011011",
  14306=>"101110010",
  14307=>"010111100",
  14308=>"000101011",
  14309=>"100001101",
  14310=>"011100010",
  14311=>"011110011",
  14312=>"110100010",
  14313=>"111100110",
  14314=>"000101001",
  14315=>"000001010",
  14316=>"111111001",
  14317=>"011101010",
  14318=>"111001001",
  14319=>"111100100",
  14320=>"000110110",
  14321=>"011011000",
  14322=>"001001000",
  14323=>"010011111",
  14324=>"010100100",
  14325=>"111101111",
  14326=>"011101001",
  14327=>"000101101",
  14328=>"011001111",
  14329=>"000110100",
  14330=>"111111000",
  14331=>"000001001",
  14332=>"101110011",
  14333=>"010011111",
  14334=>"001110110",
  14335=>"111110001",
  14336=>"011111111",
  14337=>"101001010",
  14338=>"011101111",
  14339=>"110101000",
  14340=>"001101000",
  14341=>"010011001",
  14342=>"011111111",
  14343=>"111001000",
  14344=>"101011010",
  14345=>"010010111",
  14346=>"111011101",
  14347=>"101111000",
  14348=>"010010000",
  14349=>"011111110",
  14350=>"000100010",
  14351=>"000111111",
  14352=>"011001101",
  14353=>"010001010",
  14354=>"010101110",
  14355=>"010000100",
  14356=>"011011101",
  14357=>"000000111",
  14358=>"000011100",
  14359=>"010001011",
  14360=>"001100101",
  14361=>"110001001",
  14362=>"001001110",
  14363=>"011101001",
  14364=>"000101011",
  14365=>"010110100",
  14366=>"001001000",
  14367=>"010111111",
  14368=>"110011101",
  14369=>"111000000",
  14370=>"010010010",
  14371=>"110010111",
  14372=>"110001101",
  14373=>"110010110",
  14374=>"111100101",
  14375=>"001010010",
  14376=>"011110010",
  14377=>"111111001",
  14378=>"101111011",
  14379=>"001101100",
  14380=>"010001010",
  14381=>"101110001",
  14382=>"011100010",
  14383=>"011011101",
  14384=>"100110110",
  14385=>"111111111",
  14386=>"000101111",
  14387=>"001111011",
  14388=>"000111101",
  14389=>"111010111",
  14390=>"100111011",
  14391=>"101111011",
  14392=>"001110110",
  14393=>"011101001",
  14394=>"111111100",
  14395=>"100000000",
  14396=>"110101000",
  14397=>"111000001",
  14398=>"010111100",
  14399=>"000100001",
  14400=>"011000100",
  14401=>"011011010",
  14402=>"001010110",
  14403=>"011111111",
  14404=>"110110000",
  14405=>"111010110",
  14406=>"111010110",
  14407=>"000001011",
  14408=>"011110111",
  14409=>"111110110",
  14410=>"010000001",
  14411=>"001110110",
  14412=>"000011111",
  14413=>"110110000",
  14414=>"001001001",
  14415=>"101101101",
  14416=>"000010011",
  14417=>"011000101",
  14418=>"110111000",
  14419=>"100000111",
  14420=>"001111111",
  14421=>"011101010",
  14422=>"110110101",
  14423=>"111011010",
  14424=>"110011011",
  14425=>"000000111",
  14426=>"111111001",
  14427=>"001100000",
  14428=>"110101011",
  14429=>"101100110",
  14430=>"100111001",
  14431=>"100011100",
  14432=>"000011010",
  14433=>"000010101",
  14434=>"001001001",
  14435=>"001111001",
  14436=>"000110100",
  14437=>"010101101",
  14438=>"111111011",
  14439=>"001100110",
  14440=>"111110000",
  14441=>"101101111",
  14442=>"100000000",
  14443=>"101110011",
  14444=>"010110101",
  14445=>"000111100",
  14446=>"000110000",
  14447=>"000011011",
  14448=>"000100000",
  14449=>"000000010",
  14450=>"100010010",
  14451=>"001110111",
  14452=>"010010101",
  14453=>"001001100",
  14454=>"110110010",
  14455=>"000010000",
  14456=>"110111010",
  14457=>"010001101",
  14458=>"111101011",
  14459=>"000001011",
  14460=>"001001010",
  14461=>"000000001",
  14462=>"000001010",
  14463=>"001000111",
  14464=>"010000100",
  14465=>"011100100",
  14466=>"000000000",
  14467=>"010100010",
  14468=>"011010111",
  14469=>"011110101",
  14470=>"100011111",
  14471=>"111010100",
  14472=>"110000110",
  14473=>"100001111",
  14474=>"100000001",
  14475=>"100110110",
  14476=>"100001111",
  14477=>"000111001",
  14478=>"010001010",
  14479=>"001000000",
  14480=>"110100000",
  14481=>"011011010",
  14482=>"100110100",
  14483=>"101000010",
  14484=>"101000000",
  14485=>"011000011",
  14486=>"011000000",
  14487=>"110011011",
  14488=>"010001000",
  14489=>"000011101",
  14490=>"011100111",
  14491=>"110010101",
  14492=>"101111111",
  14493=>"011011110",
  14494=>"101110000",
  14495=>"010001001",
  14496=>"100011001",
  14497=>"100010110",
  14498=>"010100000",
  14499=>"101111100",
  14500=>"100000111",
  14501=>"100011110",
  14502=>"010111000",
  14503=>"101010110",
  14504=>"001000101",
  14505=>"110100110",
  14506=>"000110000",
  14507=>"011100001",
  14508=>"000110110",
  14509=>"111010110",
  14510=>"000010000",
  14511=>"111010100",
  14512=>"101100100",
  14513=>"001101001",
  14514=>"001011101",
  14515=>"110100001",
  14516=>"111111001",
  14517=>"110000100",
  14518=>"111011101",
  14519=>"000011000",
  14520=>"101110111",
  14521=>"110001100",
  14522=>"000010000",
  14523=>"001001010",
  14524=>"010101101",
  14525=>"110100110",
  14526=>"110101011",
  14527=>"111000001",
  14528=>"001100001",
  14529=>"000000101",
  14530=>"000101011",
  14531=>"011111010",
  14532=>"110000001",
  14533=>"001000010",
  14534=>"111101111",
  14535=>"000011111",
  14536=>"010000010",
  14537=>"000111011",
  14538=>"111001000",
  14539=>"100111111",
  14540=>"010000000",
  14541=>"010111011",
  14542=>"101001001",
  14543=>"000000000",
  14544=>"011000000",
  14545=>"010010110",
  14546=>"001000101",
  14547=>"111011111",
  14548=>"010001111",
  14549=>"100011111",
  14550=>"000100001",
  14551=>"010111110",
  14552=>"101111001",
  14553=>"110101110",
  14554=>"100111100",
  14555=>"110000000",
  14556=>"000100000",
  14557=>"100100000",
  14558=>"000110111",
  14559=>"111010011",
  14560=>"110100101",
  14561=>"000110111",
  14562=>"000000101",
  14563=>"011000011",
  14564=>"110001110",
  14565=>"011001100",
  14566=>"101101000",
  14567=>"110111110",
  14568=>"101001011",
  14569=>"010010011",
  14570=>"000110111",
  14571=>"100111001",
  14572=>"001000000",
  14573=>"011101011",
  14574=>"000001101",
  14575=>"111111000",
  14576=>"101100100",
  14577=>"101010111",
  14578=>"001100110",
  14579=>"000000101",
  14580=>"110001010",
  14581=>"111111000",
  14582=>"111100010",
  14583=>"111010111",
  14584=>"000011000",
  14585=>"001010001",
  14586=>"000100111",
  14587=>"001001110",
  14588=>"000101000",
  14589=>"011100101",
  14590=>"100101001",
  14591=>"001111010",
  14592=>"001000011",
  14593=>"111000100",
  14594=>"011011011",
  14595=>"110100000",
  14596=>"110110001",
  14597=>"001000000",
  14598=>"001001000",
  14599=>"011010100",
  14600=>"011011001",
  14601=>"011101101",
  14602=>"100111000",
  14603=>"111000101",
  14604=>"101011111",
  14605=>"101100110",
  14606=>"100100110",
  14607=>"001000110",
  14608=>"111011001",
  14609=>"100111100",
  14610=>"001100000",
  14611=>"100101010",
  14612=>"110000111",
  14613=>"111111100",
  14614=>"110001100",
  14615=>"000000111",
  14616=>"111100001",
  14617=>"100110001",
  14618=>"011100011",
  14619=>"101010100",
  14620=>"111101011",
  14621=>"101011110",
  14622=>"001111011",
  14623=>"010000010",
  14624=>"010101110",
  14625=>"110110011",
  14626=>"001101101",
  14627=>"100010111",
  14628=>"000111110",
  14629=>"110110000",
  14630=>"000110111",
  14631=>"100011100",
  14632=>"011111111",
  14633=>"110010111",
  14634=>"011110000",
  14635=>"110010110",
  14636=>"001010001",
  14637=>"010010011",
  14638=>"000100100",
  14639=>"011001001",
  14640=>"111101001",
  14641=>"111000010",
  14642=>"110010101",
  14643=>"000001011",
  14644=>"110010110",
  14645=>"100110110",
  14646=>"000100110",
  14647=>"100110000",
  14648=>"111101001",
  14649=>"000010000",
  14650=>"010001100",
  14651=>"101000110",
  14652=>"101001100",
  14653=>"001111000",
  14654=>"110110001",
  14655=>"111001111",
  14656=>"010010110",
  14657=>"100110111",
  14658=>"000001100",
  14659=>"110001101",
  14660=>"001011001",
  14661=>"101110110",
  14662=>"110000010",
  14663=>"000011110",
  14664=>"111001000",
  14665=>"000001100",
  14666=>"111000101",
  14667=>"001110011",
  14668=>"111011000",
  14669=>"001101011",
  14670=>"101111011",
  14671=>"111111000",
  14672=>"011000010",
  14673=>"000110110",
  14674=>"001111110",
  14675=>"000100000",
  14676=>"110000000",
  14677=>"111101101",
  14678=>"010000110",
  14679=>"000001001",
  14680=>"110101001",
  14681=>"101101010",
  14682=>"010010001",
  14683=>"010001010",
  14684=>"010110111",
  14685=>"000101100",
  14686=>"111010000",
  14687=>"100100000",
  14688=>"111010101",
  14689=>"001100001",
  14690=>"001110000",
  14691=>"000001000",
  14692=>"010100011",
  14693=>"010001000",
  14694=>"011110100",
  14695=>"101111001",
  14696=>"100110011",
  14697=>"011001001",
  14698=>"010100011",
  14699=>"101000111",
  14700=>"111110101",
  14701=>"100101000",
  14702=>"010100010",
  14703=>"110110100",
  14704=>"000011111",
  14705=>"001011100",
  14706=>"000101110",
  14707=>"001010011",
  14708=>"001101111",
  14709=>"010011001",
  14710=>"000101000",
  14711=>"010000111",
  14712=>"000111011",
  14713=>"001001101",
  14714=>"000110010",
  14715=>"111010111",
  14716=>"111010111",
  14717=>"110101101",
  14718=>"011010010",
  14719=>"111011101",
  14720=>"110010101",
  14721=>"101000100",
  14722=>"010011011",
  14723=>"011001110",
  14724=>"011101100",
  14725=>"000000000",
  14726=>"010111110",
  14727=>"011010111",
  14728=>"100100010",
  14729=>"001010010",
  14730=>"000001010",
  14731=>"000011110",
  14732=>"010001010",
  14733=>"101101010",
  14734=>"100001101",
  14735=>"011110100",
  14736=>"000110110",
  14737=>"011010001",
  14738=>"101000000",
  14739=>"011100011",
  14740=>"001101111",
  14741=>"011111000",
  14742=>"010101001",
  14743=>"101001000",
  14744=>"110010111",
  14745=>"111110000",
  14746=>"110100011",
  14747=>"001111101",
  14748=>"000011110",
  14749=>"111011110",
  14750=>"001100100",
  14751=>"000101000",
  14752=>"101010000",
  14753=>"011010011",
  14754=>"010000111",
  14755=>"100000110",
  14756=>"111110000",
  14757=>"010011011",
  14758=>"111011111",
  14759=>"010000110",
  14760=>"000011011",
  14761=>"010100010",
  14762=>"010011101",
  14763=>"000000001",
  14764=>"111110101",
  14765=>"101000110",
  14766=>"010111010",
  14767=>"110000111",
  14768=>"111011101",
  14769=>"110110110",
  14770=>"111110101",
  14771=>"111100001",
  14772=>"001000100",
  14773=>"110100011",
  14774=>"001011101",
  14775=>"100110111",
  14776=>"110111111",
  14777=>"100011000",
  14778=>"111001100",
  14779=>"000011001",
  14780=>"111000010",
  14781=>"010111001",
  14782=>"101000000",
  14783=>"101100011",
  14784=>"010001111",
  14785=>"010100101",
  14786=>"110011111",
  14787=>"001100001",
  14788=>"101100111",
  14789=>"010010110",
  14790=>"111111010",
  14791=>"100010000",
  14792=>"000011010",
  14793=>"101001110",
  14794=>"001000001",
  14795=>"010011001",
  14796=>"010010010",
  14797=>"110100111",
  14798=>"111101001",
  14799=>"010111001",
  14800=>"001100110",
  14801=>"010111100",
  14802=>"111010000",
  14803=>"011101001",
  14804=>"111101000",
  14805=>"001010000",
  14806=>"111101011",
  14807=>"000110111",
  14808=>"011110111",
  14809=>"100011110",
  14810=>"011010011",
  14811=>"101110100",
  14812=>"111110111",
  14813=>"111101111",
  14814=>"100111011",
  14815=>"111101110",
  14816=>"110101100",
  14817=>"011100000",
  14818=>"111000001",
  14819=>"011010011",
  14820=>"101101110",
  14821=>"100010100",
  14822=>"111111100",
  14823=>"110100001",
  14824=>"111111111",
  14825=>"011101101",
  14826=>"011100011",
  14827=>"111111010",
  14828=>"000100000",
  14829=>"001111010",
  14830=>"111011010",
  14831=>"110011100",
  14832=>"101011000",
  14833=>"011010100",
  14834=>"110001010",
  14835=>"100111100",
  14836=>"001001011",
  14837=>"010101010",
  14838=>"101001101",
  14839=>"111000111",
  14840=>"111100100",
  14841=>"101100100",
  14842=>"101110101",
  14843=>"110111000",
  14844=>"001101000",
  14845=>"011110001",
  14846=>"110110101",
  14847=>"110111001",
  14848=>"011011000",
  14849=>"000001010",
  14850=>"000001111",
  14851=>"001100111",
  14852=>"010111001",
  14853=>"011110011",
  14854=>"100001001",
  14855=>"111101111",
  14856=>"101101110",
  14857=>"010011101",
  14858=>"101011011",
  14859=>"111011010",
  14860=>"101010101",
  14861=>"011000110",
  14862=>"011000010",
  14863=>"010011001",
  14864=>"011001010",
  14865=>"111000101",
  14866=>"111101001",
  14867=>"001111000",
  14868=>"011001001",
  14869=>"010000000",
  14870=>"011111001",
  14871=>"011000110",
  14872=>"010000100",
  14873=>"011010001",
  14874=>"011110100",
  14875=>"011000111",
  14876=>"110000110",
  14877=>"010010010",
  14878=>"001110101",
  14879=>"111001011",
  14880=>"010010110",
  14881=>"100110011",
  14882=>"110010111",
  14883=>"101010110",
  14884=>"011100111",
  14885=>"111000001",
  14886=>"101110111",
  14887=>"010000010",
  14888=>"011011101",
  14889=>"101110101",
  14890=>"111111111",
  14891=>"110000111",
  14892=>"100001011",
  14893=>"011110011",
  14894=>"100100001",
  14895=>"000010010",
  14896=>"010101110",
  14897=>"111100001",
  14898=>"101011001",
  14899=>"000100100",
  14900=>"110010001",
  14901=>"000110111",
  14902=>"001100111",
  14903=>"111111111",
  14904=>"111000100",
  14905=>"000010010",
  14906=>"111010000",
  14907=>"011001011",
  14908=>"110110000",
  14909=>"000000100",
  14910=>"010110101",
  14911=>"011000000",
  14912=>"111011011",
  14913=>"111000011",
  14914=>"101010111",
  14915=>"111110001",
  14916=>"111011111",
  14917=>"111101000",
  14918=>"101011001",
  14919=>"000010000",
  14920=>"110111011",
  14921=>"010010000",
  14922=>"011011111",
  14923=>"101111110",
  14924=>"101111111",
  14925=>"000000110",
  14926=>"100010011",
  14927=>"101001001",
  14928=>"110001011",
  14929=>"001001001",
  14930=>"111000101",
  14931=>"110110110",
  14932=>"101111011",
  14933=>"100001010",
  14934=>"001000110",
  14935=>"010100010",
  14936=>"011111010",
  14937=>"101001001",
  14938=>"101010000",
  14939=>"100100101",
  14940=>"001101010",
  14941=>"001000110",
  14942=>"100001101",
  14943=>"011011001",
  14944=>"011110011",
  14945=>"110100011",
  14946=>"111011010",
  14947=>"100101011",
  14948=>"101110011",
  14949=>"111010000",
  14950=>"101100010",
  14951=>"110100001",
  14952=>"100100000",
  14953=>"110111110",
  14954=>"111111000",
  14955=>"110000100",
  14956=>"001100010",
  14957=>"101000111",
  14958=>"111100110",
  14959=>"010101011",
  14960=>"111111110",
  14961=>"111110001",
  14962=>"100101011",
  14963=>"011111010",
  14964=>"001001110",
  14965=>"010111011",
  14966=>"111111001",
  14967=>"100100100",
  14968=>"000000001",
  14969=>"110110001",
  14970=>"111100101",
  14971=>"111100110",
  14972=>"001100011",
  14973=>"000101101",
  14974=>"001001011",
  14975=>"010010010",
  14976=>"000000001",
  14977=>"101100100",
  14978=>"100110110",
  14979=>"100000011",
  14980=>"111011111",
  14981=>"001000000",
  14982=>"100111100",
  14983=>"001000100",
  14984=>"111001001",
  14985=>"111000001",
  14986=>"011000110",
  14987=>"110100110",
  14988=>"001110110",
  14989=>"111100101",
  14990=>"001010100",
  14991=>"000111010",
  14992=>"100000110",
  14993=>"011111010",
  14994=>"010011010",
  14995=>"011110100",
  14996=>"110110010",
  14997=>"010101101",
  14998=>"111110101",
  14999=>"011001000",
  15000=>"100011000",
  15001=>"000110010",
  15002=>"111010101",
  15003=>"011010111",
  15004=>"011110010",
  15005=>"101111001",
  15006=>"001011110",
  15007=>"101111001",
  15008=>"110100000",
  15009=>"111100100",
  15010=>"111110010",
  15011=>"011101000",
  15012=>"001010011",
  15013=>"110111101",
  15014=>"100100101",
  15015=>"011000000",
  15016=>"010101000",
  15017=>"011011111",
  15018=>"111001011",
  15019=>"000010101",
  15020=>"011111001",
  15021=>"011110000",
  15022=>"010001100",
  15023=>"011110100",
  15024=>"110110001",
  15025=>"011110100",
  15026=>"111101011",
  15027=>"010011111",
  15028=>"101101111",
  15029=>"011111111",
  15030=>"000010100",
  15031=>"111011100",
  15032=>"000101100",
  15033=>"011110000",
  15034=>"100010111",
  15035=>"010100001",
  15036=>"010011111",
  15037=>"010000010",
  15038=>"010000000",
  15039=>"101111100",
  15040=>"111001101",
  15041=>"000000110",
  15042=>"111010000",
  15043=>"010110100",
  15044=>"010110110",
  15045=>"000000011",
  15046=>"011001100",
  15047=>"110010111",
  15048=>"000010000",
  15049=>"100111110",
  15050=>"000100011",
  15051=>"101011111",
  15052=>"100000000",
  15053=>"011010111",
  15054=>"111101001",
  15055=>"011100111",
  15056=>"010101000",
  15057=>"010011110",
  15058=>"101100101",
  15059=>"100000010",
  15060=>"101011010",
  15061=>"111000110",
  15062=>"100010110",
  15063=>"000100001",
  15064=>"101100101",
  15065=>"110001100",
  15066=>"101001011",
  15067=>"011010010",
  15068=>"000100001",
  15069=>"010100100",
  15070=>"110000001",
  15071=>"110101101",
  15072=>"000111001",
  15073=>"000110000",
  15074=>"010111101",
  15075=>"011001011",
  15076=>"100100100",
  15077=>"000100001",
  15078=>"100110100",
  15079=>"000100101",
  15080=>"110001100",
  15081=>"100101010",
  15082=>"010001011",
  15083=>"101111100",
  15084=>"000000111",
  15085=>"010000100",
  15086=>"001010000",
  15087=>"100010001",
  15088=>"101110010",
  15089=>"011011001",
  15090=>"100100100",
  15091=>"010000101",
  15092=>"001100110",
  15093=>"000011111",
  15094=>"111010011",
  15095=>"111011000",
  15096=>"100010000",
  15097=>"011111111",
  15098=>"100110000",
  15099=>"001111010",
  15100=>"101010001",
  15101=>"110000000",
  15102=>"010001001",
  15103=>"111110010",
  15104=>"001000110",
  15105=>"011110000",
  15106=>"111110110",
  15107=>"101010010",
  15108=>"100000110",
  15109=>"101000101",
  15110=>"001011010",
  15111=>"011010110",
  15112=>"100111101",
  15113=>"100000100",
  15114=>"001111111",
  15115=>"110011111",
  15116=>"001001111",
  15117=>"110101010",
  15118=>"100001100",
  15119=>"000111011",
  15120=>"010001001",
  15121=>"111011001",
  15122=>"010101110",
  15123=>"101101100",
  15124=>"110111011",
  15125=>"000000010",
  15126=>"000000111",
  15127=>"010010101",
  15128=>"110011110",
  15129=>"010110100",
  15130=>"010111000",
  15131=>"001100011",
  15132=>"001110001",
  15133=>"001100100",
  15134=>"000101001",
  15135=>"010001001",
  15136=>"001011100",
  15137=>"010000110",
  15138=>"111010000",
  15139=>"010100101",
  15140=>"001101111",
  15141=>"001000010",
  15142=>"100000101",
  15143=>"010111100",
  15144=>"001001010",
  15145=>"100010110",
  15146=>"001101000",
  15147=>"110101111",
  15148=>"100110100",
  15149=>"100000010",
  15150=>"111110001",
  15151=>"101010100",
  15152=>"100000110",
  15153=>"110010101",
  15154=>"010000000",
  15155=>"101000100",
  15156=>"101101010",
  15157=>"001110111",
  15158=>"000111000",
  15159=>"110110111",
  15160=>"011111110",
  15161=>"011011000",
  15162=>"111111101",
  15163=>"010101001",
  15164=>"110100011",
  15165=>"100011100",
  15166=>"101111111",
  15167=>"110011000",
  15168=>"110110010",
  15169=>"010000111",
  15170=>"010000011",
  15171=>"100001011",
  15172=>"101100110",
  15173=>"111000101",
  15174=>"000100010",
  15175=>"111101010",
  15176=>"011101111",
  15177=>"101000001",
  15178=>"000101010",
  15179=>"111101101",
  15180=>"000100001",
  15181=>"111100100",
  15182=>"110100100",
  15183=>"000001000",
  15184=>"011000011",
  15185=>"000101110",
  15186=>"001011010",
  15187=>"011000110",
  15188=>"010101111",
  15189=>"111110001",
  15190=>"010110110",
  15191=>"001011101",
  15192=>"001000100",
  15193=>"101000010",
  15194=>"111110001",
  15195=>"000100011",
  15196=>"101000011",
  15197=>"111111101",
  15198=>"111110001",
  15199=>"010011001",
  15200=>"011110001",
  15201=>"101001100",
  15202=>"101111010",
  15203=>"111101010",
  15204=>"101000000",
  15205=>"000001010",
  15206=>"111111001",
  15207=>"111011010",
  15208=>"000110110",
  15209=>"111101010",
  15210=>"110010010",
  15211=>"000000011",
  15212=>"110101100",
  15213=>"101110010",
  15214=>"010110111",
  15215=>"000011110",
  15216=>"001101011",
  15217=>"110011010",
  15218=>"000110111",
  15219=>"110111001",
  15220=>"111110110",
  15221=>"111001001",
  15222=>"011100000",
  15223=>"001010100",
  15224=>"011001011",
  15225=>"111111110",
  15226=>"110000100",
  15227=>"001100111",
  15228=>"011010110",
  15229=>"011010110",
  15230=>"011111011",
  15231=>"100011011",
  15232=>"111100011",
  15233=>"111101111",
  15234=>"011111000",
  15235=>"101010101",
  15236=>"000011100",
  15237=>"111111001",
  15238=>"011011000",
  15239=>"101101010",
  15240=>"011001011",
  15241=>"010111010",
  15242=>"111111110",
  15243=>"100000011",
  15244=>"011111100",
  15245=>"100010000",
  15246=>"000010000",
  15247=>"011111000",
  15248=>"011011011",
  15249=>"111111001",
  15250=>"011110111",
  15251=>"000000110",
  15252=>"101111111",
  15253=>"010000001",
  15254=>"111010101",
  15255=>"100000111",
  15256=>"001000011",
  15257=>"001000010",
  15258=>"101110110",
  15259=>"011011100",
  15260=>"011010100",
  15261=>"001101011",
  15262=>"011100000",
  15263=>"001000001",
  15264=>"001100100",
  15265=>"000011101",
  15266=>"010010101",
  15267=>"111111100",
  15268=>"110000000",
  15269=>"000000001",
  15270=>"011010111",
  15271=>"010001100",
  15272=>"111011110",
  15273=>"010000010",
  15274=>"010010000",
  15275=>"110111010",
  15276=>"100111111",
  15277=>"000001001",
  15278=>"100100101",
  15279=>"001001100",
  15280=>"010100001",
  15281=>"011111000",
  15282=>"010001110",
  15283=>"100010111",
  15284=>"011011110",
  15285=>"011001101",
  15286=>"100110011",
  15287=>"001110110",
  15288=>"100100000",
  15289=>"101111110",
  15290=>"110101000",
  15291=>"101011000",
  15292=>"010110101",
  15293=>"011101101",
  15294=>"011011100",
  15295=>"011101001",
  15296=>"101110001",
  15297=>"111000001",
  15298=>"010100101",
  15299=>"110000111",
  15300=>"011111101",
  15301=>"000011010",
  15302=>"000111100",
  15303=>"011111000",
  15304=>"000001111",
  15305=>"110101000",
  15306=>"011100010",
  15307=>"001110011",
  15308=>"011110001",
  15309=>"101110000",
  15310=>"010110110",
  15311=>"111111011",
  15312=>"010010100",
  15313=>"001100010",
  15314=>"000110100",
  15315=>"010001000",
  15316=>"101000110",
  15317=>"010010000",
  15318=>"000111110",
  15319=>"100111011",
  15320=>"110010100",
  15321=>"100011001",
  15322=>"001000000",
  15323=>"111011110",
  15324=>"010001111",
  15325=>"111010010",
  15326=>"000110001",
  15327=>"010100000",
  15328=>"101010010",
  15329=>"011101111",
  15330=>"101111001",
  15331=>"000110110",
  15332=>"111100100",
  15333=>"000001010",
  15334=>"000010010",
  15335=>"101001101",
  15336=>"010100010",
  15337=>"101001001",
  15338=>"110101111",
  15339=>"001011111",
  15340=>"110111111",
  15341=>"000000010",
  15342=>"010100010",
  15343=>"101111000",
  15344=>"010001111",
  15345=>"011101011",
  15346=>"000000010",
  15347=>"100000111",
  15348=>"110100000",
  15349=>"101110000",
  15350=>"000111100",
  15351=>"111101110",
  15352=>"000010010",
  15353=>"000000001",
  15354=>"111010100",
  15355=>"101101101",
  15356=>"010011101",
  15357=>"101100101",
  15358=>"000100011",
  15359=>"000010000",
  15360=>"000001010",
  15361=>"101110100",
  15362=>"011111110",
  15363=>"000111011",
  15364=>"001010001",
  15365=>"001000011",
  15366=>"111100011",
  15367=>"000101010",
  15368=>"010010001",
  15369=>"011011111",
  15370=>"100100010",
  15371=>"101111000",
  15372=>"101001000",
  15373=>"100000110",
  15374=>"110001000",
  15375=>"110011011",
  15376=>"000011000",
  15377=>"110011001",
  15378=>"111001110",
  15379=>"001001011",
  15380=>"110101101",
  15381=>"101000001",
  15382=>"100001111",
  15383=>"100011011",
  15384=>"000101110",
  15385=>"011101000",
  15386=>"101011110",
  15387=>"001110000",
  15388=>"001010111",
  15389=>"111010101",
  15390=>"101000001",
  15391=>"110111110",
  15392=>"111011011",
  15393=>"111010000",
  15394=>"111100101",
  15395=>"011011000",
  15396=>"111010110",
  15397=>"100011100",
  15398=>"000111000",
  15399=>"001011110",
  15400=>"010010101",
  15401=>"111100111",
  15402=>"001100011",
  15403=>"011010000",
  15404=>"110000110",
  15405=>"000110100",
  15406=>"101100100",
  15407=>"100110111",
  15408=>"010111111",
  15409=>"000100000",
  15410=>"011111100",
  15411=>"110111000",
  15412=>"010101010",
  15413=>"000100011",
  15414=>"000101110",
  15415=>"011001011",
  15416=>"101111000",
  15417=>"011100011",
  15418=>"110100000",
  15419=>"100000010",
  15420=>"111000100",
  15421=>"000100111",
  15422=>"011100110",
  15423=>"000011100",
  15424=>"000100110",
  15425=>"110101110",
  15426=>"101111111",
  15427=>"110010010",
  15428=>"100011001",
  15429=>"001111010",
  15430=>"111010110",
  15431=>"011111101",
  15432=>"110110000",
  15433=>"011111000",
  15434=>"001011100",
  15435=>"100010100",
  15436=>"110111100",
  15437=>"011110011",
  15438=>"010010100",
  15439=>"111100001",
  15440=>"000101010",
  15441=>"000000011",
  15442=>"010001100",
  15443=>"011011100",
  15444=>"011100001",
  15445=>"100101100",
  15446=>"001100010",
  15447=>"000010100",
  15448=>"111111011",
  15449=>"010100011",
  15450=>"100000111",
  15451=>"100101000",
  15452=>"000000000",
  15453=>"100001110",
  15454=>"001110100",
  15455=>"101011010",
  15456=>"101010001",
  15457=>"011010011",
  15458=>"011101001",
  15459=>"000101000",
  15460=>"011101111",
  15461=>"110111010",
  15462=>"110111111",
  15463=>"111001111",
  15464=>"110011101",
  15465=>"100100111",
  15466=>"011100100",
  15467=>"000110001",
  15468=>"001000001",
  15469=>"000011100",
  15470=>"011001101",
  15471=>"100010010",
  15472=>"100111000",
  15473=>"010000010",
  15474=>"101111100",
  15475=>"100010101",
  15476=>"110110000",
  15477=>"101101010",
  15478=>"000001010",
  15479=>"111100110",
  15480=>"101111010",
  15481=>"101000111",
  15482=>"000110100",
  15483=>"010111000",
  15484=>"010010011",
  15485=>"110100000",
  15486=>"010100111",
  15487=>"000001000",
  15488=>"110011000",
  15489=>"110101010",
  15490=>"011001110",
  15491=>"001101010",
  15492=>"101110010",
  15493=>"010000111",
  15494=>"100011010",
  15495=>"111011111",
  15496=>"110111000",
  15497=>"011000101",
  15498=>"011101001",
  15499=>"010110100",
  15500=>"110010101",
  15501=>"111100000",
  15502=>"011111011",
  15503=>"110111011",
  15504=>"000000100",
  15505=>"011111111",
  15506=>"010001000",
  15507=>"111010100",
  15508=>"001000000",
  15509=>"111001000",
  15510=>"010001101",
  15511=>"000110000",
  15512=>"111000110",
  15513=>"001000111",
  15514=>"100110000",
  15515=>"000111010",
  15516=>"110101110",
  15517=>"100000000",
  15518=>"000011100",
  15519=>"101010011",
  15520=>"000001110",
  15521=>"101100000",
  15522=>"000001101",
  15523=>"000000101",
  15524=>"101001000",
  15525=>"111100000",
  15526=>"110011000",
  15527=>"101110101",
  15528=>"000100010",
  15529=>"010001001",
  15530=>"011110000",
  15531=>"100011100",
  15532=>"110100010",
  15533=>"001111100",
  15534=>"111100111",
  15535=>"000010010",
  15536=>"001100111",
  15537=>"000101110",
  15538=>"110100100",
  15539=>"101010000",
  15540=>"100010000",
  15541=>"000111110",
  15542=>"111000111",
  15543=>"011001000",
  15544=>"110001011",
  15545=>"110101001",
  15546=>"010001010",
  15547=>"001010110",
  15548=>"010111000",
  15549=>"001000001",
  15550=>"010001000",
  15551=>"000110011",
  15552=>"111010100",
  15553=>"011111001",
  15554=>"000010111",
  15555=>"110110011",
  15556=>"000111011",
  15557=>"010101100",
  15558=>"001111001",
  15559=>"101110101",
  15560=>"010100010",
  15561=>"111111011",
  15562=>"001010100",
  15563=>"101001001",
  15564=>"100110110",
  15565=>"100011010",
  15566=>"101111101",
  15567=>"010111100",
  15568=>"011000011",
  15569=>"100110110",
  15570=>"000000011",
  15571=>"011011110",
  15572=>"101011111",
  15573=>"101011110",
  15574=>"100101010",
  15575=>"000000010",
  15576=>"001000001",
  15577=>"010111110",
  15578=>"000101110",
  15579=>"000001101",
  15580=>"111101011",
  15581=>"000001111",
  15582=>"111111011",
  15583=>"110110111",
  15584=>"010010000",
  15585=>"010000001",
  15586=>"011000100",
  15587=>"100010001",
  15588=>"011101001",
  15589=>"011000101",
  15590=>"011110010",
  15591=>"001000101",
  15592=>"110010000",
  15593=>"011001011",
  15594=>"010100001",
  15595=>"001110000",
  15596=>"000010010",
  15597=>"110001001",
  15598=>"110010110",
  15599=>"010011000",
  15600=>"000010010",
  15601=>"000010011",
  15602=>"111111011",
  15603=>"111001011",
  15604=>"010101010",
  15605=>"000001000",
  15606=>"011111001",
  15607=>"000000000",
  15608=>"010000001",
  15609=>"011010111",
  15610=>"001110111",
  15611=>"000001010",
  15612=>"000001101",
  15613=>"111111111",
  15614=>"001001001",
  15615=>"000010101",
  15616=>"010010000",
  15617=>"001110010",
  15618=>"110100001",
  15619=>"101011110",
  15620=>"010011010",
  15621=>"011111001",
  15622=>"010010011",
  15623=>"111111001",
  15624=>"101110000",
  15625=>"011000001",
  15626=>"101110110",
  15627=>"011011101",
  15628=>"110111111",
  15629=>"100110000",
  15630=>"101010101",
  15631=>"101011100",
  15632=>"110110110",
  15633=>"100000000",
  15634=>"100011000",
  15635=>"101011001",
  15636=>"101001001",
  15637=>"110101001",
  15638=>"111010011",
  15639=>"000100011",
  15640=>"011010101",
  15641=>"001100000",
  15642=>"110011111",
  15643=>"001101011",
  15644=>"000001000",
  15645=>"011100000",
  15646=>"111111000",
  15647=>"110111000",
  15648=>"100100101",
  15649=>"111011101",
  15650=>"110111001",
  15651=>"001000000",
  15652=>"111110111",
  15653=>"001100110",
  15654=>"110001001",
  15655=>"011111100",
  15656=>"110111111",
  15657=>"011001101",
  15658=>"110011101",
  15659=>"001010100",
  15660=>"111110101",
  15661=>"111110110",
  15662=>"001101111",
  15663=>"000011001",
  15664=>"100000111",
  15665=>"111111111",
  15666=>"010110100",
  15667=>"000010010",
  15668=>"111011100",
  15669=>"010011110",
  15670=>"000001011",
  15671=>"000111101",
  15672=>"110000010",
  15673=>"001100000",
  15674=>"111001010",
  15675=>"011000111",
  15676=>"101011010",
  15677=>"001011001",
  15678=>"011101001",
  15679=>"111011110",
  15680=>"100010110",
  15681=>"111010000",
  15682=>"011001010",
  15683=>"111111111",
  15684=>"000001100",
  15685=>"000111110",
  15686=>"100011010",
  15687=>"001100110",
  15688=>"111100101",
  15689=>"000111101",
  15690=>"100111101",
  15691=>"001010001",
  15692=>"000010101",
  15693=>"000011010",
  15694=>"100100111",
  15695=>"011001000",
  15696=>"011001000",
  15697=>"101000000",
  15698=>"010000100",
  15699=>"111011111",
  15700=>"100101100",
  15701=>"100010010",
  15702=>"011110111",
  15703=>"000111011",
  15704=>"111100011",
  15705=>"011111010",
  15706=>"001000100",
  15707=>"001010011",
  15708=>"000010100",
  15709=>"111101111",
  15710=>"011101011",
  15711=>"111100001",
  15712=>"000010011",
  15713=>"011010101",
  15714=>"010010000",
  15715=>"111100010",
  15716=>"101011110",
  15717=>"111010111",
  15718=>"000100100",
  15719=>"000010010",
  15720=>"111011110",
  15721=>"001110011",
  15722=>"000101110",
  15723=>"010011010",
  15724=>"110111010",
  15725=>"111000011",
  15726=>"010011000",
  15727=>"000111111",
  15728=>"100010010",
  15729=>"000101001",
  15730=>"110010100",
  15731=>"101010101",
  15732=>"101011110",
  15733=>"100000011",
  15734=>"110010010",
  15735=>"001001101",
  15736=>"110101001",
  15737=>"010111010",
  15738=>"001101011",
  15739=>"100111000",
  15740=>"111111111",
  15741=>"100010110",
  15742=>"111110111",
  15743=>"000001000",
  15744=>"000101101",
  15745=>"111001010",
  15746=>"111000010",
  15747=>"111110000",
  15748=>"001001010",
  15749=>"000111001",
  15750=>"000001001",
  15751=>"111010011",
  15752=>"000011100",
  15753=>"101101000",
  15754=>"110101001",
  15755=>"001110000",
  15756=>"100000111",
  15757=>"011110000",
  15758=>"110101000",
  15759=>"101100010",
  15760=>"101011110",
  15761=>"011000101",
  15762=>"111100101",
  15763=>"100100110",
  15764=>"011111010",
  15765=>"100110010",
  15766=>"101000000",
  15767=>"110001111",
  15768=>"110110000",
  15769=>"011100011",
  15770=>"111011011",
  15771=>"111000010",
  15772=>"110010001",
  15773=>"010100001",
  15774=>"001000100",
  15775=>"000101001",
  15776=>"000110011",
  15777=>"101000010",
  15778=>"010110101",
  15779=>"100010110",
  15780=>"111000111",
  15781=>"000101101",
  15782=>"000001010",
  15783=>"101111010",
  15784=>"110010101",
  15785=>"000011111",
  15786=>"010000011",
  15787=>"101010001",
  15788=>"110000010",
  15789=>"001100010",
  15790=>"111111011",
  15791=>"111100111",
  15792=>"111001111",
  15793=>"011111011",
  15794=>"101010101",
  15795=>"001100111",
  15796=>"010010111",
  15797=>"110111111",
  15798=>"000000101",
  15799=>"110100001",
  15800=>"001100001",
  15801=>"010011010",
  15802=>"000110001",
  15803=>"000010011",
  15804=>"101011100",
  15805=>"110101010",
  15806=>"000001001",
  15807=>"100010000",
  15808=>"000010011",
  15809=>"111101000",
  15810=>"011111000",
  15811=>"101101001",
  15812=>"100111010",
  15813=>"101111000",
  15814=>"100011001",
  15815=>"111101111",
  15816=>"111101010",
  15817=>"110100010",
  15818=>"010111101",
  15819=>"010001101",
  15820=>"110100001",
  15821=>"000010101",
  15822=>"001001111",
  15823=>"001110011",
  15824=>"001010101",
  15825=>"100011001",
  15826=>"111101101",
  15827=>"000101110",
  15828=>"101011101",
  15829=>"011010101",
  15830=>"101000101",
  15831=>"011110001",
  15832=>"000111000",
  15833=>"011001010",
  15834=>"111000010",
  15835=>"000001111",
  15836=>"011111111",
  15837=>"101110100",
  15838=>"000010011",
  15839=>"101000000",
  15840=>"111011101",
  15841=>"001010101",
  15842=>"000101101",
  15843=>"101110100",
  15844=>"101101010",
  15845=>"011011011",
  15846=>"100101001",
  15847=>"101110000",
  15848=>"101010110",
  15849=>"111110100",
  15850=>"000101101",
  15851=>"100100111",
  15852=>"011000111",
  15853=>"101000101",
  15854=>"001000011",
  15855=>"110001001",
  15856=>"100101010",
  15857=>"101011010",
  15858=>"000110111",
  15859=>"100011110",
  15860=>"001010101",
  15861=>"101111100",
  15862=>"001011100",
  15863=>"111001010",
  15864=>"000011110",
  15865=>"011011010",
  15866=>"100010101",
  15867=>"000110010",
  15868=>"111010111",
  15869=>"001010101",
  15870=>"110101100",
  15871=>"001100010",
  15872=>"111111101",
  15873=>"101101110",
  15874=>"010101101",
  15875=>"110101111",
  15876=>"101111110",
  15877=>"000111100",
  15878=>"010011011",
  15879=>"111111100",
  15880=>"101110101",
  15881=>"110000100",
  15882=>"000001110",
  15883=>"001101110",
  15884=>"100100001",
  15885=>"101111110",
  15886=>"110011111",
  15887=>"100001101",
  15888=>"101110010",
  15889=>"100001001",
  15890=>"100011010",
  15891=>"000000100",
  15892=>"001000000",
  15893=>"001101000",
  15894=>"000011011",
  15895=>"101111101",
  15896=>"100010111",
  15897=>"000101010",
  15898=>"011110000",
  15899=>"100111101",
  15900=>"100010011",
  15901=>"111011100",
  15902=>"001001111",
  15903=>"111010110",
  15904=>"111111010",
  15905=>"110111101",
  15906=>"101010101",
  15907=>"101110100",
  15908=>"001010110",
  15909=>"101011111",
  15910=>"110000100",
  15911=>"000011000",
  15912=>"000101010",
  15913=>"000000010",
  15914=>"110100000",
  15915=>"100011111",
  15916=>"100011010",
  15917=>"100100000",
  15918=>"101100110",
  15919=>"111001101",
  15920=>"110001001",
  15921=>"111100100",
  15922=>"111000110",
  15923=>"111000101",
  15924=>"110001010",
  15925=>"011010011",
  15926=>"000101001",
  15927=>"111111111",
  15928=>"111110000",
  15929=>"101110000",
  15930=>"101101101",
  15931=>"000100001",
  15932=>"000110111",
  15933=>"010010001",
  15934=>"000000011",
  15935=>"101100111",
  15936=>"011000000",
  15937=>"110011101",
  15938=>"011101110",
  15939=>"111110001",
  15940=>"001111001",
  15941=>"111110011",
  15942=>"000001001",
  15943=>"101010010",
  15944=>"010111101",
  15945=>"110001100",
  15946=>"110101111",
  15947=>"110110111",
  15948=>"100100010",
  15949=>"010000110",
  15950=>"001111110",
  15951=>"111100100",
  15952=>"100001111",
  15953=>"101000100",
  15954=>"111110111",
  15955=>"011110110",
  15956=>"000000001",
  15957=>"101110111",
  15958=>"100101111",
  15959=>"101010000",
  15960=>"000110000",
  15961=>"001111110",
  15962=>"100110110",
  15963=>"000001110",
  15964=>"001001111",
  15965=>"111101100",
  15966=>"000001110",
  15967=>"001110110",
  15968=>"100101010",
  15969=>"110010000",
  15970=>"100110000",
  15971=>"101110011",
  15972=>"010011001",
  15973=>"010100111",
  15974=>"011011111",
  15975=>"101100001",
  15976=>"010111000",
  15977=>"101100100",
  15978=>"000010111",
  15979=>"111000000",
  15980=>"001011000",
  15981=>"010101011",
  15982=>"110100010",
  15983=>"100001110",
  15984=>"000010011",
  15985=>"111000100",
  15986=>"101000111",
  15987=>"001111000",
  15988=>"110100111",
  15989=>"011001010",
  15990=>"011111001",
  15991=>"010110101",
  15992=>"100001000",
  15993=>"111110111",
  15994=>"000001011",
  15995=>"111000110",
  15996=>"001010010",
  15997=>"001011000",
  15998=>"011100100",
  15999=>"110000010",
  16000=>"010101001",
  16001=>"011110010",
  16002=>"100000101",
  16003=>"011101101",
  16004=>"110001011",
  16005=>"001100011",
  16006=>"100111001",
  16007=>"000110001",
  16008=>"010110110",
  16009=>"111010100",
  16010=>"110101011",
  16011=>"000101000",
  16012=>"010001010",
  16013=>"110101010",
  16014=>"010100100",
  16015=>"111011000",
  16016=>"110011011",
  16017=>"001100101",
  16018=>"101010101",
  16019=>"000100111",
  16020=>"000010101",
  16021=>"011101001",
  16022=>"000111100",
  16023=>"011100011",
  16024=>"101100011",
  16025=>"010100100",
  16026=>"100100111",
  16027=>"100100011",
  16028=>"001111011",
  16029=>"011101111",
  16030=>"111100010",
  16031=>"001000100",
  16032=>"001110111",
  16033=>"001010010",
  16034=>"010101101",
  16035=>"111100100",
  16036=>"011100110",
  16037=>"101000010",
  16038=>"101111111",
  16039=>"101010110",
  16040=>"000000001",
  16041=>"010111101",
  16042=>"011111010",
  16043=>"111010000",
  16044=>"111000000",
  16045=>"011010001",
  16046=>"111100100",
  16047=>"001010001",
  16048=>"110010111",
  16049=>"011011011",
  16050=>"111010100",
  16051=>"001100001",
  16052=>"011000000",
  16053=>"110011011",
  16054=>"011001110",
  16055=>"100110110",
  16056=>"010110011",
  16057=>"011101010",
  16058=>"111110111",
  16059=>"011001110",
  16060=>"101101110",
  16061=>"101111101",
  16062=>"110111001",
  16063=>"001001011",
  16064=>"011001000",
  16065=>"111110110",
  16066=>"101001101",
  16067=>"010010101",
  16068=>"101111110",
  16069=>"111001100",
  16070=>"111000110",
  16071=>"100000000",
  16072=>"101000100",
  16073=>"100110011",
  16074=>"100000010",
  16075=>"100000000",
  16076=>"111010010",
  16077=>"110011010",
  16078=>"100000110",
  16079=>"010000001",
  16080=>"111110111",
  16081=>"001001010",
  16082=>"101110010",
  16083=>"001000011",
  16084=>"110101011",
  16085=>"101011111",
  16086=>"100001111",
  16087=>"011101011",
  16088=>"101101011",
  16089=>"101001110",
  16090=>"111011011",
  16091=>"101110010",
  16092=>"010111100",
  16093=>"010001110",
  16094=>"000000110",
  16095=>"001101100",
  16096=>"100010010",
  16097=>"110010100",
  16098=>"110100110",
  16099=>"011101000",
  16100=>"110101111",
  16101=>"011001001",
  16102=>"010101011",
  16103=>"000101110",
  16104=>"110111101",
  16105=>"011101001",
  16106=>"101111001",
  16107=>"111010100",
  16108=>"110111101",
  16109=>"000100001",
  16110=>"010011011",
  16111=>"101100100",
  16112=>"100100100",
  16113=>"011001011",
  16114=>"011101010",
  16115=>"111110000",
  16116=>"111010110",
  16117=>"001001010",
  16118=>"100101100",
  16119=>"101000100",
  16120=>"101011011",
  16121=>"110110111",
  16122=>"100001101",
  16123=>"000100011",
  16124=>"110010011",
  16125=>"111011110",
  16126=>"110101111",
  16127=>"010000101",
  16128=>"110000011",
  16129=>"111110000",
  16130=>"010111001",
  16131=>"111111110",
  16132=>"110101000",
  16133=>"010110011",
  16134=>"111101000",
  16135=>"111100011",
  16136=>"111000001",
  16137=>"111010010",
  16138=>"100010011",
  16139=>"111011111",
  16140=>"011000001",
  16141=>"100101010",
  16142=>"100011110",
  16143=>"011001000",
  16144=>"011000100",
  16145=>"101111010",
  16146=>"110011000",
  16147=>"000010110",
  16148=>"111101110",
  16149=>"010011001",
  16150=>"001000101",
  16151=>"101100011",
  16152=>"110010000",
  16153=>"110011001",
  16154=>"001110000",
  16155=>"100001111",
  16156=>"101000010",
  16157=>"100001000",
  16158=>"011111110",
  16159=>"001110111",
  16160=>"111111011",
  16161=>"100000101",
  16162=>"111110111",
  16163=>"100010011",
  16164=>"101101100",
  16165=>"001110110",
  16166=>"011100000",
  16167=>"001000010",
  16168=>"011111010",
  16169=>"000000000",
  16170=>"100111101",
  16171=>"010110001",
  16172=>"010100010",
  16173=>"101110101",
  16174=>"010101001",
  16175=>"000011101",
  16176=>"101011101",
  16177=>"011011010",
  16178=>"010010100",
  16179=>"010010110",
  16180=>"011111111",
  16181=>"100101111",
  16182=>"001011000",
  16183=>"010001001",
  16184=>"101011100",
  16185=>"111100100",
  16186=>"000010100",
  16187=>"011011110",
  16188=>"011000010",
  16189=>"111010000",
  16190=>"100001110",
  16191=>"000011110",
  16192=>"001100100",
  16193=>"111101000",
  16194=>"001000101",
  16195=>"111111110",
  16196=>"100010100",
  16197=>"110010000",
  16198=>"000111000",
  16199=>"001011101",
  16200=>"101011111",
  16201=>"100001001",
  16202=>"110100110",
  16203=>"000000010",
  16204=>"101010100",
  16205=>"000110110",
  16206=>"100101001",
  16207=>"001011001",
  16208=>"001000101",
  16209=>"001110110",
  16210=>"010100100",
  16211=>"111101010",
  16212=>"010010100",
  16213=>"110010010",
  16214=>"001010001",
  16215=>"010010011",
  16216=>"110111010",
  16217=>"000011001",
  16218=>"111010110",
  16219=>"100011110",
  16220=>"000100001",
  16221=>"110000111",
  16222=>"001001011",
  16223=>"111111001",
  16224=>"110101100",
  16225=>"001010100",
  16226=>"111010001",
  16227=>"110101000",
  16228=>"010011000",
  16229=>"011010000",
  16230=>"110001100",
  16231=>"100100010",
  16232=>"110010101",
  16233=>"011000001",
  16234=>"001011100",
  16235=>"101000000",
  16236=>"000000000",
  16237=>"011011101",
  16238=>"101100101",
  16239=>"001110011",
  16240=>"000111001",
  16241=>"000110110",
  16242=>"000111100",
  16243=>"110110111",
  16244=>"110000011",
  16245=>"011110101",
  16246=>"000100111",
  16247=>"100010000",
  16248=>"010011010",
  16249=>"110010100",
  16250=>"110111010",
  16251=>"011101111",
  16252=>"111001001",
  16253=>"001110101",
  16254=>"000010111",
  16255=>"110111001",
  16256=>"000100111",
  16257=>"010011111",
  16258=>"110001001",
  16259=>"011001010",
  16260=>"010011110",
  16261=>"110010111",
  16262=>"000011101",
  16263=>"101100100",
  16264=>"100011010",
  16265=>"110011011",
  16266=>"111100000",
  16267=>"101011111",
  16268=>"111101011",
  16269=>"111001011",
  16270=>"000010101",
  16271=>"001011111",
  16272=>"110001001",
  16273=>"100100110",
  16274=>"010001100",
  16275=>"011101100",
  16276=>"111001001",
  16277=>"100101000",
  16278=>"100100100",
  16279=>"000001100",
  16280=>"010001001",
  16281=>"111101111",
  16282=>"111100000",
  16283=>"011111011",
  16284=>"010001001",
  16285=>"011110011",
  16286=>"001101010",
  16287=>"110101101",
  16288=>"010110000",
  16289=>"100001010",
  16290=>"001111010",
  16291=>"011000100",
  16292=>"011000110",
  16293=>"111110100",
  16294=>"101111101",
  16295=>"000101001",
  16296=>"100110101",
  16297=>"100110100",
  16298=>"110101111",
  16299=>"000010110",
  16300=>"001001101",
  16301=>"001001110",
  16302=>"101011011",
  16303=>"000111000",
  16304=>"001110100",
  16305=>"111100000",
  16306=>"000010000",
  16307=>"010101110",
  16308=>"110000000",
  16309=>"010000100",
  16310=>"111100010",
  16311=>"100000101",
  16312=>"100010000",
  16313=>"011010000",
  16314=>"000100011",
  16315=>"000101100",
  16316=>"110000001",
  16317=>"011111111",
  16318=>"000011000",
  16319=>"011011101",
  16320=>"100111000",
  16321=>"100100011",
  16322=>"010111001",
  16323=>"100001110",
  16324=>"001101110",
  16325=>"001101111",
  16326=>"100110000",
  16327=>"110110101",
  16328=>"100000001",
  16329=>"111110100",
  16330=>"101000100",
  16331=>"011111010",
  16332=>"110110001",
  16333=>"100001011",
  16334=>"100111000",
  16335=>"010110110",
  16336=>"111101011",
  16337=>"111101101",
  16338=>"110000011",
  16339=>"110100001",
  16340=>"000000010",
  16341=>"111000001",
  16342=>"010001100",
  16343=>"110011111",
  16344=>"000010010",
  16345=>"101110111",
  16346=>"101100000",
  16347=>"000101011",
  16348=>"000011100",
  16349=>"001110111",
  16350=>"001101110",
  16351=>"001001111",
  16352=>"010110010",
  16353=>"110010001",
  16354=>"000011111",
  16355=>"111101111",
  16356=>"100001001",
  16357=>"110111010",
  16358=>"110101111",
  16359=>"010111111",
  16360=>"110001000",
  16361=>"111011000",
  16362=>"101001111",
  16363=>"011000001",
  16364=>"001001000",
  16365=>"001101101",
  16366=>"100001001",
  16367=>"111101101",
  16368=>"001010100",
  16369=>"001111001",
  16370=>"010000000",
  16371=>"011110111",
  16372=>"100110110",
  16373=>"010111011",
  16374=>"000101000",
  16375=>"011000011",
  16376=>"100100001",
  16377=>"111111000",
  16378=>"100010010",
  16379=>"010001010",
  16380=>"111110011",
  16381=>"110001111",
  16382=>"110010000",
  16383=>"000000110",
  16384=>"111110111",
  16385=>"110010111",
  16386=>"010111011",
  16387=>"000000011",
  16388=>"111110000",
  16389=>"010000010",
  16390=>"001111001",
  16391=>"010000000",
  16392=>"100110110",
  16393=>"000001000",
  16394=>"111100011",
  16395=>"110111100",
  16396=>"000111111",
  16397=>"000101010",
  16398=>"101111110",
  16399=>"111111100",
  16400=>"010010000",
  16401=>"110110100",
  16402=>"101110000",
  16403=>"000011011",
  16404=>"100010011",
  16405=>"110000010",
  16406=>"101100101",
  16407=>"111101101",
  16408=>"111110110",
  16409=>"011111000",
  16410=>"000010000",
  16411=>"001100001",
  16412=>"001000001",
  16413=>"001011101",
  16414=>"110011101",
  16415=>"010010100",
  16416=>"010111111",
  16417=>"100101000",
  16418=>"100010001",
  16419=>"100011101",
  16420=>"101011101",
  16421=>"000101010",
  16422=>"011001101",
  16423=>"010000010",
  16424=>"000010110",
  16425=>"110100000",
  16426=>"111111110",
  16427=>"101111000",
  16428=>"011101111",
  16429=>"010110011",
  16430=>"110100100",
  16431=>"000010000",
  16432=>"010001010",
  16433=>"011011110",
  16434=>"000010000",
  16435=>"011100101",
  16436=>"110010101",
  16437=>"111100101",
  16438=>"010101001",
  16439=>"101110110",
  16440=>"101101011",
  16441=>"111010001",
  16442=>"010110101",
  16443=>"011010110",
  16444=>"000111100",
  16445=>"000001001",
  16446=>"111101101",
  16447=>"000111100",
  16448=>"100001010",
  16449=>"000110100",
  16450=>"111001110",
  16451=>"011101010",
  16452=>"101111000",
  16453=>"101111001",
  16454=>"001100001",
  16455=>"010110001",
  16456=>"110001101",
  16457=>"011001110",
  16458=>"101110110",
  16459=>"011010111",
  16460=>"011000110",
  16461=>"110010101",
  16462=>"111001110",
  16463=>"111110011",
  16464=>"111000011",
  16465=>"001011000",
  16466=>"111001001",
  16467=>"110000111",
  16468=>"110100010",
  16469=>"000000100",
  16470=>"110000100",
  16471=>"101001011",
  16472=>"110111110",
  16473=>"100011101",
  16474=>"110011011",
  16475=>"101100001",
  16476=>"010011011",
  16477=>"111101000",
  16478=>"110110001",
  16479=>"111001110",
  16480=>"011010010",
  16481=>"111001010",
  16482=>"111010010",
  16483=>"110101100",
  16484=>"101100010",
  16485=>"001111101",
  16486=>"000000000",
  16487=>"110010010",
  16488=>"111011111",
  16489=>"111000101",
  16490=>"011001000",
  16491=>"001011000",
  16492=>"001111000",
  16493=>"101010010",
  16494=>"100000010",
  16495=>"110001010",
  16496=>"001010000",
  16497=>"000001111",
  16498=>"010010110",
  16499=>"100100110",
  16500=>"111100010",
  16501=>"100000110",
  16502=>"010100110",
  16503=>"000111111",
  16504=>"101111100",
  16505=>"001000011",
  16506=>"111100110",
  16507=>"110110000",
  16508=>"110101101",
  16509=>"001110100",
  16510=>"000101110",
  16511=>"011011101",
  16512=>"011011101",
  16513=>"000111001",
  16514=>"000110011",
  16515=>"111011101",
  16516=>"100001000",
  16517=>"001110001",
  16518=>"011100110",
  16519=>"010000111",
  16520=>"000110100",
  16521=>"110110000",
  16522=>"100001011",
  16523=>"111110111",
  16524=>"100011111",
  16525=>"101011010",
  16526=>"100101110",
  16527=>"000100000",
  16528=>"111011011",
  16529=>"001110110",
  16530=>"111011011",
  16531=>"110110111",
  16532=>"100111110",
  16533=>"000011100",
  16534=>"100101100",
  16535=>"110111111",
  16536=>"010001011",
  16537=>"011100101",
  16538=>"101001010",
  16539=>"101011100",
  16540=>"110110001",
  16541=>"101010111",
  16542=>"101100100",
  16543=>"101000011",
  16544=>"110001011",
  16545=>"000101101",
  16546=>"000011111",
  16547=>"111110100",
  16548=>"001110000",
  16549=>"101001101",
  16550=>"101101011",
  16551=>"001110111",
  16552=>"110000110",
  16553=>"111001101",
  16554=>"100000110",
  16555=>"110000100",
  16556=>"000110100",
  16557=>"101010011",
  16558=>"100100011",
  16559=>"111001011",
  16560=>"001111111",
  16561=>"111011100",
  16562=>"101101101",
  16563=>"011001001",
  16564=>"000000111",
  16565=>"101100110",
  16566=>"111001011",
  16567=>"011101111",
  16568=>"100000000",
  16569=>"110011000",
  16570=>"101101001",
  16571=>"000101111",
  16572=>"011101110",
  16573=>"110100001",
  16574=>"011000110",
  16575=>"111010011",
  16576=>"000100001",
  16577=>"011001111",
  16578=>"100100100",
  16579=>"011110000",
  16580=>"001001000",
  16581=>"111010110",
  16582=>"001111000",
  16583=>"111100100",
  16584=>"011000000",
  16585=>"100011111",
  16586=>"101100111",
  16587=>"011000110",
  16588=>"001100101",
  16589=>"001011100",
  16590=>"101001100",
  16591=>"101000010",
  16592=>"110101010",
  16593=>"010111101",
  16594=>"000100111",
  16595=>"110000011",
  16596=>"101100001",
  16597=>"111000010",
  16598=>"100010110",
  16599=>"001101000",
  16600=>"010110110",
  16601=>"101100000",
  16602=>"000000011",
  16603=>"000100011",
  16604=>"001101110",
  16605=>"111110100",
  16606=>"110000111",
  16607=>"111000010",
  16608=>"101011111",
  16609=>"111000000",
  16610=>"100010100",
  16611=>"100001101",
  16612=>"100000000",
  16613=>"111011101",
  16614=>"111111010",
  16615=>"010101011",
  16616=>"011010110",
  16617=>"100011101",
  16618=>"101101000",
  16619=>"101101010",
  16620=>"110100111",
  16621=>"100010010",
  16622=>"111000000",
  16623=>"111000000",
  16624=>"010110110",
  16625=>"101000001",
  16626=>"111100001",
  16627=>"101010001",
  16628=>"001100010",
  16629=>"100111000",
  16630=>"010101010",
  16631=>"101111111",
  16632=>"110101011",
  16633=>"110101000",
  16634=>"110100000",
  16635=>"011010111",
  16636=>"101011001",
  16637=>"011000001",
  16638=>"111101011",
  16639=>"000010111",
  16640=>"000000011",
  16641=>"010001000",
  16642=>"101011011",
  16643=>"111101000",
  16644=>"011111100",
  16645=>"100001110",
  16646=>"110100010",
  16647=>"001100100",
  16648=>"110111011",
  16649=>"111011110",
  16650=>"000110110",
  16651=>"100000100",
  16652=>"010110111",
  16653=>"001110100",
  16654=>"111011000",
  16655=>"111010011",
  16656=>"000010100",
  16657=>"011111011",
  16658=>"000101101",
  16659=>"000110100",
  16660=>"100110101",
  16661=>"111111000",
  16662=>"000001111",
  16663=>"011111011",
  16664=>"101110000",
  16665=>"010010101",
  16666=>"111000010",
  16667=>"111111100",
  16668=>"111010010",
  16669=>"000001101",
  16670=>"011001100",
  16671=>"110111111",
  16672=>"111100110",
  16673=>"001001111",
  16674=>"000101101",
  16675=>"100101010",
  16676=>"010111001",
  16677=>"001010000",
  16678=>"000101111",
  16679=>"111001011",
  16680=>"101001100",
  16681=>"011011110",
  16682=>"001110000",
  16683=>"000110101",
  16684=>"100001111",
  16685=>"110100100",
  16686=>"110010000",
  16687=>"101011010",
  16688=>"011101001",
  16689=>"000001100",
  16690=>"011111110",
  16691=>"001110000",
  16692=>"111100100",
  16693=>"001101001",
  16694=>"001011011",
  16695=>"110001111",
  16696=>"110100111",
  16697=>"101100010",
  16698=>"011101011",
  16699=>"101111011",
  16700=>"111001111",
  16701=>"000000001",
  16702=>"100100110",
  16703=>"011010110",
  16704=>"110010111",
  16705=>"010000001",
  16706=>"110110101",
  16707=>"011101111",
  16708=>"010111100",
  16709=>"000001101",
  16710=>"000001110",
  16711=>"001000000",
  16712=>"000101010",
  16713=>"000000000",
  16714=>"100010010",
  16715=>"101111000",
  16716=>"001010111",
  16717=>"101010011",
  16718=>"110001100",
  16719=>"111010001",
  16720=>"000101110",
  16721=>"111111001",
  16722=>"100010010",
  16723=>"111000110",
  16724=>"001101110",
  16725=>"111010000",
  16726=>"100100110",
  16727=>"100111011",
  16728=>"111011100",
  16729=>"111011000",
  16730=>"000101111",
  16731=>"010011111",
  16732=>"011111010",
  16733=>"010001111",
  16734=>"100000111",
  16735=>"101010001",
  16736=>"110110111",
  16737=>"111011101",
  16738=>"110101110",
  16739=>"001011100",
  16740=>"000110001",
  16741=>"011111010",
  16742=>"110000000",
  16743=>"111011011",
  16744=>"100000000",
  16745=>"001101101",
  16746=>"001001101",
  16747=>"100010001",
  16748=>"110110100",
  16749=>"101000001",
  16750=>"100000100",
  16751=>"000010001",
  16752=>"100010110",
  16753=>"010111100",
  16754=>"001000100",
  16755=>"111101000",
  16756=>"001101100",
  16757=>"101001110",
  16758=>"001110000",
  16759=>"011011010",
  16760=>"100000101",
  16761=>"100101100",
  16762=>"111010000",
  16763=>"001011000",
  16764=>"111001001",
  16765=>"010011000",
  16766=>"011011001",
  16767=>"111001110",
  16768=>"010010000",
  16769=>"000110000",
  16770=>"000000000",
  16771=>"111100010",
  16772=>"110101000",
  16773=>"010000100",
  16774=>"101000111",
  16775=>"000100000",
  16776=>"000110000",
  16777=>"001100000",
  16778=>"100010101",
  16779=>"101010111",
  16780=>"100010100",
  16781=>"011010001",
  16782=>"111010000",
  16783=>"010010011",
  16784=>"101000101",
  16785=>"111111001",
  16786=>"101111010",
  16787=>"000010111",
  16788=>"111110100",
  16789=>"010011111",
  16790=>"110100010",
  16791=>"001001110",
  16792=>"001010110",
  16793=>"111000101",
  16794=>"101010010",
  16795=>"110011101",
  16796=>"001010111",
  16797=>"111111011",
  16798=>"011100101",
  16799=>"110100001",
  16800=>"011010001",
  16801=>"001111001",
  16802=>"001111001",
  16803=>"010101111",
  16804=>"101011000",
  16805=>"101001100",
  16806=>"100100000",
  16807=>"101011000",
  16808=>"100010111",
  16809=>"011100010",
  16810=>"101011001",
  16811=>"001101110",
  16812=>"000110111",
  16813=>"111011111",
  16814=>"101010110",
  16815=>"101111001",
  16816=>"100010011",
  16817=>"011100101",
  16818=>"111000101",
  16819=>"100000110",
  16820=>"111110110",
  16821=>"110110011",
  16822=>"000111000",
  16823=>"011100000",
  16824=>"110100011",
  16825=>"110101001",
  16826=>"001011000",
  16827=>"100011110",
  16828=>"001001100",
  16829=>"000100111",
  16830=>"110111111",
  16831=>"100001011",
  16832=>"101000011",
  16833=>"100111100",
  16834=>"010111011",
  16835=>"010011010",
  16836=>"000100000",
  16837=>"010010110",
  16838=>"011001001",
  16839=>"101111000",
  16840=>"000001111",
  16841=>"100110111",
  16842=>"101111010",
  16843=>"101010010",
  16844=>"000011100",
  16845=>"000010100",
  16846=>"000010111",
  16847=>"101011010",
  16848=>"011001000",
  16849=>"110111110",
  16850=>"000001100",
  16851=>"010111000",
  16852=>"110000101",
  16853=>"001010100",
  16854=>"011000100",
  16855=>"101100101",
  16856=>"001100011",
  16857=>"101111001",
  16858=>"110010101",
  16859=>"100100000",
  16860=>"011011110",
  16861=>"010000000",
  16862=>"100001000",
  16863=>"110001101",
  16864=>"110101010",
  16865=>"111100010",
  16866=>"011000101",
  16867=>"000110110",
  16868=>"101000001",
  16869=>"011010011",
  16870=>"110110100",
  16871=>"101001100",
  16872=>"000011001",
  16873=>"010001010",
  16874=>"110111011",
  16875=>"001010000",
  16876=>"100010110",
  16877=>"100011000",
  16878=>"110011011",
  16879=>"001000001",
  16880=>"001111010",
  16881=>"110010111",
  16882=>"011001010",
  16883=>"001101001",
  16884=>"000000101",
  16885=>"100100010",
  16886=>"011011110",
  16887=>"100001101",
  16888=>"000100011",
  16889=>"000010100",
  16890=>"111011101",
  16891=>"010110111",
  16892=>"111110101",
  16893=>"011011100",
  16894=>"110100111",
  16895=>"010110001",
  16896=>"101001011",
  16897=>"111001111",
  16898=>"101111001",
  16899=>"001111101",
  16900=>"100010010",
  16901=>"011000111",
  16902=>"110011010",
  16903=>"010001110",
  16904=>"000101101",
  16905=>"101110010",
  16906=>"100100010",
  16907=>"111011101",
  16908=>"010001101",
  16909=>"001111111",
  16910=>"101110100",
  16911=>"010010111",
  16912=>"010110000",
  16913=>"101101011",
  16914=>"100011101",
  16915=>"100010001",
  16916=>"010010001",
  16917=>"010110110",
  16918=>"111000101",
  16919=>"111110100",
  16920=>"000000101",
  16921=>"001010000",
  16922=>"101001010",
  16923=>"110011000",
  16924=>"000001011",
  16925=>"101101111",
  16926=>"100000000",
  16927=>"000011101",
  16928=>"111010110",
  16929=>"011001010",
  16930=>"100101010",
  16931=>"011000111",
  16932=>"001110011",
  16933=>"100000101",
  16934=>"111011111",
  16935=>"000111000",
  16936=>"110011111",
  16937=>"111101010",
  16938=>"100101011",
  16939=>"011101110",
  16940=>"111000011",
  16941=>"100001101",
  16942=>"001100101",
  16943=>"101010101",
  16944=>"110001110",
  16945=>"000010110",
  16946=>"010101110",
  16947=>"100000100",
  16948=>"110111110",
  16949=>"010011111",
  16950=>"000101011",
  16951=>"000101011",
  16952=>"100011111",
  16953=>"001110011",
  16954=>"010101001",
  16955=>"111011110",
  16956=>"100001001",
  16957=>"000011100",
  16958=>"000001110",
  16959=>"100110001",
  16960=>"101010001",
  16961=>"011001110",
  16962=>"110000000",
  16963=>"100001000",
  16964=>"001011100",
  16965=>"101011000",
  16966=>"111110110",
  16967=>"010001110",
  16968=>"001111111",
  16969=>"011001010",
  16970=>"011001100",
  16971=>"011010001",
  16972=>"111101110",
  16973=>"011011011",
  16974=>"011001010",
  16975=>"011011111",
  16976=>"110111101",
  16977=>"000100111",
  16978=>"100000001",
  16979=>"101001011",
  16980=>"001110011",
  16981=>"011101010",
  16982=>"000110111",
  16983=>"101000011",
  16984=>"011011110",
  16985=>"010010111",
  16986=>"010101011",
  16987=>"010010011",
  16988=>"010001011",
  16989=>"101100001",
  16990=>"110000100",
  16991=>"010011011",
  16992=>"010001110",
  16993=>"000011101",
  16994=>"110101110",
  16995=>"110001100",
  16996=>"100110011",
  16997=>"001001000",
  16998=>"110010111",
  16999=>"010100101",
  17000=>"100001010",
  17001=>"110110111",
  17002=>"100000110",
  17003=>"110111100",
  17004=>"100100111",
  17005=>"111111101",
  17006=>"110011000",
  17007=>"000000111",
  17008=>"010010001",
  17009=>"000000000",
  17010=>"010101101",
  17011=>"001000100",
  17012=>"110111000",
  17013=>"001011101",
  17014=>"100000110",
  17015=>"001001111",
  17016=>"011100011",
  17017=>"010110101",
  17018=>"001101010",
  17019=>"001111100",
  17020=>"000110001",
  17021=>"110110000",
  17022=>"000010011",
  17023=>"001000100",
  17024=>"011000011",
  17025=>"010011100",
  17026=>"001110101",
  17027=>"110111001",
  17028=>"000000011",
  17029=>"101000000",
  17030=>"001010000",
  17031=>"000010011",
  17032=>"010110011",
  17033=>"100100000",
  17034=>"110011110",
  17035=>"001111000",
  17036=>"000110011",
  17037=>"000101101",
  17038=>"100101011",
  17039=>"001110010",
  17040=>"110101110",
  17041=>"010001111",
  17042=>"101000011",
  17043=>"111010111",
  17044=>"011000101",
  17045=>"100011011",
  17046=>"011011010",
  17047=>"000001111",
  17048=>"110110101",
  17049=>"001011000",
  17050=>"000010111",
  17051=>"101101110",
  17052=>"010001010",
  17053=>"101011000",
  17054=>"100111001",
  17055=>"011011101",
  17056=>"001110001",
  17057=>"001001011",
  17058=>"000001111",
  17059=>"010011011",
  17060=>"101000000",
  17061=>"011111010",
  17062=>"111000010",
  17063=>"010100110",
  17064=>"111011011",
  17065=>"011000000",
  17066=>"100000101",
  17067=>"110010010",
  17068=>"110011000",
  17069=>"011111010",
  17070=>"000001111",
  17071=>"110010000",
  17072=>"100000110",
  17073=>"110100101",
  17074=>"111000110",
  17075=>"110110010",
  17076=>"011100001",
  17077=>"110110011",
  17078=>"000011110",
  17079=>"000011010",
  17080=>"110111101",
  17081=>"100010101",
  17082=>"001101111",
  17083=>"011000001",
  17084=>"010100101",
  17085=>"000000100",
  17086=>"110100010",
  17087=>"001010010",
  17088=>"110110111",
  17089=>"011111101",
  17090=>"001000011",
  17091=>"111000010",
  17092=>"111011000",
  17093=>"110100000",
  17094=>"100111000",
  17095=>"000001001",
  17096=>"101101110",
  17097=>"000011001",
  17098=>"111100110",
  17099=>"101010010",
  17100=>"111010101",
  17101=>"010100100",
  17102=>"101011101",
  17103=>"101000111",
  17104=>"000001000",
  17105=>"010110110",
  17106=>"011010110",
  17107=>"011010111",
  17108=>"001011100",
  17109=>"010101000",
  17110=>"110010000",
  17111=>"001111000",
  17112=>"011001000",
  17113=>"111010110",
  17114=>"000101000",
  17115=>"110010001",
  17116=>"111101101",
  17117=>"100001000",
  17118=>"101100000",
  17119=>"000100101",
  17120=>"010110001",
  17121=>"110100010",
  17122=>"111000100",
  17123=>"011100010",
  17124=>"110011111",
  17125=>"101001100",
  17126=>"010100000",
  17127=>"000000101",
  17128=>"111011011",
  17129=>"111111001",
  17130=>"010100001",
  17131=>"011000110",
  17132=>"010111111",
  17133=>"010000100",
  17134=>"101000001",
  17135=>"110000010",
  17136=>"011101010",
  17137=>"000111000",
  17138=>"111111011",
  17139=>"011110110",
  17140=>"100011110",
  17141=>"001110111",
  17142=>"011011101",
  17143=>"000111000",
  17144=>"110000010",
  17145=>"101100101",
  17146=>"101000001",
  17147=>"011101101",
  17148=>"100100111",
  17149=>"101101000",
  17150=>"010000011",
  17151=>"101000110",
  17152=>"110000011",
  17153=>"111101000",
  17154=>"000100011",
  17155=>"101100001",
  17156=>"100000111",
  17157=>"000101000",
  17158=>"111101101",
  17159=>"100101101",
  17160=>"011101110",
  17161=>"101100111",
  17162=>"010000101",
  17163=>"010000010",
  17164=>"010111011",
  17165=>"010000010",
  17166=>"110000111",
  17167=>"011000000",
  17168=>"010010111",
  17169=>"001110011",
  17170=>"111110001",
  17171=>"111110000",
  17172=>"000000110",
  17173=>"010011000",
  17174=>"101000010",
  17175=>"101011010",
  17176=>"111101001",
  17177=>"110010100",
  17178=>"100100101",
  17179=>"111110111",
  17180=>"011100000",
  17181=>"110111111",
  17182=>"110100111",
  17183=>"010100101",
  17184=>"010101101",
  17185=>"110111111",
  17186=>"101000100",
  17187=>"011101111",
  17188=>"111001101",
  17189=>"110011001",
  17190=>"110010111",
  17191=>"000110101",
  17192=>"000000111",
  17193=>"011011011",
  17194=>"010111011",
  17195=>"001101000",
  17196=>"110100001",
  17197=>"011000100",
  17198=>"001110100",
  17199=>"000010000",
  17200=>"010011110",
  17201=>"011011100",
  17202=>"000111111",
  17203=>"010001000",
  17204=>"011010010",
  17205=>"010000001",
  17206=>"101111110",
  17207=>"111000111",
  17208=>"111111101",
  17209=>"000001110",
  17210=>"000000000",
  17211=>"011010100",
  17212=>"100001101",
  17213=>"100010010",
  17214=>"000001011",
  17215=>"000010100",
  17216=>"011100010",
  17217=>"010000101",
  17218=>"111011001",
  17219=>"111100101",
  17220=>"110000100",
  17221=>"001010111",
  17222=>"100011110",
  17223=>"100001110",
  17224=>"111111110",
  17225=>"110100100",
  17226=>"011110101",
  17227=>"110100001",
  17228=>"011000011",
  17229=>"100111101",
  17230=>"101100001",
  17231=>"001011110",
  17232=>"011100101",
  17233=>"111010000",
  17234=>"110001011",
  17235=>"001001000",
  17236=>"010110100",
  17237=>"100000111",
  17238=>"000000111",
  17239=>"111101001",
  17240=>"011010011",
  17241=>"100011011",
  17242=>"101111011",
  17243=>"001101001",
  17244=>"101111001",
  17245=>"100101011",
  17246=>"111011010",
  17247=>"100101011",
  17248=>"010111010",
  17249=>"011010100",
  17250=>"101100010",
  17251=>"101001110",
  17252=>"101111010",
  17253=>"111001000",
  17254=>"010010011",
  17255=>"100010011",
  17256=>"110000110",
  17257=>"001100011",
  17258=>"111111011",
  17259=>"010110110",
  17260=>"001000000",
  17261=>"001111010",
  17262=>"011101010",
  17263=>"011011001",
  17264=>"101101100",
  17265=>"010011010",
  17266=>"110111001",
  17267=>"001101100",
  17268=>"011101101",
  17269=>"100001001",
  17270=>"111100001",
  17271=>"100011110",
  17272=>"100000000",
  17273=>"001100111",
  17274=>"011011010",
  17275=>"011001101",
  17276=>"110011110",
  17277=>"010101101",
  17278=>"011110011",
  17279=>"011100000",
  17280=>"100100100",
  17281=>"110100001",
  17282=>"001000100",
  17283=>"111101011",
  17284=>"011101111",
  17285=>"111100000",
  17286=>"101110010",
  17287=>"010001110",
  17288=>"101100101",
  17289=>"100010110",
  17290=>"100111010",
  17291=>"111100011",
  17292=>"001100000",
  17293=>"011110111",
  17294=>"000100100",
  17295=>"010011110",
  17296=>"011000001",
  17297=>"000011110",
  17298=>"100010111",
  17299=>"111111000",
  17300=>"101011110",
  17301=>"110111001",
  17302=>"011001101",
  17303=>"101111111",
  17304=>"010000101",
  17305=>"001001100",
  17306=>"000110011",
  17307=>"001100011",
  17308=>"111010000",
  17309=>"111101110",
  17310=>"000100101",
  17311=>"001110111",
  17312=>"111001001",
  17313=>"101011001",
  17314=>"111110011",
  17315=>"011111010",
  17316=>"011110111",
  17317=>"001101111",
  17318=>"101100011",
  17319=>"101001011",
  17320=>"001101101",
  17321=>"010011000",
  17322=>"011111110",
  17323=>"010100011",
  17324=>"010001111",
  17325=>"100111100",
  17326=>"110110110",
  17327=>"000100100",
  17328=>"110000100",
  17329=>"010100111",
  17330=>"011111010",
  17331=>"010110001",
  17332=>"111100001",
  17333=>"011010100",
  17334=>"101110011",
  17335=>"010111001",
  17336=>"111010010",
  17337=>"010111000",
  17338=>"100100101",
  17339=>"110001010",
  17340=>"110100111",
  17341=>"100100000",
  17342=>"010110111",
  17343=>"101111011",
  17344=>"001010011",
  17345=>"010010110",
  17346=>"001100001",
  17347=>"100110010",
  17348=>"101011101",
  17349=>"000001010",
  17350=>"000000010",
  17351=>"100100101",
  17352=>"111000101",
  17353=>"110101101",
  17354=>"000101101",
  17355=>"000011100",
  17356=>"010000100",
  17357=>"010001100",
  17358=>"001001001",
  17359=>"001001110",
  17360=>"110000100",
  17361=>"011001101",
  17362=>"000010011",
  17363=>"100100010",
  17364=>"011101101",
  17365=>"010001011",
  17366=>"110011010",
  17367=>"000111011",
  17368=>"100100001",
  17369=>"110000111",
  17370=>"011100010",
  17371=>"101111110",
  17372=>"010110000",
  17373=>"110100000",
  17374=>"000000011",
  17375=>"011000110",
  17376=>"101010100",
  17377=>"110011001",
  17378=>"011011111",
  17379=>"111101010",
  17380=>"101101010",
  17381=>"111100001",
  17382=>"101010011",
  17383=>"100011010",
  17384=>"111011111",
  17385=>"000001011",
  17386=>"110000110",
  17387=>"011111111",
  17388=>"010101011",
  17389=>"110000111",
  17390=>"100000111",
  17391=>"100110011",
  17392=>"010010101",
  17393=>"110010010",
  17394=>"100011100",
  17395=>"001011000",
  17396=>"011111110",
  17397=>"000111100",
  17398=>"111101101",
  17399=>"011001110",
  17400=>"011010001",
  17401=>"001111010",
  17402=>"110000100",
  17403=>"000001011",
  17404=>"000010100",
  17405=>"101111001",
  17406=>"110000100",
  17407=>"010001000",
  17408=>"000110110",
  17409=>"001001011",
  17410=>"010101101",
  17411=>"001010010",
  17412=>"111010110",
  17413=>"011101111",
  17414=>"110000010",
  17415=>"011110011",
  17416=>"111111011",
  17417=>"001001011",
  17418=>"111101000",
  17419=>"111101001",
  17420=>"110101101",
  17421=>"110100000",
  17422=>"011001000",
  17423=>"100000110",
  17424=>"001000111",
  17425=>"001110001",
  17426=>"010011111",
  17427=>"110110101",
  17428=>"100101010",
  17429=>"101000010",
  17430=>"100111111",
  17431=>"001001010",
  17432=>"011001010",
  17433=>"111111101",
  17434=>"000111110",
  17435=>"111111101",
  17436=>"000010000",
  17437=>"100111000",
  17438=>"100111100",
  17439=>"010100000",
  17440=>"111101010",
  17441=>"001011111",
  17442=>"001111101",
  17443=>"010101101",
  17444=>"111111101",
  17445=>"010111000",
  17446=>"001010011",
  17447=>"101111100",
  17448=>"010001101",
  17449=>"010000000",
  17450=>"101001010",
  17451=>"101100010",
  17452=>"101101111",
  17453=>"011010010",
  17454=>"001111010",
  17455=>"111011000",
  17456=>"001101101",
  17457=>"100010010",
  17458=>"111001101",
  17459=>"101100111",
  17460=>"111000011",
  17461=>"111110111",
  17462=>"110110100",
  17463=>"110101000",
  17464=>"010001100",
  17465=>"000100100",
  17466=>"001001110",
  17467=>"011100101",
  17468=>"000000001",
  17469=>"000000111",
  17470=>"010110100",
  17471=>"100110101",
  17472=>"010010010",
  17473=>"000101110",
  17474=>"001011110",
  17475=>"000010000",
  17476=>"000111001",
  17477=>"001001111",
  17478=>"110111001",
  17479=>"101100100",
  17480=>"111010111",
  17481=>"111000101",
  17482=>"011100101",
  17483=>"101111110",
  17484=>"100101010",
  17485=>"010001000",
  17486=>"000010100",
  17487=>"101101011",
  17488=>"000000111",
  17489=>"111111101",
  17490=>"011000000",
  17491=>"100010100",
  17492=>"011100000",
  17493=>"011100101",
  17494=>"000101111",
  17495=>"000110001",
  17496=>"011101001",
  17497=>"111110111",
  17498=>"101110100",
  17499=>"000110000",
  17500=>"010010000",
  17501=>"001100111",
  17502=>"010011110",
  17503=>"110011000",
  17504=>"101001100",
  17505=>"011001001",
  17506=>"110000000",
  17507=>"010110000",
  17508=>"010010010",
  17509=>"011110001",
  17510=>"110110101",
  17511=>"010000011",
  17512=>"110000101",
  17513=>"100111100",
  17514=>"100110000",
  17515=>"010110010",
  17516=>"000001000",
  17517=>"111010101",
  17518=>"011110110",
  17519=>"011000001",
  17520=>"111111111",
  17521=>"100100101",
  17522=>"001001011",
  17523=>"100010001",
  17524=>"101001100",
  17525=>"111011001",
  17526=>"100111000",
  17527=>"001110010",
  17528=>"001110000",
  17529=>"100001000",
  17530=>"000011001",
  17531=>"010100010",
  17532=>"110111010",
  17533=>"111011010",
  17534=>"010100110",
  17535=>"000111100",
  17536=>"100001100",
  17537=>"011011101",
  17538=>"000011000",
  17539=>"111010010",
  17540=>"000001010",
  17541=>"011000111",
  17542=>"101101101",
  17543=>"110111100",
  17544=>"000110010",
  17545=>"101000000",
  17546=>"110001101",
  17547=>"101111010",
  17548=>"000001101",
  17549=>"001000111",
  17550=>"010100000",
  17551=>"000111110",
  17552=>"111010011",
  17553=>"001001110",
  17554=>"000011010",
  17555=>"111101110",
  17556=>"111101111",
  17557=>"000001101",
  17558=>"010011000",
  17559=>"111110100",
  17560=>"011101001",
  17561=>"010100011",
  17562=>"100010111",
  17563=>"010100010",
  17564=>"000100100",
  17565=>"111101000",
  17566=>"001010010",
  17567=>"010101110",
  17568=>"111010001",
  17569=>"000111010",
  17570=>"101011001",
  17571=>"101000111",
  17572=>"111011111",
  17573=>"010000010",
  17574=>"000100001",
  17575=>"110011101",
  17576=>"110000111",
  17577=>"101001001",
  17578=>"010100001",
  17579=>"100110010",
  17580=>"000000100",
  17581=>"011000100",
  17582=>"101101111",
  17583=>"100010010",
  17584=>"011001010",
  17585=>"110001100",
  17586=>"011110000",
  17587=>"000111000",
  17588=>"011000110",
  17589=>"101101101",
  17590=>"100100100",
  17591=>"111101010",
  17592=>"101011100",
  17593=>"010000101",
  17594=>"101111000",
  17595=>"011010010",
  17596=>"010010001",
  17597=>"101011010",
  17598=>"101001111",
  17599=>"011010100",
  17600=>"101010111",
  17601=>"110011101",
  17602=>"001011111",
  17603=>"000101111",
  17604=>"110100101",
  17605=>"010001101",
  17606=>"000111010",
  17607=>"110001111",
  17608=>"010010110",
  17609=>"001100111",
  17610=>"001000101",
  17611=>"101001100",
  17612=>"100001101",
  17613=>"011101001",
  17614=>"100111101",
  17615=>"110000011",
  17616=>"111110010",
  17617=>"011010001",
  17618=>"010110101",
  17619=>"011101011",
  17620=>"100001001",
  17621=>"000001011",
  17622=>"010110000",
  17623=>"010100101",
  17624=>"100010010",
  17625=>"010001010",
  17626=>"001100101",
  17627=>"011010111",
  17628=>"001110111",
  17629=>"010001100",
  17630=>"000100011",
  17631=>"011111111",
  17632=>"110001101",
  17633=>"111110001",
  17634=>"110001100",
  17635=>"010001011",
  17636=>"010100101",
  17637=>"111011101",
  17638=>"111100101",
  17639=>"011010111",
  17640=>"100000010",
  17641=>"010000010",
  17642=>"110100111",
  17643=>"011110101",
  17644=>"000100100",
  17645=>"010010000",
  17646=>"000000010",
  17647=>"010001000",
  17648=>"011010000",
  17649=>"111101001",
  17650=>"001111111",
  17651=>"011101011",
  17652=>"101110101",
  17653=>"000010100",
  17654=>"001011000",
  17655=>"111001000",
  17656=>"111001001",
  17657=>"101010011",
  17658=>"110001000",
  17659=>"001001001",
  17660=>"100000111",
  17661=>"111011101",
  17662=>"001110010",
  17663=>"111110100",
  17664=>"010000010",
  17665=>"110100011",
  17666=>"000010011",
  17667=>"000111010",
  17668=>"111111101",
  17669=>"001111001",
  17670=>"010011010",
  17671=>"000110001",
  17672=>"110111010",
  17673=>"010100011",
  17674=>"101011010",
  17675=>"010010001",
  17676=>"100010100",
  17677=>"110100010",
  17678=>"111111000",
  17679=>"010001100",
  17680=>"000111110",
  17681=>"011100100",
  17682=>"000000000",
  17683=>"100100011",
  17684=>"100010111",
  17685=>"000100101",
  17686=>"110100010",
  17687=>"110111100",
  17688=>"010000011",
  17689=>"011000011",
  17690=>"010100010",
  17691=>"010000011",
  17692=>"110101101",
  17693=>"000101101",
  17694=>"001011111",
  17695=>"100001001",
  17696=>"001100010",
  17697=>"010010100",
  17698=>"101010101",
  17699=>"000000100",
  17700=>"110111001",
  17701=>"011001011",
  17702=>"000010011",
  17703=>"010100100",
  17704=>"000100100",
  17705=>"111110111",
  17706=>"011000111",
  17707=>"111000001",
  17708=>"010110100",
  17709=>"011011110",
  17710=>"010101101",
  17711=>"011111111",
  17712=>"000110010",
  17713=>"010010111",
  17714=>"001010010",
  17715=>"001110000",
  17716=>"111000010",
  17717=>"111011001",
  17718=>"100111111",
  17719=>"011010011",
  17720=>"000111101",
  17721=>"001010110",
  17722=>"111111001",
  17723=>"001011110",
  17724=>"111101001",
  17725=>"001000010",
  17726=>"000011111",
  17727=>"000000100",
  17728=>"111110011",
  17729=>"000110011",
  17730=>"101110011",
  17731=>"011101100",
  17732=>"100000010",
  17733=>"101100110",
  17734=>"010011101",
  17735=>"000111111",
  17736=>"001001000",
  17737=>"011010110",
  17738=>"011000001",
  17739=>"101110000",
  17740=>"101110111",
  17741=>"001111011",
  17742=>"111010001",
  17743=>"101000111",
  17744=>"100110100",
  17745=>"001000000",
  17746=>"010000010",
  17747=>"000001110",
  17748=>"000000100",
  17749=>"011000000",
  17750=>"011110100",
  17751=>"010111000",
  17752=>"010010101",
  17753=>"000110001",
  17754=>"111111110",
  17755=>"011001001",
  17756=>"001110101",
  17757=>"111010110",
  17758=>"000111001",
  17759=>"000010001",
  17760=>"001110010",
  17761=>"011100100",
  17762=>"010011100",
  17763=>"000101101",
  17764=>"011010000",
  17765=>"000001101",
  17766=>"111111110",
  17767=>"110011101",
  17768=>"101011000",
  17769=>"000110110",
  17770=>"100111001",
  17771=>"011010111",
  17772=>"101101000",
  17773=>"011110111",
  17774=>"100001110",
  17775=>"100111011",
  17776=>"100000000",
  17777=>"011011011",
  17778=>"001101001",
  17779=>"100101010",
  17780=>"110000100",
  17781=>"001011111",
  17782=>"100010110",
  17783=>"010000011",
  17784=>"001110000",
  17785=>"001001001",
  17786=>"100010111",
  17787=>"110000000",
  17788=>"110110101",
  17789=>"110000101",
  17790=>"111011000",
  17791=>"110001101",
  17792=>"010101101",
  17793=>"011011010",
  17794=>"111010111",
  17795=>"001010000",
  17796=>"101101110",
  17797=>"100010110",
  17798=>"101000101",
  17799=>"011010000",
  17800=>"101100000",
  17801=>"001111000",
  17802=>"100000011",
  17803=>"010100101",
  17804=>"000000010",
  17805=>"001111100",
  17806=>"101111111",
  17807=>"100100101",
  17808=>"110010000",
  17809=>"111001101",
  17810=>"011111100",
  17811=>"111010111",
  17812=>"100010101",
  17813=>"001000000",
  17814=>"000100001",
  17815=>"001001001",
  17816=>"010011100",
  17817=>"001010110",
  17818=>"001001011",
  17819=>"111010110",
  17820=>"110000000",
  17821=>"000010101",
  17822=>"100011001",
  17823=>"101000111",
  17824=>"110010001",
  17825=>"101000100",
  17826=>"100011001",
  17827=>"010000010",
  17828=>"100101100",
  17829=>"010100010",
  17830=>"011110011",
  17831=>"101011100",
  17832=>"001110011",
  17833=>"000100000",
  17834=>"100000110",
  17835=>"110010110",
  17836=>"010100000",
  17837=>"010111010",
  17838=>"110011011",
  17839=>"010110110",
  17840=>"100010011",
  17841=>"101011010",
  17842=>"111100110",
  17843=>"100000100",
  17844=>"000100101",
  17845=>"000000111",
  17846=>"110110010",
  17847=>"000111100",
  17848=>"001100101",
  17849=>"100010001",
  17850=>"111011100",
  17851=>"110111011",
  17852=>"100000100",
  17853=>"111100111",
  17854=>"001010110",
  17855=>"100000100",
  17856=>"001101010",
  17857=>"000000110",
  17858=>"011100011",
  17859=>"111011011",
  17860=>"100111110",
  17861=>"110101100",
  17862=>"000111001",
  17863=>"101010100",
  17864=>"000111110",
  17865=>"010010110",
  17866=>"011101110",
  17867=>"001101111",
  17868=>"000110000",
  17869=>"101011100",
  17870=>"001001000",
  17871=>"010001101",
  17872=>"000010011",
  17873=>"100000011",
  17874=>"011011111",
  17875=>"000110111",
  17876=>"001110101",
  17877=>"110000010",
  17878=>"100101110",
  17879=>"110111100",
  17880=>"101001010",
  17881=>"111111101",
  17882=>"001100001",
  17883=>"110010110",
  17884=>"101101111",
  17885=>"001010100",
  17886=>"110100111",
  17887=>"000000000",
  17888=>"111100000",
  17889=>"001110111",
  17890=>"101010010",
  17891=>"000010000",
  17892=>"001010000",
  17893=>"000010000",
  17894=>"001100010",
  17895=>"100111001",
  17896=>"000110001",
  17897=>"000011010",
  17898=>"001011111",
  17899=>"001001011",
  17900=>"000000110",
  17901=>"001010010",
  17902=>"010110100",
  17903=>"000000011",
  17904=>"101111111",
  17905=>"101000101",
  17906=>"011000000",
  17907=>"110101100",
  17908=>"100100011",
  17909=>"011010001",
  17910=>"010101010",
  17911=>"111011010",
  17912=>"000101101",
  17913=>"011110000",
  17914=>"110011111",
  17915=>"111101110",
  17916=>"101010011",
  17917=>"010111100",
  17918=>"011001101",
  17919=>"111110001",
  17920=>"010000010",
  17921=>"000100000",
  17922=>"100110011",
  17923=>"001110010",
  17924=>"100000110",
  17925=>"101101011",
  17926=>"011011011",
  17927=>"100001011",
  17928=>"001001100",
  17929=>"111101001",
  17930=>"011100101",
  17931=>"011000100",
  17932=>"100111111",
  17933=>"101000010",
  17934=>"011110111",
  17935=>"111100101",
  17936=>"001011100",
  17937=>"101011011",
  17938=>"000010001",
  17939=>"010010010",
  17940=>"000000010",
  17941=>"101001100",
  17942=>"100111111",
  17943=>"011000000",
  17944=>"111101000",
  17945=>"011110111",
  17946=>"101001100",
  17947=>"001110110",
  17948=>"111100000",
  17949=>"000111101",
  17950=>"100100000",
  17951=>"101101011",
  17952=>"010010000",
  17953=>"100001001",
  17954=>"100000110",
  17955=>"011111110",
  17956=>"001010110",
  17957=>"101000001",
  17958=>"101001010",
  17959=>"010010001",
  17960=>"001110010",
  17961=>"001111101",
  17962=>"101101111",
  17963=>"011100101",
  17964=>"100100100",
  17965=>"010001001",
  17966=>"111001001",
  17967=>"011100000",
  17968=>"010100011",
  17969=>"111111111",
  17970=>"111101101",
  17971=>"100011110",
  17972=>"001101100",
  17973=>"010001000",
  17974=>"110011111",
  17975=>"000101001",
  17976=>"011000001",
  17977=>"011001110",
  17978=>"001110000",
  17979=>"111110000",
  17980=>"101000010",
  17981=>"111111110",
  17982=>"111010100",
  17983=>"010100011",
  17984=>"111100000",
  17985=>"001101001",
  17986=>"100100101",
  17987=>"000010111",
  17988=>"111101011",
  17989=>"001011010",
  17990=>"100101111",
  17991=>"010111111",
  17992=>"001100101",
  17993=>"000111000",
  17994=>"101000010",
  17995=>"001101111",
  17996=>"101100011",
  17997=>"101001100",
  17998=>"011011100",
  17999=>"001001001",
  18000=>"111111111",
  18001=>"100101000",
  18002=>"000111011",
  18003=>"010111111",
  18004=>"000100100",
  18005=>"111010011",
  18006=>"100100100",
  18007=>"111010000",
  18008=>"101010000",
  18009=>"111001110",
  18010=>"110101000",
  18011=>"100011101",
  18012=>"101010110",
  18013=>"100100100",
  18014=>"010000111",
  18015=>"110111010",
  18016=>"000010111",
  18017=>"101001011",
  18018=>"011000011",
  18019=>"000001010",
  18020=>"111000000",
  18021=>"000000010",
  18022=>"000000111",
  18023=>"001000000",
  18024=>"001111101",
  18025=>"010110101",
  18026=>"111101010",
  18027=>"100111100",
  18028=>"010000010",
  18029=>"100000011",
  18030=>"100011000",
  18031=>"100001110",
  18032=>"111010000",
  18033=>"000000101",
  18034=>"010100101",
  18035=>"100110110",
  18036=>"100001111",
  18037=>"110111100",
  18038=>"001111011",
  18039=>"101110101",
  18040=>"010011100",
  18041=>"101100101",
  18042=>"010001011",
  18043=>"011101100",
  18044=>"001110100",
  18045=>"101110001",
  18046=>"101111101",
  18047=>"000111110",
  18048=>"100010010",
  18049=>"100101010",
  18050=>"101011100",
  18051=>"100110100",
  18052=>"011111000",
  18053=>"110001100",
  18054=>"101011000",
  18055=>"101010001",
  18056=>"101110101",
  18057=>"010110010",
  18058=>"101111001",
  18059=>"101000100",
  18060=>"100111100",
  18061=>"000000100",
  18062=>"100011011",
  18063=>"001001010",
  18064=>"111110111",
  18065=>"101001001",
  18066=>"000111101",
  18067=>"101000110",
  18068=>"110000011",
  18069=>"001100001",
  18070=>"100011011",
  18071=>"011010100",
  18072=>"010010011",
  18073=>"010010000",
  18074=>"110111000",
  18075=>"110000001",
  18076=>"101011010",
  18077=>"100101110",
  18078=>"001100000",
  18079=>"011001111",
  18080=>"100101101",
  18081=>"101010110",
  18082=>"001111111",
  18083=>"110001010",
  18084=>"010101110",
  18085=>"110111010",
  18086=>"010100010",
  18087=>"100010001",
  18088=>"110001100",
  18089=>"000001010",
  18090=>"010110011",
  18091=>"001000001",
  18092=>"000000110",
  18093=>"100110110",
  18094=>"010100011",
  18095=>"100011100",
  18096=>"111001001",
  18097=>"110000101",
  18098=>"100001000",
  18099=>"100010101",
  18100=>"100011100",
  18101=>"110001001",
  18102=>"100001100",
  18103=>"000001011",
  18104=>"001011110",
  18105=>"000001100",
  18106=>"010011111",
  18107=>"100011110",
  18108=>"000110011",
  18109=>"101000010",
  18110=>"000001000",
  18111=>"000010100",
  18112=>"011000101",
  18113=>"011101111",
  18114=>"000100110",
  18115=>"110011001",
  18116=>"010000111",
  18117=>"000010001",
  18118=>"111110011",
  18119=>"111101011",
  18120=>"001010010",
  18121=>"111111110",
  18122=>"110001111",
  18123=>"000000000",
  18124=>"011111111",
  18125=>"001010011",
  18126=>"000000010",
  18127=>"011100110",
  18128=>"010110101",
  18129=>"111000001",
  18130=>"101101011",
  18131=>"110000010",
  18132=>"101110000",
  18133=>"101111010",
  18134=>"101001011",
  18135=>"010010110",
  18136=>"101111001",
  18137=>"001000011",
  18138=>"111101001",
  18139=>"101111011",
  18140=>"110011111",
  18141=>"100101111",
  18142=>"000010100",
  18143=>"101000101",
  18144=>"010011001",
  18145=>"001111111",
  18146=>"010100010",
  18147=>"111001101",
  18148=>"111000011",
  18149=>"011001010",
  18150=>"001001000",
  18151=>"101001010",
  18152=>"001011010",
  18153=>"101010110",
  18154=>"011100000",
  18155=>"000010010",
  18156=>"000010111",
  18157=>"011100000",
  18158=>"111111100",
  18159=>"000110110",
  18160=>"110110110",
  18161=>"111000100",
  18162=>"111111100",
  18163=>"010011111",
  18164=>"001011100",
  18165=>"001011101",
  18166=>"111001011",
  18167=>"110010010",
  18168=>"011011000",
  18169=>"100110100",
  18170=>"101001010",
  18171=>"110010001",
  18172=>"000000010",
  18173=>"100111011",
  18174=>"000000101",
  18175=>"111111101",
  18176=>"111001001",
  18177=>"111110110",
  18178=>"010001101",
  18179=>"111110011",
  18180=>"000111110",
  18181=>"110101100",
  18182=>"100000010",
  18183=>"101101101",
  18184=>"111101000",
  18185=>"000011101",
  18186=>"011011010",
  18187=>"000010111",
  18188=>"111111000",
  18189=>"101111010",
  18190=>"001100100",
  18191=>"001001111",
  18192=>"110010011",
  18193=>"111000111",
  18194=>"110101100",
  18195=>"010110000",
  18196=>"001001101",
  18197=>"000010110",
  18198=>"000010010",
  18199=>"110101001",
  18200=>"100000000",
  18201=>"001110000",
  18202=>"111001010",
  18203=>"001000010",
  18204=>"101111101",
  18205=>"101110000",
  18206=>"010000001",
  18207=>"111011010",
  18208=>"000011100",
  18209=>"101110111",
  18210=>"001001100",
  18211=>"101110011",
  18212=>"111001000",
  18213=>"101100100",
  18214=>"001001001",
  18215=>"111000010",
  18216=>"100110111",
  18217=>"100010100",
  18218=>"101010100",
  18219=>"100000000",
  18220=>"111000111",
  18221=>"011100011",
  18222=>"011100000",
  18223=>"010110001",
  18224=>"101010001",
  18225=>"000011010",
  18226=>"011101011",
  18227=>"101011100",
  18228=>"111100111",
  18229=>"010011010",
  18230=>"101111011",
  18231=>"011111011",
  18232=>"001001010",
  18233=>"011010001",
  18234=>"001100110",
  18235=>"100010010",
  18236=>"101111111",
  18237=>"101110111",
  18238=>"000111010",
  18239=>"000110101",
  18240=>"100011000",
  18241=>"000011110",
  18242=>"010100100",
  18243=>"100011101",
  18244=>"001000000",
  18245=>"101011111",
  18246=>"100100010",
  18247=>"011111000",
  18248=>"111101110",
  18249=>"001100100",
  18250=>"010110001",
  18251=>"010011100",
  18252=>"101001010",
  18253=>"010001010",
  18254=>"101000000",
  18255=>"001001000",
  18256=>"010010110",
  18257=>"000100111",
  18258=>"111100101",
  18259=>"010111001",
  18260=>"011000011",
  18261=>"100000000",
  18262=>"011100100",
  18263=>"101000000",
  18264=>"111010111",
  18265=>"011100011",
  18266=>"111011100",
  18267=>"111111010",
  18268=>"100011101",
  18269=>"011101000",
  18270=>"010001011",
  18271=>"001111100",
  18272=>"010011110",
  18273=>"101111100",
  18274=>"010111011",
  18275=>"001010110",
  18276=>"111111110",
  18277=>"100101001",
  18278=>"100000110",
  18279=>"110001101",
  18280=>"011011001",
  18281=>"001100101",
  18282=>"000101001",
  18283=>"110011000",
  18284=>"111010000",
  18285=>"101001111",
  18286=>"111110101",
  18287=>"101100100",
  18288=>"111101111",
  18289=>"001001101",
  18290=>"111010100",
  18291=>"011010101",
  18292=>"000101000",
  18293=>"000110010",
  18294=>"011111000",
  18295=>"001010101",
  18296=>"111100011",
  18297=>"001111011",
  18298=>"101011000",
  18299=>"001010010",
  18300=>"110101011",
  18301=>"000110100",
  18302=>"001101010",
  18303=>"100010010",
  18304=>"101110100",
  18305=>"110000101",
  18306=>"011001000",
  18307=>"110110101",
  18308=>"110110010",
  18309=>"111110111",
  18310=>"110101011",
  18311=>"000001101",
  18312=>"101000111",
  18313=>"000100100",
  18314=>"100011001",
  18315=>"111010011",
  18316=>"010000111",
  18317=>"110000011",
  18318=>"001011100",
  18319=>"000010110",
  18320=>"111010110",
  18321=>"111001111",
  18322=>"011000110",
  18323=>"101100000",
  18324=>"011101000",
  18325=>"010101111",
  18326=>"000011101",
  18327=>"011111100",
  18328=>"011010000",
  18329=>"101101011",
  18330=>"101011010",
  18331=>"100011110",
  18332=>"001001000",
  18333=>"001010001",
  18334=>"001101100",
  18335=>"010100011",
  18336=>"011111100",
  18337=>"000001011",
  18338=>"010100110",
  18339=>"101000100",
  18340=>"111011010",
  18341=>"011101111",
  18342=>"111101010",
  18343=>"110101101",
  18344=>"010010001",
  18345=>"100100000",
  18346=>"110101100",
  18347=>"101000111",
  18348=>"111110000",
  18349=>"111100011",
  18350=>"010100011",
  18351=>"100110110",
  18352=>"011001100",
  18353=>"001000011",
  18354=>"100010010",
  18355=>"111111011",
  18356=>"111010100",
  18357=>"000001100",
  18358=>"101010110",
  18359=>"111111111",
  18360=>"111000110",
  18361=>"000101001",
  18362=>"000111101",
  18363=>"010101111",
  18364=>"111111001",
  18365=>"011101111",
  18366=>"011010100",
  18367=>"010010110",
  18368=>"111010000",
  18369=>"010111000",
  18370=>"111101110",
  18371=>"011010010",
  18372=>"111010110",
  18373=>"001110011",
  18374=>"011011100",
  18375=>"011101101",
  18376=>"001111001",
  18377=>"010010110",
  18378=>"010000010",
  18379=>"001011100",
  18380=>"101010101",
  18381=>"101111001",
  18382=>"010011010",
  18383=>"101101011",
  18384=>"101101111",
  18385=>"001100010",
  18386=>"001110110",
  18387=>"101010110",
  18388=>"100100001",
  18389=>"011011011",
  18390=>"101011011",
  18391=>"110110101",
  18392=>"011011010",
  18393=>"000111110",
  18394=>"010001010",
  18395=>"110000000",
  18396=>"101001100",
  18397=>"010100100",
  18398=>"010110000",
  18399=>"011011000",
  18400=>"110001111",
  18401=>"100011001",
  18402=>"111101000",
  18403=>"100000000",
  18404=>"101010001",
  18405=>"111001010",
  18406=>"000110010",
  18407=>"001111111",
  18408=>"100111011",
  18409=>"111111111",
  18410=>"011100011",
  18411=>"000001111",
  18412=>"001001000",
  18413=>"101100001",
  18414=>"110011101",
  18415=>"111001100",
  18416=>"110111101",
  18417=>"111010110",
  18418=>"011000101",
  18419=>"000101111",
  18420=>"001111000",
  18421=>"100100001",
  18422=>"101100100",
  18423=>"001010011",
  18424=>"000000000",
  18425=>"000000101",
  18426=>"100110100",
  18427=>"100111011",
  18428=>"001110010",
  18429=>"001101001",
  18430=>"100111001",
  18431=>"100001101",
  18432=>"100000001",
  18433=>"000010011",
  18434=>"001111010",
  18435=>"011111000",
  18436=>"000011001",
  18437=>"010011010",
  18438=>"110111111",
  18439=>"101100001",
  18440=>"101010110",
  18441=>"011011101",
  18442=>"011110111",
  18443=>"111001000",
  18444=>"110010001",
  18445=>"110011011",
  18446=>"101010100",
  18447=>"011101010",
  18448=>"000001001",
  18449=>"010001001",
  18450=>"100011010",
  18451=>"100101000",
  18452=>"011110101",
  18453=>"011001011",
  18454=>"110000101",
  18455=>"011011111",
  18456=>"101010001",
  18457=>"000101000",
  18458=>"011100100",
  18459=>"001010010",
  18460=>"000000001",
  18461=>"000010110",
  18462=>"111111111",
  18463=>"010000001",
  18464=>"100101010",
  18465=>"111100001",
  18466=>"001100000",
  18467=>"111110010",
  18468=>"110001100",
  18469=>"101101001",
  18470=>"110101001",
  18471=>"100010100",
  18472=>"001000100",
  18473=>"001000011",
  18474=>"001110100",
  18475=>"110001001",
  18476=>"100110111",
  18477=>"001000000",
  18478=>"010010100",
  18479=>"111110111",
  18480=>"110101000",
  18481=>"000100110",
  18482=>"000011001",
  18483=>"011010110",
  18484=>"101111100",
  18485=>"001000000",
  18486=>"011001100",
  18487=>"010000110",
  18488=>"010110110",
  18489=>"001011110",
  18490=>"110100001",
  18491=>"010000100",
  18492=>"010100000",
  18493=>"001011111",
  18494=>"111000011",
  18495=>"000100010",
  18496=>"101000011",
  18497=>"000000010",
  18498=>"000101011",
  18499=>"001100111",
  18500=>"110001100",
  18501=>"000100101",
  18502=>"001011000",
  18503=>"101011001",
  18504=>"001100100",
  18505=>"111000111",
  18506=>"101111110",
  18507=>"001101110",
  18508=>"100000101",
  18509=>"000111011",
  18510=>"001101000",
  18511=>"011010010",
  18512=>"011111010",
  18513=>"101100011",
  18514=>"101101110",
  18515=>"010100000",
  18516=>"111000010",
  18517=>"011111111",
  18518=>"000100111",
  18519=>"011000111",
  18520=>"110111101",
  18521=>"101101000",
  18522=>"001100101",
  18523=>"000100101",
  18524=>"110010101",
  18525=>"101111110",
  18526=>"110100010",
  18527=>"111101000",
  18528=>"101000000",
  18529=>"010001101",
  18530=>"001100101",
  18531=>"001000010",
  18532=>"100111000",
  18533=>"100101101",
  18534=>"110001011",
  18535=>"010101100",
  18536=>"100000000",
  18537=>"010010010",
  18538=>"011001110",
  18539=>"000001100",
  18540=>"101000101",
  18541=>"001110000",
  18542=>"110001110",
  18543=>"000111111",
  18544=>"110110000",
  18545=>"101000001",
  18546=>"010001101",
  18547=>"110111100",
  18548=>"110000111",
  18549=>"100000101",
  18550=>"011111101",
  18551=>"110101110",
  18552=>"000100010",
  18553=>"000101100",
  18554=>"100111000",
  18555=>"001100101",
  18556=>"000000101",
  18557=>"110100100",
  18558=>"110110101",
  18559=>"001100011",
  18560=>"001000110",
  18561=>"011111010",
  18562=>"101010000",
  18563=>"010001110",
  18564=>"010000101",
  18565=>"010101110",
  18566=>"101010111",
  18567=>"110110000",
  18568=>"000100101",
  18569=>"111111000",
  18570=>"010111001",
  18571=>"010010110",
  18572=>"010100011",
  18573=>"111011100",
  18574=>"011010000",
  18575=>"100101011",
  18576=>"000111101",
  18577=>"010101001",
  18578=>"110010001",
  18579=>"111100010",
  18580=>"000011101",
  18581=>"110110111",
  18582=>"101010111",
  18583=>"111100111",
  18584=>"101111100",
  18585=>"100000010",
  18586=>"101000011",
  18587=>"010111101",
  18588=>"001011100",
  18589=>"111100100",
  18590=>"110011110",
  18591=>"000000010",
  18592=>"001010100",
  18593=>"011010000",
  18594=>"001010011",
  18595=>"111001101",
  18596=>"010100001",
  18597=>"011110101",
  18598=>"101011011",
  18599=>"011101011",
  18600=>"010001001",
  18601=>"011100111",
  18602=>"011111111",
  18603=>"110101100",
  18604=>"111010111",
  18605=>"100101001",
  18606=>"011101111",
  18607=>"100011111",
  18608=>"100100000",
  18609=>"000111000",
  18610=>"111111111",
  18611=>"100010011",
  18612=>"111110001",
  18613=>"011110011",
  18614=>"000110001",
  18615=>"110110101",
  18616=>"110000000",
  18617=>"010101001",
  18618=>"000010111",
  18619=>"101101011",
  18620=>"101111001",
  18621=>"101000110",
  18622=>"100101011",
  18623=>"000110101",
  18624=>"010110101",
  18625=>"110111101",
  18626=>"111011010",
  18627=>"101100100",
  18628=>"100100001",
  18629=>"000100001",
  18630=>"101111101",
  18631=>"100010111",
  18632=>"111111100",
  18633=>"111101001",
  18634=>"100110100",
  18635=>"001000100",
  18636=>"101100110",
  18637=>"101001110",
  18638=>"111000000",
  18639=>"100111011",
  18640=>"111011111",
  18641=>"001001010",
  18642=>"010101100",
  18643=>"010011011",
  18644=>"101101100",
  18645=>"101111010",
  18646=>"111001000",
  18647=>"000001101",
  18648=>"111100100",
  18649=>"101010100",
  18650=>"110011011",
  18651=>"100010010",
  18652=>"111011011",
  18653=>"111011010",
  18654=>"101110100",
  18655=>"100100011",
  18656=>"101110101",
  18657=>"011101011",
  18658=>"111110001",
  18659=>"000101000",
  18660=>"111100010",
  18661=>"000110111",
  18662=>"110111010",
  18663=>"100000010",
  18664=>"000000111",
  18665=>"100110001",
  18666=>"100001001",
  18667=>"110011000",
  18668=>"010011111",
  18669=>"110110001",
  18670=>"011010111",
  18671=>"110000000",
  18672=>"001101111",
  18673=>"001011111",
  18674=>"111110000",
  18675=>"011010000",
  18676=>"010100101",
  18677=>"111111110",
  18678=>"010011000",
  18679=>"011110100",
  18680=>"011111000",
  18681=>"100101011",
  18682=>"000100000",
  18683=>"101100100",
  18684=>"011100000",
  18685=>"100111111",
  18686=>"001100000",
  18687=>"111001100",
  18688=>"000111111",
  18689=>"000100110",
  18690=>"101001000",
  18691=>"100100000",
  18692=>"100111100",
  18693=>"000000111",
  18694=>"010011001",
  18695=>"110101011",
  18696=>"000011011",
  18697=>"000000011",
  18698=>"000111110",
  18699=>"011010101",
  18700=>"001010110",
  18701=>"000000110",
  18702=>"001111110",
  18703=>"011111011",
  18704=>"110001100",
  18705=>"010001000",
  18706=>"110011110",
  18707=>"000101001",
  18708=>"000000011",
  18709=>"011000110",
  18710=>"000110111",
  18711=>"010010101",
  18712=>"010110101",
  18713=>"000011001",
  18714=>"110101111",
  18715=>"010011001",
  18716=>"110011100",
  18717=>"110011000",
  18718=>"001111010",
  18719=>"000110010",
  18720=>"111110111",
  18721=>"100101100",
  18722=>"000001100",
  18723=>"100110000",
  18724=>"000000111",
  18725=>"011110010",
  18726=>"101001011",
  18727=>"100101011",
  18728=>"101010001",
  18729=>"001111000",
  18730=>"001100011",
  18731=>"101110011",
  18732=>"101000100",
  18733=>"110111110",
  18734=>"001111111",
  18735=>"111101110",
  18736=>"010101001",
  18737=>"101111111",
  18738=>"100010101",
  18739=>"010101010",
  18740=>"011010101",
  18741=>"010110110",
  18742=>"110001011",
  18743=>"101001100",
  18744=>"001111010",
  18745=>"010001101",
  18746=>"011011010",
  18747=>"010100111",
  18748=>"110100101",
  18749=>"010100001",
  18750=>"011111101",
  18751=>"000000100",
  18752=>"011101011",
  18753=>"000010111",
  18754=>"011010111",
  18755=>"100001001",
  18756=>"111110111",
  18757=>"110110011",
  18758=>"001001010",
  18759=>"010100011",
  18760=>"110110011",
  18761=>"011100001",
  18762=>"010111010",
  18763=>"010100111",
  18764=>"101101001",
  18765=>"100010101",
  18766=>"001100001",
  18767=>"011001110",
  18768=>"110011110",
  18769=>"111101000",
  18770=>"001101011",
  18771=>"001011000",
  18772=>"000101011",
  18773=>"111111001",
  18774=>"110100000",
  18775=>"111110100",
  18776=>"110011111",
  18777=>"101001011",
  18778=>"100000000",
  18779=>"011101110",
  18780=>"110000101",
  18781=>"101111100",
  18782=>"100011100",
  18783=>"000011001",
  18784=>"001111000",
  18785=>"001000001",
  18786=>"010100100",
  18787=>"100000010",
  18788=>"000001111",
  18789=>"001100000",
  18790=>"101111011",
  18791=>"100110011",
  18792=>"111011110",
  18793=>"101011110",
  18794=>"100110111",
  18795=>"011101001",
  18796=>"001011100",
  18797=>"000110101",
  18798=>"100100000",
  18799=>"100001110",
  18800=>"100011001",
  18801=>"001000111",
  18802=>"110000101",
  18803=>"010001000",
  18804=>"011100001",
  18805=>"100100010",
  18806=>"101000111",
  18807=>"000001111",
  18808=>"000100010",
  18809=>"011111100",
  18810=>"010110100",
  18811=>"110000010",
  18812=>"000000001",
  18813=>"010111111",
  18814=>"001001101",
  18815=>"101011000",
  18816=>"000010001",
  18817=>"000000111",
  18818=>"000001001",
  18819=>"111011100",
  18820=>"011011111",
  18821=>"110100001",
  18822=>"010110111",
  18823=>"011000101",
  18824=>"001010101",
  18825=>"110111100",
  18826=>"100001111",
  18827=>"111111101",
  18828=>"000111100",
  18829=>"011101111",
  18830=>"100001101",
  18831=>"101010000",
  18832=>"100001100",
  18833=>"110111100",
  18834=>"111011010",
  18835=>"000011100",
  18836=>"110101100",
  18837=>"000110001",
  18838=>"000111001",
  18839=>"101100011",
  18840=>"110000001",
  18841=>"010011110",
  18842=>"000000000",
  18843=>"100000000",
  18844=>"111001011",
  18845=>"111000111",
  18846=>"110000000",
  18847=>"011100000",
  18848=>"010100011",
  18849=>"010100111",
  18850=>"000001000",
  18851=>"111001001",
  18852=>"101100111",
  18853=>"000010001",
  18854=>"010100011",
  18855=>"101101011",
  18856=>"001111110",
  18857=>"010101010",
  18858=>"000110100",
  18859=>"010010001",
  18860=>"101001001",
  18861=>"000100000",
  18862=>"010001011",
  18863=>"110110001",
  18864=>"111011000",
  18865=>"110101000",
  18866=>"001101110",
  18867=>"010111011",
  18868=>"000111110",
  18869=>"010111011",
  18870=>"101110010",
  18871=>"000110010",
  18872=>"001000100",
  18873=>"101100001",
  18874=>"100111110",
  18875=>"001010011",
  18876=>"110011111",
  18877=>"001110111",
  18878=>"001001010",
  18879=>"000001000",
  18880=>"110000100",
  18881=>"011011100",
  18882=>"000110100",
  18883=>"010100110",
  18884=>"011011111",
  18885=>"000101111",
  18886=>"111110001",
  18887=>"000100000",
  18888=>"011100111",
  18889=>"110001110",
  18890=>"011100111",
  18891=>"001101101",
  18892=>"001111111",
  18893=>"010111010",
  18894=>"001110100",
  18895=>"111111000",
  18896=>"100011001",
  18897=>"010011010",
  18898=>"010110000",
  18899=>"111001001",
  18900=>"000011001",
  18901=>"100010010",
  18902=>"111110111",
  18903=>"101011011",
  18904=>"011110111",
  18905=>"100101100",
  18906=>"110100001",
  18907=>"000100100",
  18908=>"111010011",
  18909=>"000110100",
  18910=>"010001111",
  18911=>"101101100",
  18912=>"011101001",
  18913=>"000000010",
  18914=>"101100100",
  18915=>"011001011",
  18916=>"010100001",
  18917=>"010000000",
  18918=>"011111001",
  18919=>"000000000",
  18920=>"011110001",
  18921=>"110001101",
  18922=>"000001100",
  18923=>"011111111",
  18924=>"110110110",
  18925=>"101011010",
  18926=>"111010110",
  18927=>"000000001",
  18928=>"010111001",
  18929=>"011110111",
  18930=>"101001001",
  18931=>"001111001",
  18932=>"111000111",
  18933=>"101100001",
  18934=>"110100010",
  18935=>"100001100",
  18936=>"000100000",
  18937=>"111110100",
  18938=>"100000111",
  18939=>"010000011",
  18940=>"100011100",
  18941=>"011000111",
  18942=>"001101000",
  18943=>"010011010",
  18944=>"110011100",
  18945=>"100000001",
  18946=>"100010100",
  18947=>"011010010",
  18948=>"000010101",
  18949=>"010001000",
  18950=>"111110101",
  18951=>"010011001",
  18952=>"111100101",
  18953=>"011101100",
  18954=>"000100010",
  18955=>"100001000",
  18956=>"110001000",
  18957=>"111011111",
  18958=>"010001110",
  18959=>"110110100",
  18960=>"001111001",
  18961=>"000111010",
  18962=>"110001101",
  18963=>"110001111",
  18964=>"101100001",
  18965=>"101000001",
  18966=>"011101101",
  18967=>"101011010",
  18968=>"110011101",
  18969=>"101111011",
  18970=>"111111001",
  18971=>"010100011",
  18972=>"101100110",
  18973=>"011010000",
  18974=>"111000111",
  18975=>"001000010",
  18976=>"111111000",
  18977=>"111101001",
  18978=>"001100110",
  18979=>"110111111",
  18980=>"100011100",
  18981=>"100010000",
  18982=>"011001100",
  18983=>"110100101",
  18984=>"111110001",
  18985=>"001001010",
  18986=>"100000001",
  18987=>"010101100",
  18988=>"001111110",
  18989=>"111000001",
  18990=>"011000001",
  18991=>"000100001",
  18992=>"000010001",
  18993=>"000010111",
  18994=>"001000000",
  18995=>"000001110",
  18996=>"110001101",
  18997=>"001110111",
  18998=>"001110001",
  18999=>"011000111",
  19000=>"110010001",
  19001=>"010100100",
  19002=>"101110111",
  19003=>"100101111",
  19004=>"011110100",
  19005=>"001100001",
  19006=>"101010101",
  19007=>"100101101",
  19008=>"101111000",
  19009=>"110111010",
  19010=>"110000000",
  19011=>"110010101",
  19012=>"110100101",
  19013=>"001110101",
  19014=>"111111100",
  19015=>"001010001",
  19016=>"101010110",
  19017=>"000111001",
  19018=>"100000111",
  19019=>"011011011",
  19020=>"111011111",
  19021=>"110110110",
  19022=>"110100000",
  19023=>"110010100",
  19024=>"111101111",
  19025=>"001001001",
  19026=>"010110100",
  19027=>"010100100",
  19028=>"100010001",
  19029=>"101011110",
  19030=>"101010010",
  19031=>"000000010",
  19032=>"111111100",
  19033=>"001000011",
  19034=>"111100111",
  19035=>"001000010",
  19036=>"110111100",
  19037=>"000001000",
  19038=>"111011000",
  19039=>"110101101",
  19040=>"110101111",
  19041=>"100010100",
  19042=>"100110100",
  19043=>"001000011",
  19044=>"111011110",
  19045=>"010001100",
  19046=>"101010100",
  19047=>"000101001",
  19048=>"001001100",
  19049=>"101111111",
  19050=>"111111111",
  19051=>"101101010",
  19052=>"111101001",
  19053=>"110001110",
  19054=>"100110001",
  19055=>"111110100",
  19056=>"010101010",
  19057=>"101000110",
  19058=>"001100011",
  19059=>"000011111",
  19060=>"010111101",
  19061=>"011001011",
  19062=>"101000111",
  19063=>"000110011",
  19064=>"100100010",
  19065=>"000110101",
  19066=>"100101001",
  19067=>"111001010",
  19068=>"100100100",
  19069=>"000101010",
  19070=>"000111000",
  19071=>"010100101",
  19072=>"100100101",
  19073=>"001001101",
  19074=>"011111111",
  19075=>"110000010",
  19076=>"101000101",
  19077=>"000011101",
  19078=>"100010110",
  19079=>"100011001",
  19080=>"010100001",
  19081=>"000000001",
  19082=>"011001111",
  19083=>"011010111",
  19084=>"011101000",
  19085=>"000110011",
  19086=>"011110100",
  19087=>"110010011",
  19088=>"011100010",
  19089=>"111000111",
  19090=>"001101110",
  19091=>"111000010",
  19092=>"101010000",
  19093=>"000100110",
  19094=>"001111011",
  19095=>"111011101",
  19096=>"101001001",
  19097=>"001101001",
  19098=>"000001001",
  19099=>"100000101",
  19100=>"110110011",
  19101=>"001100001",
  19102=>"011100100",
  19103=>"011000010",
  19104=>"111011011",
  19105=>"010000011",
  19106=>"010001101",
  19107=>"011010100",
  19108=>"001011001",
  19109=>"001101011",
  19110=>"110110010",
  19111=>"111111011",
  19112=>"111111010",
  19113=>"111011100",
  19114=>"010010100",
  19115=>"011010100",
  19116=>"101011000",
  19117=>"101100100",
  19118=>"101110011",
  19119=>"111011111",
  19120=>"110101101",
  19121=>"011000100",
  19122=>"010111011",
  19123=>"010001100",
  19124=>"010110100",
  19125=>"101001100",
  19126=>"011100001",
  19127=>"111110011",
  19128=>"000011000",
  19129=>"010001001",
  19130=>"100000101",
  19131=>"100111110",
  19132=>"101101111",
  19133=>"110111011",
  19134=>"000110010",
  19135=>"101111000",
  19136=>"101101110",
  19137=>"011001011",
  19138=>"000001110",
  19139=>"111011101",
  19140=>"111111001",
  19141=>"000000110",
  19142=>"011011110",
  19143=>"111110010",
  19144=>"100001000",
  19145=>"010111101",
  19146=>"001010101",
  19147=>"000000011",
  19148=>"111011100",
  19149=>"111001111",
  19150=>"010111011",
  19151=>"000000000",
  19152=>"111001001",
  19153=>"100101001",
  19154=>"100111000",
  19155=>"011111100",
  19156=>"001000000",
  19157=>"000011101",
  19158=>"010101111",
  19159=>"001011110",
  19160=>"000100011",
  19161=>"100100100",
  19162=>"011001010",
  19163=>"110010001",
  19164=>"000001110",
  19165=>"111001011",
  19166=>"010111111",
  19167=>"110111000",
  19168=>"011111000",
  19169=>"101100000",
  19170=>"011011001",
  19171=>"101101111",
  19172=>"001100001",
  19173=>"001000000",
  19174=>"100011011",
  19175=>"111000000",
  19176=>"111111000",
  19177=>"100100000",
  19178=>"110011000",
  19179=>"010100010",
  19180=>"100001010",
  19181=>"111010010",
  19182=>"000001110",
  19183=>"001010000",
  19184=>"010100101",
  19185=>"000000011",
  19186=>"011011111",
  19187=>"011010000",
  19188=>"011111000",
  19189=>"101001100",
  19190=>"100000101",
  19191=>"010101101",
  19192=>"101010010",
  19193=>"111100100",
  19194=>"000000010",
  19195=>"010111101",
  19196=>"101110101",
  19197=>"100001000",
  19198=>"010110000",
  19199=>"010110001",
  19200=>"100010010",
  19201=>"001000101",
  19202=>"110110111",
  19203=>"000110001",
  19204=>"111111000",
  19205=>"011110100",
  19206=>"011111111",
  19207=>"110110000",
  19208=>"100000101",
  19209=>"100101101",
  19210=>"010100001",
  19211=>"100000101",
  19212=>"000100001",
  19213=>"011100011",
  19214=>"001100010",
  19215=>"011010010",
  19216=>"110101010",
  19217=>"011000010",
  19218=>"111001010",
  19219=>"010010100",
  19220=>"100110110",
  19221=>"001111010",
  19222=>"111001000",
  19223=>"100100110",
  19224=>"000100111",
  19225=>"100110100",
  19226=>"010000010",
  19227=>"010111100",
  19228=>"101110011",
  19229=>"110011001",
  19230=>"101001010",
  19231=>"111001011",
  19232=>"011010110",
  19233=>"001101101",
  19234=>"001000110",
  19235=>"011100111",
  19236=>"111110010",
  19237=>"100101011",
  19238=>"100111111",
  19239=>"100110100",
  19240=>"110111100",
  19241=>"010001100",
  19242=>"010010110",
  19243=>"011111100",
  19244=>"100100111",
  19245=>"111000011",
  19246=>"100010101",
  19247=>"010000100",
  19248=>"100110010",
  19249=>"101010111",
  19250=>"111111000",
  19251=>"100001010",
  19252=>"010100111",
  19253=>"101110100",
  19254=>"111101100",
  19255=>"111100101",
  19256=>"110110000",
  19257=>"110101010",
  19258=>"110000010",
  19259=>"110000101",
  19260=>"010000101",
  19261=>"010010100",
  19262=>"100000000",
  19263=>"000001001",
  19264=>"011000110",
  19265=>"111000111",
  19266=>"111100000",
  19267=>"110100100",
  19268=>"011010011",
  19269=>"111010011",
  19270=>"010011100",
  19271=>"010010001",
  19272=>"110110010",
  19273=>"001000000",
  19274=>"011001100",
  19275=>"111000110",
  19276=>"100010101",
  19277=>"110111011",
  19278=>"110001100",
  19279=>"010010111",
  19280=>"110100111",
  19281=>"100101001",
  19282=>"111001011",
  19283=>"101010011",
  19284=>"101001001",
  19285=>"001101101",
  19286=>"101000110",
  19287=>"000100001",
  19288=>"010010010",
  19289=>"100111010",
  19290=>"110000110",
  19291=>"011010011",
  19292=>"000100001",
  19293=>"111001011",
  19294=>"001110011",
  19295=>"000011001",
  19296=>"111000100",
  19297=>"011111100",
  19298=>"000000100",
  19299=>"100001011",
  19300=>"001100001",
  19301=>"100011111",
  19302=>"011000011",
  19303=>"010111110",
  19304=>"111010010",
  19305=>"010011110",
  19306=>"001100000",
  19307=>"101011000",
  19308=>"100101101",
  19309=>"101101100",
  19310=>"001111101",
  19311=>"001110011",
  19312=>"010101101",
  19313=>"000101000",
  19314=>"111000100",
  19315=>"001110101",
  19316=>"111001100",
  19317=>"010110010",
  19318=>"111111010",
  19319=>"111000000",
  19320=>"111100111",
  19321=>"001110111",
  19322=>"101110100",
  19323=>"101001001",
  19324=>"000011001",
  19325=>"111001101",
  19326=>"011110000",
  19327=>"011010111",
  19328=>"101111100",
  19329=>"101110111",
  19330=>"100000000",
  19331=>"000111111",
  19332=>"011111001",
  19333=>"010011001",
  19334=>"100010010",
  19335=>"101010101",
  19336=>"000100011",
  19337=>"100111010",
  19338=>"110110110",
  19339=>"011010001",
  19340=>"111011110",
  19341=>"010010011",
  19342=>"001100001",
  19343=>"100101011",
  19344=>"000100100",
  19345=>"010010100",
  19346=>"111110100",
  19347=>"110010001",
  19348=>"001101000",
  19349=>"001101111",
  19350=>"001100100",
  19351=>"001111111",
  19352=>"010110110",
  19353=>"110011001",
  19354=>"000101011",
  19355=>"100111111",
  19356=>"101001000",
  19357=>"011001000",
  19358=>"100101110",
  19359=>"111010000",
  19360=>"111010011",
  19361=>"111000000",
  19362=>"000000001",
  19363=>"011000011",
  19364=>"110010101",
  19365=>"010110101",
  19366=>"100111101",
  19367=>"100100000",
  19368=>"101101110",
  19369=>"011001001",
  19370=>"001100010",
  19371=>"001101010",
  19372=>"111001100",
  19373=>"110001010",
  19374=>"011000100",
  19375=>"100101101",
  19376=>"010110110",
  19377=>"001101110",
  19378=>"100101111",
  19379=>"111101110",
  19380=>"001000010",
  19381=>"000000100",
  19382=>"001110100",
  19383=>"001000010",
  19384=>"000101100",
  19385=>"100000100",
  19386=>"010010010",
  19387=>"101001010",
  19388=>"000001110",
  19389=>"110110001",
  19390=>"101101111",
  19391=>"111110101",
  19392=>"011000101",
  19393=>"001001001",
  19394=>"000011110",
  19395=>"001000100",
  19396=>"111100100",
  19397=>"010111000",
  19398=>"100000110",
  19399=>"100100000",
  19400=>"011010110",
  19401=>"000101001",
  19402=>"000111001",
  19403=>"001111000",
  19404=>"100110010",
  19405=>"111001111",
  19406=>"101010000",
  19407=>"110000000",
  19408=>"111000110",
  19409=>"110000000",
  19410=>"101110000",
  19411=>"000001000",
  19412=>"001001001",
  19413=>"101010110",
  19414=>"110001111",
  19415=>"000101111",
  19416=>"000111100",
  19417=>"010010110",
  19418=>"111101110",
  19419=>"011011111",
  19420=>"111101000",
  19421=>"001110000",
  19422=>"100111001",
  19423=>"011101101",
  19424=>"100000110",
  19425=>"001111110",
  19426=>"100100001",
  19427=>"001111101",
  19428=>"001101011",
  19429=>"010111001",
  19430=>"000111100",
  19431=>"001111100",
  19432=>"011011000",
  19433=>"110111010",
  19434=>"101101001",
  19435=>"010001011",
  19436=>"101011011",
  19437=>"011101000",
  19438=>"000110110",
  19439=>"100111101",
  19440=>"110110111",
  19441=>"010101000",
  19442=>"100110000",
  19443=>"011100011",
  19444=>"101111101",
  19445=>"110100000",
  19446=>"111001100",
  19447=>"110000100",
  19448=>"110001000",
  19449=>"001010101",
  19450=>"101100001",
  19451=>"101110001",
  19452=>"000011101",
  19453=>"001010110",
  19454=>"111010100",
  19455=>"000111010",
  19456=>"110100100",
  19457=>"111011001",
  19458=>"011000111",
  19459=>"111100001",
  19460=>"010110111",
  19461=>"001001111",
  19462=>"001100000",
  19463=>"100110101",
  19464=>"111101100",
  19465=>"001100010",
  19466=>"000000110",
  19467=>"010000111",
  19468=>"101010111",
  19469=>"000001011",
  19470=>"011001100",
  19471=>"001101100",
  19472=>"101100001",
  19473=>"001001111",
  19474=>"110010100",
  19475=>"011101001",
  19476=>"101010000",
  19477=>"001101100",
  19478=>"000100000",
  19479=>"111010000",
  19480=>"110001101",
  19481=>"000000101",
  19482=>"001111001",
  19483=>"000000000",
  19484=>"100111100",
  19485=>"100000010",
  19486=>"100111111",
  19487=>"011010100",
  19488=>"101111101",
  19489=>"001101001",
  19490=>"111101111",
  19491=>"100110001",
  19492=>"110101011",
  19493=>"111111011",
  19494=>"110011010",
  19495=>"101010001",
  19496=>"011001011",
  19497=>"111101001",
  19498=>"111101101",
  19499=>"010001101",
  19500=>"000010000",
  19501=>"111111101",
  19502=>"000000010",
  19503=>"100110110",
  19504=>"001101101",
  19505=>"011000010",
  19506=>"110010010",
  19507=>"100011001",
  19508=>"111111111",
  19509=>"110000001",
  19510=>"111100011",
  19511=>"001000010",
  19512=>"111101000",
  19513=>"000001100",
  19514=>"001110110",
  19515=>"000101001",
  19516=>"010011101",
  19517=>"011001110",
  19518=>"100010110",
  19519=>"100101010",
  19520=>"001111011",
  19521=>"000010010",
  19522=>"011100100",
  19523=>"100001000",
  19524=>"111111000",
  19525=>"000101101",
  19526=>"010100011",
  19527=>"110110101",
  19528=>"010101011",
  19529=>"100111010",
  19530=>"101011100",
  19531=>"100110000",
  19532=>"000001001",
  19533=>"001111001",
  19534=>"110011000",
  19535=>"101010111",
  19536=>"111001011",
  19537=>"001111010",
  19538=>"101001111",
  19539=>"000010000",
  19540=>"000000100",
  19541=>"100110011",
  19542=>"010011100",
  19543=>"111011000",
  19544=>"010010000",
  19545=>"011000011",
  19546=>"000010111",
  19547=>"111001010",
  19548=>"101001101",
  19549=>"111111100",
  19550=>"000111110",
  19551=>"101011010",
  19552=>"100100011",
  19553=>"111011011",
  19554=>"001010011",
  19555=>"101001000",
  19556=>"001001100",
  19557=>"101100111",
  19558=>"111101000",
  19559=>"110110000",
  19560=>"101001110",
  19561=>"001010001",
  19562=>"101010001",
  19563=>"001100100",
  19564=>"101110100",
  19565=>"001101001",
  19566=>"101000010",
  19567=>"001010011",
  19568=>"001001101",
  19569=>"011001111",
  19570=>"110000110",
  19571=>"111011000",
  19572=>"000001000",
  19573=>"101100101",
  19574=>"000001011",
  19575=>"011011110",
  19576=>"111111101",
  19577=>"000010010",
  19578=>"101101111",
  19579=>"100110011",
  19580=>"010000000",
  19581=>"100000110",
  19582=>"001000100",
  19583=>"111111111",
  19584=>"011000001",
  19585=>"001110111",
  19586=>"110110111",
  19587=>"001000100",
  19588=>"011101110",
  19589=>"110000001",
  19590=>"001100111",
  19591=>"010010100",
  19592=>"111100011",
  19593=>"011011010",
  19594=>"101010111",
  19595=>"110111101",
  19596=>"001100000",
  19597=>"110101111",
  19598=>"100100111",
  19599=>"110001010",
  19600=>"111100010",
  19601=>"100001111",
  19602=>"111000110",
  19603=>"000111010",
  19604=>"111001110",
  19605=>"001111100",
  19606=>"011101111",
  19607=>"100100001",
  19608=>"100100110",
  19609=>"010110111",
  19610=>"100000100",
  19611=>"111001101",
  19612=>"111100010",
  19613=>"111000000",
  19614=>"110100111",
  19615=>"001101010",
  19616=>"000111011",
  19617=>"010101000",
  19618=>"000110100",
  19619=>"100110010",
  19620=>"101101100",
  19621=>"101101100",
  19622=>"000010110",
  19623=>"111011110",
  19624=>"100010111",
  19625=>"111111001",
  19626=>"110110111",
  19627=>"110111110",
  19628=>"000111011",
  19629=>"111000011",
  19630=>"101110011",
  19631=>"110011100",
  19632=>"011111010",
  19633=>"000110000",
  19634=>"000001111",
  19635=>"001000000",
  19636=>"010011100",
  19637=>"100010010",
  19638=>"111111101",
  19639=>"001011000",
  19640=>"110011010",
  19641=>"100001000",
  19642=>"011000000",
  19643=>"011000101",
  19644=>"001111110",
  19645=>"111011101",
  19646=>"001101110",
  19647=>"001000011",
  19648=>"010001000",
  19649=>"101101010",
  19650=>"010010011",
  19651=>"111010010",
  19652=>"011001111",
  19653=>"111100000",
  19654=>"100100100",
  19655=>"100011100",
  19656=>"011011011",
  19657=>"010111101",
  19658=>"001011000",
  19659=>"100110111",
  19660=>"111100000",
  19661=>"001001001",
  19662=>"110011010",
  19663=>"110100000",
  19664=>"111011011",
  19665=>"000000100",
  19666=>"011010111",
  19667=>"110011110",
  19668=>"010000100",
  19669=>"011011100",
  19670=>"001001000",
  19671=>"011101110",
  19672=>"011110010",
  19673=>"110001001",
  19674=>"101001000",
  19675=>"011000110",
  19676=>"011111101",
  19677=>"110000011",
  19678=>"111011101",
  19679=>"010100000",
  19680=>"011001100",
  19681=>"111111001",
  19682=>"101111101",
  19683=>"000010010",
  19684=>"001100011",
  19685=>"011010101",
  19686=>"101110111",
  19687=>"000011111",
  19688=>"001111010",
  19689=>"111110100",
  19690=>"100100001",
  19691=>"000001000",
  19692=>"011000001",
  19693=>"110110101",
  19694=>"001110001",
  19695=>"011111000",
  19696=>"110100101",
  19697=>"111000000",
  19698=>"000010010",
  19699=>"101010001",
  19700=>"100100000",
  19701=>"111001011",
  19702=>"010110010",
  19703=>"100110100",
  19704=>"111010001",
  19705=>"001111000",
  19706=>"100001001",
  19707=>"110010011",
  19708=>"000000001",
  19709=>"001110001",
  19710=>"011001100",
  19711=>"000010111",
  19712=>"101011001",
  19713=>"110001001",
  19714=>"000110100",
  19715=>"010110000",
  19716=>"001000000",
  19717=>"001101101",
  19718=>"001000010",
  19719=>"100011111",
  19720=>"010011001",
  19721=>"011101111",
  19722=>"100000000",
  19723=>"111001000",
  19724=>"111110110",
  19725=>"101101000",
  19726=>"100100100",
  19727=>"011010110",
  19728=>"001011010",
  19729=>"010001100",
  19730=>"111011111",
  19731=>"000011101",
  19732=>"110100110",
  19733=>"000000000",
  19734=>"011100001",
  19735=>"100011110",
  19736=>"101000010",
  19737=>"000101001",
  19738=>"001001000",
  19739=>"010000111",
  19740=>"011000010",
  19741=>"100001111",
  19742=>"110011110",
  19743=>"000011101",
  19744=>"001011101",
  19745=>"000011100",
  19746=>"010111010",
  19747=>"111011101",
  19748=>"000010101",
  19749=>"110001001",
  19750=>"100000000",
  19751=>"000111101",
  19752=>"001111010",
  19753=>"100101011",
  19754=>"011010100",
  19755=>"100000000",
  19756=>"101100010",
  19757=>"011100111",
  19758=>"000000100",
  19759=>"010001000",
  19760=>"000000110",
  19761=>"110101011",
  19762=>"110111010",
  19763=>"110011010",
  19764=>"010110110",
  19765=>"010101011",
  19766=>"010111011",
  19767=>"001000010",
  19768=>"001100110",
  19769=>"110000111",
  19770=>"101001100",
  19771=>"010000010",
  19772=>"011101111",
  19773=>"001111110",
  19774=>"111011111",
  19775=>"100010111",
  19776=>"011010011",
  19777=>"011011010",
  19778=>"101100000",
  19779=>"000011101",
  19780=>"011010001",
  19781=>"100110111",
  19782=>"010001010",
  19783=>"000010111",
  19784=>"011100001",
  19785=>"100000111",
  19786=>"100001101",
  19787=>"101100001",
  19788=>"000000101",
  19789=>"101001001",
  19790=>"001111000",
  19791=>"110001101",
  19792=>"010000010",
  19793=>"001110110",
  19794=>"111101010",
  19795=>"101110110",
  19796=>"110000100",
  19797=>"011101111",
  19798=>"000010101",
  19799=>"111100100",
  19800=>"001100101",
  19801=>"001001110",
  19802=>"110001110",
  19803=>"011100011",
  19804=>"101001100",
  19805=>"000010100",
  19806=>"110110110",
  19807=>"111000001",
  19808=>"010110001",
  19809=>"011101001",
  19810=>"110101110",
  19811=>"000000110",
  19812=>"100000001",
  19813=>"010000010",
  19814=>"010011110",
  19815=>"001000110",
  19816=>"001100010",
  19817=>"111101000",
  19818=>"001001010",
  19819=>"001101001",
  19820=>"010000010",
  19821=>"111110011",
  19822=>"010000111",
  19823=>"101000001",
  19824=>"110011111",
  19825=>"011111111",
  19826=>"111001010",
  19827=>"101000101",
  19828=>"001001111",
  19829=>"000000001",
  19830=>"011010010",
  19831=>"100110010",
  19832=>"010100010",
  19833=>"010001111",
  19834=>"110011000",
  19835=>"100001000",
  19836=>"000100110",
  19837=>"110011010",
  19838=>"001111100",
  19839=>"101111000",
  19840=>"101001000",
  19841=>"001010110",
  19842=>"100000110",
  19843=>"011101110",
  19844=>"010011001",
  19845=>"000100100",
  19846=>"001011100",
  19847=>"110001011",
  19848=>"000110001",
  19849=>"011000001",
  19850=>"000100100",
  19851=>"010110110",
  19852=>"010101111",
  19853=>"111001111",
  19854=>"110101111",
  19855=>"010101011",
  19856=>"010100111",
  19857=>"001101001",
  19858=>"101010111",
  19859=>"110000101",
  19860=>"000001101",
  19861=>"001100010",
  19862=>"100111101",
  19863=>"100010010",
  19864=>"011010001",
  19865=>"100101101",
  19866=>"100110100",
  19867=>"111011010",
  19868=>"100010110",
  19869=>"011111011",
  19870=>"011101110",
  19871=>"010110111",
  19872=>"101001101",
  19873=>"001110111",
  19874=>"110100100",
  19875=>"000001100",
  19876=>"011010100",
  19877=>"001101111",
  19878=>"010111001",
  19879=>"011001000",
  19880=>"010111011",
  19881=>"101010111",
  19882=>"011100000",
  19883=>"010100010",
  19884=>"010110100",
  19885=>"010110000",
  19886=>"010010100",
  19887=>"111110110",
  19888=>"000101110",
  19889=>"101111100",
  19890=>"100111100",
  19891=>"001111011",
  19892=>"111001101",
  19893=>"010010100",
  19894=>"011001000",
  19895=>"100101001",
  19896=>"011001010",
  19897=>"100110000",
  19898=>"100001111",
  19899=>"100011010",
  19900=>"110011001",
  19901=>"111110000",
  19902=>"101101110",
  19903=>"111011011",
  19904=>"000011011",
  19905=>"111110111",
  19906=>"100101111",
  19907=>"110000110",
  19908=>"101111110",
  19909=>"101100011",
  19910=>"111001010",
  19911=>"111111001",
  19912=>"110000001",
  19913=>"000101100",
  19914=>"011111010",
  19915=>"001100100",
  19916=>"101111001",
  19917=>"100100101",
  19918=>"111011111",
  19919=>"100010110",
  19920=>"111101100",
  19921=>"101111011",
  19922=>"001001111",
  19923=>"010001100",
  19924=>"110010110",
  19925=>"001000010",
  19926=>"000011000",
  19927=>"000010111",
  19928=>"001011000",
  19929=>"111011000",
  19930=>"011001001",
  19931=>"100111001",
  19932=>"001001010",
  19933=>"110001110",
  19934=>"100011100",
  19935=>"100011100",
  19936=>"101101111",
  19937=>"100110001",
  19938=>"110111110",
  19939=>"000010111",
  19940=>"110000000",
  19941=>"111100101",
  19942=>"011111000",
  19943=>"101110110",
  19944=>"000100110",
  19945=>"010000111",
  19946=>"000110001",
  19947=>"111111100",
  19948=>"101001111",
  19949=>"111101111",
  19950=>"001111011",
  19951=>"000100101",
  19952=>"001000000",
  19953=>"001100101",
  19954=>"110001101",
  19955=>"110001101",
  19956=>"011001001",
  19957=>"010111110",
  19958=>"000011001",
  19959=>"000101110",
  19960=>"001011110",
  19961=>"000110110",
  19962=>"110100001",
  19963=>"111001111",
  19964=>"000000010",
  19965=>"110111100",
  19966=>"011101011",
  19967=>"010111111",
  19968=>"010000100",
  19969=>"001110011",
  19970=>"101110010",
  19971=>"111010101",
  19972=>"010111000",
  19973=>"111111000",
  19974=>"000010110",
  19975=>"010100011",
  19976=>"100111110",
  19977=>"011101111",
  19978=>"100110010",
  19979=>"111001111",
  19980=>"100011001",
  19981=>"101010011",
  19982=>"101010010",
  19983=>"010000000",
  19984=>"111101011",
  19985=>"010001111",
  19986=>"100010010",
  19987=>"111100101",
  19988=>"110000011",
  19989=>"101000001",
  19990=>"001010010",
  19991=>"110101010",
  19992=>"011011101",
  19993=>"100100010",
  19994=>"010111101",
  19995=>"100110111",
  19996=>"001101010",
  19997=>"001001110",
  19998=>"000011111",
  19999=>"100000001",
  20000=>"101011001",
  20001=>"110010010",
  20002=>"001111100",
  20003=>"000001100",
  20004=>"010101010",
  20005=>"000101011",
  20006=>"001010110",
  20007=>"001010101",
  20008=>"000111011",
  20009=>"010101101",
  20010=>"101010111",
  20011=>"010101011",
  20012=>"010110000",
  20013=>"010111110",
  20014=>"010111011",
  20015=>"101000110",
  20016=>"110110011",
  20017=>"111010000",
  20018=>"001101110",
  20019=>"101101111",
  20020=>"111010011",
  20021=>"000111101",
  20022=>"110111111",
  20023=>"000000010",
  20024=>"010110101",
  20025=>"111011101",
  20026=>"001111000",
  20027=>"111001000",
  20028=>"111101010",
  20029=>"001001101",
  20030=>"011101111",
  20031=>"010100000",
  20032=>"101010110",
  20033=>"000100111",
  20034=>"000011101",
  20035=>"111010110",
  20036=>"001010111",
  20037=>"110001000",
  20038=>"001110100",
  20039=>"100100110",
  20040=>"000000010",
  20041=>"111001111",
  20042=>"101111111",
  20043=>"011100100",
  20044=>"101001110",
  20045=>"111001101",
  20046=>"110010110",
  20047=>"101000001",
  20048=>"111001100",
  20049=>"010101011",
  20050=>"110111110",
  20051=>"100100000",
  20052=>"011001000",
  20053=>"001011100",
  20054=>"000110110",
  20055=>"000100010",
  20056=>"001011001",
  20057=>"110010000",
  20058=>"101001110",
  20059=>"101001110",
  20060=>"010010001",
  20061=>"110001111",
  20062=>"001010000",
  20063=>"000001111",
  20064=>"001001001",
  20065=>"011101111",
  20066=>"101000011",
  20067=>"010010000",
  20068=>"110010011",
  20069=>"000001011",
  20070=>"010100100",
  20071=>"011110101",
  20072=>"001100001",
  20073=>"110010110",
  20074=>"111000111",
  20075=>"000001000",
  20076=>"000111001",
  20077=>"001001001",
  20078=>"000000001",
  20079=>"011010111",
  20080=>"110111101",
  20081=>"111110010",
  20082=>"100101001",
  20083=>"100111110",
  20084=>"001001100",
  20085=>"000000110",
  20086=>"100010100",
  20087=>"001101010",
  20088=>"010111111",
  20089=>"011101110",
  20090=>"100010100",
  20091=>"110001111",
  20092=>"001000000",
  20093=>"100001000",
  20094=>"101011111",
  20095=>"000010110",
  20096=>"110100111",
  20097=>"100100100",
  20098=>"011101101",
  20099=>"010000101",
  20100=>"100111011",
  20101=>"100101001",
  20102=>"101001110",
  20103=>"011111001",
  20104=>"100100100",
  20105=>"110000010",
  20106=>"111111101",
  20107=>"001100100",
  20108=>"010001110",
  20109=>"111010101",
  20110=>"100101101",
  20111=>"000101111",
  20112=>"100100101",
  20113=>"001010010",
  20114=>"111111100",
  20115=>"110010111",
  20116=>"101100100",
  20117=>"111011000",
  20118=>"100000000",
  20119=>"000001010",
  20120=>"011000001",
  20121=>"000000110",
  20122=>"101110101",
  20123=>"001110000",
  20124=>"011011010",
  20125=>"101101111",
  20126=>"000111011",
  20127=>"011001000",
  20128=>"111100100",
  20129=>"000000111",
  20130=>"110010000",
  20131=>"011001011",
  20132=>"010000001",
  20133=>"000010100",
  20134=>"100011010",
  20135=>"100101001",
  20136=>"010110000",
  20137=>"010100011",
  20138=>"001011010",
  20139=>"011000110",
  20140=>"100011110",
  20141=>"111111001",
  20142=>"111110000",
  20143=>"100001101",
  20144=>"110011011",
  20145=>"000101101",
  20146=>"111010111",
  20147=>"101101100",
  20148=>"100000001",
  20149=>"011000111",
  20150=>"000110100",
  20151=>"011101110",
  20152=>"000101000",
  20153=>"101110100",
  20154=>"111011001",
  20155=>"100100001",
  20156=>"110100101",
  20157=>"011011000",
  20158=>"101101101",
  20159=>"011011001",
  20160=>"000000101",
  20161=>"111010100",
  20162=>"001011011",
  20163=>"111101100",
  20164=>"110010011",
  20165=>"001011000",
  20166=>"001100110",
  20167=>"000100011",
  20168=>"001011111",
  20169=>"100110001",
  20170=>"100001010",
  20171=>"100100001",
  20172=>"001010011",
  20173=>"000011001",
  20174=>"011101100",
  20175=>"100111010",
  20176=>"110101010",
  20177=>"110111010",
  20178=>"100101000",
  20179=>"111011101",
  20180=>"101100110",
  20181=>"110111101",
  20182=>"011111100",
  20183=>"110010001",
  20184=>"100010011",
  20185=>"110111111",
  20186=>"111101000",
  20187=>"100011001",
  20188=>"101011001",
  20189=>"000000000",
  20190=>"110001101",
  20191=>"111110011",
  20192=>"010111100",
  20193=>"101000100",
  20194=>"110000011",
  20195=>"001001011",
  20196=>"101011000",
  20197=>"100001110",
  20198=>"100000100",
  20199=>"110001100",
  20200=>"111111000",
  20201=>"010001011",
  20202=>"100010111",
  20203=>"001001000",
  20204=>"001000111",
  20205=>"110001000",
  20206=>"110011000",
  20207=>"100000010",
  20208=>"110000101",
  20209=>"101000010",
  20210=>"110011010",
  20211=>"110110110",
  20212=>"001100111",
  20213=>"011111010",
  20214=>"110010111",
  20215=>"000111111",
  20216=>"111010001",
  20217=>"100000010",
  20218=>"001111011",
  20219=>"100101011",
  20220=>"010010001",
  20221=>"000010100",
  20222=>"111000101",
  20223=>"110111101",
  20224=>"111110011",
  20225=>"111101111",
  20226=>"000111010",
  20227=>"000000111",
  20228=>"111000000",
  20229=>"000000011",
  20230=>"001010000",
  20231=>"101100001",
  20232=>"100001101",
  20233=>"000110101",
  20234=>"111100100",
  20235=>"010000010",
  20236=>"100001111",
  20237=>"101100110",
  20238=>"100000001",
  20239=>"011110010",
  20240=>"100010000",
  20241=>"110110101",
  20242=>"110110011",
  20243=>"110101111",
  20244=>"000110101",
  20245=>"000001010",
  20246=>"100011111",
  20247=>"010010101",
  20248=>"100100100",
  20249=>"010100001",
  20250=>"110001011",
  20251=>"111011110",
  20252=>"111001000",
  20253=>"101001111",
  20254=>"011011100",
  20255=>"111110100",
  20256=>"100100100",
  20257=>"111001111",
  20258=>"111101101",
  20259=>"111111010",
  20260=>"100010101",
  20261=>"101010011",
  20262=>"101011110",
  20263=>"111101110",
  20264=>"100100101",
  20265=>"111011011",
  20266=>"110000001",
  20267=>"000100001",
  20268=>"010101001",
  20269=>"101001000",
  20270=>"100011111",
  20271=>"110111110",
  20272=>"000011101",
  20273=>"110110010",
  20274=>"101100110",
  20275=>"100010000",
  20276=>"000111010",
  20277=>"000110011",
  20278=>"100101110",
  20279=>"011111011",
  20280=>"001011101",
  20281=>"010101000",
  20282=>"001111001",
  20283=>"001101110",
  20284=>"111100010",
  20285=>"000111100",
  20286=>"111010000",
  20287=>"000111010",
  20288=>"011111011",
  20289=>"000101111",
  20290=>"000101000",
  20291=>"100111100",
  20292=>"101010100",
  20293=>"010000101",
  20294=>"000111110",
  20295=>"100001000",
  20296=>"001110110",
  20297=>"000011010",
  20298=>"010001110",
  20299=>"111001110",
  20300=>"011100000",
  20301=>"001001011",
  20302=>"011000110",
  20303=>"000110000",
  20304=>"110101111",
  20305=>"110001010",
  20306=>"011100010",
  20307=>"000000000",
  20308=>"010100100",
  20309=>"100111101",
  20310=>"001001000",
  20311=>"110110011",
  20312=>"110101000",
  20313=>"111110100",
  20314=>"110111101",
  20315=>"110001100",
  20316=>"100101001",
  20317=>"011101011",
  20318=>"011100001",
  20319=>"001011011",
  20320=>"111000001",
  20321=>"010100010",
  20322=>"001100001",
  20323=>"100000111",
  20324=>"000101011",
  20325=>"000101101",
  20326=>"110111011",
  20327=>"011011010",
  20328=>"101011111",
  20329=>"000001000",
  20330=>"110011011",
  20331=>"111101101",
  20332=>"100111011",
  20333=>"110001011",
  20334=>"010110011",
  20335=>"110101001",
  20336=>"100000101",
  20337=>"001110010",
  20338=>"001110110",
  20339=>"111001011",
  20340=>"100001000",
  20341=>"110100001",
  20342=>"100110101",
  20343=>"000000110",
  20344=>"011101110",
  20345=>"101110110",
  20346=>"100111001",
  20347=>"110010101",
  20348=>"100001010",
  20349=>"010011000",
  20350=>"110101001",
  20351=>"000100000",
  20352=>"100001010",
  20353=>"111110100",
  20354=>"101001001",
  20355=>"010100111",
  20356=>"011101000",
  20357=>"000011000",
  20358=>"101110001",
  20359=>"010001100",
  20360=>"011011101",
  20361=>"111110101",
  20362=>"000111110",
  20363=>"000111011",
  20364=>"010101100",
  20365=>"110111111",
  20366=>"100011000",
  20367=>"000001101",
  20368=>"000101001",
  20369=>"010110011",
  20370=>"000011000",
  20371=>"000001010",
  20372=>"010100011",
  20373=>"001000101",
  20374=>"010001101",
  20375=>"111111011",
  20376=>"000011101",
  20377=>"110111100",
  20378=>"101000001",
  20379=>"100101001",
  20380=>"101000110",
  20381=>"010111101",
  20382=>"001101100",
  20383=>"101000110",
  20384=>"000011001",
  20385=>"101000001",
  20386=>"000011010",
  20387=>"111001100",
  20388=>"100111111",
  20389=>"111011111",
  20390=>"001111001",
  20391=>"111110010",
  20392=>"111110011",
  20393=>"111011101",
  20394=>"001010010",
  20395=>"001010101",
  20396=>"110001100",
  20397=>"100011010",
  20398=>"100100010",
  20399=>"111101111",
  20400=>"110010111",
  20401=>"001111010",
  20402=>"001000001",
  20403=>"111101000",
  20404=>"000001000",
  20405=>"100110111",
  20406=>"000011010",
  20407=>"111000011",
  20408=>"111011001",
  20409=>"100000000",
  20410=>"010001010",
  20411=>"001110011",
  20412=>"000111000",
  20413=>"101010001",
  20414=>"001111111",
  20415=>"100111000",
  20416=>"101000101",
  20417=>"010001110",
  20418=>"000100101",
  20419=>"011010010",
  20420=>"000111001",
  20421=>"000001110",
  20422=>"111110011",
  20423=>"110101010",
  20424=>"101001100",
  20425=>"100110000",
  20426=>"110000100",
  20427=>"100100111",
  20428=>"111111010",
  20429=>"011010111",
  20430=>"110000000",
  20431=>"110100110",
  20432=>"100100111",
  20433=>"110010010",
  20434=>"110000010",
  20435=>"010100101",
  20436=>"111111000",
  20437=>"000110111",
  20438=>"101000001",
  20439=>"110101110",
  20440=>"111001101",
  20441=>"101101000",
  20442=>"111000111",
  20443=>"010010100",
  20444=>"101100110",
  20445=>"101000000",
  20446=>"010010100",
  20447=>"110011001",
  20448=>"110011100",
  20449=>"001011010",
  20450=>"111101010",
  20451=>"000110010",
  20452=>"111011110",
  20453=>"010111001",
  20454=>"111001010",
  20455=>"010011110",
  20456=>"000011000",
  20457=>"111111011",
  20458=>"111000110",
  20459=>"001110011",
  20460=>"000011011",
  20461=>"010110001",
  20462=>"010101001",
  20463=>"000101101",
  20464=>"100001101",
  20465=>"101001110",
  20466=>"000001110",
  20467=>"110001110",
  20468=>"100011011",
  20469=>"000111110",
  20470=>"001110001",
  20471=>"101111111",
  20472=>"010011000",
  20473=>"001010100",
  20474=>"000100110",
  20475=>"110101011",
  20476=>"101001100",
  20477=>"001000000",
  20478=>"110100101",
  20479=>"100001001",
  20480=>"110010100",
  20481=>"001111011",
  20482=>"010110101",
  20483=>"000001000",
  20484=>"100011101",
  20485=>"100100100",
  20486=>"010101101",
  20487=>"000000001",
  20488=>"000000111",
  20489=>"000000011",
  20490=>"111101111",
  20491=>"110110111",
  20492=>"010010010",
  20493=>"100000010",
  20494=>"100100101",
  20495=>"011101000",
  20496=>"010100111",
  20497=>"010011001",
  20498=>"001011101",
  20499=>"001110111",
  20500=>"000111110",
  20501=>"001011000",
  20502=>"101100011",
  20503=>"111111100",
  20504=>"000101000",
  20505=>"111111001",
  20506=>"011010100",
  20507=>"110000111",
  20508=>"010011110",
  20509=>"000010011",
  20510=>"110101110",
  20511=>"001001101",
  20512=>"000111000",
  20513=>"000011000",
  20514=>"001101010",
  20515=>"010000001",
  20516=>"110101010",
  20517=>"101011001",
  20518=>"011000100",
  20519=>"110100100",
  20520=>"001100101",
  20521=>"010110011",
  20522=>"111100001",
  20523=>"100111110",
  20524=>"101110010",
  20525=>"111011111",
  20526=>"001010101",
  20527=>"010110111",
  20528=>"110110111",
  20529=>"000000001",
  20530=>"000110111",
  20531=>"110110011",
  20532=>"000100000",
  20533=>"101111100",
  20534=>"100110011",
  20535=>"100110001",
  20536=>"011001100",
  20537=>"010010000",
  20538=>"010100011",
  20539=>"000101100",
  20540=>"001010100",
  20541=>"001101101",
  20542=>"001001001",
  20543=>"000001111",
  20544=>"011110011",
  20545=>"001000001",
  20546=>"100111000",
  20547=>"010001011",
  20548=>"000111101",
  20549=>"011011000",
  20550=>"010000001",
  20551=>"100110100",
  20552=>"101100001",
  20553=>"110011100",
  20554=>"100001110",
  20555=>"101010110",
  20556=>"111100100",
  20557=>"100110001",
  20558=>"110100101",
  20559=>"100111100",
  20560=>"111001001",
  20561=>"101000001",
  20562=>"101011010",
  20563=>"001001000",
  20564=>"110111011",
  20565=>"110100011",
  20566=>"101101111",
  20567=>"010001001",
  20568=>"111100111",
  20569=>"010000100",
  20570=>"010111001",
  20571=>"001110100",
  20572=>"100101100",
  20573=>"010111011",
  20574=>"111101010",
  20575=>"110010001",
  20576=>"101011000",
  20577=>"000100111",
  20578=>"001010010",
  20579=>"100001000",
  20580=>"000101000",
  20581=>"001110110",
  20582=>"100010100",
  20583=>"000011110",
  20584=>"111100000",
  20585=>"110110110",
  20586=>"101101000",
  20587=>"100011100",
  20588=>"111000001",
  20589=>"111111110",
  20590=>"001111101",
  20591=>"101110000",
  20592=>"110101011",
  20593=>"011001010",
  20594=>"001101101",
  20595=>"111101011",
  20596=>"001000111",
  20597=>"000101000",
  20598=>"100011001",
  20599=>"011011100",
  20600=>"010010111",
  20601=>"100111001",
  20602=>"111111010",
  20603=>"110000001",
  20604=>"100110011",
  20605=>"111011001",
  20606=>"000100000",
  20607=>"010000000",
  20608=>"001111000",
  20609=>"100011100",
  20610=>"011111111",
  20611=>"001010011",
  20612=>"000110111",
  20613=>"100001100",
  20614=>"000000010",
  20615=>"001000011",
  20616=>"011000000",
  20617=>"000000011",
  20618=>"011011110",
  20619=>"101101111",
  20620=>"011001100",
  20621=>"000000100",
  20622=>"100100111",
  20623=>"110111001",
  20624=>"010101001",
  20625=>"100011111",
  20626=>"011110110",
  20627=>"110100100",
  20628=>"001101111",
  20629=>"001111011",
  20630=>"110110110",
  20631=>"100101000",
  20632=>"010100000",
  20633=>"000110011",
  20634=>"000110011",
  20635=>"001101110",
  20636=>"000001100",
  20637=>"111101111",
  20638=>"101011000",
  20639=>"100000011",
  20640=>"000001110",
  20641=>"110100011",
  20642=>"010110111",
  20643=>"001110001",
  20644=>"000000010",
  20645=>"001011100",
  20646=>"000010000",
  20647=>"000000011",
  20648=>"000111101",
  20649=>"011101011",
  20650=>"011100000",
  20651=>"111001110",
  20652=>"001111001",
  20653=>"000111111",
  20654=>"100011101",
  20655=>"111001111",
  20656=>"011110100",
  20657=>"010010010",
  20658=>"010110110",
  20659=>"101001000",
  20660=>"111101001",
  20661=>"011010000",
  20662=>"001110100",
  20663=>"000110011",
  20664=>"011101010",
  20665=>"111010010",
  20666=>"100101011",
  20667=>"100010111",
  20668=>"010111000",
  20669=>"100101000",
  20670=>"110001100",
  20671=>"000010000",
  20672=>"111011000",
  20673=>"000100110",
  20674=>"011101000",
  20675=>"111000111",
  20676=>"100101000",
  20677=>"011111111",
  20678=>"101111101",
  20679=>"100110101",
  20680=>"011111100",
  20681=>"001101111",
  20682=>"111101111",
  20683=>"001111100",
  20684=>"111110010",
  20685=>"110000000",
  20686=>"000100100",
  20687=>"000000000",
  20688=>"111101001",
  20689=>"111001110",
  20690=>"101000000",
  20691=>"000110111",
  20692=>"000001111",
  20693=>"001000101",
  20694=>"000110001",
  20695=>"001100001",
  20696=>"000011101",
  20697=>"001010000",
  20698=>"111111010",
  20699=>"111000101",
  20700=>"000000100",
  20701=>"101110100",
  20702=>"100010100",
  20703=>"011001100",
  20704=>"001001001",
  20705=>"111100010",
  20706=>"010000110",
  20707=>"111100111",
  20708=>"010111110",
  20709=>"011001100",
  20710=>"101101001",
  20711=>"110010111",
  20712=>"010010010",
  20713=>"001101100",
  20714=>"001011001",
  20715=>"110100111",
  20716=>"011000000",
  20717=>"010101101",
  20718=>"001111000",
  20719=>"001001110",
  20720=>"111010000",
  20721=>"011110001",
  20722=>"011011010",
  20723=>"011100010",
  20724=>"111001110",
  20725=>"001110100",
  20726=>"100111100",
  20727=>"011001011",
  20728=>"101110001",
  20729=>"100100000",
  20730=>"111011100",
  20731=>"101101110",
  20732=>"111101101",
  20733=>"101101000",
  20734=>"001000110",
  20735=>"100001011",
  20736=>"010001001",
  20737=>"010011101",
  20738=>"010111011",
  20739=>"100110011",
  20740=>"011000010",
  20741=>"110000111",
  20742=>"011111000",
  20743=>"110100011",
  20744=>"001001011",
  20745=>"100000101",
  20746=>"111111101",
  20747=>"111110000",
  20748=>"111111011",
  20749=>"010110111",
  20750=>"100100111",
  20751=>"100011000",
  20752=>"111111000",
  20753=>"001000010",
  20754=>"000000011",
  20755=>"000001010",
  20756=>"001001001",
  20757=>"101010000",
  20758=>"001111000",
  20759=>"111110101",
  20760=>"010001010",
  20761=>"110011111",
  20762=>"111101101",
  20763=>"100110101",
  20764=>"111110110",
  20765=>"101000010",
  20766=>"110000110",
  20767=>"000001110",
  20768=>"011000101",
  20769=>"110111100",
  20770=>"011111111",
  20771=>"111010010",
  20772=>"011101010",
  20773=>"111000111",
  20774=>"011011010",
  20775=>"000010111",
  20776=>"110010110",
  20777=>"010001101",
  20778=>"110111010",
  20779=>"010001101",
  20780=>"101000001",
  20781=>"001100001",
  20782=>"000000001",
  20783=>"010000110",
  20784=>"010001010",
  20785=>"001011000",
  20786=>"110110111",
  20787=>"100000110",
  20788=>"010000111",
  20789=>"111000101",
  20790=>"110111000",
  20791=>"011101011",
  20792=>"110011110",
  20793=>"000100001",
  20794=>"101001011",
  20795=>"111110011",
  20796=>"110111011",
  20797=>"011111110",
  20798=>"010000000",
  20799=>"001101101",
  20800=>"000000001",
  20801=>"000010101",
  20802=>"101011000",
  20803=>"110101010",
  20804=>"001000111",
  20805=>"101000101",
  20806=>"101101011",
  20807=>"011100100",
  20808=>"111000000",
  20809=>"101100010",
  20810=>"110110000",
  20811=>"001010001",
  20812=>"010101001",
  20813=>"001101100",
  20814=>"111000100",
  20815=>"010100010",
  20816=>"110101111",
  20817=>"010111010",
  20818=>"001010100",
  20819=>"110011000",
  20820=>"010011000",
  20821=>"011011100",
  20822=>"011110110",
  20823=>"011111110",
  20824=>"011110100",
  20825=>"010010101",
  20826=>"001010101",
  20827=>"011100110",
  20828=>"001010010",
  20829=>"000010000",
  20830=>"101110011",
  20831=>"100011110",
  20832=>"000110000",
  20833=>"010011001",
  20834=>"110010111",
  20835=>"010001001",
  20836=>"010101010",
  20837=>"011101000",
  20838=>"000011100",
  20839=>"011001001",
  20840=>"010111000",
  20841=>"101001000",
  20842=>"000110011",
  20843=>"111010101",
  20844=>"110110011",
  20845=>"001101011",
  20846=>"000010000",
  20847=>"001000010",
  20848=>"100111110",
  20849=>"010110011",
  20850=>"010100000",
  20851=>"001010111",
  20852=>"101101100",
  20853=>"111101111",
  20854=>"001101011",
  20855=>"010100001",
  20856=>"110111101",
  20857=>"111000001",
  20858=>"111001011",
  20859=>"110010111",
  20860=>"111101001",
  20861=>"111101001",
  20862=>"110110100",
  20863=>"001110000",
  20864=>"110011111",
  20865=>"000001111",
  20866=>"111111010",
  20867=>"101000001",
  20868=>"001111010",
  20869=>"000101001",
  20870=>"110011100",
  20871=>"000110110",
  20872=>"010011001",
  20873=>"101011100",
  20874=>"100101100",
  20875=>"100100110",
  20876=>"110000100",
  20877=>"010111101",
  20878=>"001000010",
  20879=>"010100100",
  20880=>"001011100",
  20881=>"001100110",
  20882=>"011001001",
  20883=>"001000111",
  20884=>"000000000",
  20885=>"001010011",
  20886=>"100110111",
  20887=>"100101110",
  20888=>"101010111",
  20889=>"011001010",
  20890=>"111000100",
  20891=>"111011101",
  20892=>"101000010",
  20893=>"110011000",
  20894=>"010111011",
  20895=>"111000010",
  20896=>"110101010",
  20897=>"000100110",
  20898=>"100111111",
  20899=>"101011011",
  20900=>"010000001",
  20901=>"000101100",
  20902=>"000000111",
  20903=>"111010101",
  20904=>"001110010",
  20905=>"101101111",
  20906=>"110100101",
  20907=>"110011000",
  20908=>"111000001",
  20909=>"101011110",
  20910=>"010010000",
  20911=>"111001011",
  20912=>"111001001",
  20913=>"110100110",
  20914=>"100001101",
  20915=>"111101000",
  20916=>"111101010",
  20917=>"000100001",
  20918=>"110111100",
  20919=>"001100110",
  20920=>"010100100",
  20921=>"001101110",
  20922=>"111111001",
  20923=>"111101101",
  20924=>"000110000",
  20925=>"101100011",
  20926=>"000110101",
  20927=>"101100101",
  20928=>"010101001",
  20929=>"111111110",
  20930=>"111011010",
  20931=>"110000010",
  20932=>"000010000",
  20933=>"101111101",
  20934=>"000010100",
  20935=>"010000100",
  20936=>"011001001",
  20937=>"001110000",
  20938=>"010100110",
  20939=>"011101010",
  20940=>"101001100",
  20941=>"100110000",
  20942=>"001101011",
  20943=>"110100111",
  20944=>"110011100",
  20945=>"011001010",
  20946=>"101011010",
  20947=>"101100101",
  20948=>"010101001",
  20949=>"111101101",
  20950=>"011110000",
  20951=>"101111111",
  20952=>"001000100",
  20953=>"011111100",
  20954=>"101100010",
  20955=>"101111100",
  20956=>"001110010",
  20957=>"110001111",
  20958=>"010011111",
  20959=>"101101010",
  20960=>"001111101",
  20961=>"011001100",
  20962=>"001011110",
  20963=>"011100010",
  20964=>"100100110",
  20965=>"001111011",
  20966=>"010000010",
  20967=>"000011011",
  20968=>"000011100",
  20969=>"101010011",
  20970=>"010100000",
  20971=>"101110001",
  20972=>"100111100",
  20973=>"000110000",
  20974=>"100100111",
  20975=>"100110010",
  20976=>"110001100",
  20977=>"100010111",
  20978=>"101101101",
  20979=>"000000000",
  20980=>"110001001",
  20981=>"000110100",
  20982=>"100101010",
  20983=>"101101000",
  20984=>"001101001",
  20985=>"100111001",
  20986=>"100011011",
  20987=>"100001111",
  20988=>"101110110",
  20989=>"000011100",
  20990=>"001001101",
  20991=>"101111001",
  20992=>"001001100",
  20993=>"001010000",
  20994=>"011010110",
  20995=>"110100001",
  20996=>"010011001",
  20997=>"010111111",
  20998=>"010110001",
  20999=>"111000100",
  21000=>"101000101",
  21001=>"101011101",
  21002=>"100001110",
  21003=>"011101001",
  21004=>"110111000",
  21005=>"010011101",
  21006=>"010100011",
  21007=>"001011000",
  21008=>"111101110",
  21009=>"100000000",
  21010=>"000000111",
  21011=>"110001110",
  21012=>"011101100",
  21013=>"011011001",
  21014=>"101010111",
  21015=>"111100010",
  21016=>"010111001",
  21017=>"111100001",
  21018=>"111001111",
  21019=>"001001001",
  21020=>"100000001",
  21021=>"011001011",
  21022=>"111000001",
  21023=>"001110111",
  21024=>"101000011",
  21025=>"110100110",
  21026=>"101101000",
  21027=>"100010001",
  21028=>"110111100",
  21029=>"000000110",
  21030=>"100100110",
  21031=>"011010001",
  21032=>"010100100",
  21033=>"001000100",
  21034=>"001011110",
  21035=>"100100100",
  21036=>"101111110",
  21037=>"111111110",
  21038=>"010100001",
  21039=>"010110101",
  21040=>"001010110",
  21041=>"100011110",
  21042=>"111100100",
  21043=>"100010100",
  21044=>"001010010",
  21045=>"001111000",
  21046=>"110110100",
  21047=>"100100100",
  21048=>"010011001",
  21049=>"001000010",
  21050=>"011001110",
  21051=>"001010010",
  21052=>"111111010",
  21053=>"010101011",
  21054=>"111110001",
  21055=>"101001110",
  21056=>"000100101",
  21057=>"010000110",
  21058=>"100111111",
  21059=>"110000001",
  21060=>"101011110",
  21061=>"100100110",
  21062=>"110000010",
  21063=>"000010011",
  21064=>"001000101",
  21065=>"000111110",
  21066=>"101011001",
  21067=>"100110111",
  21068=>"101000101",
  21069=>"011111111",
  21070=>"000101011",
  21071=>"110111010",
  21072=>"101001111",
  21073=>"001000000",
  21074=>"110101111",
  21075=>"111101000",
  21076=>"011001000",
  21077=>"000011100",
  21078=>"111111111",
  21079=>"100101111",
  21080=>"100010000",
  21081=>"000000011",
  21082=>"111110111",
  21083=>"000001100",
  21084=>"111011100",
  21085=>"100110011",
  21086=>"001100010",
  21087=>"100000110",
  21088=>"100000110",
  21089=>"101110111",
  21090=>"110111010",
  21091=>"110101111",
  21092=>"101000101",
  21093=>"001101010",
  21094=>"101010000",
  21095=>"101111000",
  21096=>"000001101",
  21097=>"001001111",
  21098=>"110010000",
  21099=>"011011100",
  21100=>"000001100",
  21101=>"111011011",
  21102=>"101101011",
  21103=>"001010111",
  21104=>"111100011",
  21105=>"101101100",
  21106=>"110011110",
  21107=>"111101110",
  21108=>"110000011",
  21109=>"111110111",
  21110=>"011001001",
  21111=>"100001000",
  21112=>"111011110",
  21113=>"010001000",
  21114=>"111000000",
  21115=>"011100111",
  21116=>"010110110",
  21117=>"101010111",
  21118=>"110011101",
  21119=>"001110011",
  21120=>"111101011",
  21121=>"101001000",
  21122=>"111111011",
  21123=>"110110100",
  21124=>"001100100",
  21125=>"000100000",
  21126=>"101111000",
  21127=>"010110110",
  21128=>"101010101",
  21129=>"100101011",
  21130=>"111000110",
  21131=>"001001100",
  21132=>"111001011",
  21133=>"001111101",
  21134=>"100101110",
  21135=>"000100110",
  21136=>"000111000",
  21137=>"001101000",
  21138=>"111100001",
  21139=>"010101100",
  21140=>"011110000",
  21141=>"011000001",
  21142=>"001111001",
  21143=>"111101100",
  21144=>"111110100",
  21145=>"011110011",
  21146=>"011001000",
  21147=>"010110000",
  21148=>"000100010",
  21149=>"111011001",
  21150=>"001111101",
  21151=>"011001111",
  21152=>"101010110",
  21153=>"101001010",
  21154=>"111011101",
  21155=>"111011011",
  21156=>"011111101",
  21157=>"101011100",
  21158=>"010100010",
  21159=>"111000111",
  21160=>"011011101",
  21161=>"111110111",
  21162=>"101110111",
  21163=>"001111001",
  21164=>"001111011",
  21165=>"100001001",
  21166=>"101000111",
  21167=>"000001000",
  21168=>"110101111",
  21169=>"110000001",
  21170=>"111011100",
  21171=>"001100011",
  21172=>"110100111",
  21173=>"000111001",
  21174=>"011010110",
  21175=>"111101100",
  21176=>"111011011",
  21177=>"001111111",
  21178=>"100101010",
  21179=>"000000000",
  21180=>"011001100",
  21181=>"010011011",
  21182=>"011011010",
  21183=>"111110111",
  21184=>"110100001",
  21185=>"011011101",
  21186=>"111111111",
  21187=>"101000000",
  21188=>"111111100",
  21189=>"001011010",
  21190=>"001011101",
  21191=>"011101100",
  21192=>"101101111",
  21193=>"010000001",
  21194=>"111110010",
  21195=>"111000011",
  21196=>"000010011",
  21197=>"111101101",
  21198=>"110011000",
  21199=>"000100000",
  21200=>"011011111",
  21201=>"011111001",
  21202=>"001000010",
  21203=>"101111111",
  21204=>"101000100",
  21205=>"000111110",
  21206=>"100110011",
  21207=>"000101100",
  21208=>"100011100",
  21209=>"110110100",
  21210=>"001110000",
  21211=>"001010001",
  21212=>"111011000",
  21213=>"000101001",
  21214=>"111011001",
  21215=>"001101001",
  21216=>"010001111",
  21217=>"000111011",
  21218=>"011100110",
  21219=>"101101111",
  21220=>"001001000",
  21221=>"100100000",
  21222=>"100100101",
  21223=>"000000001",
  21224=>"100111100",
  21225=>"101111111",
  21226=>"011001111",
  21227=>"100101101",
  21228=>"110101001",
  21229=>"110101000",
  21230=>"110110110",
  21231=>"000010000",
  21232=>"000100101",
  21233=>"110111101",
  21234=>"100010101",
  21235=>"010010001",
  21236=>"101110011",
  21237=>"110000000",
  21238=>"110110110",
  21239=>"001000011",
  21240=>"101110111",
  21241=>"100100011",
  21242=>"000010001",
  21243=>"011011100",
  21244=>"010100001",
  21245=>"101010101",
  21246=>"110011000",
  21247=>"010000100",
  21248=>"101110000",
  21249=>"100111111",
  21250=>"101011101",
  21251=>"000000100",
  21252=>"000000001",
  21253=>"101010001",
  21254=>"111100110",
  21255=>"100111011",
  21256=>"010000010",
  21257=>"010010101",
  21258=>"000011001",
  21259=>"011100100",
  21260=>"010001100",
  21261=>"010100001",
  21262=>"010111011",
  21263=>"000010000",
  21264=>"010100110",
  21265=>"010011001",
  21266=>"010011111",
  21267=>"101101011",
  21268=>"010100101",
  21269=>"111100000",
  21270=>"010100000",
  21271=>"000111111",
  21272=>"010100010",
  21273=>"110000000",
  21274=>"000111100",
  21275=>"111101010",
  21276=>"001000100",
  21277=>"111010011",
  21278=>"001101101",
  21279=>"001010111",
  21280=>"010101111",
  21281=>"110011000",
  21282=>"011111101",
  21283=>"100000101",
  21284=>"010111110",
  21285=>"100001111",
  21286=>"111011010",
  21287=>"100011100",
  21288=>"000000000",
  21289=>"100000000",
  21290=>"111110011",
  21291=>"000000111",
  21292=>"001011100",
  21293=>"001011010",
  21294=>"011110101",
  21295=>"111011101",
  21296=>"111101001",
  21297=>"101100100",
  21298=>"001000000",
  21299=>"100001000",
  21300=>"000000101",
  21301=>"100110110",
  21302=>"101010011",
  21303=>"100001000",
  21304=>"100000000",
  21305=>"011011111",
  21306=>"000101001",
  21307=>"011001111",
  21308=>"110110110",
  21309=>"110010010",
  21310=>"111110101",
  21311=>"110101101",
  21312=>"111100100",
  21313=>"010101001",
  21314=>"010100110",
  21315=>"111100001",
  21316=>"100011001",
  21317=>"000100010",
  21318=>"110010101",
  21319=>"101011010",
  21320=>"011110010",
  21321=>"110111100",
  21322=>"100001000",
  21323=>"000001001",
  21324=>"101111001",
  21325=>"111010101",
  21326=>"100101110",
  21327=>"000011010",
  21328=>"110000101",
  21329=>"011000010",
  21330=>"100110001",
  21331=>"100000101",
  21332=>"001001101",
  21333=>"001100101",
  21334=>"100000110",
  21335=>"001101100",
  21336=>"101101010",
  21337=>"100001010",
  21338=>"101110111",
  21339=>"001110111",
  21340=>"101000111",
  21341=>"001110111",
  21342=>"110010000",
  21343=>"001111010",
  21344=>"000100011",
  21345=>"111001011",
  21346=>"110100111",
  21347=>"101110000",
  21348=>"010001110",
  21349=>"101111111",
  21350=>"101100101",
  21351=>"000001110",
  21352=>"110111010",
  21353=>"111111001",
  21354=>"111001010",
  21355=>"001111001",
  21356=>"111100101",
  21357=>"010100010",
  21358=>"111011011",
  21359=>"110000011",
  21360=>"101111101",
  21361=>"001000100",
  21362=>"111000111",
  21363=>"001110111",
  21364=>"011010110",
  21365=>"101000111",
  21366=>"010011101",
  21367=>"000101111",
  21368=>"101000011",
  21369=>"001111000",
  21370=>"101101000",
  21371=>"111010110",
  21372=>"010001001",
  21373=>"111111110",
  21374=>"100011100",
  21375=>"000100001",
  21376=>"001100100",
  21377=>"110110110",
  21378=>"100001000",
  21379=>"100111001",
  21380=>"101111110",
  21381=>"001010000",
  21382=>"010000111",
  21383=>"001011110",
  21384=>"111110000",
  21385=>"111111010",
  21386=>"110101100",
  21387=>"000111111",
  21388=>"000000101",
  21389=>"101010000",
  21390=>"001101111",
  21391=>"010110001",
  21392=>"001010101",
  21393=>"110011111",
  21394=>"101111000",
  21395=>"111001001",
  21396=>"001011101",
  21397=>"100111010",
  21398=>"100001111",
  21399=>"000100110",
  21400=>"010011010",
  21401=>"001000100",
  21402=>"110101000",
  21403=>"010101101",
  21404=>"111001000",
  21405=>"100111000",
  21406=>"110001010",
  21407=>"010001010",
  21408=>"010000101",
  21409=>"110001100",
  21410=>"100111110",
  21411=>"110101011",
  21412=>"000000001",
  21413=>"110100000",
  21414=>"001011111",
  21415=>"010011110",
  21416=>"000010110",
  21417=>"100001000",
  21418=>"111101000",
  21419=>"101111001",
  21420=>"011100111",
  21421=>"011101010",
  21422=>"001111001",
  21423=>"001100001",
  21424=>"100101101",
  21425=>"111010011",
  21426=>"101100001",
  21427=>"100100111",
  21428=>"101110000",
  21429=>"101000100",
  21430=>"000101100",
  21431=>"000111100",
  21432=>"111010111",
  21433=>"010010011",
  21434=>"111011010",
  21435=>"101001000",
  21436=>"011000010",
  21437=>"011111111",
  21438=>"000100100",
  21439=>"100000101",
  21440=>"100001111",
  21441=>"100010010",
  21442=>"111100001",
  21443=>"111011010",
  21444=>"010000100",
  21445=>"000011010",
  21446=>"000000100",
  21447=>"101110101",
  21448=>"011010100",
  21449=>"100100000",
  21450=>"101100011",
  21451=>"111011000",
  21452=>"010111110",
  21453=>"011100010",
  21454=>"110111111",
  21455=>"011001100",
  21456=>"111100010",
  21457=>"101101010",
  21458=>"101011000",
  21459=>"100000000",
  21460=>"111000010",
  21461=>"010011000",
  21462=>"001001100",
  21463=>"110010101",
  21464=>"000010011",
  21465=>"100001010",
  21466=>"000000101",
  21467=>"000001110",
  21468=>"110010110",
  21469=>"101100011",
  21470=>"010010001",
  21471=>"110010011",
  21472=>"111111011",
  21473=>"010100100",
  21474=>"011010011",
  21475=>"000000100",
  21476=>"010010110",
  21477=>"000010010",
  21478=>"101000010",
  21479=>"100110111",
  21480=>"001001100",
  21481=>"111111110",
  21482=>"110101000",
  21483=>"000000001",
  21484=>"011101001",
  21485=>"001000000",
  21486=>"010001000",
  21487=>"111000010",
  21488=>"101111011",
  21489=>"000111010",
  21490=>"101110000",
  21491=>"100111100",
  21492=>"110001010",
  21493=>"011010111",
  21494=>"011110111",
  21495=>"000111011",
  21496=>"101001010",
  21497=>"011101100",
  21498=>"111111111",
  21499=>"111011110",
  21500=>"110011100",
  21501=>"101101101",
  21502=>"010101111",
  21503=>"011000000",
  21504=>"001000101",
  21505=>"001011100",
  21506=>"000011110",
  21507=>"110111100",
  21508=>"001000010",
  21509=>"000010010",
  21510=>"010000100",
  21511=>"101001001",
  21512=>"011111011",
  21513=>"000000100",
  21514=>"001011000",
  21515=>"101110101",
  21516=>"001011000",
  21517=>"101100010",
  21518=>"010011010",
  21519=>"000110011",
  21520=>"000001111",
  21521=>"110000110",
  21522=>"100000100",
  21523=>"101110010",
  21524=>"101101010",
  21525=>"011110100",
  21526=>"000010111",
  21527=>"001010111",
  21528=>"111100100",
  21529=>"001111011",
  21530=>"111011001",
  21531=>"010000101",
  21532=>"011100000",
  21533=>"001001110",
  21534=>"000000010",
  21535=>"110010011",
  21536=>"100100101",
  21537=>"101011100",
  21538=>"000001001",
  21539=>"100000001",
  21540=>"100011111",
  21541=>"111100011",
  21542=>"101000111",
  21543=>"010000100",
  21544=>"100011010",
  21545=>"101111111",
  21546=>"000100000",
  21547=>"001000110",
  21548=>"011010001",
  21549=>"010111111",
  21550=>"010101011",
  21551=>"000101110",
  21552=>"011101111",
  21553=>"110010111",
  21554=>"011101110",
  21555=>"101011111",
  21556=>"011111011",
  21557=>"101001011",
  21558=>"110101000",
  21559=>"100100001",
  21560=>"001110101",
  21561=>"000010100",
  21562=>"011011100",
  21563=>"101100000",
  21564=>"010101000",
  21565=>"011100000",
  21566=>"001010100",
  21567=>"000010111",
  21568=>"011001000",
  21569=>"110100000",
  21570=>"101010001",
  21571=>"101000000",
  21572=>"100000110",
  21573=>"000001100",
  21574=>"110111000",
  21575=>"000000011",
  21576=>"011011100",
  21577=>"110101000",
  21578=>"100111111",
  21579=>"111101010",
  21580=>"101010011",
  21581=>"011010100",
  21582=>"001011110",
  21583=>"001110101",
  21584=>"011010000",
  21585=>"001000000",
  21586=>"101100100",
  21587=>"100000000",
  21588=>"000101011",
  21589=>"111110110",
  21590=>"101011000",
  21591=>"101101000",
  21592=>"111101110",
  21593=>"100000001",
  21594=>"001000110",
  21595=>"001001010",
  21596=>"101101011",
  21597=>"101000101",
  21598=>"011001001",
  21599=>"011001110",
  21600=>"101101101",
  21601=>"001101010",
  21602=>"001010111",
  21603=>"011101001",
  21604=>"100000001",
  21605=>"011001100",
  21606=>"001110111",
  21607=>"110010111",
  21608=>"101010101",
  21609=>"111110110",
  21610=>"101111000",
  21611=>"101000101",
  21612=>"001111101",
  21613=>"110011100",
  21614=>"101111010",
  21615=>"111011110",
  21616=>"101101001",
  21617=>"000111010",
  21618=>"000011111",
  21619=>"000010000",
  21620=>"101100010",
  21621=>"101001000",
  21622=>"001101011",
  21623=>"110011011",
  21624=>"011111010",
  21625=>"011011111",
  21626=>"111111111",
  21627=>"000101010",
  21628=>"000001011",
  21629=>"101101010",
  21630=>"010110010",
  21631=>"100011000",
  21632=>"000101100",
  21633=>"000011001",
  21634=>"100101000",
  21635=>"111010110",
  21636=>"101011000",
  21637=>"011000101",
  21638=>"001101011",
  21639=>"011110111",
  21640=>"100111111",
  21641=>"111000010",
  21642=>"111000011",
  21643=>"000010111",
  21644=>"000010011",
  21645=>"010010000",
  21646=>"001010100",
  21647=>"111111111",
  21648=>"001101110",
  21649=>"011000011",
  21650=>"111111000",
  21651=>"000100110",
  21652=>"111111101",
  21653=>"100110101",
  21654=>"100000001",
  21655=>"111011111",
  21656=>"101110111",
  21657=>"001000000",
  21658=>"111100101",
  21659=>"011111101",
  21660=>"000000110",
  21661=>"111110100",
  21662=>"111101010",
  21663=>"101101111",
  21664=>"011110011",
  21665=>"100000110",
  21666=>"100100000",
  21667=>"100100111",
  21668=>"001110010",
  21669=>"110000000",
  21670=>"001100111",
  21671=>"011011110",
  21672=>"100011001",
  21673=>"001010000",
  21674=>"000010100",
  21675=>"000100000",
  21676=>"100111100",
  21677=>"000111011",
  21678=>"101110110",
  21679=>"010011100",
  21680=>"001101110",
  21681=>"110110100",
  21682=>"001101010",
  21683=>"001111001",
  21684=>"000100111",
  21685=>"010001000",
  21686=>"100001100",
  21687=>"011011110",
  21688=>"110111011",
  21689=>"111000111",
  21690=>"101010010",
  21691=>"100011010",
  21692=>"100001000",
  21693=>"001100111",
  21694=>"010110110",
  21695=>"010000010",
  21696=>"010101100",
  21697=>"101101100",
  21698=>"111100100",
  21699=>"010010101",
  21700=>"111111100",
  21701=>"100100101",
  21702=>"011101000",
  21703=>"101110110",
  21704=>"110100001",
  21705=>"110010110",
  21706=>"111001000",
  21707=>"101010111",
  21708=>"101110100",
  21709=>"011011100",
  21710=>"000000000",
  21711=>"100100001",
  21712=>"100100111",
  21713=>"101100010",
  21714=>"100010001",
  21715=>"010000111",
  21716=>"110000011",
  21717=>"001011001",
  21718=>"000110000",
  21719=>"111000010",
  21720=>"100101111",
  21721=>"000001010",
  21722=>"100110011",
  21723=>"001101001",
  21724=>"111001000",
  21725=>"010111010",
  21726=>"010000101",
  21727=>"101000101",
  21728=>"010000110",
  21729=>"100111010",
  21730=>"110001011",
  21731=>"110100000",
  21732=>"100111110",
  21733=>"110011111",
  21734=>"001001111",
  21735=>"110010001",
  21736=>"000000101",
  21737=>"001000100",
  21738=>"111111110",
  21739=>"101101000",
  21740=>"110100010",
  21741=>"110100111",
  21742=>"010000000",
  21743=>"111001011",
  21744=>"011011110",
  21745=>"101000000",
  21746=>"101100100",
  21747=>"100111001",
  21748=>"010000011",
  21749=>"101010110",
  21750=>"100011010",
  21751=>"010100111",
  21752=>"010011000",
  21753=>"000000100",
  21754=>"011111101",
  21755=>"100110110",
  21756=>"000011100",
  21757=>"111110101",
  21758=>"100001110",
  21759=>"110110000",
  21760=>"010111111",
  21761=>"010101011",
  21762=>"111011011",
  21763=>"101101000",
  21764=>"100100000",
  21765=>"000000100",
  21766=>"100100100",
  21767=>"100001101",
  21768=>"101010100",
  21769=>"101000011",
  21770=>"000011101",
  21771=>"001101101",
  21772=>"111011111",
  21773=>"111101001",
  21774=>"001101101",
  21775=>"000001001",
  21776=>"100110010",
  21777=>"111010011",
  21778=>"000000010",
  21779=>"011111110",
  21780=>"111011100",
  21781=>"100111110",
  21782=>"110010111",
  21783=>"101101100",
  21784=>"000001000",
  21785=>"101101101",
  21786=>"001010110",
  21787=>"000110011",
  21788=>"100010011",
  21789=>"111001000",
  21790=>"001010101",
  21791=>"001001111",
  21792=>"010110001",
  21793=>"000111110",
  21794=>"101110111",
  21795=>"010010111",
  21796=>"100000101",
  21797=>"101010110",
  21798=>"101010000",
  21799=>"011010110",
  21800=>"111101101",
  21801=>"001001001",
  21802=>"011111100",
  21803=>"010010110",
  21804=>"101000000",
  21805=>"011001010",
  21806=>"101000101",
  21807=>"101001011",
  21808=>"000101011",
  21809=>"111110011",
  21810=>"001010110",
  21811=>"101110111",
  21812=>"000001110",
  21813=>"011110101",
  21814=>"111110101",
  21815=>"101000000",
  21816=>"000001000",
  21817=>"010000000",
  21818=>"110011100",
  21819=>"111010101",
  21820=>"111001111",
  21821=>"001001000",
  21822=>"000010011",
  21823=>"000101001",
  21824=>"010010101",
  21825=>"111011101",
  21826=>"100101001",
  21827=>"110110000",
  21828=>"110110011",
  21829=>"100000101",
  21830=>"101101101",
  21831=>"000000110",
  21832=>"111110101",
  21833=>"101010000",
  21834=>"010111001",
  21835=>"010110000",
  21836=>"110011100",
  21837=>"010011101",
  21838=>"011101010",
  21839=>"101100000",
  21840=>"101001001",
  21841=>"000111101",
  21842=>"011100000",
  21843=>"100111100",
  21844=>"001110001",
  21845=>"111101101",
  21846=>"111000101",
  21847=>"111100001",
  21848=>"100010110",
  21849=>"100101111",
  21850=>"000011001",
  21851=>"011001001",
  21852=>"111001110",
  21853=>"110111000",
  21854=>"011001000",
  21855=>"001110111",
  21856=>"001010100",
  21857=>"001010000",
  21858=>"001101101",
  21859=>"000011101",
  21860=>"101010101",
  21861=>"011010000",
  21862=>"100011101",
  21863=>"000110011",
  21864=>"010011001",
  21865=>"001010100",
  21866=>"010001011",
  21867=>"011000100",
  21868=>"100000010",
  21869=>"011101101",
  21870=>"001010111",
  21871=>"001010111",
  21872=>"001011111",
  21873=>"010110000",
  21874=>"011100101",
  21875=>"110001011",
  21876=>"100101001",
  21877=>"111111011",
  21878=>"100101000",
  21879=>"101001100",
  21880=>"000010110",
  21881=>"101011110",
  21882=>"010101110",
  21883=>"101011011",
  21884=>"110100011",
  21885=>"000010110",
  21886=>"001100101",
  21887=>"011000010",
  21888=>"101100011",
  21889=>"000111111",
  21890=>"110101101",
  21891=>"011010011",
  21892=>"110110000",
  21893=>"111111101",
  21894=>"100101011",
  21895=>"000110000",
  21896=>"001001010",
  21897=>"110100111",
  21898=>"110000001",
  21899=>"100110101",
  21900=>"000001001",
  21901=>"101000101",
  21902=>"000011010",
  21903=>"000101010",
  21904=>"101111000",
  21905=>"101000101",
  21906=>"010100011",
  21907=>"010110010",
  21908=>"010001000",
  21909=>"001110000",
  21910=>"010000111",
  21911=>"100110011",
  21912=>"011101010",
  21913=>"001101111",
  21914=>"001011010",
  21915=>"100000010",
  21916=>"100010001",
  21917=>"100101010",
  21918=>"011001000",
  21919=>"110110010",
  21920=>"001111010",
  21921=>"111011101",
  21922=>"111110101",
  21923=>"000011111",
  21924=>"101101001",
  21925=>"100110001",
  21926=>"000010000",
  21927=>"011100100",
  21928=>"000000000",
  21929=>"111000110",
  21930=>"100110111",
  21931=>"101010101",
  21932=>"110001111",
  21933=>"100100000",
  21934=>"101011101",
  21935=>"010011010",
  21936=>"100101010",
  21937=>"100100110",
  21938=>"000110011",
  21939=>"010011101",
  21940=>"001000100",
  21941=>"111110010",
  21942=>"010010111",
  21943=>"110111001",
  21944=>"111101101",
  21945=>"010000011",
  21946=>"001010100",
  21947=>"010100101",
  21948=>"000100111",
  21949=>"000110111",
  21950=>"000100100",
  21951=>"011001111",
  21952=>"011011000",
  21953=>"010110001",
  21954=>"101101011",
  21955=>"111111000",
  21956=>"100001001",
  21957=>"111011000",
  21958=>"111100001",
  21959=>"110000010",
  21960=>"001101111",
  21961=>"010111011",
  21962=>"011011000",
  21963=>"000000100",
  21964=>"000000111",
  21965=>"010110101",
  21966=>"100101101",
  21967=>"111101111",
  21968=>"101000100",
  21969=>"100110110",
  21970=>"000000011",
  21971=>"100011000",
  21972=>"101001100",
  21973=>"111000010",
  21974=>"100111010",
  21975=>"101011000",
  21976=>"010111011",
  21977=>"100100000",
  21978=>"110110100",
  21979=>"101100101",
  21980=>"110011111",
  21981=>"000011110",
  21982=>"101001110",
  21983=>"111001111",
  21984=>"011111001",
  21985=>"110011011",
  21986=>"001110101",
  21987=>"111100000",
  21988=>"100001101",
  21989=>"000011101",
  21990=>"001011111",
  21991=>"000010100",
  21992=>"110011110",
  21993=>"111011011",
  21994=>"110101111",
  21995=>"100010101",
  21996=>"111100110",
  21997=>"000101100",
  21998=>"101101000",
  21999=>"011000101",
  22000=>"110111111",
  22001=>"111100101",
  22002=>"111001101",
  22003=>"010001001",
  22004=>"000001000",
  22005=>"010101011",
  22006=>"100110100",
  22007=>"110101010",
  22008=>"011111111",
  22009=>"011011101",
  22010=>"001001100",
  22011=>"000111011",
  22012=>"100111110",
  22013=>"001011010",
  22014=>"110000011",
  22015=>"001000001",
  22016=>"011100001",
  22017=>"001100110",
  22018=>"100110111",
  22019=>"101100001",
  22020=>"111100010",
  22021=>"100000010",
  22022=>"111001111",
  22023=>"001101111",
  22024=>"101011001",
  22025=>"001110011",
  22026=>"011100100",
  22027=>"001011111",
  22028=>"101010001",
  22029=>"111001100",
  22030=>"110100111",
  22031=>"000000101",
  22032=>"100111110",
  22033=>"110100000",
  22034=>"000011111",
  22035=>"110111001",
  22036=>"001010000",
  22037=>"100000011",
  22038=>"001111000",
  22039=>"111110010",
  22040=>"100111110",
  22041=>"001000001",
  22042=>"100101010",
  22043=>"110111011",
  22044=>"000111101",
  22045=>"100110000",
  22046=>"011111101",
  22047=>"110011101",
  22048=>"011000001",
  22049=>"110010101",
  22050=>"100001101",
  22051=>"001110000",
  22052=>"011011011",
  22053=>"110100100",
  22054=>"011111110",
  22055=>"010010011",
  22056=>"101001011",
  22057=>"111001001",
  22058=>"110001111",
  22059=>"100001001",
  22060=>"111001011",
  22061=>"100001111",
  22062=>"111101011",
  22063=>"111101111",
  22064=>"011010011",
  22065=>"110100001",
  22066=>"100001010",
  22067=>"101111011",
  22068=>"111111000",
  22069=>"100001111",
  22070=>"011110001",
  22071=>"010110111",
  22072=>"000010100",
  22073=>"111001010",
  22074=>"101110110",
  22075=>"001010111",
  22076=>"100001111",
  22077=>"001111101",
  22078=>"001000010",
  22079=>"111001001",
  22080=>"111101000",
  22081=>"011111100",
  22082=>"101010101",
  22083=>"000001001",
  22084=>"110011101",
  22085=>"101100000",
  22086=>"010101000",
  22087=>"010001001",
  22088=>"100100011",
  22089=>"101111001",
  22090=>"000011110",
  22091=>"011010100",
  22092=>"110100101",
  22093=>"110010100",
  22094=>"101101111",
  22095=>"010011101",
  22096=>"110101101",
  22097=>"000110111",
  22098=>"001100000",
  22099=>"101101111",
  22100=>"010001010",
  22101=>"101001000",
  22102=>"001000010",
  22103=>"100111101",
  22104=>"000011101",
  22105=>"100100111",
  22106=>"110011001",
  22107=>"001100111",
  22108=>"110110101",
  22109=>"001001100",
  22110=>"101001010",
  22111=>"000011010",
  22112=>"011010111",
  22113=>"101010100",
  22114=>"001001001",
  22115=>"001110111",
  22116=>"111010110",
  22117=>"100111000",
  22118=>"010101111",
  22119=>"001001100",
  22120=>"000101010",
  22121=>"100100000",
  22122=>"011100100",
  22123=>"010000001",
  22124=>"101001111",
  22125=>"100011100",
  22126=>"101000010",
  22127=>"110001111",
  22128=>"111001000",
  22129=>"001100000",
  22130=>"111001110",
  22131=>"001010011",
  22132=>"000110101",
  22133=>"011100111",
  22134=>"000011001",
  22135=>"000010001",
  22136=>"110100111",
  22137=>"010110100",
  22138=>"000001000",
  22139=>"011010000",
  22140=>"010111111",
  22141=>"011100001",
  22142=>"011111010",
  22143=>"111001011",
  22144=>"000111100",
  22145=>"000111100",
  22146=>"000100100",
  22147=>"011010000",
  22148=>"000010101",
  22149=>"000111101",
  22150=>"110101101",
  22151=>"011010101",
  22152=>"111101110",
  22153=>"000000111",
  22154=>"111100010",
  22155=>"001010110",
  22156=>"000001100",
  22157=>"110010100",
  22158=>"001001101",
  22159=>"010101010",
  22160=>"101000000",
  22161=>"111111000",
  22162=>"100110011",
  22163=>"101100101",
  22164=>"110011010",
  22165=>"010110111",
  22166=>"111010000",
  22167=>"101000000",
  22168=>"111101111",
  22169=>"100100111",
  22170=>"110010011",
  22171=>"010000010",
  22172=>"010110111",
  22173=>"010110100",
  22174=>"000011000",
  22175=>"110001001",
  22176=>"100110111",
  22177=>"011110101",
  22178=>"100110010",
  22179=>"110101101",
  22180=>"100101000",
  22181=>"100101110",
  22182=>"101001110",
  22183=>"100011011",
  22184=>"100110100",
  22185=>"010110010",
  22186=>"100110011",
  22187=>"000011010",
  22188=>"100110000",
  22189=>"101010011",
  22190=>"111001101",
  22191=>"010101000",
  22192=>"100101000",
  22193=>"100001001",
  22194=>"000101101",
  22195=>"000000110",
  22196=>"101011001",
  22197=>"000110011",
  22198=>"101110000",
  22199=>"000101101",
  22200=>"110111110",
  22201=>"001000000",
  22202=>"111100010",
  22203=>"001111101",
  22204=>"001101110",
  22205=>"011010010",
  22206=>"001101011",
  22207=>"010100100",
  22208=>"001110101",
  22209=>"001101010",
  22210=>"101001111",
  22211=>"100111100",
  22212=>"011001001",
  22213=>"001001011",
  22214=>"111101100",
  22215=>"010100111",
  22216=>"100111011",
  22217=>"011010100",
  22218=>"101001101",
  22219=>"110000101",
  22220=>"111101101",
  22221=>"101001110",
  22222=>"101100011",
  22223=>"010000100",
  22224=>"111001110",
  22225=>"111000110",
  22226=>"000001100",
  22227=>"101110011",
  22228=>"010001110",
  22229=>"110010001",
  22230=>"111010100",
  22231=>"110011000",
  22232=>"010011111",
  22233=>"101111001",
  22234=>"001001101",
  22235=>"001111101",
  22236=>"101101100",
  22237=>"100010000",
  22238=>"111110111",
  22239=>"100011111",
  22240=>"011101011",
  22241=>"011010110",
  22242=>"101111111",
  22243=>"000011111",
  22244=>"101000110",
  22245=>"011011100",
  22246=>"110001001",
  22247=>"110110011",
  22248=>"111100101",
  22249=>"001100101",
  22250=>"011011111",
  22251=>"100110010",
  22252=>"101111001",
  22253=>"000000011",
  22254=>"101011110",
  22255=>"000011100",
  22256=>"001111000",
  22257=>"000000110",
  22258=>"111110011",
  22259=>"101001111",
  22260=>"111000001",
  22261=>"100101100",
  22262=>"111110011",
  22263=>"011001011",
  22264=>"011111100",
  22265=>"101000111",
  22266=>"100101010",
  22267=>"111000111",
  22268=>"100110001",
  22269=>"010010111",
  22270=>"010001110",
  22271=>"001110010",
  22272=>"010100010",
  22273=>"111000100",
  22274=>"001000010",
  22275=>"010000001",
  22276=>"110100000",
  22277=>"111101011",
  22278=>"101111100",
  22279=>"101110110",
  22280=>"011011010",
  22281=>"111100101",
  22282=>"110011101",
  22283=>"000110111",
  22284=>"011010011",
  22285=>"001001001",
  22286=>"111010011",
  22287=>"001000010",
  22288=>"011000010",
  22289=>"110000010",
  22290=>"011101010",
  22291=>"110000110",
  22292=>"011111111",
  22293=>"001010001",
  22294=>"010000000",
  22295=>"100101101",
  22296=>"001000111",
  22297=>"010101010",
  22298=>"001010111",
  22299=>"111011010",
  22300=>"111111010",
  22301=>"111011101",
  22302=>"010101101",
  22303=>"111110110",
  22304=>"111110011",
  22305=>"000100010",
  22306=>"001111010",
  22307=>"110101011",
  22308=>"000001001",
  22309=>"000111111",
  22310=>"011100010",
  22311=>"000110101",
  22312=>"101110010",
  22313=>"100000101",
  22314=>"011011000",
  22315=>"101001111",
  22316=>"101011100",
  22317=>"011100011",
  22318=>"000111011",
  22319=>"011101001",
  22320=>"000000011",
  22321=>"110111110",
  22322=>"000011001",
  22323=>"100110101",
  22324=>"000110100",
  22325=>"001100111",
  22326=>"010011000",
  22327=>"100001010",
  22328=>"011001111",
  22329=>"010110101",
  22330=>"010101001",
  22331=>"001110101",
  22332=>"101000010",
  22333=>"000001111",
  22334=>"100100000",
  22335=>"110101111",
  22336=>"111101001",
  22337=>"110111100",
  22338=>"011011000",
  22339=>"111111110",
  22340=>"001110011",
  22341=>"110010101",
  22342=>"000110111",
  22343=>"001101101",
  22344=>"000001001",
  22345=>"101010000",
  22346=>"011010100",
  22347=>"100001101",
  22348=>"010001110",
  22349=>"111110110",
  22350=>"100011111",
  22351=>"000011000",
  22352=>"110110010",
  22353=>"010001110",
  22354=>"010111011",
  22355=>"100111101",
  22356=>"000110011",
  22357=>"111110111",
  22358=>"011110011",
  22359=>"100110010",
  22360=>"001101010",
  22361=>"000000100",
  22362=>"111010010",
  22363=>"000100100",
  22364=>"000100000",
  22365=>"011000000",
  22366=>"000000011",
  22367=>"001000101",
  22368=>"100001010",
  22369=>"000110000",
  22370=>"010100111",
  22371=>"010110101",
  22372=>"101110101",
  22373=>"110111100",
  22374=>"001001000",
  22375=>"111101000",
  22376=>"010000001",
  22377=>"000011010",
  22378=>"001100100",
  22379=>"011000101",
  22380=>"111101101",
  22381=>"000110110",
  22382=>"100111000",
  22383=>"111011011",
  22384=>"111000010",
  22385=>"101000001",
  22386=>"010000011",
  22387=>"011110111",
  22388=>"000001011",
  22389=>"000011000",
  22390=>"011010011",
  22391=>"011101100",
  22392=>"101110011",
  22393=>"101111000",
  22394=>"100011101",
  22395=>"101001000",
  22396=>"000011100",
  22397=>"110101000",
  22398=>"100000011",
  22399=>"110001000",
  22400=>"001110111",
  22401=>"000001110",
  22402=>"111011111",
  22403=>"101011101",
  22404=>"110111100",
  22405=>"000010011",
  22406=>"011010011",
  22407=>"001101010",
  22408=>"101001010",
  22409=>"001000000",
  22410=>"000010010",
  22411=>"010110011",
  22412=>"000101011",
  22413=>"000010010",
  22414=>"101011001",
  22415=>"100110111",
  22416=>"111001111",
  22417=>"011000001",
  22418=>"000010110",
  22419=>"100110101",
  22420=>"011010001",
  22421=>"000001010",
  22422=>"101100111",
  22423=>"111001010",
  22424=>"101011000",
  22425=>"000101100",
  22426=>"011111011",
  22427=>"100010111",
  22428=>"100011000",
  22429=>"100100101",
  22430=>"101101101",
  22431=>"001011010",
  22432=>"101010000",
  22433=>"101100000",
  22434=>"011101101",
  22435=>"001001000",
  22436=>"010010100",
  22437=>"110001101",
  22438=>"001011100",
  22439=>"010100101",
  22440=>"000101011",
  22441=>"100111001",
  22442=>"011001101",
  22443=>"110001111",
  22444=>"000001001",
  22445=>"001001110",
  22446=>"000001110",
  22447=>"001010100",
  22448=>"000010100",
  22449=>"111110111",
  22450=>"110110110",
  22451=>"100011110",
  22452=>"010001001",
  22453=>"111010001",
  22454=>"111010111",
  22455=>"001111010",
  22456=>"100110011",
  22457=>"010011101",
  22458=>"100101111",
  22459=>"010011110",
  22460=>"111011000",
  22461=>"111010000",
  22462=>"010101011",
  22463=>"100010000",
  22464=>"000001100",
  22465=>"110000010",
  22466=>"011101011",
  22467=>"011011111",
  22468=>"010110110",
  22469=>"001101001",
  22470=>"010010100",
  22471=>"110111100",
  22472=>"001000001",
  22473=>"100001101",
  22474=>"100111111",
  22475=>"110100011",
  22476=>"110111101",
  22477=>"111111101",
  22478=>"110111100",
  22479=>"010001000",
  22480=>"001110110",
  22481=>"100001011",
  22482=>"111000011",
  22483=>"001100111",
  22484=>"000011100",
  22485=>"000000110",
  22486=>"110110110",
  22487=>"101110111",
  22488=>"111001110",
  22489=>"101101111",
  22490=>"100011000",
  22491=>"000101000",
  22492=>"011100100",
  22493=>"000111010",
  22494=>"011001100",
  22495=>"000011000",
  22496=>"110000100",
  22497=>"000110101",
  22498=>"011011111",
  22499=>"111101001",
  22500=>"011100110",
  22501=>"010111001",
  22502=>"010100100",
  22503=>"101011001",
  22504=>"111100001",
  22505=>"000011000",
  22506=>"000111001",
  22507=>"000011111",
  22508=>"011010010",
  22509=>"101001100",
  22510=>"011010110",
  22511=>"011110110",
  22512=>"110010111",
  22513=>"111000100",
  22514=>"111001100",
  22515=>"010000100",
  22516=>"100111011",
  22517=>"100001101",
  22518=>"000111001",
  22519=>"000000001",
  22520=>"101110101",
  22521=>"001010001",
  22522=>"011111101",
  22523=>"101100011",
  22524=>"110101110",
  22525=>"001000010",
  22526=>"010001001",
  22527=>"001011111",
  22528=>"010000110",
  22529=>"010000001",
  22530=>"000110100",
  22531=>"011101010",
  22532=>"011111011",
  22533=>"000101011",
  22534=>"001111110",
  22535=>"010001010",
  22536=>"100001000",
  22537=>"100011011",
  22538=>"000011010",
  22539=>"100010100",
  22540=>"010001110",
  22541=>"101000101",
  22542=>"011011010",
  22543=>"000101000",
  22544=>"100010001",
  22545=>"011011110",
  22546=>"001110010",
  22547=>"011010100",
  22548=>"000111101",
  22549=>"010000001",
  22550=>"101011101",
  22551=>"011010000",
  22552=>"000011100",
  22553=>"100101000",
  22554=>"000101111",
  22555=>"110101100",
  22556=>"100101001",
  22557=>"101100101",
  22558=>"110000000",
  22559=>"000011011",
  22560=>"101010111",
  22561=>"000000101",
  22562=>"001100101",
  22563=>"001101000",
  22564=>"100111111",
  22565=>"010110110",
  22566=>"100011011",
  22567=>"000110100",
  22568=>"000011000",
  22569=>"010011100",
  22570=>"111011110",
  22571=>"010011011",
  22572=>"110010001",
  22573=>"011101110",
  22574=>"001110011",
  22575=>"111111101",
  22576=>"101001000",
  22577=>"111000101",
  22578=>"000111101",
  22579=>"011110101",
  22580=>"001001000",
  22581=>"001001001",
  22582=>"011101101",
  22583=>"100111101",
  22584=>"000110011",
  22585=>"000110110",
  22586=>"100111110",
  22587=>"000000100",
  22588=>"000111010",
  22589=>"001000110",
  22590=>"101101010",
  22591=>"001000101",
  22592=>"001101110",
  22593=>"111101101",
  22594=>"001111010",
  22595=>"111010111",
  22596=>"100101100",
  22597=>"010000111",
  22598=>"101010100",
  22599=>"011111110",
  22600=>"100010010",
  22601=>"110111010",
  22602=>"010010010",
  22603=>"001000001",
  22604=>"000100111",
  22605=>"111100011",
  22606=>"111011010",
  22607=>"000110000",
  22608=>"001111001",
  22609=>"001110000",
  22610=>"100001110",
  22611=>"101101000",
  22612=>"110101010",
  22613=>"110111011",
  22614=>"101110111",
  22615=>"011011100",
  22616=>"110111011",
  22617=>"111101111",
  22618=>"110001011",
  22619=>"000000001",
  22620=>"000001100",
  22621=>"001011100",
  22622=>"001000000",
  22623=>"010001000",
  22624=>"011101010",
  22625=>"001000010",
  22626=>"010101110",
  22627=>"010110001",
  22628=>"100000011",
  22629=>"000110101",
  22630=>"010101101",
  22631=>"000100111",
  22632=>"011111000",
  22633=>"001111100",
  22634=>"100001011",
  22635=>"110110101",
  22636=>"110011010",
  22637=>"111000000",
  22638=>"000111011",
  22639=>"000011110",
  22640=>"010111000",
  22641=>"010111010",
  22642=>"000100010",
  22643=>"110010110",
  22644=>"000110011",
  22645=>"101011110",
  22646=>"010001001",
  22647=>"010100111",
  22648=>"010111110",
  22649=>"011111111",
  22650=>"000111011",
  22651=>"001000000",
  22652=>"100111110",
  22653=>"001000000",
  22654=>"010001100",
  22655=>"001011011",
  22656=>"110100111",
  22657=>"000000011",
  22658=>"111110110",
  22659=>"101001010",
  22660=>"110110011",
  22661=>"101010011",
  22662=>"001010000",
  22663=>"110001111",
  22664=>"101110000",
  22665=>"001000100",
  22666=>"100001000",
  22667=>"010110110",
  22668=>"110110100",
  22669=>"101110100",
  22670=>"101001001",
  22671=>"010101000",
  22672=>"011111001",
  22673=>"101101100",
  22674=>"000101111",
  22675=>"111001111",
  22676=>"001000100",
  22677=>"111101110",
  22678=>"111001001",
  22679=>"101011110",
  22680=>"111000100",
  22681=>"100111100",
  22682=>"101010101",
  22683=>"011010000",
  22684=>"011111100",
  22685=>"100001001",
  22686=>"010001111",
  22687=>"010100001",
  22688=>"100010001",
  22689=>"101101100",
  22690=>"100101110",
  22691=>"100110100",
  22692=>"001101110",
  22693=>"011110111",
  22694=>"001101001",
  22695=>"000100011",
  22696=>"111011010",
  22697=>"100011000",
  22698=>"111001111",
  22699=>"011110100",
  22700=>"011101111",
  22701=>"110101100",
  22702=>"001001101",
  22703=>"111101011",
  22704=>"011101000",
  22705=>"010011011",
  22706=>"110110110",
  22707=>"000101000",
  22708=>"000011111",
  22709=>"011011000",
  22710=>"011111110",
  22711=>"010111100",
  22712=>"101001000",
  22713=>"110100101",
  22714=>"010001111",
  22715=>"011101100",
  22716=>"101101000",
  22717=>"011110101",
  22718=>"111100101",
  22719=>"101100100",
  22720=>"100001101",
  22721=>"100101010",
  22722=>"111001101",
  22723=>"001010110",
  22724=>"111001010",
  22725=>"001100110",
  22726=>"111011110",
  22727=>"110001110",
  22728=>"100110111",
  22729=>"101010111",
  22730=>"110100000",
  22731=>"101000011",
  22732=>"110100110",
  22733=>"011100011",
  22734=>"010110010",
  22735=>"000011000",
  22736=>"101001110",
  22737=>"000010101",
  22738=>"101001110",
  22739=>"000111111",
  22740=>"010100011",
  22741=>"001000101",
  22742=>"100111000",
  22743=>"110010111",
  22744=>"010001001",
  22745=>"000010111",
  22746=>"010111001",
  22747=>"100011110",
  22748=>"011000011",
  22749=>"111110110",
  22750=>"011001010",
  22751=>"001111010",
  22752=>"001011110",
  22753=>"010000100",
  22754=>"000100110",
  22755=>"011000011",
  22756=>"101000000",
  22757=>"000100111",
  22758=>"001010101",
  22759=>"100110100",
  22760=>"101011000",
  22761=>"100001100",
  22762=>"000101101",
  22763=>"111111111",
  22764=>"011100110",
  22765=>"001101100",
  22766=>"010011100",
  22767=>"001011010",
  22768=>"001110001",
  22769=>"001011111",
  22770=>"000001101",
  22771=>"100111100",
  22772=>"101010000",
  22773=>"001010010",
  22774=>"111001111",
  22775=>"001100110",
  22776=>"101101110",
  22777=>"001110000",
  22778=>"000001101",
  22779=>"010000000",
  22780=>"101000100",
  22781=>"000101000",
  22782=>"000100111",
  22783=>"111111110",
  22784=>"010011111",
  22785=>"100100000",
  22786=>"000100101",
  22787=>"001001000",
  22788=>"000110010",
  22789=>"001000100",
  22790=>"101100110",
  22791=>"000101100",
  22792=>"101000011",
  22793=>"000101110",
  22794=>"101101001",
  22795=>"110010000",
  22796=>"001000000",
  22797=>"110101100",
  22798=>"100101101",
  22799=>"000010111",
  22800=>"101011011",
  22801=>"110000111",
  22802=>"010100000",
  22803=>"000000000",
  22804=>"110111111",
  22805=>"001101101",
  22806=>"010101101",
  22807=>"000101101",
  22808=>"011001000",
  22809=>"101111101",
  22810=>"101110101",
  22811=>"111101111",
  22812=>"100101110",
  22813=>"011101111",
  22814=>"011111100",
  22815=>"000011011",
  22816=>"000100011",
  22817=>"000111011",
  22818=>"001001110",
  22819=>"110100001",
  22820=>"000100101",
  22821=>"100111010",
  22822=>"001101110",
  22823=>"101101100",
  22824=>"100101111",
  22825=>"000000010",
  22826=>"100000111",
  22827=>"101000010",
  22828=>"010000010",
  22829=>"110010111",
  22830=>"101000011",
  22831=>"011011001",
  22832=>"100100101",
  22833=>"010000000",
  22834=>"111010100",
  22835=>"010001111",
  22836=>"100000101",
  22837=>"100011110",
  22838=>"001001100",
  22839=>"101011100",
  22840=>"011110111",
  22841=>"011110000",
  22842=>"100111000",
  22843=>"010000010",
  22844=>"011001110",
  22845=>"101101011",
  22846=>"001111011",
  22847=>"101110110",
  22848=>"011100100",
  22849=>"110100110",
  22850=>"110110100",
  22851=>"000001000",
  22852=>"001100100",
  22853=>"000010001",
  22854=>"010100111",
  22855=>"100110001",
  22856=>"101000001",
  22857=>"011001000",
  22858=>"101010111",
  22859=>"100000001",
  22860=>"010110111",
  22861=>"111101010",
  22862=>"000000010",
  22863=>"101111110",
  22864=>"100000101",
  22865=>"011100111",
  22866=>"001000011",
  22867=>"100110110",
  22868=>"000010101",
  22869=>"000001111",
  22870=>"111111000",
  22871=>"100111010",
  22872=>"011011001",
  22873=>"010010111",
  22874=>"011111111",
  22875=>"010001101",
  22876=>"101011100",
  22877=>"111001010",
  22878=>"011111110",
  22879=>"111110101",
  22880=>"011111101",
  22881=>"000011000",
  22882=>"100110111",
  22883=>"001001100",
  22884=>"011011100",
  22885=>"001111011",
  22886=>"010011101",
  22887=>"111100110",
  22888=>"000111011",
  22889=>"010100100",
  22890=>"010000000",
  22891=>"111000011",
  22892=>"000100100",
  22893=>"000100011",
  22894=>"010111110",
  22895=>"101010101",
  22896=>"010101111",
  22897=>"101101110",
  22898=>"000011000",
  22899=>"111100001",
  22900=>"110111111",
  22901=>"101100101",
  22902=>"100011110",
  22903=>"000101001",
  22904=>"100110011",
  22905=>"001010010",
  22906=>"010010011",
  22907=>"111010101",
  22908=>"101111100",
  22909=>"110011010",
  22910=>"100011101",
  22911=>"111000100",
  22912=>"010001100",
  22913=>"000100100",
  22914=>"100011010",
  22915=>"000101110",
  22916=>"001110101",
  22917=>"001011100",
  22918=>"100110101",
  22919=>"111000110",
  22920=>"011011000",
  22921=>"000110111",
  22922=>"000000000",
  22923=>"000101111",
  22924=>"010110110",
  22925=>"001000011",
  22926=>"010100110",
  22927=>"101010100",
  22928=>"001000001",
  22929=>"000000001",
  22930=>"010001001",
  22931=>"110000110",
  22932=>"010000000",
  22933=>"010011001",
  22934=>"011001001",
  22935=>"000001110",
  22936=>"001110111",
  22937=>"000101001",
  22938=>"111010000",
  22939=>"000111010",
  22940=>"011101010",
  22941=>"100010010",
  22942=>"000110000",
  22943=>"111010111",
  22944=>"111101000",
  22945=>"110010010",
  22946=>"001000000",
  22947=>"010111010",
  22948=>"011000010",
  22949=>"100000000",
  22950=>"110010001",
  22951=>"010011000",
  22952=>"100110101",
  22953=>"010001111",
  22954=>"001101111",
  22955=>"110000100",
  22956=>"100101100",
  22957=>"011110100",
  22958=>"010011010",
  22959=>"001100011",
  22960=>"101000100",
  22961=>"000000111",
  22962=>"101110000",
  22963=>"111110001",
  22964=>"100100011",
  22965=>"001011000",
  22966=>"011111110",
  22967=>"101111111",
  22968=>"011101001",
  22969=>"010001110",
  22970=>"100100010",
  22971=>"000010110",
  22972=>"111101111",
  22973=>"100001001",
  22974=>"100011000",
  22975=>"111010101",
  22976=>"110001111",
  22977=>"111010100",
  22978=>"110000101",
  22979=>"000110001",
  22980=>"110100100",
  22981=>"010111111",
  22982=>"110110010",
  22983=>"010110010",
  22984=>"111110101",
  22985=>"101010111",
  22986=>"111001101",
  22987=>"000111111",
  22988=>"100110100",
  22989=>"111011011",
  22990=>"001110000",
  22991=>"111111111",
  22992=>"100110111",
  22993=>"011001110",
  22994=>"011011101",
  22995=>"101111111",
  22996=>"010110110",
  22997=>"111101100",
  22998=>"101001011",
  22999=>"111010110",
  23000=>"110100110",
  23001=>"110001101",
  23002=>"111111000",
  23003=>"110101111",
  23004=>"111100011",
  23005=>"111101010",
  23006=>"101011101",
  23007=>"001010100",
  23008=>"010111101",
  23009=>"111010111",
  23010=>"000011110",
  23011=>"011100100",
  23012=>"001010111",
  23013=>"111100001",
  23014=>"000100010",
  23015=>"111111010",
  23016=>"010011000",
  23017=>"011101010",
  23018=>"010011011",
  23019=>"111000010",
  23020=>"011000010",
  23021=>"101010110",
  23022=>"110011110",
  23023=>"010010100",
  23024=>"100100110",
  23025=>"000111100",
  23026=>"101000010",
  23027=>"011110111",
  23028=>"000010100",
  23029=>"000010011",
  23030=>"001100000",
  23031=>"111010001",
  23032=>"110100011",
  23033=>"111001110",
  23034=>"000001001",
  23035=>"101011010",
  23036=>"011011111",
  23037=>"011000110",
  23038=>"010000010",
  23039=>"010000101",
  23040=>"010000100",
  23041=>"011001111",
  23042=>"011110001",
  23043=>"011101000",
  23044=>"000000011",
  23045=>"100110110",
  23046=>"110010011",
  23047=>"100000111",
  23048=>"000111010",
  23049=>"000111011",
  23050=>"011101110",
  23051=>"001100000",
  23052=>"101011011",
  23053=>"010100000",
  23054=>"101011000",
  23055=>"011011001",
  23056=>"011111001",
  23057=>"010110011",
  23058=>"010011101",
  23059=>"101100101",
  23060=>"000111101",
  23061=>"000000011",
  23062=>"110110010",
  23063=>"110000110",
  23064=>"010101000",
  23065=>"001001000",
  23066=>"011101101",
  23067=>"011000110",
  23068=>"000001010",
  23069=>"000000000",
  23070=>"101100010",
  23071=>"100110101",
  23072=>"001111010",
  23073=>"011110001",
  23074=>"000101000",
  23075=>"100011100",
  23076=>"110110001",
  23077=>"000000001",
  23078=>"000111100",
  23079=>"110001001",
  23080=>"100001010",
  23081=>"100001110",
  23082=>"110100011",
  23083=>"101111010",
  23084=>"111001101",
  23085=>"001011110",
  23086=>"011101000",
  23087=>"000001001",
  23088=>"110111101",
  23089=>"001000101",
  23090=>"100010000",
  23091=>"001111011",
  23092=>"100000001",
  23093=>"001100110",
  23094=>"010111011",
  23095=>"000111101",
  23096=>"010101000",
  23097=>"100100110",
  23098=>"000110010",
  23099=>"011010001",
  23100=>"111110100",
  23101=>"010011010",
  23102=>"000101000",
  23103=>"011000111",
  23104=>"110011111",
  23105=>"001111101",
  23106=>"010001100",
  23107=>"001000001",
  23108=>"011100000",
  23109=>"011010010",
  23110=>"001010010",
  23111=>"001001001",
  23112=>"011011111",
  23113=>"000101110",
  23114=>"110010100",
  23115=>"101110001",
  23116=>"001101000",
  23117=>"101111110",
  23118=>"111100111",
  23119=>"000000111",
  23120=>"101011111",
  23121=>"101100111",
  23122=>"010010011",
  23123=>"011110110",
  23124=>"111001010",
  23125=>"101000010",
  23126=>"000110110",
  23127=>"001011111",
  23128=>"100101110",
  23129=>"101101010",
  23130=>"011011011",
  23131=>"100001101",
  23132=>"000010000",
  23133=>"010000011",
  23134=>"001011100",
  23135=>"010101100",
  23136=>"011011101",
  23137=>"111101101",
  23138=>"110110100",
  23139=>"001111101",
  23140=>"011011111",
  23141=>"111000011",
  23142=>"000101110",
  23143=>"000100101",
  23144=>"001110100",
  23145=>"011000110",
  23146=>"001100111",
  23147=>"010110011",
  23148=>"000010001",
  23149=>"010101110",
  23150=>"110010110",
  23151=>"101100110",
  23152=>"010100010",
  23153=>"101101100",
  23154=>"110100110",
  23155=>"010010111",
  23156=>"011010011",
  23157=>"111010011",
  23158=>"000000110",
  23159=>"011111010",
  23160=>"100001101",
  23161=>"000110001",
  23162=>"111110100",
  23163=>"000110100",
  23164=>"001100101",
  23165=>"010101010",
  23166=>"100001001",
  23167=>"010100101",
  23168=>"101101001",
  23169=>"111010011",
  23170=>"011001001",
  23171=>"111011000",
  23172=>"101110110",
  23173=>"101111010",
  23174=>"001000011",
  23175=>"011010111",
  23176=>"011010011",
  23177=>"101001100",
  23178=>"010111101",
  23179=>"101101111",
  23180=>"110110001",
  23181=>"010110110",
  23182=>"111001000",
  23183=>"111111101",
  23184=>"000010100",
  23185=>"111010111",
  23186=>"011011000",
  23187=>"100011111",
  23188=>"101111111",
  23189=>"000111111",
  23190=>"001011110",
  23191=>"110001000",
  23192=>"010111110",
  23193=>"000100001",
  23194=>"101000000",
  23195=>"011110101",
  23196=>"010101110",
  23197=>"111101001",
  23198=>"110010111",
  23199=>"000001011",
  23200=>"001101001",
  23201=>"011111010",
  23202=>"011100100",
  23203=>"111100101",
  23204=>"001000101",
  23205=>"011111111",
  23206=>"000000011",
  23207=>"001100001",
  23208=>"010000000",
  23209=>"010111011",
  23210=>"101111111",
  23211=>"111101110",
  23212=>"011010011",
  23213=>"101111111",
  23214=>"001000010",
  23215=>"110000110",
  23216=>"110110001",
  23217=>"010000100",
  23218=>"000101100",
  23219=>"011011000",
  23220=>"101011011",
  23221=>"010101111",
  23222=>"010010011",
  23223=>"000001010",
  23224=>"100100100",
  23225=>"111101110",
  23226=>"011010001",
  23227=>"111000001",
  23228=>"001111101",
  23229=>"000010010",
  23230=>"001000100",
  23231=>"000100110",
  23232=>"101011110",
  23233=>"100010110",
  23234=>"001100000",
  23235=>"101000111",
  23236=>"001101001",
  23237=>"010101001",
  23238=>"010010011",
  23239=>"000101101",
  23240=>"001100001",
  23241=>"000001000",
  23242=>"010111011",
  23243=>"001001100",
  23244=>"000001011",
  23245=>"110011111",
  23246=>"010100111",
  23247=>"001101010",
  23248=>"110111111",
  23249=>"100101000",
  23250=>"011101000",
  23251=>"011011001",
  23252=>"000111110",
  23253=>"010110110",
  23254=>"011110101",
  23255=>"111010101",
  23256=>"010100000",
  23257=>"011110010",
  23258=>"000010001",
  23259=>"001111111",
  23260=>"110001111",
  23261=>"010111010",
  23262=>"010101101",
  23263=>"010000100",
  23264=>"001100110",
  23265=>"100000110",
  23266=>"010101110",
  23267=>"001101000",
  23268=>"110100110",
  23269=>"000011110",
  23270=>"001111000",
  23271=>"000010011",
  23272=>"010111001",
  23273=>"010000111",
  23274=>"101100000",
  23275=>"010001101",
  23276=>"000100010",
  23277=>"101001000",
  23278=>"101110111",
  23279=>"111000101",
  23280=>"100011101",
  23281=>"111100011",
  23282=>"111101001",
  23283=>"101011011",
  23284=>"111000010",
  23285=>"000010000",
  23286=>"111001101",
  23287=>"101000011",
  23288=>"100010110",
  23289=>"111010010",
  23290=>"101101000",
  23291=>"011000111",
  23292=>"000010001",
  23293=>"000101010",
  23294=>"011000001",
  23295=>"000100010",
  23296=>"111001110",
  23297=>"111111011",
  23298=>"101101101",
  23299=>"001111001",
  23300=>"010110110",
  23301=>"000010100",
  23302=>"011001111",
  23303=>"111011110",
  23304=>"100100011",
  23305=>"001101001",
  23306=>"001111011",
  23307=>"001001110",
  23308=>"001010000",
  23309=>"111001100",
  23310=>"110111010",
  23311=>"001010001",
  23312=>"000110101",
  23313=>"011110101",
  23314=>"001110000",
  23315=>"100111100",
  23316=>"011001010",
  23317=>"010010001",
  23318=>"101110101",
  23319=>"000000101",
  23320=>"000000100",
  23321=>"111011010",
  23322=>"101100001",
  23323=>"110010101",
  23324=>"011010100",
  23325=>"010110000",
  23326=>"000100000",
  23327=>"111010010",
  23328=>"111010011",
  23329=>"111000101",
  23330=>"101010010",
  23331=>"100011111",
  23332=>"111001001",
  23333=>"111010111",
  23334=>"011001000",
  23335=>"000111001",
  23336=>"000100101",
  23337=>"101100001",
  23338=>"000101110",
  23339=>"100101101",
  23340=>"110011010",
  23341=>"101011101",
  23342=>"000111000",
  23343=>"111111000",
  23344=>"101110101",
  23345=>"110000100",
  23346=>"101100000",
  23347=>"100000100",
  23348=>"010100011",
  23349=>"101100100",
  23350=>"010001001",
  23351=>"100110000",
  23352=>"001110111",
  23353=>"110011100",
  23354=>"011000011",
  23355=>"111110110",
  23356=>"000001000",
  23357=>"010010101",
  23358=>"111100010",
  23359=>"011110101",
  23360=>"001100010",
  23361=>"010101110",
  23362=>"101001011",
  23363=>"001011100",
  23364=>"001000101",
  23365=>"111111100",
  23366=>"000111110",
  23367=>"000111110",
  23368=>"010101111",
  23369=>"111111011",
  23370=>"101110011",
  23371=>"100101100",
  23372=>"111111110",
  23373=>"110000101",
  23374=>"110000101",
  23375=>"100100111",
  23376=>"000111100",
  23377=>"111110010",
  23378=>"011001001",
  23379=>"011000011",
  23380=>"000101011",
  23381=>"111100111",
  23382=>"001001011",
  23383=>"011010100",
  23384=>"011111010",
  23385=>"001111110",
  23386=>"111101011",
  23387=>"101100100",
  23388=>"000011111",
  23389=>"111001111",
  23390=>"101001110",
  23391=>"000101001",
  23392=>"010001001",
  23393=>"101111010",
  23394=>"100110110",
  23395=>"001100010",
  23396=>"100100010",
  23397=>"111010010",
  23398=>"101000000",
  23399=>"000110011",
  23400=>"110010011",
  23401=>"011011001",
  23402=>"010110100",
  23403=>"011111101",
  23404=>"011111100",
  23405=>"000011001",
  23406=>"100111101",
  23407=>"000101001",
  23408=>"111100000",
  23409=>"011101010",
  23410=>"101011110",
  23411=>"101001001",
  23412=>"000111010",
  23413=>"110011111",
  23414=>"100011011",
  23415=>"100111000",
  23416=>"100000001",
  23417=>"000011001",
  23418=>"001101100",
  23419=>"000101101",
  23420=>"001110011",
  23421=>"110101101",
  23422=>"101101101",
  23423=>"010010100",
  23424=>"110111000",
  23425=>"100010001",
  23426=>"100100111",
  23427=>"010110111",
  23428=>"111101011",
  23429=>"001010011",
  23430=>"111100110",
  23431=>"011101110",
  23432=>"000000010",
  23433=>"001001101",
  23434=>"001000111",
  23435=>"001111100",
  23436=>"100111111",
  23437=>"100110000",
  23438=>"101111111",
  23439=>"001000101",
  23440=>"101010101",
  23441=>"010001100",
  23442=>"000010000",
  23443=>"111111100",
  23444=>"110010101",
  23445=>"000111100",
  23446=>"110000100",
  23447=>"011000110",
  23448=>"010100011",
  23449=>"110011100",
  23450=>"110111001",
  23451=>"000000101",
  23452=>"100100111",
  23453=>"111111001",
  23454=>"101100110",
  23455=>"001111000",
  23456=>"001010010",
  23457=>"110000001",
  23458=>"000111010",
  23459=>"000011101",
  23460=>"000010001",
  23461=>"101110101",
  23462=>"001000110",
  23463=>"010111000",
  23464=>"010111100",
  23465=>"101000101",
  23466=>"110001101",
  23467=>"000010110",
  23468=>"000100001",
  23469=>"000000110",
  23470=>"110011000",
  23471=>"110100001",
  23472=>"101100101",
  23473=>"111000111",
  23474=>"001101101",
  23475=>"011000111",
  23476=>"011001110",
  23477=>"101100111",
  23478=>"101101100",
  23479=>"010111100",
  23480=>"101111100",
  23481=>"110010110",
  23482=>"101100101",
  23483=>"100010000",
  23484=>"011111111",
  23485=>"111100001",
  23486=>"110110111",
  23487=>"100100001",
  23488=>"011010011",
  23489=>"000000100",
  23490=>"110110101",
  23491=>"110101001",
  23492=>"010000111",
  23493=>"010101011",
  23494=>"010010000",
  23495=>"001110001",
  23496=>"010001010",
  23497=>"000101110",
  23498=>"110101001",
  23499=>"100000111",
  23500=>"111101011",
  23501=>"100000111",
  23502=>"001111010",
  23503=>"110001110",
  23504=>"110111101",
  23505=>"010110101",
  23506=>"101111110",
  23507=>"101001001",
  23508=>"011100110",
  23509=>"110001100",
  23510=>"110111110",
  23511=>"100100000",
  23512=>"100011001",
  23513=>"001101101",
  23514=>"101101011",
  23515=>"000001001",
  23516=>"111110101",
  23517=>"100010010",
  23518=>"110111011",
  23519=>"100101111",
  23520=>"101100110",
  23521=>"111011110",
  23522=>"010111001",
  23523=>"110111100",
  23524=>"010110110",
  23525=>"000101001",
  23526=>"100100011",
  23527=>"000000101",
  23528=>"110001010",
  23529=>"000101010",
  23530=>"010011100",
  23531=>"110011010",
  23532=>"110010110",
  23533=>"100010001",
  23534=>"011001010",
  23535=>"000011001",
  23536=>"110011110",
  23537=>"110111000",
  23538=>"000110110",
  23539=>"110010111",
  23540=>"001110100",
  23541=>"010101010",
  23542=>"011111000",
  23543=>"101111100",
  23544=>"010000100",
  23545=>"001011000",
  23546=>"100001010",
  23547=>"011000001",
  23548=>"001101110",
  23549=>"000101000",
  23550=>"001010011",
  23551=>"100010011",
  23552=>"001000101",
  23553=>"111011011",
  23554=>"000011001",
  23555=>"010100011",
  23556=>"110000001",
  23557=>"011000101",
  23558=>"001000101",
  23559=>"111000011",
  23560=>"100101110",
  23561=>"110000110",
  23562=>"111011110",
  23563=>"110110111",
  23564=>"011100001",
  23565=>"011110011",
  23566=>"011111101",
  23567=>"111110101",
  23568=>"000110111",
  23569=>"101110100",
  23570=>"010000011",
  23571=>"110010011",
  23572=>"011001001",
  23573=>"000100011",
  23574=>"111111110",
  23575=>"100101010",
  23576=>"101000001",
  23577=>"110000111",
  23578=>"110100001",
  23579=>"001101111",
  23580=>"111011001",
  23581=>"001000001",
  23582=>"000000001",
  23583=>"110101101",
  23584=>"011001000",
  23585=>"101000101",
  23586=>"111010110",
  23587=>"001000110",
  23588=>"111000010",
  23589=>"001000000",
  23590=>"000110110",
  23591=>"111011000",
  23592=>"000100111",
  23593=>"010001001",
  23594=>"010000111",
  23595=>"101110101",
  23596=>"000010110",
  23597=>"100001011",
  23598=>"111101101",
  23599=>"010001000",
  23600=>"101111010",
  23601=>"101111111",
  23602=>"101001110",
  23603=>"000111010",
  23604=>"111000000",
  23605=>"101111000",
  23606=>"110110000",
  23607=>"101000010",
  23608=>"110111010",
  23609=>"100010011",
  23610=>"000101000",
  23611=>"001111000",
  23612=>"000100011",
  23613=>"000000010",
  23614=>"001111001",
  23615=>"011101101",
  23616=>"000111111",
  23617=>"001111001",
  23618=>"001010100",
  23619=>"011111000",
  23620=>"100010011",
  23621=>"001111110",
  23622=>"000100001",
  23623=>"001111001",
  23624=>"010010011",
  23625=>"111111100",
  23626=>"011101000",
  23627=>"011100000",
  23628=>"100011010",
  23629=>"010111110",
  23630=>"001100000",
  23631=>"100011010",
  23632=>"000011100",
  23633=>"001111110",
  23634=>"111111001",
  23635=>"110010011",
  23636=>"110100001",
  23637=>"000111011",
  23638=>"110011110",
  23639=>"100101100",
  23640=>"110101111",
  23641=>"110000111",
  23642=>"000001111",
  23643=>"110101101",
  23644=>"001111001",
  23645=>"111110000",
  23646=>"110111101",
  23647=>"011001100",
  23648=>"001010010",
  23649=>"010011100",
  23650=>"010110100",
  23651=>"101100011",
  23652=>"100100101",
  23653=>"111111011",
  23654=>"011011001",
  23655=>"111111111",
  23656=>"011100000",
  23657=>"101011000",
  23658=>"000000010",
  23659=>"110010010",
  23660=>"001000001",
  23661=>"100001011",
  23662=>"011111001",
  23663=>"000001011",
  23664=>"111010101",
  23665=>"001010000",
  23666=>"100101011",
  23667=>"111100110",
  23668=>"011001110",
  23669=>"100000101",
  23670=>"100110110",
  23671=>"101111010",
  23672=>"111110001",
  23673=>"111110111",
  23674=>"101010011",
  23675=>"101000001",
  23676=>"100001001",
  23677=>"000000000",
  23678=>"111110010",
  23679=>"100010000",
  23680=>"101010000",
  23681=>"111110101",
  23682=>"010100110",
  23683=>"010101001",
  23684=>"111100010",
  23685=>"100011010",
  23686=>"110111011",
  23687=>"101110011",
  23688=>"100111001",
  23689=>"110000001",
  23690=>"100001011",
  23691=>"101011011",
  23692=>"011110001",
  23693=>"110010101",
  23694=>"001010010",
  23695=>"100111100",
  23696=>"011001000",
  23697=>"100011100",
  23698=>"000000010",
  23699=>"011110101",
  23700=>"011000111",
  23701=>"001000110",
  23702=>"001010100",
  23703=>"000101111",
  23704=>"101011010",
  23705=>"001110100",
  23706=>"110001110",
  23707=>"110001110",
  23708=>"000110100",
  23709=>"110100000",
  23710=>"101010100",
  23711=>"010000010",
  23712=>"100011111",
  23713=>"010110010",
  23714=>"000100100",
  23715=>"011011111",
  23716=>"101100100",
  23717=>"001010010",
  23718=>"000111001",
  23719=>"010100011",
  23720=>"110100100",
  23721=>"111000011",
  23722=>"000101001",
  23723=>"001001111",
  23724=>"100100000",
  23725=>"110101010",
  23726=>"010001100",
  23727=>"001010011",
  23728=>"010111000",
  23729=>"111011010",
  23730=>"011001011",
  23731=>"010000001",
  23732=>"001001001",
  23733=>"111110001",
  23734=>"001110011",
  23735=>"111110100",
  23736=>"000101011",
  23737=>"101010101",
  23738=>"010110100",
  23739=>"110101011",
  23740=>"001010101",
  23741=>"100100111",
  23742=>"101110011",
  23743=>"100001000",
  23744=>"001101010",
  23745=>"001000101",
  23746=>"001001111",
  23747=>"010110010",
  23748=>"111101010",
  23749=>"000001010",
  23750=>"110101100",
  23751=>"001110101",
  23752=>"101110011",
  23753=>"111111001",
  23754=>"001100100",
  23755=>"001111111",
  23756=>"110001010",
  23757=>"101001110",
  23758=>"001001101",
  23759=>"111010101",
  23760=>"101111110",
  23761=>"010010000",
  23762=>"111111010",
  23763=>"111101010",
  23764=>"000001011",
  23765=>"111001000",
  23766=>"100001011",
  23767=>"011011000",
  23768=>"011101110",
  23769=>"010010011",
  23770=>"000100100",
  23771=>"111110111",
  23772=>"000000111",
  23773=>"000111001",
  23774=>"001110001",
  23775=>"010011111",
  23776=>"000111001",
  23777=>"100111110",
  23778=>"010000100",
  23779=>"000111110",
  23780=>"001011011",
  23781=>"100100010",
  23782=>"101010101",
  23783=>"011101001",
  23784=>"000001100",
  23785=>"101011100",
  23786=>"011001111",
  23787=>"101110111",
  23788=>"000011100",
  23789=>"100000010",
  23790=>"100010001",
  23791=>"010000000",
  23792=>"001111100",
  23793=>"001000000",
  23794=>"100000110",
  23795=>"001101011",
  23796=>"001000011",
  23797=>"101001011",
  23798=>"001111001",
  23799=>"100111100",
  23800=>"101000000",
  23801=>"111100000",
  23802=>"101000100",
  23803=>"001000001",
  23804=>"010000001",
  23805=>"111011110",
  23806=>"010111010",
  23807=>"111010101",
  23808=>"110011110",
  23809=>"110111101",
  23810=>"101010101",
  23811=>"110111110",
  23812=>"000011110",
  23813=>"011000001",
  23814=>"000000101",
  23815=>"111101101",
  23816=>"001111010",
  23817=>"001001111",
  23818=>"101111000",
  23819=>"011100110",
  23820=>"010011011",
  23821=>"000111011",
  23822=>"100001011",
  23823=>"011110110",
  23824=>"101100111",
  23825=>"001011001",
  23826=>"001000100",
  23827=>"111011010",
  23828=>"010000000",
  23829=>"010001100",
  23830=>"010110011",
  23831=>"011000001",
  23832=>"011111011",
  23833=>"111111011",
  23834=>"111010101",
  23835=>"000111100",
  23836=>"010110110",
  23837=>"111000111",
  23838=>"001101101",
  23839=>"000011011",
  23840=>"100010101",
  23841=>"110001110",
  23842=>"110111011",
  23843=>"000010110",
  23844=>"010000110",
  23845=>"010010001",
  23846=>"100010001",
  23847=>"111111110",
  23848=>"010001100",
  23849=>"010111110",
  23850=>"100100111",
  23851=>"110110100",
  23852=>"100100011",
  23853=>"011110110",
  23854=>"000101100",
  23855=>"101011111",
  23856=>"111011100",
  23857=>"000101110",
  23858=>"011101000",
  23859=>"100011011",
  23860=>"110110000",
  23861=>"000011000",
  23862=>"101001110",
  23863=>"100000010",
  23864=>"101100111",
  23865=>"010111000",
  23866=>"010100010",
  23867=>"000111100",
  23868=>"111001000",
  23869=>"101011010",
  23870=>"110110101",
  23871=>"111011000",
  23872=>"000101110",
  23873=>"001100100",
  23874=>"000110100",
  23875=>"101001011",
  23876=>"000011011",
  23877=>"010010111",
  23878=>"011000111",
  23879=>"101101111",
  23880=>"001000000",
  23881=>"110000010",
  23882=>"110011101",
  23883=>"101110001",
  23884=>"101001011",
  23885=>"101110010",
  23886=>"100111001",
  23887=>"011000110",
  23888=>"011010101",
  23889=>"000001011",
  23890=>"000001110",
  23891=>"111011000",
  23892=>"001100000",
  23893=>"001011011",
  23894=>"010111111",
  23895=>"011111010",
  23896=>"101101000",
  23897=>"110001010",
  23898=>"000111101",
  23899=>"111101001",
  23900=>"110000110",
  23901=>"100101000",
  23902=>"110001100",
  23903=>"110010101",
  23904=>"110010000",
  23905=>"001100010",
  23906=>"011001110",
  23907=>"101101101",
  23908=>"110001001",
  23909=>"101000001",
  23910=>"100011001",
  23911=>"111100100",
  23912=>"000011011",
  23913=>"100110110",
  23914=>"010110100",
  23915=>"101000011",
  23916=>"101011001",
  23917=>"101011111",
  23918=>"100000011",
  23919=>"010011110",
  23920=>"101100111",
  23921=>"101111111",
  23922=>"101001100",
  23923=>"001000011",
  23924=>"111000111",
  23925=>"001001110",
  23926=>"100000010",
  23927=>"001101100",
  23928=>"010101001",
  23929=>"100111101",
  23930=>"111011110",
  23931=>"111111111",
  23932=>"001001110",
  23933=>"011010010",
  23934=>"010101101",
  23935=>"011000110",
  23936=>"111110010",
  23937=>"001111101",
  23938=>"101111110",
  23939=>"001100101",
  23940=>"011001011",
  23941=>"100001010",
  23942=>"101110111",
  23943=>"010001101",
  23944=>"011000111",
  23945=>"011001001",
  23946=>"000100111",
  23947=>"000001000",
  23948=>"000001110",
  23949=>"001010011",
  23950=>"100101111",
  23951=>"010100001",
  23952=>"001100011",
  23953=>"111101110",
  23954=>"001010011",
  23955=>"100000011",
  23956=>"001000101",
  23957=>"000111001",
  23958=>"101001010",
  23959=>"111001100",
  23960=>"101110011",
  23961=>"001100101",
  23962=>"110100101",
  23963=>"110010000",
  23964=>"000100111",
  23965=>"000101001",
  23966=>"111011100",
  23967=>"011110101",
  23968=>"100100100",
  23969=>"011100000",
  23970=>"110010101",
  23971=>"011100111",
  23972=>"101000110",
  23973=>"000000110",
  23974=>"111110001",
  23975=>"011101000",
  23976=>"010100111",
  23977=>"100101000",
  23978=>"111110000",
  23979=>"110001000",
  23980=>"111101101",
  23981=>"111100010",
  23982=>"000000000",
  23983=>"010001000",
  23984=>"000111000",
  23985=>"100100000",
  23986=>"101110001",
  23987=>"011011001",
  23988=>"110111001",
  23989=>"110000101",
  23990=>"001010111",
  23991=>"111100111",
  23992=>"001100010",
  23993=>"010111111",
  23994=>"001100010",
  23995=>"000111000",
  23996=>"110110010",
  23997=>"011110101",
  23998=>"110000011",
  23999=>"100011111",
  24000=>"111100100",
  24001=>"011110010",
  24002=>"110010101",
  24003=>"011010001",
  24004=>"010000110",
  24005=>"011111100",
  24006=>"000010000",
  24007=>"101010000",
  24008=>"101101001",
  24009=>"011100000",
  24010=>"011101011",
  24011=>"011101010",
  24012=>"000000000",
  24013=>"000101100",
  24014=>"111011111",
  24015=>"101100101",
  24016=>"101100001",
  24017=>"111001100",
  24018=>"001011001",
  24019=>"100011011",
  24020=>"101110101",
  24021=>"000110000",
  24022=>"100011001",
  24023=>"100100000",
  24024=>"101100100",
  24025=>"000011101",
  24026=>"011110101",
  24027=>"111001100",
  24028=>"000000011",
  24029=>"000111011",
  24030=>"000111100",
  24031=>"110011100",
  24032=>"001110100",
  24033=>"110010010",
  24034=>"000000100",
  24035=>"110111101",
  24036=>"111100100",
  24037=>"011010110",
  24038=>"110110110",
  24039=>"101110110",
  24040=>"011010011",
  24041=>"001101110",
  24042=>"100000100",
  24043=>"010001000",
  24044=>"010000010",
  24045=>"010001000",
  24046=>"101000011",
  24047=>"110001011",
  24048=>"010111000",
  24049=>"111010111",
  24050=>"000010000",
  24051=>"100011011",
  24052=>"010111000",
  24053=>"101011011",
  24054=>"111000011",
  24055=>"011001010",
  24056=>"000111100",
  24057=>"011011011",
  24058=>"001000110",
  24059=>"001100010",
  24060=>"100000001",
  24061=>"110010010",
  24062=>"011100001",
  24063=>"111110111",
  24064=>"100001001",
  24065=>"101111101",
  24066=>"000101001",
  24067=>"010001010",
  24068=>"010000001",
  24069=>"100101100",
  24070=>"110100110",
  24071=>"100110111",
  24072=>"010000011",
  24073=>"110111011",
  24074=>"010101011",
  24075=>"000100000",
  24076=>"111100101",
  24077=>"111110010",
  24078=>"000100101",
  24079=>"000001010",
  24080=>"100011001",
  24081=>"111111110",
  24082=>"001110000",
  24083=>"111101010",
  24084=>"111100000",
  24085=>"011000101",
  24086=>"100101000",
  24087=>"010110000",
  24088=>"000111111",
  24089=>"010111000",
  24090=>"001000000",
  24091=>"010100001",
  24092=>"101001000",
  24093=>"101001100",
  24094=>"010011110",
  24095=>"110100110",
  24096=>"000001001",
  24097=>"010010101",
  24098=>"000011111",
  24099=>"101100001",
  24100=>"010101000",
  24101=>"011011001",
  24102=>"000101011",
  24103=>"000100000",
  24104=>"111111100",
  24105=>"111001111",
  24106=>"001100000",
  24107=>"001010110",
  24108=>"100111101",
  24109=>"111011010",
  24110=>"110010000",
  24111=>"101110110",
  24112=>"100111011",
  24113=>"011011010",
  24114=>"000001000",
  24115=>"000110100",
  24116=>"111011010",
  24117=>"000000111",
  24118=>"111001111",
  24119=>"000111101",
  24120=>"000010011",
  24121=>"000000110",
  24122=>"101111101",
  24123=>"011111010",
  24124=>"000011110",
  24125=>"111110001",
  24126=>"000101001",
  24127=>"011101001",
  24128=>"011010001",
  24129=>"110000011",
  24130=>"000111111",
  24131=>"010010111",
  24132=>"101100110",
  24133=>"100100001",
  24134=>"111101011",
  24135=>"001001110",
  24136=>"111010000",
  24137=>"111100001",
  24138=>"000010010",
  24139=>"100000011",
  24140=>"011110000",
  24141=>"111010001",
  24142=>"001000000",
  24143=>"101100011",
  24144=>"111101101",
  24145=>"011001101",
  24146=>"010010011",
  24147=>"101110101",
  24148=>"100000101",
  24149=>"100010110",
  24150=>"100110101",
  24151=>"000111001",
  24152=>"010100011",
  24153=>"101011101",
  24154=>"100101001",
  24155=>"110010110",
  24156=>"001001001",
  24157=>"111110110",
  24158=>"011101010",
  24159=>"010110001",
  24160=>"101101111",
  24161=>"110011111",
  24162=>"011110100",
  24163=>"000000010",
  24164=>"010101100",
  24165=>"110101000",
  24166=>"101100111",
  24167=>"100001000",
  24168=>"110010001",
  24169=>"111001110",
  24170=>"111000110",
  24171=>"111110001",
  24172=>"000001010",
  24173=>"110011010",
  24174=>"011111101",
  24175=>"111100000",
  24176=>"110001011",
  24177=>"110000000",
  24178=>"011110011",
  24179=>"111111101",
  24180=>"110110010",
  24181=>"010111101",
  24182=>"010001110",
  24183=>"110001000",
  24184=>"100011011",
  24185=>"000111111",
  24186=>"011100101",
  24187=>"011111111",
  24188=>"000001011",
  24189=>"010000110",
  24190=>"101110101",
  24191=>"001010101",
  24192=>"000100000",
  24193=>"001000111",
  24194=>"100100110",
  24195=>"101101110",
  24196=>"001010011",
  24197=>"111001000",
  24198=>"010100011",
  24199=>"111010011",
  24200=>"000001110",
  24201=>"010111110",
  24202=>"011100111",
  24203=>"111001100",
  24204=>"011000111",
  24205=>"010100011",
  24206=>"000000100",
  24207=>"110000110",
  24208=>"100110100",
  24209=>"011100001",
  24210=>"001011110",
  24211=>"001011111",
  24212=>"100110111",
  24213=>"001011001",
  24214=>"100101111",
  24215=>"010011101",
  24216=>"000101010",
  24217=>"011111101",
  24218=>"100000011",
  24219=>"110101111",
  24220=>"000000110",
  24221=>"111110110",
  24222=>"100011100",
  24223=>"001011110",
  24224=>"010001000",
  24225=>"000110001",
  24226=>"000011101",
  24227=>"101110100",
  24228=>"101011001",
  24229=>"010011011",
  24230=>"010101000",
  24231=>"100101100",
  24232=>"000001111",
  24233=>"100111110",
  24234=>"000011000",
  24235=>"001110111",
  24236=>"100000111",
  24237=>"011010100",
  24238=>"011111001",
  24239=>"100001101",
  24240=>"111000100",
  24241=>"000110110",
  24242=>"101010110",
  24243=>"011100001",
  24244=>"101111111",
  24245=>"010111100",
  24246=>"110001100",
  24247=>"010101001",
  24248=>"011111001",
  24249=>"111010011",
  24250=>"000010110",
  24251=>"011001010",
  24252=>"100010110",
  24253=>"000001011",
  24254=>"100000110",
  24255=>"110111111",
  24256=>"010111111",
  24257=>"101011111",
  24258=>"110001111",
  24259=>"011100010",
  24260=>"000100001",
  24261=>"011010001",
  24262=>"001111110",
  24263=>"111011101",
  24264=>"111111001",
  24265=>"100100001",
  24266=>"001001000",
  24267=>"111110100",
  24268=>"000011000",
  24269=>"011010010",
  24270=>"111001100",
  24271=>"111001011",
  24272=>"100011101",
  24273=>"100000101",
  24274=>"110111000",
  24275=>"001000000",
  24276=>"000101101",
  24277=>"101111111",
  24278=>"101010010",
  24279=>"010000001",
  24280=>"000110101",
  24281=>"111100101",
  24282=>"100100000",
  24283=>"101100101",
  24284=>"100100010",
  24285=>"101011000",
  24286=>"100110010",
  24287=>"111000000",
  24288=>"110110110",
  24289=>"110100100",
  24290=>"111001000",
  24291=>"010101100",
  24292=>"111101110",
  24293=>"111100000",
  24294=>"011010000",
  24295=>"110110000",
  24296=>"110011101",
  24297=>"110001101",
  24298=>"000111100",
  24299=>"110010001",
  24300=>"100111011",
  24301=>"110110100",
  24302=>"001001100",
  24303=>"101111100",
  24304=>"101000100",
  24305=>"010101110",
  24306=>"101001011",
  24307=>"010101110",
  24308=>"110110000",
  24309=>"101001000",
  24310=>"001111100",
  24311=>"011110110",
  24312=>"111101101",
  24313=>"110101100",
  24314=>"011001010",
  24315=>"111001101",
  24316=>"110100010",
  24317=>"100100111",
  24318=>"111110111",
  24319=>"011010001",
  24320=>"100111010",
  24321=>"001011011",
  24322=>"000011110",
  24323=>"010001111",
  24324=>"100101111",
  24325=>"100111000",
  24326=>"101011011",
  24327=>"001101001",
  24328=>"011101000",
  24329=>"001010010",
  24330=>"100000000",
  24331=>"001101001",
  24332=>"110011101",
  24333=>"111000011",
  24334=>"101100001",
  24335=>"101001100",
  24336=>"001001101",
  24337=>"111101100",
  24338=>"111000001",
  24339=>"110000101",
  24340=>"000001111",
  24341=>"101010100",
  24342=>"101111101",
  24343=>"001100110",
  24344=>"001000000",
  24345=>"100000010",
  24346=>"101100101",
  24347=>"110100110",
  24348=>"101100010",
  24349=>"100011000",
  24350=>"100110111",
  24351=>"001111110",
  24352=>"111001101",
  24353=>"010010011",
  24354=>"100001000",
  24355=>"010010000",
  24356=>"011101000",
  24357=>"000000110",
  24358=>"001001100",
  24359=>"101001001",
  24360=>"111001100",
  24361=>"100110010",
  24362=>"111111011",
  24363=>"110011001",
  24364=>"010010100",
  24365=>"101000111",
  24366=>"000011000",
  24367=>"110110101",
  24368=>"110011011",
  24369=>"001111011",
  24370=>"000111000",
  24371=>"000010010",
  24372=>"101111011",
  24373=>"011101001",
  24374=>"100100111",
  24375=>"111011011",
  24376=>"110111010",
  24377=>"010000000",
  24378=>"111111111",
  24379=>"111010010",
  24380=>"010000011",
  24381=>"101011001",
  24382=>"000010000",
  24383=>"111010001",
  24384=>"011010011",
  24385=>"101101110",
  24386=>"011010011",
  24387=>"101111010",
  24388=>"110010000",
  24389=>"001101110",
  24390=>"000111100",
  24391=>"001111101",
  24392=>"101111100",
  24393=>"000100000",
  24394=>"001111001",
  24395=>"011110001",
  24396=>"011100000",
  24397=>"011110001",
  24398=>"101011000",
  24399=>"001001000",
  24400=>"000111000",
  24401=>"100001011",
  24402=>"110000001",
  24403=>"010111111",
  24404=>"011100110",
  24405=>"110000011",
  24406=>"000101011",
  24407=>"110000101",
  24408=>"111001100",
  24409=>"100010011",
  24410=>"011100011",
  24411=>"000010001",
  24412=>"011101000",
  24413=>"001100001",
  24414=>"100010110",
  24415=>"000101011",
  24416=>"010010100",
  24417=>"010011011",
  24418=>"111011110",
  24419=>"010010011",
  24420=>"100100011",
  24421=>"011110100",
  24422=>"011111001",
  24423=>"000100001",
  24424=>"010010010",
  24425=>"100111001",
  24426=>"001110011",
  24427=>"110011111",
  24428=>"110001010",
  24429=>"001111010",
  24430=>"101111110",
  24431=>"000010000",
  24432=>"010101011",
  24433=>"101010000",
  24434=>"011000101",
  24435=>"010101001",
  24436=>"001100001",
  24437=>"100100010",
  24438=>"101101101",
  24439=>"101101111",
  24440=>"110101010",
  24441=>"010101101",
  24442=>"101100001",
  24443=>"111000000",
  24444=>"000001000",
  24445=>"001111111",
  24446=>"111111100",
  24447=>"110010111",
  24448=>"011111011",
  24449=>"000100111",
  24450=>"111001011",
  24451=>"100011100",
  24452=>"000110111",
  24453=>"010110101",
  24454=>"101010011",
  24455=>"110101010",
  24456=>"111011110",
  24457=>"111110001",
  24458=>"001101111",
  24459=>"101000010",
  24460=>"110101101",
  24461=>"101100001",
  24462=>"101110111",
  24463=>"010101100",
  24464=>"100001110",
  24465=>"011101101",
  24466=>"000111111",
  24467=>"100111011",
  24468=>"011001100",
  24469=>"100001111",
  24470=>"000100010",
  24471=>"100000110",
  24472=>"110001010",
  24473=>"000001001",
  24474=>"111100100",
  24475=>"000011010",
  24476=>"000001110",
  24477=>"000110000",
  24478=>"111001011",
  24479=>"101110001",
  24480=>"001101111",
  24481=>"100011010",
  24482=>"100011011",
  24483=>"011010010",
  24484=>"101100011",
  24485=>"011101101",
  24486=>"011101001",
  24487=>"101001011",
  24488=>"010011101",
  24489=>"111001111",
  24490=>"110100001",
  24491=>"001000100",
  24492=>"001111001",
  24493=>"000111110",
  24494=>"100001110",
  24495=>"001001101",
  24496=>"110000101",
  24497=>"110000101",
  24498=>"001001011",
  24499=>"011101101",
  24500=>"101111110",
  24501=>"001011100",
  24502=>"010011110",
  24503=>"001000000",
  24504=>"001010111",
  24505=>"100101100",
  24506=>"100101100",
  24507=>"000000100",
  24508=>"001111010",
  24509=>"111101101",
  24510=>"010100000",
  24511=>"001100001",
  24512=>"010111001",
  24513=>"000110100",
  24514=>"001101110",
  24515=>"101100101",
  24516=>"110111111",
  24517=>"101110000",
  24518=>"111111010",
  24519=>"011000010",
  24520=>"000010011",
  24521=>"001011000",
  24522=>"010001100",
  24523=>"101101111",
  24524=>"011011101",
  24525=>"100010111",
  24526=>"000000100",
  24527=>"101011011",
  24528=>"111000010",
  24529=>"100001110",
  24530=>"110000000",
  24531=>"011101010",
  24532=>"011001111",
  24533=>"000100110",
  24534=>"011011000",
  24535=>"101101110",
  24536=>"001010101",
  24537=>"110110110",
  24538=>"111101101",
  24539=>"010000001",
  24540=>"000111011",
  24541=>"010001000",
  24542=>"111100010",
  24543=>"111101101",
  24544=>"100111001",
  24545=>"001101011",
  24546=>"101110011",
  24547=>"001111001",
  24548=>"110001011",
  24549=>"000111001",
  24550=>"110000110",
  24551=>"100010100",
  24552=>"001000100",
  24553=>"011001011",
  24554=>"101110101",
  24555=>"111000101",
  24556=>"011100100",
  24557=>"001101001",
  24558=>"110001011",
  24559=>"000011001",
  24560=>"100111101",
  24561=>"011100111",
  24562=>"000010110",
  24563=>"010010110",
  24564=>"010000110",
  24565=>"000001001",
  24566=>"000000111",
  24567=>"001110010",
  24568=>"110011111",
  24569=>"010100101",
  24570=>"111110111",
  24571=>"010101111",
  24572=>"010010111",
  24573=>"010011111",
  24574=>"100000111",
  24575=>"100011101",
  24576=>"111101101",
  24577=>"110010101",
  24578=>"010110110",
  24579=>"101101010",
  24580=>"011011100",
  24581=>"100101110",
  24582=>"011100010",
  24583=>"110000111",
  24584=>"000110000",
  24585=>"100101010",
  24586=>"111111011",
  24587=>"000010000",
  24588=>"001111011",
  24589=>"001011000",
  24590=>"111110011",
  24591=>"101111011",
  24592=>"010001100",
  24593=>"111100100",
  24594=>"100110111",
  24595=>"110000100",
  24596=>"111110111",
  24597=>"111010001",
  24598=>"110100011",
  24599=>"011010010",
  24600=>"111010010",
  24601=>"010000101",
  24602=>"100001001",
  24603=>"100111101",
  24604=>"000110111",
  24605=>"101001010",
  24606=>"000101101",
  24607=>"101010111",
  24608=>"110111101",
  24609=>"001110000",
  24610=>"011110010",
  24611=>"011011100",
  24612=>"110000001",
  24613=>"110110001",
  24614=>"111100101",
  24615=>"100100010",
  24616=>"101000101",
  24617=>"100001000",
  24618=>"111101100",
  24619=>"110000111",
  24620=>"011110001",
  24621=>"000010101",
  24622=>"011100111",
  24623=>"110110111",
  24624=>"111010111",
  24625=>"010101110",
  24626=>"110100101",
  24627=>"110011011",
  24628=>"011000010",
  24629=>"000111110",
  24630=>"010001011",
  24631=>"000100010",
  24632=>"110010001",
  24633=>"111100101",
  24634=>"101011110",
  24635=>"001010110",
  24636=>"010111001",
  24637=>"101000111",
  24638=>"001111111",
  24639=>"010110011",
  24640=>"110010100",
  24641=>"110101010",
  24642=>"110001001",
  24643=>"101011010",
  24644=>"111110001",
  24645=>"100100111",
  24646=>"111001001",
  24647=>"000110011",
  24648=>"111000101",
  24649=>"001001111",
  24650=>"111000110",
  24651=>"101011000",
  24652=>"101001001",
  24653=>"100010000",
  24654=>"110111101",
  24655=>"101111001",
  24656=>"000110100",
  24657=>"010100001",
  24658=>"101010111",
  24659=>"100110100",
  24660=>"111101110",
  24661=>"100010001",
  24662=>"000011010",
  24663=>"111010001",
  24664=>"101111101",
  24665=>"101001111",
  24666=>"111010010",
  24667=>"011101000",
  24668=>"001101110",
  24669=>"010001101",
  24670=>"111010111",
  24671=>"011110110",
  24672=>"000000010",
  24673=>"011110011",
  24674=>"100010010",
  24675=>"001101100",
  24676=>"001100001",
  24677=>"000000110",
  24678=>"010101001",
  24679=>"011011000",
  24680=>"111001111",
  24681=>"010010101",
  24682=>"001110000",
  24683=>"101010111",
  24684=>"010001011",
  24685=>"110011001",
  24686=>"101100001",
  24687=>"101000011",
  24688=>"001010001",
  24689=>"101011100",
  24690=>"101111100",
  24691=>"111100000",
  24692=>"100000100",
  24693=>"100001100",
  24694=>"011111000",
  24695=>"111101110",
  24696=>"001100001",
  24697=>"101111100",
  24698=>"111111100",
  24699=>"101110101",
  24700=>"000111110",
  24701=>"111011011",
  24702=>"111110010",
  24703=>"010111111",
  24704=>"000100001",
  24705=>"100101100",
  24706=>"000011001",
  24707=>"010001101",
  24708=>"000110010",
  24709=>"000001000",
  24710=>"010110001",
  24711=>"001000001",
  24712=>"000010111",
  24713=>"000100000",
  24714=>"100001000",
  24715=>"000011010",
  24716=>"110111111",
  24717=>"111001110",
  24718=>"001100001",
  24719=>"101000110",
  24720=>"010111010",
  24721=>"000110101",
  24722=>"101101100",
  24723=>"001000011",
  24724=>"100000000",
  24725=>"010110100",
  24726=>"101111011",
  24727=>"111111100",
  24728=>"100110101",
  24729=>"010011000",
  24730=>"100100110",
  24731=>"111101010",
  24732=>"011010100",
  24733=>"000101000",
  24734=>"011100011",
  24735=>"011010110",
  24736=>"000001000",
  24737=>"101110011",
  24738=>"100100001",
  24739=>"000101011",
  24740=>"110011101",
  24741=>"110110100",
  24742=>"101110101",
  24743=>"011000010",
  24744=>"111000111",
  24745=>"011110001",
  24746=>"010101101",
  24747=>"100100011",
  24748=>"110010001",
  24749=>"011000101",
  24750=>"001100101",
  24751=>"001001110",
  24752=>"111010001",
  24753=>"111010011",
  24754=>"111110000",
  24755=>"110010100",
  24756=>"010101111",
  24757=>"100101011",
  24758=>"001111001",
  24759=>"000111110",
  24760=>"101000110",
  24761=>"011001011",
  24762=>"010100111",
  24763=>"001101101",
  24764=>"010101111",
  24765=>"011010111",
  24766=>"110001011",
  24767=>"100110111",
  24768=>"001011101",
  24769=>"011100011",
  24770=>"100100001",
  24771=>"010100100",
  24772=>"010101010",
  24773=>"000111110",
  24774=>"010000010",
  24775=>"110110110",
  24776=>"110000000",
  24777=>"001001101",
  24778=>"110000001",
  24779=>"101110111",
  24780=>"001011000",
  24781=>"110110110",
  24782=>"100110010",
  24783=>"100001010",
  24784=>"011011100",
  24785=>"110111010",
  24786=>"100111000",
  24787=>"010111010",
  24788=>"100010110",
  24789=>"101011011",
  24790=>"001000011",
  24791=>"011110010",
  24792=>"011110000",
  24793=>"011111110",
  24794=>"011000111",
  24795=>"101111100",
  24796=>"010010110",
  24797=>"101111011",
  24798=>"111101011",
  24799=>"001100100",
  24800=>"100000101",
  24801=>"011111111",
  24802=>"111000111",
  24803=>"110111110",
  24804=>"000000100",
  24805=>"011100111",
  24806=>"100010001",
  24807=>"101001010",
  24808=>"101111010",
  24809=>"101110001",
  24810=>"000001101",
  24811=>"110011110",
  24812=>"011110001",
  24813=>"100011110",
  24814=>"111111100",
  24815=>"010110100",
  24816=>"111101111",
  24817=>"111100110",
  24818=>"100010101",
  24819=>"001111111",
  24820=>"101010100",
  24821=>"001010101",
  24822=>"000001010",
  24823=>"110111110",
  24824=>"100011000",
  24825=>"100011001",
  24826=>"101011000",
  24827=>"110011100",
  24828=>"111000010",
  24829=>"010010110",
  24830=>"101101011",
  24831=>"101010101",
  24832=>"110110011",
  24833=>"010010000",
  24834=>"111001111",
  24835=>"111010110",
  24836=>"110000101",
  24837=>"010001000",
  24838=>"101101110",
  24839=>"101110100",
  24840=>"001000101",
  24841=>"001001011",
  24842=>"100010110",
  24843=>"011111111",
  24844=>"000111100",
  24845=>"111010110",
  24846=>"111101111",
  24847=>"010111010",
  24848=>"110100111",
  24849=>"110000100",
  24850=>"100001111",
  24851=>"100111011",
  24852=>"111000101",
  24853=>"000110101",
  24854=>"101000010",
  24855=>"011000100",
  24856=>"101000100",
  24857=>"111010010",
  24858=>"000010000",
  24859=>"011111110",
  24860=>"000100111",
  24861=>"110101011",
  24862=>"001110101",
  24863=>"101110010",
  24864=>"100010111",
  24865=>"110101010",
  24866=>"101000010",
  24867=>"001110111",
  24868=>"101000011",
  24869=>"001110000",
  24870=>"100100011",
  24871=>"011000011",
  24872=>"101101100",
  24873=>"110001010",
  24874=>"101101000",
  24875=>"111011100",
  24876=>"010111110",
  24877=>"000001011",
  24878=>"100101001",
  24879=>"001011111",
  24880=>"010101101",
  24881=>"011110100",
  24882=>"111011000",
  24883=>"011101011",
  24884=>"100110001",
  24885=>"001101010",
  24886=>"111011100",
  24887=>"011011100",
  24888=>"111011000",
  24889=>"101001000",
  24890=>"100001010",
  24891=>"111110000",
  24892=>"000011100",
  24893=>"000000001",
  24894=>"100011001",
  24895=>"011110111",
  24896=>"110100000",
  24897=>"101101011",
  24898=>"111100111",
  24899=>"110110100",
  24900=>"110000011",
  24901=>"100100111",
  24902=>"100100011",
  24903=>"010110111",
  24904=>"000110100",
  24905=>"110001101",
  24906=>"011011000",
  24907=>"100000010",
  24908=>"110010010",
  24909=>"111110111",
  24910=>"000100100",
  24911=>"100101000",
  24912=>"000101111",
  24913=>"111110100",
  24914=>"010011001",
  24915=>"110101101",
  24916=>"010100100",
  24917=>"110000111",
  24918=>"000001001",
  24919=>"011101100",
  24920=>"110110010",
  24921=>"011001001",
  24922=>"000010000",
  24923=>"101110011",
  24924=>"000010010",
  24925=>"111001101",
  24926=>"001000100",
  24927=>"111110111",
  24928=>"110010100",
  24929=>"111010100",
  24930=>"001000001",
  24931=>"011100010",
  24932=>"000010010",
  24933=>"010100110",
  24934=>"101110011",
  24935=>"110110000",
  24936=>"000101100",
  24937=>"111111010",
  24938=>"100011010",
  24939=>"111101110",
  24940=>"111000000",
  24941=>"000101111",
  24942=>"101010101",
  24943=>"110001110",
  24944=>"100011111",
  24945=>"101001101",
  24946=>"011100001",
  24947=>"000111101",
  24948=>"100111011",
  24949=>"110111011",
  24950=>"010100000",
  24951=>"000110100",
  24952=>"101010100",
  24953=>"011110010",
  24954=>"101101001",
  24955=>"110101111",
  24956=>"010011111",
  24957=>"010000001",
  24958=>"011101000",
  24959=>"111010011",
  24960=>"010100111",
  24961=>"001100011",
  24962=>"100101101",
  24963=>"100101010",
  24964=>"010110111",
  24965=>"011011001",
  24966=>"100001111",
  24967=>"010010010",
  24968=>"001011010",
  24969=>"111100010",
  24970=>"101001101",
  24971=>"111001000",
  24972=>"001101100",
  24973=>"111100111",
  24974=>"011010001",
  24975=>"010110011",
  24976=>"101110111",
  24977=>"010011010",
  24978=>"101100100",
  24979=>"000000110",
  24980=>"011110100",
  24981=>"001000101",
  24982=>"001010000",
  24983=>"000110101",
  24984=>"100101100",
  24985=>"000110110",
  24986=>"010100011",
  24987=>"000101101",
  24988=>"111100011",
  24989=>"011110011",
  24990=>"000111010",
  24991=>"110100110",
  24992=>"110000100",
  24993=>"001000000",
  24994=>"001111101",
  24995=>"000000001",
  24996=>"001001000",
  24997=>"100000000",
  24998=>"010000110",
  24999=>"111000011",
  25000=>"001110000",
  25001=>"000110010",
  25002=>"000001011",
  25003=>"001001001",
  25004=>"101111101",
  25005=>"000000001",
  25006=>"010000101",
  25007=>"101010111",
  25008=>"110011100",
  25009=>"011010010",
  25010=>"000001001",
  25011=>"000011001",
  25012=>"101010111",
  25013=>"101110010",
  25014=>"110101101",
  25015=>"101001100",
  25016=>"011110010",
  25017=>"011111101",
  25018=>"101110100",
  25019=>"101101011",
  25020=>"100010101",
  25021=>"100000110",
  25022=>"000010011",
  25023=>"100011010",
  25024=>"111001110",
  25025=>"111111001",
  25026=>"100001110",
  25027=>"000111000",
  25028=>"111111010",
  25029=>"110111110",
  25030=>"010100110",
  25031=>"101010111",
  25032=>"111110001",
  25033=>"001011101",
  25034=>"011011011",
  25035=>"010001110",
  25036=>"010001000",
  25037=>"110010101",
  25038=>"100011001",
  25039=>"001101111",
  25040=>"110100110",
  25041=>"000101000",
  25042=>"010011100",
  25043=>"111001000",
  25044=>"000000100",
  25045=>"001000110",
  25046=>"000010000",
  25047=>"011011101",
  25048=>"100010111",
  25049=>"000011111",
  25050=>"110011101",
  25051=>"010110110",
  25052=>"110110000",
  25053=>"011001111",
  25054=>"011001010",
  25055=>"111110101",
  25056=>"000101000",
  25057=>"011000000",
  25058=>"101011010",
  25059=>"111101001",
  25060=>"011011001",
  25061=>"001110111",
  25062=>"001101011",
  25063=>"000111100",
  25064=>"000111100",
  25065=>"110101011",
  25066=>"001001001",
  25067=>"111111010",
  25068=>"101001011",
  25069=>"001100000",
  25070=>"111000100",
  25071=>"101010010",
  25072=>"101101100",
  25073=>"110101010",
  25074=>"000001010",
  25075=>"111100101",
  25076=>"011011100",
  25077=>"101110110",
  25078=>"000011000",
  25079=>"110011001",
  25080=>"101001111",
  25081=>"110100000",
  25082=>"010001101",
  25083=>"000000101",
  25084=>"111010010",
  25085=>"011100101",
  25086=>"101110110",
  25087=>"010110111",
  25088=>"010100001",
  25089=>"100100110",
  25090=>"101011110",
  25091=>"110100011",
  25092=>"111000000",
  25093=>"111100100",
  25094=>"001110010",
  25095=>"000111100",
  25096=>"111100001",
  25097=>"000000100",
  25098=>"001110100",
  25099=>"100001100",
  25100=>"010111111",
  25101=>"010110001",
  25102=>"000000110",
  25103=>"011110010",
  25104=>"111101101",
  25105=>"110001110",
  25106=>"101010111",
  25107=>"110100100",
  25108=>"110110101",
  25109=>"010011010",
  25110=>"001000000",
  25111=>"110100011",
  25112=>"000110011",
  25113=>"111100111",
  25114=>"011000101",
  25115=>"000111011",
  25116=>"010100100",
  25117=>"111100011",
  25118=>"111010111",
  25119=>"011011111",
  25120=>"111101010",
  25121=>"101110011",
  25122=>"110000010",
  25123=>"001011011",
  25124=>"010011000",
  25125=>"010001111",
  25126=>"110001111",
  25127=>"010011001",
  25128=>"101111010",
  25129=>"111111110",
  25130=>"100011011",
  25131=>"000100111",
  25132=>"111110101",
  25133=>"000000000",
  25134=>"011010000",
  25135=>"000000111",
  25136=>"010001101",
  25137=>"111110110",
  25138=>"111100100",
  25139=>"010101000",
  25140=>"111111111",
  25141=>"100011011",
  25142=>"110010000",
  25143=>"110110000",
  25144=>"011110110",
  25145=>"101001100",
  25146=>"100100011",
  25147=>"001101110",
  25148=>"101100110",
  25149=>"001010100",
  25150=>"111011010",
  25151=>"101111111",
  25152=>"000100111",
  25153=>"100101101",
  25154=>"011111011",
  25155=>"110011001",
  25156=>"110101011",
  25157=>"111100011",
  25158=>"101010001",
  25159=>"110101000",
  25160=>"000111011",
  25161=>"010010100",
  25162=>"101100101",
  25163=>"111111111",
  25164=>"111100110",
  25165=>"110111100",
  25166=>"110101011",
  25167=>"110110011",
  25168=>"010100001",
  25169=>"111100011",
  25170=>"011111011",
  25171=>"001010101",
  25172=>"111100000",
  25173=>"110010111",
  25174=>"000011010",
  25175=>"111000001",
  25176=>"111111000",
  25177=>"000100011",
  25178=>"111000111",
  25179=>"011001101",
  25180=>"001100101",
  25181=>"000100101",
  25182=>"101110011",
  25183=>"101111110",
  25184=>"110011111",
  25185=>"101001100",
  25186=>"011110000",
  25187=>"001110100",
  25188=>"100011001",
  25189=>"110011010",
  25190=>"111101011",
  25191=>"110100110",
  25192=>"011110101",
  25193=>"000111101",
  25194=>"000001010",
  25195=>"001011101",
  25196=>"101110010",
  25197=>"101110000",
  25198=>"100101010",
  25199=>"001100100",
  25200=>"111010110",
  25201=>"110111001",
  25202=>"110001000",
  25203=>"010000110",
  25204=>"101111010",
  25205=>"011110101",
  25206=>"011010001",
  25207=>"110101110",
  25208=>"000000111",
  25209=>"101010100",
  25210=>"000111011",
  25211=>"100111001",
  25212=>"000100110",
  25213=>"010011111",
  25214=>"111110001",
  25215=>"101010011",
  25216=>"111010111",
  25217=>"000010001",
  25218=>"110001001",
  25219=>"111011111",
  25220=>"011000101",
  25221=>"110101100",
  25222=>"000010111",
  25223=>"011010010",
  25224=>"011000010",
  25225=>"001000111",
  25226=>"001011100",
  25227=>"001010110",
  25228=>"000001011",
  25229=>"010001001",
  25230=>"101110111",
  25231=>"010110001",
  25232=>"011101011",
  25233=>"110000001",
  25234=>"000011001",
  25235=>"111010000",
  25236=>"101101111",
  25237=>"110001100",
  25238=>"011000111",
  25239=>"011000000",
  25240=>"101001110",
  25241=>"001100101",
  25242=>"111110111",
  25243=>"101000110",
  25244=>"100101100",
  25245=>"111111011",
  25246=>"001100001",
  25247=>"000111111",
  25248=>"001000000",
  25249=>"101001111",
  25250=>"000111010",
  25251=>"100101110",
  25252=>"000110011",
  25253=>"011001101",
  25254=>"001000011",
  25255=>"110011010",
  25256=>"110000000",
  25257=>"011111110",
  25258=>"011111011",
  25259=>"100010100",
  25260=>"111001100",
  25261=>"111101101",
  25262=>"000000010",
  25263=>"111111110",
  25264=>"010011111",
  25265=>"011010111",
  25266=>"001110101",
  25267=>"111010100",
  25268=>"111100100",
  25269=>"110110001",
  25270=>"000101001",
  25271=>"000010000",
  25272=>"011111101",
  25273=>"011011011",
  25274=>"010110011",
  25275=>"010101111",
  25276=>"011111001",
  25277=>"000001010",
  25278=>"110100110",
  25279=>"100111001",
  25280=>"111000100",
  25281=>"111011101",
  25282=>"101000011",
  25283=>"011111111",
  25284=>"010010011",
  25285=>"100100011",
  25286=>"010010010",
  25287=>"100001100",
  25288=>"110110100",
  25289=>"010101101",
  25290=>"000000111",
  25291=>"100011100",
  25292=>"010010010",
  25293=>"111010100",
  25294=>"111110101",
  25295=>"110100100",
  25296=>"111110100",
  25297=>"110110100",
  25298=>"110111000",
  25299=>"001000011",
  25300=>"111111110",
  25301=>"011000001",
  25302=>"001110000",
  25303=>"111111110",
  25304=>"001011110",
  25305=>"101001011",
  25306=>"001001011",
  25307=>"110111000",
  25308=>"010100011",
  25309=>"001000110",
  25310=>"111110010",
  25311=>"000110101",
  25312=>"000000111",
  25313=>"100000010",
  25314=>"101101011",
  25315=>"011101001",
  25316=>"100011111",
  25317=>"111111111",
  25318=>"111110100",
  25319=>"101011110",
  25320=>"101101001",
  25321=>"110001101",
  25322=>"101010111",
  25323=>"111010100",
  25324=>"111000101",
  25325=>"100000101",
  25326=>"101101000",
  25327=>"111010101",
  25328=>"010010011",
  25329=>"100101101",
  25330=>"010000011",
  25331=>"001111110",
  25332=>"010111000",
  25333=>"111111101",
  25334=>"110011110",
  25335=>"110001010",
  25336=>"100110011",
  25337=>"001110000",
  25338=>"100011010",
  25339=>"110110001",
  25340=>"000110111",
  25341=>"011001101",
  25342=>"110100100",
  25343=>"101001000",
  25344=>"001001101",
  25345=>"110100000",
  25346=>"111110001",
  25347=>"000101001",
  25348=>"100101010",
  25349=>"011111110",
  25350=>"110100111",
  25351=>"010011001",
  25352=>"000010000",
  25353=>"010110101",
  25354=>"101011110",
  25355=>"110101110",
  25356=>"011011111",
  25357=>"000110101",
  25358=>"010100010",
  25359=>"011010000",
  25360=>"111101011",
  25361=>"111101111",
  25362=>"011010001",
  25363=>"101101101",
  25364=>"111000010",
  25365=>"000010000",
  25366=>"010100101",
  25367=>"011000110",
  25368=>"010111100",
  25369=>"101100001",
  25370=>"101100111",
  25371=>"111001010",
  25372=>"100001010",
  25373=>"110001100",
  25374=>"111001011",
  25375=>"110111001",
  25376=>"011001101",
  25377=>"010101110",
  25378=>"000011111",
  25379=>"001000110",
  25380=>"010101010",
  25381=>"100000111",
  25382=>"000011110",
  25383=>"011111011",
  25384=>"010010011",
  25385=>"101111011",
  25386=>"111110111",
  25387=>"010110100",
  25388=>"011110001",
  25389=>"011110010",
  25390=>"101001111",
  25391=>"010010011",
  25392=>"100111011",
  25393=>"010100011",
  25394=>"010000100",
  25395=>"110001010",
  25396=>"001111000",
  25397=>"111010101",
  25398=>"101000011",
  25399=>"101011100",
  25400=>"000110001",
  25401=>"011110011",
  25402=>"000101001",
  25403=>"101010110",
  25404=>"110011000",
  25405=>"010101011",
  25406=>"111100001",
  25407=>"110101001",
  25408=>"111011111",
  25409=>"001100110",
  25410=>"101101101",
  25411=>"110001011",
  25412=>"101100000",
  25413=>"010111000",
  25414=>"100111110",
  25415=>"111010000",
  25416=>"010100111",
  25417=>"100100011",
  25418=>"110100110",
  25419=>"110010100",
  25420=>"101101111",
  25421=>"111110010",
  25422=>"100111011",
  25423=>"010011101",
  25424=>"101101110",
  25425=>"101011111",
  25426=>"001100101",
  25427=>"110001001",
  25428=>"011111011",
  25429=>"001000101",
  25430=>"000010001",
  25431=>"100011001",
  25432=>"000101110",
  25433=>"100000010",
  25434=>"010111001",
  25435=>"000110001",
  25436=>"010011101",
  25437=>"000000001",
  25438=>"110011000",
  25439=>"101111111",
  25440=>"010011011",
  25441=>"111101010",
  25442=>"100011000",
  25443=>"110111111",
  25444=>"100000000",
  25445=>"100000000",
  25446=>"011110100",
  25447=>"000110001",
  25448=>"011100000",
  25449=>"111100110",
  25450=>"100010000",
  25451=>"010010011",
  25452=>"010000000",
  25453=>"111110111",
  25454=>"011001110",
  25455=>"010111100",
  25456=>"100010101",
  25457=>"101000010",
  25458=>"111011010",
  25459=>"010011011",
  25460=>"000000011",
  25461=>"101000000",
  25462=>"010111001",
  25463=>"010100101",
  25464=>"001111110",
  25465=>"010011101",
  25466=>"111011100",
  25467=>"111101101",
  25468=>"110110001",
  25469=>"011101100",
  25470=>"110111011",
  25471=>"011110101",
  25472=>"110011011",
  25473=>"010100001",
  25474=>"000000100",
  25475=>"011010000",
  25476=>"011111001",
  25477=>"110001000",
  25478=>"000000011",
  25479=>"000001001",
  25480=>"100101101",
  25481=>"010101011",
  25482=>"111011000",
  25483=>"000111001",
  25484=>"110001111",
  25485=>"100110100",
  25486=>"110111110",
  25487=>"110010001",
  25488=>"010010010",
  25489=>"110101101",
  25490=>"001000110",
  25491=>"000000100",
  25492=>"100011000",
  25493=>"000110111",
  25494=>"101010101",
  25495=>"010110110",
  25496=>"101001100",
  25497=>"111100101",
  25498=>"110001011",
  25499=>"110110011",
  25500=>"010111100",
  25501=>"101110000",
  25502=>"110011101",
  25503=>"010001010",
  25504=>"001001111",
  25505=>"000100011",
  25506=>"000110010",
  25507=>"000000001",
  25508=>"001110001",
  25509=>"000000010",
  25510=>"100100111",
  25511=>"010110001",
  25512=>"011111100",
  25513=>"000000010",
  25514=>"101100101",
  25515=>"100110110",
  25516=>"000001110",
  25517=>"101100011",
  25518=>"101100011",
  25519=>"100111100",
  25520=>"111110100",
  25521=>"110110001",
  25522=>"001010101",
  25523=>"000001010",
  25524=>"011101110",
  25525=>"100001011",
  25526=>"000010001",
  25527=>"000001000",
  25528=>"100010011",
  25529=>"010101100",
  25530=>"001001110",
  25531=>"100000100",
  25532=>"111011101",
  25533=>"010000111",
  25534=>"001100100",
  25535=>"111010101",
  25536=>"010111001",
  25537=>"000111110",
  25538=>"100000100",
  25539=>"110101111",
  25540=>"011110011",
  25541=>"011111011",
  25542=>"001111101",
  25543=>"011100110",
  25544=>"111110101",
  25545=>"100111101",
  25546=>"101001001",
  25547=>"101110111",
  25548=>"000101000",
  25549=>"111001010",
  25550=>"000000110",
  25551=>"010000011",
  25552=>"101001110",
  25553=>"100000000",
  25554=>"000010110",
  25555=>"110111011",
  25556=>"000001101",
  25557=>"010011100",
  25558=>"101111010",
  25559=>"111010000",
  25560=>"101100000",
  25561=>"111011011",
  25562=>"110100000",
  25563=>"000111011",
  25564=>"110010101",
  25565=>"000000011",
  25566=>"101111111",
  25567=>"000011101",
  25568=>"011000110",
  25569=>"110000000",
  25570=>"110100010",
  25571=>"000110011",
  25572=>"010100111",
  25573=>"011001000",
  25574=>"110111011",
  25575=>"101011000",
  25576=>"011010000",
  25577=>"110110000",
  25578=>"010100001",
  25579=>"011000001",
  25580=>"110001101",
  25581=>"110101010",
  25582=>"000001110",
  25583=>"100011011",
  25584=>"110101111",
  25585=>"101111010",
  25586=>"111001111",
  25587=>"011010010",
  25588=>"010000101",
  25589=>"101100100",
  25590=>"000000000",
  25591=>"011111111",
  25592=>"111111001",
  25593=>"001011000",
  25594=>"000100110",
  25595=>"001100011",
  25596=>"010001011",
  25597=>"110100001",
  25598=>"011010011",
  25599=>"100100010",
  25600=>"111101111",
  25601=>"011011011",
  25602=>"000001010",
  25603=>"101000111",
  25604=>"110110001",
  25605=>"101011111",
  25606=>"101111010",
  25607=>"111011110",
  25608=>"001101010",
  25609=>"010000110",
  25610=>"101111100",
  25611=>"000100001",
  25612=>"110011010",
  25613=>"010110110",
  25614=>"101111001",
  25615=>"101000010",
  25616=>"010011001",
  25617=>"111100001",
  25618=>"001111110",
  25619=>"001101100",
  25620=>"010101100",
  25621=>"010011000",
  25622=>"101010100",
  25623=>"000000000",
  25624=>"001100001",
  25625=>"000110110",
  25626=>"100011111",
  25627=>"101101110",
  25628=>"000011000",
  25629=>"111000001",
  25630=>"111110100",
  25631=>"000110001",
  25632=>"100001000",
  25633=>"111110110",
  25634=>"010101001",
  25635=>"001101111",
  25636=>"110111010",
  25637=>"000101111",
  25638=>"100110100",
  25639=>"001111111",
  25640=>"010101011",
  25641=>"111111100",
  25642=>"011111010",
  25643=>"100011100",
  25644=>"111100111",
  25645=>"011110000",
  25646=>"010010000",
  25647=>"001010011",
  25648=>"111101100",
  25649=>"011111100",
  25650=>"111110000",
  25651=>"111111111",
  25652=>"001011010",
  25653=>"000000110",
  25654=>"111101100",
  25655=>"111011000",
  25656=>"000011101",
  25657=>"010111010",
  25658=>"100000110",
  25659=>"010101010",
  25660=>"000010001",
  25661=>"111110000",
  25662=>"011000110",
  25663=>"101100011",
  25664=>"001010101",
  25665=>"000110000",
  25666=>"010110101",
  25667=>"111011010",
  25668=>"111110100",
  25669=>"100001000",
  25670=>"011111010",
  25671=>"101111110",
  25672=>"101001010",
  25673=>"000000101",
  25674=>"000001011",
  25675=>"101101000",
  25676=>"011100000",
  25677=>"101011010",
  25678=>"111000100",
  25679=>"101100101",
  25680=>"100000110",
  25681=>"011111011",
  25682=>"011111100",
  25683=>"000111010",
  25684=>"111100001",
  25685=>"011100100",
  25686=>"100111010",
  25687=>"000001111",
  25688=>"100110010",
  25689=>"101111010",
  25690=>"110111010",
  25691=>"011110000",
  25692=>"000011100",
  25693=>"111011010",
  25694=>"010011110",
  25695=>"010001111",
  25696=>"111100101",
  25697=>"001011010",
  25698=>"001110010",
  25699=>"111001010",
  25700=>"010000001",
  25701=>"110101011",
  25702=>"011110010",
  25703=>"000111101",
  25704=>"110111010",
  25705=>"001111000",
  25706=>"111100111",
  25707=>"000001100",
  25708=>"001000001",
  25709=>"101011011",
  25710=>"000111010",
  25711=>"100011101",
  25712=>"101100111",
  25713=>"010111010",
  25714=>"110011011",
  25715=>"111110100",
  25716=>"111111010",
  25717=>"010011111",
  25718=>"000100101",
  25719=>"010111000",
  25720=>"010010001",
  25721=>"001111000",
  25722=>"010000011",
  25723=>"001101110",
  25724=>"100101011",
  25725=>"100111101",
  25726=>"101100111",
  25727=>"000000100",
  25728=>"110101110",
  25729=>"111111101",
  25730=>"011001110",
  25731=>"110010010",
  25732=>"100100100",
  25733=>"011010010",
  25734=>"001000000",
  25735=>"011100100",
  25736=>"001011110",
  25737=>"000111011",
  25738=>"111101010",
  25739=>"111111110",
  25740=>"000011011",
  25741=>"100110010",
  25742=>"001010111",
  25743=>"101101011",
  25744=>"000110100",
  25745=>"011010100",
  25746=>"000010111",
  25747=>"010011000",
  25748=>"100100101",
  25749=>"000110011",
  25750=>"000010010",
  25751=>"000100101",
  25752=>"011101010",
  25753=>"001110000",
  25754=>"111111001",
  25755=>"001101001",
  25756=>"001101101",
  25757=>"101000100",
  25758=>"000010100",
  25759=>"110000010",
  25760=>"001101111",
  25761=>"000001110",
  25762=>"111010000",
  25763=>"100011010",
  25764=>"111110100",
  25765=>"010011011",
  25766=>"001100000",
  25767=>"011010111",
  25768=>"011011100",
  25769=>"001010010",
  25770=>"000000011",
  25771=>"011101111",
  25772=>"011100100",
  25773=>"110011100",
  25774=>"001000001",
  25775=>"001011001",
  25776=>"010111001",
  25777=>"111100111",
  25778=>"001001000",
  25779=>"101111111",
  25780=>"011110001",
  25781=>"110011100",
  25782=>"100001111",
  25783=>"111010011",
  25784=>"100000100",
  25785=>"100011101",
  25786=>"000010111",
  25787=>"101100010",
  25788=>"111001111",
  25789=>"001011111",
  25790=>"000101001",
  25791=>"001100010",
  25792=>"111110011",
  25793=>"001100111",
  25794=>"010011111",
  25795=>"000011001",
  25796=>"001010100",
  25797=>"101001111",
  25798=>"101110101",
  25799=>"100101111",
  25800=>"110010100",
  25801=>"101001001",
  25802=>"100101100",
  25803=>"110011001",
  25804=>"001110010",
  25805=>"011110001",
  25806=>"010000110",
  25807=>"101110101",
  25808=>"000010001",
  25809=>"001101010",
  25810=>"011010011",
  25811=>"000001010",
  25812=>"110100111",
  25813=>"000110011",
  25814=>"010011000",
  25815=>"101011001",
  25816=>"101011100",
  25817=>"000010110",
  25818=>"100101100",
  25819=>"000100011",
  25820=>"110010010",
  25821=>"111101111",
  25822=>"010111111",
  25823=>"100100111",
  25824=>"011010010",
  25825=>"000110110",
  25826=>"101001111",
  25827=>"100111100",
  25828=>"110111010",
  25829=>"011100001",
  25830=>"000000010",
  25831=>"001000111",
  25832=>"010001011",
  25833=>"010000100",
  25834=>"111010100",
  25835=>"111111111",
  25836=>"000010010",
  25837=>"000001011",
  25838=>"001011000",
  25839=>"000001110",
  25840=>"100110001",
  25841=>"010000010",
  25842=>"100001110",
  25843=>"001010011",
  25844=>"100111111",
  25845=>"100011100",
  25846=>"011001111",
  25847=>"101100011",
  25848=>"011011011",
  25849=>"001101011",
  25850=>"011001000",
  25851=>"000011100",
  25852=>"101100111",
  25853=>"010111000",
  25854=>"101000001",
  25855=>"011111101",
  25856=>"111000010",
  25857=>"000011111",
  25858=>"001100011",
  25859=>"101010011",
  25860=>"010111110",
  25861=>"010000110",
  25862=>"000000101",
  25863=>"001110101",
  25864=>"111101101",
  25865=>"000111000",
  25866=>"110101111",
  25867=>"111001011",
  25868=>"110110110",
  25869=>"110110000",
  25870=>"111011101",
  25871=>"111001011",
  25872=>"011001110",
  25873=>"101110010",
  25874=>"001010010",
  25875=>"110001010",
  25876=>"100100101",
  25877=>"011000101",
  25878=>"101001001",
  25879=>"100010011",
  25880=>"101001111",
  25881=>"010110100",
  25882=>"101111101",
  25883=>"011101100",
  25884=>"000011010",
  25885=>"101100111",
  25886=>"010011110",
  25887=>"111000010",
  25888=>"011001110",
  25889=>"001111011",
  25890=>"110111110",
  25891=>"010011100",
  25892=>"111110111",
  25893=>"111110011",
  25894=>"011010111",
  25895=>"101101101",
  25896=>"101000100",
  25897=>"001010011",
  25898=>"110100011",
  25899=>"011101000",
  25900=>"111000111",
  25901=>"001100100",
  25902=>"001101100",
  25903=>"001100111",
  25904=>"101110100",
  25905=>"101101100",
  25906=>"110001110",
  25907=>"101110001",
  25908=>"110110100",
  25909=>"010110010",
  25910=>"110111001",
  25911=>"010101001",
  25912=>"001101101",
  25913=>"100101110",
  25914=>"010100011",
  25915=>"110000001",
  25916=>"100000010",
  25917=>"011100010",
  25918=>"010110000",
  25919=>"110101110",
  25920=>"101011101",
  25921=>"101101101",
  25922=>"101100011",
  25923=>"010110101",
  25924=>"011001010",
  25925=>"110001001",
  25926=>"000010001",
  25927=>"100101010",
  25928=>"010011010",
  25929=>"010100100",
  25930=>"101111100",
  25931=>"101000001",
  25932=>"010010111",
  25933=>"010111110",
  25934=>"000000001",
  25935=>"010010011",
  25936=>"111100011",
  25937=>"111110001",
  25938=>"000000111",
  25939=>"101111011",
  25940=>"110001111",
  25941=>"001101000",
  25942=>"000101111",
  25943=>"110111010",
  25944=>"011110100",
  25945=>"110010011",
  25946=>"101000011",
  25947=>"000110010",
  25948=>"111000011",
  25949=>"101000001",
  25950=>"010111001",
  25951=>"010011110",
  25952=>"101101111",
  25953=>"110011111",
  25954=>"000001010",
  25955=>"111111110",
  25956=>"111001111",
  25957=>"010101110",
  25958=>"100011001",
  25959=>"100110111",
  25960=>"000110101",
  25961=>"100111110",
  25962=>"100111011",
  25963=>"101101000",
  25964=>"000001010",
  25965=>"000101110",
  25966=>"111101110",
  25967=>"100011111",
  25968=>"111110001",
  25969=>"100111101",
  25970=>"000010111",
  25971=>"100010001",
  25972=>"110000001",
  25973=>"111001111",
  25974=>"011100011",
  25975=>"100110101",
  25976=>"101010000",
  25977=>"010010110",
  25978=>"000010110",
  25979=>"100111001",
  25980=>"111100010",
  25981=>"001011011",
  25982=>"110010110",
  25983=>"100010110",
  25984=>"010001001",
  25985=>"011010010",
  25986=>"101101011",
  25987=>"000110000",
  25988=>"011111011",
  25989=>"101111100",
  25990=>"111010110",
  25991=>"010000000",
  25992=>"110111000",
  25993=>"001010000",
  25994=>"011001001",
  25995=>"001101010",
  25996=>"100011100",
  25997=>"000011101",
  25998=>"000010101",
  25999=>"011011111",
  26000=>"111011000",
  26001=>"010001010",
  26002=>"101000111",
  26003=>"111101100",
  26004=>"101011111",
  26005=>"000111001",
  26006=>"000101011",
  26007=>"011100001",
  26008=>"101110000",
  26009=>"010101011",
  26010=>"100001011",
  26011=>"000000011",
  26012=>"000001101",
  26013=>"001001000",
  26014=>"011000010",
  26015=>"101110110",
  26016=>"110110000",
  26017=>"111011111",
  26018=>"000000010",
  26019=>"011101111",
  26020=>"111010010",
  26021=>"110011001",
  26022=>"111010100",
  26023=>"111010100",
  26024=>"011001010",
  26025=>"100000011",
  26026=>"001011100",
  26027=>"010010100",
  26028=>"010111010",
  26029=>"000001001",
  26030=>"101001001",
  26031=>"000111110",
  26032=>"011000100",
  26033=>"100101111",
  26034=>"010010000",
  26035=>"001111111",
  26036=>"111100010",
  26037=>"101111111",
  26038=>"011011000",
  26039=>"111011111",
  26040=>"110011000",
  26041=>"111001010",
  26042=>"011011010",
  26043=>"111001110",
  26044=>"110110110",
  26045=>"001101000",
  26046=>"111001101",
  26047=>"001011010",
  26048=>"000110110",
  26049=>"000110100",
  26050=>"011001010",
  26051=>"000111101",
  26052=>"101011111",
  26053=>"100110001",
  26054=>"000010011",
  26055=>"000100111",
  26056=>"001101111",
  26057=>"110110100",
  26058=>"001100101",
  26059=>"000000000",
  26060=>"111011011",
  26061=>"111110000",
  26062=>"000101000",
  26063=>"000110000",
  26064=>"001100111",
  26065=>"100010111",
  26066=>"010101000",
  26067=>"100011010",
  26068=>"011000010",
  26069=>"011001110",
  26070=>"110001101",
  26071=>"000011000",
  26072=>"111111101",
  26073=>"110111010",
  26074=>"101000110",
  26075=>"000010011",
  26076=>"110000001",
  26077=>"001111011",
  26078=>"010000010",
  26079=>"101010111",
  26080=>"000001111",
  26081=>"001111000",
  26082=>"001010000",
  26083=>"111010101",
  26084=>"011001000",
  26085=>"111110111",
  26086=>"011001011",
  26087=>"011101010",
  26088=>"011000100",
  26089=>"011111101",
  26090=>"101010010",
  26091=>"101000110",
  26092=>"001110011",
  26093=>"110001000",
  26094=>"110111001",
  26095=>"110011000",
  26096=>"010001011",
  26097=>"000011000",
  26098=>"110010111",
  26099=>"010100100",
  26100=>"010001000",
  26101=>"111100011",
  26102=>"101111110",
  26103=>"000111101",
  26104=>"101101010",
  26105=>"001010001",
  26106=>"101101011",
  26107=>"011000010",
  26108=>"111101100",
  26109=>"101100000",
  26110=>"100011101",
  26111=>"111100100",
  26112=>"111010010",
  26113=>"000011111",
  26114=>"011010111",
  26115=>"011001011",
  26116=>"001101010",
  26117=>"110110000",
  26118=>"101100011",
  26119=>"011011100",
  26120=>"100001011",
  26121=>"100100111",
  26122=>"001011110",
  26123=>"101110000",
  26124=>"111101001",
  26125=>"101011110",
  26126=>"111010000",
  26127=>"110111101",
  26128=>"011000011",
  26129=>"000010001",
  26130=>"110101110",
  26131=>"010101101",
  26132=>"111111001",
  26133=>"110001011",
  26134=>"111110011",
  26135=>"101101001",
  26136=>"001101111",
  26137=>"010010010",
  26138=>"001011001",
  26139=>"110011010",
  26140=>"101011000",
  26141=>"010001000",
  26142=>"001000000",
  26143=>"011010000",
  26144=>"001110110",
  26145=>"000111111",
  26146=>"000101010",
  26147=>"100100010",
  26148=>"110100001",
  26149=>"010011000",
  26150=>"010111101",
  26151=>"010110110",
  26152=>"100010010",
  26153=>"110000000",
  26154=>"000110001",
  26155=>"110111000",
  26156=>"000001101",
  26157=>"100101100",
  26158=>"111101101",
  26159=>"000100111",
  26160=>"100100100",
  26161=>"110001110",
  26162=>"010001000",
  26163=>"101010111",
  26164=>"011000101",
  26165=>"001001100",
  26166=>"000011010",
  26167=>"100101111",
  26168=>"000010100",
  26169=>"100101011",
  26170=>"000011010",
  26171=>"111100110",
  26172=>"101001110",
  26173=>"110000011",
  26174=>"101100111",
  26175=>"010011101",
  26176=>"011100111",
  26177=>"110111011",
  26178=>"100000111",
  26179=>"111101010",
  26180=>"111001110",
  26181=>"100000010",
  26182=>"011000110",
  26183=>"110100111",
  26184=>"011101111",
  26185=>"001010011",
  26186=>"000111110",
  26187=>"000111100",
  26188=>"001001110",
  26189=>"001100000",
  26190=>"101100101",
  26191=>"010100100",
  26192=>"101100111",
  26193=>"001010010",
  26194=>"101011011",
  26195=>"101010110",
  26196=>"000110111",
  26197=>"100011000",
  26198=>"010000010",
  26199=>"011011011",
  26200=>"001000110",
  26201=>"010101110",
  26202=>"011010011",
  26203=>"101110010",
  26204=>"110110010",
  26205=>"000010001",
  26206=>"111000111",
  26207=>"101000100",
  26208=>"101000110",
  26209=>"000011100",
  26210=>"011110111",
  26211=>"110001100",
  26212=>"001111011",
  26213=>"111011111",
  26214=>"000101000",
  26215=>"001011001",
  26216=>"000101001",
  26217=>"000001011",
  26218=>"011110000",
  26219=>"010011000",
  26220=>"110110000",
  26221=>"010000000",
  26222=>"011110011",
  26223=>"000000110",
  26224=>"110010111",
  26225=>"100001001",
  26226=>"110111001",
  26227=>"011010000",
  26228=>"110110111",
  26229=>"001100010",
  26230=>"010000001",
  26231=>"110110011",
  26232=>"001110111",
  26233=>"110100010",
  26234=>"011110101",
  26235=>"010011111",
  26236=>"000000101",
  26237=>"001000000",
  26238=>"001000000",
  26239=>"000111010",
  26240=>"100101010",
  26241=>"010001001",
  26242=>"111000000",
  26243=>"110101001",
  26244=>"000011101",
  26245=>"000100101",
  26246=>"111100110",
  26247=>"000000111",
  26248=>"011010110",
  26249=>"010110000",
  26250=>"000100000",
  26251=>"011001000",
  26252=>"000100010",
  26253=>"010100111",
  26254=>"000000010",
  26255=>"100111000",
  26256=>"111001111",
  26257=>"010010000",
  26258=>"001001010",
  26259=>"011001011",
  26260=>"011101100",
  26261=>"001000010",
  26262=>"100000001",
  26263=>"111111111",
  26264=>"001000011",
  26265=>"010000111",
  26266=>"000111111",
  26267=>"001100101",
  26268=>"011110001",
  26269=>"101011011",
  26270=>"101000101",
  26271=>"100100000",
  26272=>"000011000",
  26273=>"000010011",
  26274=>"110111101",
  26275=>"001010100",
  26276=>"010111111",
  26277=>"001000011",
  26278=>"111110011",
  26279=>"100111010",
  26280=>"111111111",
  26281=>"101010001",
  26282=>"010001001",
  26283=>"000011001",
  26284=>"011001000",
  26285=>"111111010",
  26286=>"010111110",
  26287=>"000010111",
  26288=>"001100111",
  26289=>"101001101",
  26290=>"000101000",
  26291=>"110101101",
  26292=>"110101100",
  26293=>"001100000",
  26294=>"011111111",
  26295=>"011011111",
  26296=>"100010001",
  26297=>"001100001",
  26298=>"111000000",
  26299=>"110000111",
  26300=>"100001010",
  26301=>"110110010",
  26302=>"100100011",
  26303=>"110101110",
  26304=>"110111001",
  26305=>"001111110",
  26306=>"011100000",
  26307=>"000010000",
  26308=>"110111001",
  26309=>"000000001",
  26310=>"101001000",
  26311=>"111110000",
  26312=>"101101110",
  26313=>"111011010",
  26314=>"100010011",
  26315=>"111010100",
  26316=>"110110011",
  26317=>"010010101",
  26318=>"110110111",
  26319=>"101000001",
  26320=>"000000100",
  26321=>"001100010",
  26322=>"011010110",
  26323=>"000001000",
  26324=>"100110101",
  26325=>"010001100",
  26326=>"010101010",
  26327=>"011101100",
  26328=>"001011111",
  26329=>"111011110",
  26330=>"111101111",
  26331=>"011110110",
  26332=>"101011000",
  26333=>"001010010",
  26334=>"100010111",
  26335=>"010010000",
  26336=>"100000110",
  26337=>"010111011",
  26338=>"000000010",
  26339=>"010111111",
  26340=>"001110110",
  26341=>"110000011",
  26342=>"100010011",
  26343=>"110101011",
  26344=>"110110111",
  26345=>"100011101",
  26346=>"111111001",
  26347=>"110010111",
  26348=>"000010000",
  26349=>"110101101",
  26350=>"001001100",
  26351=>"111111111",
  26352=>"001110111",
  26353=>"111100000",
  26354=>"001101110",
  26355=>"111001111",
  26356=>"011110010",
  26357=>"101101000",
  26358=>"011111111",
  26359=>"110110000",
  26360=>"000111010",
  26361=>"010010001",
  26362=>"111010100",
  26363=>"101011111",
  26364=>"111101001",
  26365=>"111111100",
  26366=>"111010111",
  26367=>"111100100",
  26368=>"000011010",
  26369=>"101101000",
  26370=>"010001010",
  26371=>"100101000",
  26372=>"010010001",
  26373=>"101000001",
  26374=>"010000101",
  26375=>"010011001",
  26376=>"111001101",
  26377=>"111110111",
  26378=>"111001001",
  26379=>"001110001",
  26380=>"111101010",
  26381=>"000111101",
  26382=>"101010001",
  26383=>"010001100",
  26384=>"001110110",
  26385=>"110001010",
  26386=>"010001000",
  26387=>"000010000",
  26388=>"001101100",
  26389=>"011111000",
  26390=>"100011110",
  26391=>"111100100",
  26392=>"000111111",
  26393=>"010000110",
  26394=>"111101110",
  26395=>"000100110",
  26396=>"101111110",
  26397=>"011000101",
  26398=>"111110010",
  26399=>"111001110",
  26400=>"110110010",
  26401=>"110000000",
  26402=>"001000011",
  26403=>"001110111",
  26404=>"110010010",
  26405=>"101100101",
  26406=>"101100000",
  26407=>"000000100",
  26408=>"011001110",
  26409=>"111001011",
  26410=>"000011001",
  26411=>"100001110",
  26412=>"100000011",
  26413=>"011100011",
  26414=>"010010000",
  26415=>"000110100",
  26416=>"011111111",
  26417=>"111111100",
  26418=>"111001111",
  26419=>"001000100",
  26420=>"001001110",
  26421=>"000100010",
  26422=>"101000001",
  26423=>"000111001",
  26424=>"110101001",
  26425=>"001001011",
  26426=>"010000010",
  26427=>"100111110",
  26428=>"010010101",
  26429=>"100110111",
  26430=>"001001011",
  26431=>"010010111",
  26432=>"011100011",
  26433=>"100100100",
  26434=>"010111000",
  26435=>"000011011",
  26436=>"001111010",
  26437=>"101000000",
  26438=>"101110110",
  26439=>"000001101",
  26440=>"100010101",
  26441=>"001110010",
  26442=>"111101010",
  26443=>"000001101",
  26444=>"001110110",
  26445=>"001011011",
  26446=>"000001100",
  26447=>"111101100",
  26448=>"110000001",
  26449=>"000011101",
  26450=>"100000110",
  26451=>"000110010",
  26452=>"011001110",
  26453=>"011000010",
  26454=>"110101000",
  26455=>"000111111",
  26456=>"000110010",
  26457=>"010101101",
  26458=>"110000011",
  26459=>"000011110",
  26460=>"111001010",
  26461=>"111100000",
  26462=>"110011101",
  26463=>"000000000",
  26464=>"000101111",
  26465=>"100011111",
  26466=>"110110111",
  26467=>"101101010",
  26468=>"000100111",
  26469=>"001000010",
  26470=>"101111010",
  26471=>"011111101",
  26472=>"010001001",
  26473=>"100110110",
  26474=>"111110100",
  26475=>"000110010",
  26476=>"100101001",
  26477=>"001110110",
  26478=>"111111000",
  26479=>"011000000",
  26480=>"001111110",
  26481=>"100111011",
  26482=>"111010011",
  26483=>"000110110",
  26484=>"000110111",
  26485=>"001110100",
  26486=>"100000110",
  26487=>"011001011",
  26488=>"010000000",
  26489=>"101111100",
  26490=>"011011001",
  26491=>"011101010",
  26492=>"100011100",
  26493=>"010000011",
  26494=>"100110100",
  26495=>"010000111",
  26496=>"000000110",
  26497=>"100100010",
  26498=>"011111011",
  26499=>"000010100",
  26500=>"110000101",
  26501=>"011010101",
  26502=>"000111101",
  26503=>"011101100",
  26504=>"001000111",
  26505=>"111000101",
  26506=>"101001011",
  26507=>"010001000",
  26508=>"010101100",
  26509=>"100100010",
  26510=>"000011111",
  26511=>"110101110",
  26512=>"111111011",
  26513=>"001110111",
  26514=>"100100110",
  26515=>"010101000",
  26516=>"001110101",
  26517=>"100100010",
  26518=>"011100100",
  26519=>"111011000",
  26520=>"011111001",
  26521=>"000010010",
  26522=>"011001000",
  26523=>"011111010",
  26524=>"101110000",
  26525=>"001100000",
  26526=>"111000000",
  26527=>"111111011",
  26528=>"111100010",
  26529=>"010010000",
  26530=>"111110101",
  26531=>"100110100",
  26532=>"000000010",
  26533=>"101110011",
  26534=>"101001010",
  26535=>"101101000",
  26536=>"010111100",
  26537=>"100101001",
  26538=>"001101011",
  26539=>"001001011",
  26540=>"010011101",
  26541=>"111111011",
  26542=>"110100001",
  26543=>"001101000",
  26544=>"111010000",
  26545=>"001101001",
  26546=>"100000000",
  26547=>"111001101",
  26548=>"110101110",
  26549=>"100111100",
  26550=>"000100000",
  26551=>"001110010",
  26552=>"100000011",
  26553=>"010001110",
  26554=>"101001111",
  26555=>"110111011",
  26556=>"001000010",
  26557=>"110010010",
  26558=>"110100101",
  26559=>"001010100",
  26560=>"010000011",
  26561=>"011110101",
  26562=>"100101110",
  26563=>"100001110",
  26564=>"100100101",
  26565=>"100110101",
  26566=>"100111010",
  26567=>"111010111",
  26568=>"100100001",
  26569=>"000111011",
  26570=>"100101110",
  26571=>"111111100",
  26572=>"000011100",
  26573=>"111100101",
  26574=>"010111010",
  26575=>"101110001",
  26576=>"000110001",
  26577=>"010111100",
  26578=>"110100000",
  26579=>"100011100",
  26580=>"111111111",
  26581=>"101100100",
  26582=>"001010101",
  26583=>"001101010",
  26584=>"111000111",
  26585=>"100001111",
  26586=>"000100111",
  26587=>"110110000",
  26588=>"111010000",
  26589=>"010000111",
  26590=>"111001101",
  26591=>"111011010",
  26592=>"001101111",
  26593=>"100111110",
  26594=>"000100101",
  26595=>"101000110",
  26596=>"011111011",
  26597=>"111110010",
  26598=>"000011010",
  26599=>"000101000",
  26600=>"000010100",
  26601=>"111001001",
  26602=>"000011000",
  26603=>"011000101",
  26604=>"100111100",
  26605=>"000001010",
  26606=>"001001001",
  26607=>"001011011",
  26608=>"001010110",
  26609=>"100101111",
  26610=>"010110101",
  26611=>"000011011",
  26612=>"100100010",
  26613=>"101000000",
  26614=>"111101011",
  26615=>"010111111",
  26616=>"011100011",
  26617=>"101011111",
  26618=>"010111010",
  26619=>"011011100",
  26620=>"010110110",
  26621=>"011010110",
  26622=>"001000000",
  26623=>"101101000",
  26624=>"010001101",
  26625=>"000010111",
  26626=>"011011110",
  26627=>"001100110",
  26628=>"011101010",
  26629=>"111011100",
  26630=>"100000100",
  26631=>"010111110",
  26632=>"111010110",
  26633=>"010100111",
  26634=>"111110000",
  26635=>"100011000",
  26636=>"100101010",
  26637=>"000101010",
  26638=>"111011111",
  26639=>"101111110",
  26640=>"011111110",
  26641=>"001101010",
  26642=>"011101111",
  26643=>"110111011",
  26644=>"001010111",
  26645=>"100010100",
  26646=>"010101111",
  26647=>"100111010",
  26648=>"111001100",
  26649=>"110000110",
  26650=>"011110000",
  26651=>"011101110",
  26652=>"001100011",
  26653=>"010000001",
  26654=>"001110101",
  26655=>"001001100",
  26656=>"001000000",
  26657=>"111100011",
  26658=>"111110111",
  26659=>"001000111",
  26660=>"010010100",
  26661=>"010001100",
  26662=>"011100101",
  26663=>"001110010",
  26664=>"010111010",
  26665=>"000000000",
  26666=>"001001111",
  26667=>"001000101",
  26668=>"001111100",
  26669=>"100011101",
  26670=>"011001000",
  26671=>"000000100",
  26672=>"110011011",
  26673=>"001010101",
  26674=>"110000111",
  26675=>"111011011",
  26676=>"001101001",
  26677=>"001001001",
  26678=>"011010000",
  26679=>"111111000",
  26680=>"111111110",
  26681=>"001011101",
  26682=>"000101010",
  26683=>"010010101",
  26684=>"011110111",
  26685=>"001111001",
  26686=>"010010111",
  26687=>"010101110",
  26688=>"000011011",
  26689=>"111100100",
  26690=>"110011001",
  26691=>"010101001",
  26692=>"110000100",
  26693=>"111011000",
  26694=>"010011110",
  26695=>"000000010",
  26696=>"101101110",
  26697=>"010010010",
  26698=>"001010110",
  26699=>"100011010",
  26700=>"101101101",
  26701=>"011111101",
  26702=>"110010100",
  26703=>"100110011",
  26704=>"101011101",
  26705=>"110011100",
  26706=>"101011000",
  26707=>"011101110",
  26708=>"000100001",
  26709=>"110010111",
  26710=>"010101001",
  26711=>"011000111",
  26712=>"000100001",
  26713=>"111011111",
  26714=>"110101110",
  26715=>"101000000",
  26716=>"000000100",
  26717=>"110011010",
  26718=>"001100111",
  26719=>"011100000",
  26720=>"010101101",
  26721=>"010101111",
  26722=>"001111100",
  26723=>"101100000",
  26724=>"111001001",
  26725=>"101101101",
  26726=>"011010010",
  26727=>"010101001",
  26728=>"010010000",
  26729=>"110000011",
  26730=>"011100111",
  26731=>"110110000",
  26732=>"100100000",
  26733=>"011000110",
  26734=>"010001111",
  26735=>"101001101",
  26736=>"100101101",
  26737=>"101000111",
  26738=>"000101101",
  26739=>"010000000",
  26740=>"110110110",
  26741=>"010111111",
  26742=>"110111110",
  26743=>"110111000",
  26744=>"000101111",
  26745=>"100010001",
  26746=>"000001000",
  26747=>"000101101",
  26748=>"001100010",
  26749=>"100001101",
  26750=>"110110101",
  26751=>"011011110",
  26752=>"001000110",
  26753=>"011001010",
  26754=>"100000101",
  26755=>"101000100",
  26756=>"111000111",
  26757=>"010110000",
  26758=>"001011011",
  26759=>"011011001",
  26760=>"101000000",
  26761=>"000110010",
  26762=>"110000011",
  26763=>"011101100",
  26764=>"011101101",
  26765=>"101110001",
  26766=>"010011100",
  26767=>"101001110",
  26768=>"100110110",
  26769=>"010111110",
  26770=>"111011000",
  26771=>"011010000",
  26772=>"101100000",
  26773=>"000001001",
  26774=>"011001000",
  26775=>"001001010",
  26776=>"000001001",
  26777=>"000110000",
  26778=>"000111000",
  26779=>"011100001",
  26780=>"101110100",
  26781=>"100111000",
  26782=>"000011000",
  26783=>"000011000",
  26784=>"000111111",
  26785=>"101101001",
  26786=>"001110110",
  26787=>"011001111",
  26788=>"110010100",
  26789=>"011000111",
  26790=>"010000111",
  26791=>"110100001",
  26792=>"100010011",
  26793=>"011010000",
  26794=>"111010010",
  26795=>"101011101",
  26796=>"001101000",
  26797=>"110110100",
  26798=>"100110010",
  26799=>"011101100",
  26800=>"011100001",
  26801=>"000111101",
  26802=>"000010110",
  26803=>"100001100",
  26804=>"110001111",
  26805=>"101100011",
  26806=>"011110111",
  26807=>"111101100",
  26808=>"100011110",
  26809=>"001111111",
  26810=>"111000010",
  26811=>"111101100",
  26812=>"000000001",
  26813=>"111010111",
  26814=>"111100001",
  26815=>"101010111",
  26816=>"000011110",
  26817=>"001101000",
  26818=>"000100101",
  26819=>"011001001",
  26820=>"101000011",
  26821=>"110001011",
  26822=>"110010110",
  26823=>"100111000",
  26824=>"001101101",
  26825=>"111110000",
  26826=>"001001011",
  26827=>"010001011",
  26828=>"111011001",
  26829=>"100100110",
  26830=>"100000100",
  26831=>"110001110",
  26832=>"111100101",
  26833=>"000101100",
  26834=>"111011001",
  26835=>"101111111",
  26836=>"111010111",
  26837=>"001000010",
  26838=>"000000100",
  26839=>"000001011",
  26840=>"000000011",
  26841=>"110101010",
  26842=>"111011011",
  26843=>"100111110",
  26844=>"010011110",
  26845=>"011100100",
  26846=>"110010001",
  26847=>"000000010",
  26848=>"001111110",
  26849=>"101000000",
  26850=>"111001100",
  26851=>"001110111",
  26852=>"000011001",
  26853=>"110000010",
  26854=>"000010010",
  26855=>"101111110",
  26856=>"101100110",
  26857=>"111110001",
  26858=>"001011000",
  26859=>"100010110",
  26860=>"001001110",
  26861=>"100111001",
  26862=>"000000000",
  26863=>"111000010",
  26864=>"100100010",
  26865=>"101010000",
  26866=>"010111110",
  26867=>"110101001",
  26868=>"001000011",
  26869=>"000110001",
  26870=>"000010111",
  26871=>"010000010",
  26872=>"100111111",
  26873=>"100100010",
  26874=>"111101111",
  26875=>"001110000",
  26876=>"001001000",
  26877=>"000001000",
  26878=>"100100110",
  26879=>"111111111",
  26880=>"111001001",
  26881=>"010010001",
  26882=>"001011111",
  26883=>"110001000",
  26884=>"101111101",
  26885=>"011011101",
  26886=>"011101101",
  26887=>"100000110",
  26888=>"010001001",
  26889=>"111110011",
  26890=>"111111101",
  26891=>"001111001",
  26892=>"101000110",
  26893=>"010111110",
  26894=>"001000010",
  26895=>"100010100",
  26896=>"001101100",
  26897=>"100110101",
  26898=>"101111111",
  26899=>"011001010",
  26900=>"111101100",
  26901=>"010111111",
  26902=>"010010000",
  26903=>"001101111",
  26904=>"110010001",
  26905=>"010000011",
  26906=>"011111000",
  26907=>"101010101",
  26908=>"010010001",
  26909=>"010110110",
  26910=>"010011010",
  26911=>"101110110",
  26912=>"001100101",
  26913=>"000011110",
  26914=>"000110110",
  26915=>"111110000",
  26916=>"001000111",
  26917=>"001110110",
  26918=>"100100101",
  26919=>"010000101",
  26920=>"001011101",
  26921=>"000011111",
  26922=>"101000010",
  26923=>"111110011",
  26924=>"011111010",
  26925=>"011111110",
  26926=>"001100110",
  26927=>"101101000",
  26928=>"010011011",
  26929=>"110011111",
  26930=>"000000111",
  26931=>"001100111",
  26932=>"010111011",
  26933=>"111111010",
  26934=>"011000010",
  26935=>"111110010",
  26936=>"000101011",
  26937=>"011100111",
  26938=>"111011110",
  26939=>"110110010",
  26940=>"100000000",
  26941=>"100001100",
  26942=>"010111111",
  26943=>"011111000",
  26944=>"100101100",
  26945=>"100100110",
  26946=>"100111011",
  26947=>"011100100",
  26948=>"101111010",
  26949=>"110101000",
  26950=>"100111000",
  26951=>"110010110",
  26952=>"111010011",
  26953=>"111010001",
  26954=>"011001010",
  26955=>"101101000",
  26956=>"101100001",
  26957=>"110011100",
  26958=>"011101100",
  26959=>"010011001",
  26960=>"010000011",
  26961=>"100101010",
  26962=>"000001100",
  26963=>"001010101",
  26964=>"101101101",
  26965=>"011001010",
  26966=>"111001111",
  26967=>"001101010",
  26968=>"110100101",
  26969=>"010011010",
  26970=>"111111011",
  26971=>"011011101",
  26972=>"010101111",
  26973=>"110110101",
  26974=>"011010101",
  26975=>"001001110",
  26976=>"011111010",
  26977=>"101100010",
  26978=>"000110100",
  26979=>"000110011",
  26980=>"000110001",
  26981=>"110101110",
  26982=>"011011101",
  26983=>"010011111",
  26984=>"010101001",
  26985=>"101000110",
  26986=>"001010100",
  26987=>"111110011",
  26988=>"011000110",
  26989=>"000110000",
  26990=>"100110000",
  26991=>"001111110",
  26992=>"101010011",
  26993=>"011111110",
  26994=>"011000111",
  26995=>"110101111",
  26996=>"110100111",
  26997=>"010010010",
  26998=>"110011100",
  26999=>"001111111",
  27000=>"101100010",
  27001=>"010000001",
  27002=>"001001011",
  27003=>"111111001",
  27004=>"111011001",
  27005=>"110010000",
  27006=>"011011101",
  27007=>"010011110",
  27008=>"011000001",
  27009=>"110110111",
  27010=>"000011011",
  27011=>"111110110",
  27012=>"000010101",
  27013=>"011110111",
  27014=>"101101001",
  27015=>"110110100",
  27016=>"001001001",
  27017=>"001001110",
  27018=>"100111001",
  27019=>"110100011",
  27020=>"101111111",
  27021=>"001011000",
  27022=>"011100101",
  27023=>"111111111",
  27024=>"010111010",
  27025=>"111110111",
  27026=>"111111010",
  27027=>"011110101",
  27028=>"011000100",
  27029=>"000111101",
  27030=>"100101000",
  27031=>"011011100",
  27032=>"011101100",
  27033=>"001100001",
  27034=>"110101101",
  27035=>"001101111",
  27036=>"000100101",
  27037=>"110101111",
  27038=>"110001111",
  27039=>"001001011",
  27040=>"101101110",
  27041=>"010101001",
  27042=>"101001000",
  27043=>"011000010",
  27044=>"110101100",
  27045=>"101111001",
  27046=>"000000001",
  27047=>"100111100",
  27048=>"110110001",
  27049=>"110101010",
  27050=>"000110111",
  27051=>"111101101",
  27052=>"001001011",
  27053=>"100100100",
  27054=>"010111110",
  27055=>"100001101",
  27056=>"001101000",
  27057=>"100100101",
  27058=>"000111001",
  27059=>"100101100",
  27060=>"100101010",
  27061=>"011011000",
  27062=>"110100000",
  27063=>"100011111",
  27064=>"011111010",
  27065=>"111000101",
  27066=>"100110110",
  27067=>"111111101",
  27068=>"001000000",
  27069=>"100010100",
  27070=>"001000010",
  27071=>"011100010",
  27072=>"001011000",
  27073=>"001000010",
  27074=>"100001111",
  27075=>"111011011",
  27076=>"001100110",
  27077=>"010110011",
  27078=>"000100000",
  27079=>"011100110",
  27080=>"100000110",
  27081=>"000001100",
  27082=>"110110110",
  27083=>"110000000",
  27084=>"011101001",
  27085=>"011011010",
  27086=>"100111101",
  27087=>"001111111",
  27088=>"110010011",
  27089=>"100110100",
  27090=>"100101100",
  27091=>"011111000",
  27092=>"000111010",
  27093=>"001011110",
  27094=>"000100001",
  27095=>"101100010",
  27096=>"111010101",
  27097=>"101101010",
  27098=>"101011000",
  27099=>"011000110",
  27100=>"001101100",
  27101=>"101101001",
  27102=>"111111000",
  27103=>"111101101",
  27104=>"010101101",
  27105=>"100001101",
  27106=>"100101000",
  27107=>"011000001",
  27108=>"111100010",
  27109=>"100011110",
  27110=>"111010111",
  27111=>"001110111",
  27112=>"010111010",
  27113=>"011001100",
  27114=>"000110100",
  27115=>"100010001",
  27116=>"101000111",
  27117=>"000100100",
  27118=>"010010000",
  27119=>"011011110",
  27120=>"010000111",
  27121=>"110000000",
  27122=>"111111001",
  27123=>"011100001",
  27124=>"110110001",
  27125=>"100110000",
  27126=>"011110001",
  27127=>"011101000",
  27128=>"111111110",
  27129=>"011110001",
  27130=>"111110111",
  27131=>"111100101",
  27132=>"100110110",
  27133=>"010100100",
  27134=>"111001100",
  27135=>"011001001",
  27136=>"111100001",
  27137=>"111101110",
  27138=>"001111111",
  27139=>"110001111",
  27140=>"001110101",
  27141=>"000011000",
  27142=>"110101101",
  27143=>"111110011",
  27144=>"000111000",
  27145=>"110110110",
  27146=>"010010100",
  27147=>"111110000",
  27148=>"111110000",
  27149=>"110110101",
  27150=>"011010011",
  27151=>"000011110",
  27152=>"101010110",
  27153=>"100010010",
  27154=>"111000011",
  27155=>"001100000",
  27156=>"001110101",
  27157=>"111101100",
  27158=>"100111101",
  27159=>"110100110",
  27160=>"001110111",
  27161=>"100110001",
  27162=>"101100010",
  27163=>"100100000",
  27164=>"101011001",
  27165=>"010011100",
  27166=>"110110111",
  27167=>"011001001",
  27168=>"010100100",
  27169=>"110001000",
  27170=>"010111110",
  27171=>"101000100",
  27172=>"011001011",
  27173=>"001111010",
  27174=>"000001110",
  27175=>"000110011",
  27176=>"100101101",
  27177=>"000001110",
  27178=>"110101010",
  27179=>"111010101",
  27180=>"011110001",
  27181=>"000010110",
  27182=>"111001010",
  27183=>"001000100",
  27184=>"111011101",
  27185=>"110010001",
  27186=>"110111010",
  27187=>"010101001",
  27188=>"001110101",
  27189=>"000111001",
  27190=>"100110001",
  27191=>"100000101",
  27192=>"100101110",
  27193=>"011100001",
  27194=>"111111110",
  27195=>"011110000",
  27196=>"100010101",
  27197=>"010011111",
  27198=>"010001100",
  27199=>"011000101",
  27200=>"100101000",
  27201=>"110000000",
  27202=>"001101111",
  27203=>"100110011",
  27204=>"111011111",
  27205=>"111011011",
  27206=>"101000100",
  27207=>"101001100",
  27208=>"001100000",
  27209=>"000011101",
  27210=>"011001001",
  27211=>"100100100",
  27212=>"010101011",
  27213=>"101111001",
  27214=>"000100000",
  27215=>"101001001",
  27216=>"101110101",
  27217=>"001000000",
  27218=>"001101110",
  27219=>"000111101",
  27220=>"111100001",
  27221=>"111111011",
  27222=>"000101101",
  27223=>"110111100",
  27224=>"111000011",
  27225=>"101101111",
  27226=>"001010000",
  27227=>"000011100",
  27228=>"100100011",
  27229=>"110101111",
  27230=>"110110110",
  27231=>"110101100",
  27232=>"000111001",
  27233=>"101100110",
  27234=>"110101000",
  27235=>"101011011",
  27236=>"110110101",
  27237=>"111010111",
  27238=>"110010110",
  27239=>"111110111",
  27240=>"000001010",
  27241=>"111001000",
  27242=>"111111001",
  27243=>"111111110",
  27244=>"001110000",
  27245=>"000000010",
  27246=>"000111101",
  27247=>"010000010",
  27248=>"100111011",
  27249=>"111111011",
  27250=>"001111011",
  27251=>"101111100",
  27252=>"100011111",
  27253=>"011100011",
  27254=>"101111100",
  27255=>"101001011",
  27256=>"101100001",
  27257=>"001101110",
  27258=>"110110111",
  27259=>"010000001",
  27260=>"010100001",
  27261=>"101110111",
  27262=>"001110101",
  27263=>"110111111",
  27264=>"010001110",
  27265=>"010001101",
  27266=>"101101101",
  27267=>"000001100",
  27268=>"010110010",
  27269=>"110001110",
  27270=>"110101111",
  27271=>"011101101",
  27272=>"111001001",
  27273=>"000110110",
  27274=>"100111100",
  27275=>"001101001",
  27276=>"110101011",
  27277=>"011000001",
  27278=>"010010110",
  27279=>"110110100",
  27280=>"011110111",
  27281=>"111111101",
  27282=>"100010101",
  27283=>"100001001",
  27284=>"100100110",
  27285=>"000100010",
  27286=>"000100011",
  27287=>"110001111",
  27288=>"100000101",
  27289=>"000111110",
  27290=>"011011011",
  27291=>"111111010",
  27292=>"100110001",
  27293=>"110000001",
  27294=>"101000110",
  27295=>"000010000",
  27296=>"010110110",
  27297=>"110100000",
  27298=>"101011001",
  27299=>"100010111",
  27300=>"101101100",
  27301=>"111111111",
  27302=>"111111100",
  27303=>"110111000",
  27304=>"000001100",
  27305=>"111010001",
  27306=>"111111010",
  27307=>"100101010",
  27308=>"100110111",
  27309=>"111101111",
  27310=>"010010110",
  27311=>"111111010",
  27312=>"000110111",
  27313=>"000110101",
  27314=>"111011110",
  27315=>"101011111",
  27316=>"001100010",
  27317=>"001000100",
  27318=>"000111110",
  27319=>"100110110",
  27320=>"110001101",
  27321=>"000110110",
  27322=>"001000101",
  27323=>"111000111",
  27324=>"001010011",
  27325=>"100100101",
  27326=>"110111010",
  27327=>"100110110",
  27328=>"000111011",
  27329=>"000010010",
  27330=>"111111111",
  27331=>"100110000",
  27332=>"101111001",
  27333=>"000110111",
  27334=>"010101100",
  27335=>"001011011",
  27336=>"111110001",
  27337=>"011010111",
  27338=>"011111111",
  27339=>"010111111",
  27340=>"111100000",
  27341=>"111000110",
  27342=>"100010100",
  27343=>"111011010",
  27344=>"110100000",
  27345=>"010101110",
  27346=>"100100100",
  27347=>"000001110",
  27348=>"111010111",
  27349=>"110111011",
  27350=>"100101001",
  27351=>"001000010",
  27352=>"101100100",
  27353=>"010101001",
  27354=>"100111101",
  27355=>"000001001",
  27356=>"110011011",
  27357=>"110011011",
  27358=>"111111000",
  27359=>"111101100",
  27360=>"011001100",
  27361=>"011000111",
  27362=>"100111011",
  27363=>"010011000",
  27364=>"111100010",
  27365=>"010001010",
  27366=>"111110000",
  27367=>"001011111",
  27368=>"000101011",
  27369=>"101111111",
  27370=>"011010000",
  27371=>"101101110",
  27372=>"101100001",
  27373=>"111000100",
  27374=>"011010100",
  27375=>"100100111",
  27376=>"100110010",
  27377=>"011111011",
  27378=>"010100011",
  27379=>"110001110",
  27380=>"110111001",
  27381=>"111010011",
  27382=>"011100010",
  27383=>"100111110",
  27384=>"111000010",
  27385=>"111011101",
  27386=>"101011001",
  27387=>"001100111",
  27388=>"101110011",
  27389=>"011011101",
  27390=>"110101000",
  27391=>"111111001",
  27392=>"010100001",
  27393=>"001111110",
  27394=>"110100010",
  27395=>"011101001",
  27396=>"100000000",
  27397=>"001010100",
  27398=>"110000000",
  27399=>"011101100",
  27400=>"010010101",
  27401=>"010010101",
  27402=>"010101000",
  27403=>"110110100",
  27404=>"000000011",
  27405=>"000011000",
  27406=>"011101011",
  27407=>"111101001",
  27408=>"000000100",
  27409=>"011101000",
  27410=>"010101000",
  27411=>"110011101",
  27412=>"010000100",
  27413=>"110110100",
  27414=>"000101111",
  27415=>"000000110",
  27416=>"000010011",
  27417=>"000100011",
  27418=>"110001000",
  27419=>"101110000",
  27420=>"011000010",
  27421=>"101011111",
  27422=>"110000010",
  27423=>"010001100",
  27424=>"111010111",
  27425=>"011010000",
  27426=>"000001100",
  27427=>"101100101",
  27428=>"101110111",
  27429=>"111111110",
  27430=>"111001111",
  27431=>"011111110",
  27432=>"100111000",
  27433=>"010101000",
  27434=>"110101010",
  27435=>"011000111",
  27436=>"010000111",
  27437=>"111111101",
  27438=>"101001111",
  27439=>"100110100",
  27440=>"001100111",
  27441=>"111111110",
  27442=>"000100101",
  27443=>"000101001",
  27444=>"110010100",
  27445=>"110011001",
  27446=>"000010011",
  27447=>"111111111",
  27448=>"111111110",
  27449=>"110011111",
  27450=>"001110000",
  27451=>"010011110",
  27452=>"001100000",
  27453=>"111111001",
  27454=>"001110110",
  27455=>"010100000",
  27456=>"101000101",
  27457=>"010111011",
  27458=>"011101111",
  27459=>"001100111",
  27460=>"100011111",
  27461=>"010111000",
  27462=>"101100101",
  27463=>"110101110",
  27464=>"001001001",
  27465=>"010011001",
  27466=>"011010101",
  27467=>"000110111",
  27468=>"111000101",
  27469=>"010100010",
  27470=>"110000110",
  27471=>"111001111",
  27472=>"100100101",
  27473=>"011011110",
  27474=>"000111100",
  27475=>"011010100",
  27476=>"010001111",
  27477=>"010100000",
  27478=>"010001011",
  27479=>"011010101",
  27480=>"111000011",
  27481=>"111111100",
  27482=>"110011101",
  27483=>"100100001",
  27484=>"111100010",
  27485=>"010000011",
  27486=>"010000110",
  27487=>"101010110",
  27488=>"100100011",
  27489=>"100100111",
  27490=>"111111110",
  27491=>"100100001",
  27492=>"010000111",
  27493=>"000100111",
  27494=>"010110110",
  27495=>"001110010",
  27496=>"000000000",
  27497=>"110001001",
  27498=>"000101000",
  27499=>"110001001",
  27500=>"110000000",
  27501=>"010100011",
  27502=>"100101111",
  27503=>"010011011",
  27504=>"110100010",
  27505=>"000001101",
  27506=>"110111111",
  27507=>"011001010",
  27508=>"010100111",
  27509=>"001100011",
  27510=>"000010000",
  27511=>"000011100",
  27512=>"100001001",
  27513=>"101000111",
  27514=>"000000110",
  27515=>"111101100",
  27516=>"000010110",
  27517=>"010010011",
  27518=>"101111110",
  27519=>"001011000",
  27520=>"110001000",
  27521=>"000001011",
  27522=>"000101010",
  27523=>"000000100",
  27524=>"111100000",
  27525=>"011101001",
  27526=>"110011111",
  27527=>"100001110",
  27528=>"111110111",
  27529=>"011010111",
  27530=>"111100111",
  27531=>"110011110",
  27532=>"010100111",
  27533=>"101100001",
  27534=>"000110011",
  27535=>"110000001",
  27536=>"110110111",
  27537=>"011101000",
  27538=>"010011010",
  27539=>"101101110",
  27540=>"001000000",
  27541=>"111000100",
  27542=>"101100010",
  27543=>"001000001",
  27544=>"101010100",
  27545=>"010101010",
  27546=>"001111110",
  27547=>"110001000",
  27548=>"101010101",
  27549=>"111111011",
  27550=>"111010000",
  27551=>"100010011",
  27552=>"001010100",
  27553=>"010010110",
  27554=>"000001011",
  27555=>"010001101",
  27556=>"010000001",
  27557=>"101100010",
  27558=>"101010110",
  27559=>"110110001",
  27560=>"000000101",
  27561=>"100001110",
  27562=>"000001111",
  27563=>"010001101",
  27564=>"001100000",
  27565=>"001000100",
  27566=>"100001011",
  27567=>"110110010",
  27568=>"011011000",
  27569=>"101111011",
  27570=>"011011000",
  27571=>"111011100",
  27572=>"111101001",
  27573=>"100100101",
  27574=>"010100001",
  27575=>"000110111",
  27576=>"111010011",
  27577=>"010011110",
  27578=>"101100110",
  27579=>"011101000",
  27580=>"000100000",
  27581=>"001011000",
  27582=>"001110000",
  27583=>"100111100",
  27584=>"110010100",
  27585=>"111100111",
  27586=>"001101000",
  27587=>"010111010",
  27588=>"011011001",
  27589=>"000100100",
  27590=>"011111111",
  27591=>"110000111",
  27592=>"010100111",
  27593=>"001111011",
  27594=>"011100110",
  27595=>"000111100",
  27596=>"000100010",
  27597=>"011011111",
  27598=>"110011010",
  27599=>"001011000",
  27600=>"110110111",
  27601=>"000000001",
  27602=>"110101001",
  27603=>"110111111",
  27604=>"111101111",
  27605=>"011110010",
  27606=>"000101111",
  27607=>"000000110",
  27608=>"010110010",
  27609=>"101100011",
  27610=>"000111110",
  27611=>"110110110",
  27612=>"111101101",
  27613=>"111001001",
  27614=>"011100100",
  27615=>"111111110",
  27616=>"001000000",
  27617=>"110010110",
  27618=>"101011100",
  27619=>"011100000",
  27620=>"111100110",
  27621=>"001100000",
  27622=>"111111101",
  27623=>"001011010",
  27624=>"010101111",
  27625=>"111001100",
  27626=>"000001010",
  27627=>"111101011",
  27628=>"111110010",
  27629=>"110101111",
  27630=>"111110101",
  27631=>"010011000",
  27632=>"001110000",
  27633=>"001110010",
  27634=>"111011010",
  27635=>"000010001",
  27636=>"010110110",
  27637=>"000110010",
  27638=>"100001010",
  27639=>"011001010",
  27640=>"110001000",
  27641=>"101000001",
  27642=>"110111011",
  27643=>"101010000",
  27644=>"100100101",
  27645=>"010000100",
  27646=>"110010011",
  27647=>"010010001",
  27648=>"110110101",
  27649=>"001010001",
  27650=>"100101111",
  27651=>"010011001",
  27652=>"011101111",
  27653=>"100100101",
  27654=>"010000001",
  27655=>"000110010",
  27656=>"101011000",
  27657=>"101101111",
  27658=>"100100000",
  27659=>"011100110",
  27660=>"100100110",
  27661=>"000011000",
  27662=>"110010100",
  27663=>"110100100",
  27664=>"111100000",
  27665=>"110110101",
  27666=>"010110000",
  27667=>"100011111",
  27668=>"010100011",
  27669=>"011110001",
  27670=>"011011011",
  27671=>"100101111",
  27672=>"101000010",
  27673=>"110110100",
  27674=>"110000011",
  27675=>"101100101",
  27676=>"101101001",
  27677=>"001011011",
  27678=>"100000101",
  27679=>"010101100",
  27680=>"011011011",
  27681=>"101101100",
  27682=>"111110011",
  27683=>"001101010",
  27684=>"001101110",
  27685=>"111100011",
  27686=>"111011101",
  27687=>"111110101",
  27688=>"000010111",
  27689=>"110101101",
  27690=>"011100110",
  27691=>"111011101",
  27692=>"110010000",
  27693=>"010110111",
  27694=>"100001010",
  27695=>"011000111",
  27696=>"001010001",
  27697=>"101011110",
  27698=>"001111000",
  27699=>"000100011",
  27700=>"000010010",
  27701=>"010011000",
  27702=>"100100011",
  27703=>"000010101",
  27704=>"001100110",
  27705=>"010011010",
  27706=>"100110100",
  27707=>"111111101",
  27708=>"110100011",
  27709=>"010000101",
  27710=>"110011100",
  27711=>"011011111",
  27712=>"011011000",
  27713=>"100000111",
  27714=>"111000010",
  27715=>"000110110",
  27716=>"110110010",
  27717=>"001100101",
  27718=>"000001100",
  27719=>"000000110",
  27720=>"111000100",
  27721=>"011111010",
  27722=>"100011001",
  27723=>"101001101",
  27724=>"101001101",
  27725=>"111100001",
  27726=>"101110110",
  27727=>"010010011",
  27728=>"110000101",
  27729=>"111100101",
  27730=>"111111001",
  27731=>"101011000",
  27732=>"110111100",
  27733=>"011000000",
  27734=>"000001001",
  27735=>"000000000",
  27736=>"110000011",
  27737=>"110111010",
  27738=>"111101111",
  27739=>"000010110",
  27740=>"011001001",
  27741=>"100100010",
  27742=>"111010000",
  27743=>"001110111",
  27744=>"001010100",
  27745=>"100110100",
  27746=>"000010110",
  27747=>"110011100",
  27748=>"001111011",
  27749=>"011011001",
  27750=>"100101000",
  27751=>"111010110",
  27752=>"011110100",
  27753=>"111000000",
  27754=>"001101100",
  27755=>"111101101",
  27756=>"001110000",
  27757=>"101101001",
  27758=>"110001101",
  27759=>"111110110",
  27760=>"010001000",
  27761=>"000001000",
  27762=>"110100100",
  27763=>"101011111",
  27764=>"000000100",
  27765=>"110110001",
  27766=>"110110001",
  27767=>"111011001",
  27768=>"010100101",
  27769=>"001101001",
  27770=>"110101011",
  27771=>"100110101",
  27772=>"001100101",
  27773=>"111101111",
  27774=>"110011011",
  27775=>"110010010",
  27776=>"110100100",
  27777=>"000000001",
  27778=>"010101101",
  27779=>"011010001",
  27780=>"010001001",
  27781=>"010111011",
  27782=>"000101000",
  27783=>"001111011",
  27784=>"110001001",
  27785=>"100000001",
  27786=>"000100001",
  27787=>"100010001",
  27788=>"011011000",
  27789=>"111011111",
  27790=>"110101111",
  27791=>"110001001",
  27792=>"100010100",
  27793=>"011000111",
  27794=>"101000000",
  27795=>"111100110",
  27796=>"100000110",
  27797=>"010000110",
  27798=>"000101100",
  27799=>"001100100",
  27800=>"100101110",
  27801=>"011111110",
  27802=>"100100010",
  27803=>"111001001",
  27804=>"100111001",
  27805=>"001101101",
  27806=>"111011110",
  27807=>"100111101",
  27808=>"110110001",
  27809=>"011011101",
  27810=>"111111110",
  27811=>"010011011",
  27812=>"100110110",
  27813=>"011011101",
  27814=>"101101001",
  27815=>"010111000",
  27816=>"100101011",
  27817=>"100110010",
  27818=>"101110100",
  27819=>"001111111",
  27820=>"100001101",
  27821=>"100110101",
  27822=>"011010100",
  27823=>"101000100",
  27824=>"010100000",
  27825=>"100110111",
  27826=>"110101011",
  27827=>"100100001",
  27828=>"100110101",
  27829=>"111110100",
  27830=>"001001110",
  27831=>"000111011",
  27832=>"100111110",
  27833=>"101010100",
  27834=>"000100000",
  27835=>"110111100",
  27836=>"100011110",
  27837=>"111000111",
  27838=>"100000111",
  27839=>"000100100",
  27840=>"001111001",
  27841=>"100100100",
  27842=>"010110100",
  27843=>"010000000",
  27844=>"110101000",
  27845=>"100000110",
  27846=>"110000001",
  27847=>"100110111",
  27848=>"111111011",
  27849=>"001001111",
  27850=>"101111111",
  27851=>"001101101",
  27852=>"100001011",
  27853=>"100101100",
  27854=>"100100100",
  27855=>"000111100",
  27856=>"111110100",
  27857=>"011111100",
  27858=>"000100101",
  27859=>"110111110",
  27860=>"000000010",
  27861=>"110010101",
  27862=>"100100110",
  27863=>"101001010",
  27864=>"110011100",
  27865=>"111001110",
  27866=>"010000111",
  27867=>"111111100",
  27868=>"111011101",
  27869=>"011010111",
  27870=>"111001000",
  27871=>"111001000",
  27872=>"101100001",
  27873=>"101110100",
  27874=>"111000001",
  27875=>"110100110",
  27876=>"111001001",
  27877=>"101010101",
  27878=>"000100100",
  27879=>"110010011",
  27880=>"001101111",
  27881=>"000111001",
  27882=>"100010001",
  27883=>"101100000",
  27884=>"111010010",
  27885=>"110110000",
  27886=>"100011001",
  27887=>"001101111",
  27888=>"010010000",
  27889=>"100001111",
  27890=>"100100101",
  27891=>"010100101",
  27892=>"010010011",
  27893=>"001101101",
  27894=>"011011100",
  27895=>"100100010",
  27896=>"010110110",
  27897=>"100011110",
  27898=>"000100011",
  27899=>"111111111",
  27900=>"110011001",
  27901=>"010110110",
  27902=>"111110000",
  27903=>"110110001",
  27904=>"001111111",
  27905=>"110010001",
  27906=>"000001001",
  27907=>"001000000",
  27908=>"101101100",
  27909=>"101111000",
  27910=>"101001100",
  27911=>"011010110",
  27912=>"010011001",
  27913=>"111000100",
  27914=>"101000010",
  27915=>"011010101",
  27916=>"000101001",
  27917=>"000010000",
  27918=>"001100011",
  27919=>"101111100",
  27920=>"010010000",
  27921=>"100100001",
  27922=>"110001110",
  27923=>"101110010",
  27924=>"111001001",
  27925=>"101010010",
  27926=>"011111011",
  27927=>"000111110",
  27928=>"000010010",
  27929=>"110110001",
  27930=>"101011010",
  27931=>"100110110",
  27932=>"001011111",
  27933=>"101110110",
  27934=>"001110010",
  27935=>"010001010",
  27936=>"100010100",
  27937=>"100000000",
  27938=>"000010110",
  27939=>"100011010",
  27940=>"101101110",
  27941=>"010011000",
  27942=>"000110100",
  27943=>"000010001",
  27944=>"000001111",
  27945=>"111101011",
  27946=>"001000001",
  27947=>"100011101",
  27948=>"010010111",
  27949=>"101100010",
  27950=>"010001101",
  27951=>"001011100",
  27952=>"111010100",
  27953=>"111010000",
  27954=>"011010100",
  27955=>"110100111",
  27956=>"101100100",
  27957=>"100010110",
  27958=>"110001011",
  27959=>"011001011",
  27960=>"101101000",
  27961=>"000001001",
  27962=>"111110111",
  27963=>"110000010",
  27964=>"100100111",
  27965=>"110111110",
  27966=>"101110111",
  27967=>"011001000",
  27968=>"001101011",
  27969=>"011111110",
  27970=>"101011111",
  27971=>"100100110",
  27972=>"110000101",
  27973=>"011000000",
  27974=>"000010010",
  27975=>"110100111",
  27976=>"100110100",
  27977=>"001101001",
  27978=>"001000101",
  27979=>"110010100",
  27980=>"110100100",
  27981=>"000001001",
  27982=>"110110101",
  27983=>"010100000",
  27984=>"001011000",
  27985=>"000100011",
  27986=>"001011010",
  27987=>"000111011",
  27988=>"001000110",
  27989=>"000111111",
  27990=>"000111110",
  27991=>"000101010",
  27992=>"010010011",
  27993=>"001010011",
  27994=>"111011111",
  27995=>"011010110",
  27996=>"111000001",
  27997=>"110110011",
  27998=>"111110010",
  27999=>"001011111",
  28000=>"110101110",
  28001=>"010101000",
  28002=>"110110100",
  28003=>"001110000",
  28004=>"001000100",
  28005=>"110010011",
  28006=>"001100000",
  28007=>"111111101",
  28008=>"000011110",
  28009=>"101100100",
  28010=>"001100010",
  28011=>"111001011",
  28012=>"000100101",
  28013=>"110001001",
  28014=>"110100110",
  28015=>"001000101",
  28016=>"001001111",
  28017=>"010100001",
  28018=>"101000111",
  28019=>"000110110",
  28020=>"101001100",
  28021=>"001101101",
  28022=>"100101110",
  28023=>"001010000",
  28024=>"010111110",
  28025=>"010010001",
  28026=>"010010001",
  28027=>"101101001",
  28028=>"011000000",
  28029=>"111110101",
  28030=>"101110100",
  28031=>"100001101",
  28032=>"010110101",
  28033=>"110010100",
  28034=>"100010010",
  28035=>"010000011",
  28036=>"000011010",
  28037=>"110100001",
  28038=>"011101001",
  28039=>"011110110",
  28040=>"111011000",
  28041=>"111101101",
  28042=>"001000101",
  28043=>"001001001",
  28044=>"110110100",
  28045=>"111001000",
  28046=>"111010111",
  28047=>"101011000",
  28048=>"011001001",
  28049=>"101110110",
  28050=>"110000011",
  28051=>"011101011",
  28052=>"101000001",
  28053=>"111111110",
  28054=>"110111110",
  28055=>"111001010",
  28056=>"000011000",
  28057=>"011001101",
  28058=>"100111111",
  28059=>"100010000",
  28060=>"101100111",
  28061=>"100110101",
  28062=>"110111001",
  28063=>"011100001",
  28064=>"111101111",
  28065=>"111010110",
  28066=>"101000000",
  28067=>"000110001",
  28068=>"111110000",
  28069=>"011111000",
  28070=>"100001001",
  28071=>"100001011",
  28072=>"011001010",
  28073=>"000110011",
  28074=>"000100011",
  28075=>"001101011",
  28076=>"111111101",
  28077=>"001100000",
  28078=>"100110101",
  28079=>"110001011",
  28080=>"100100001",
  28081=>"100101110",
  28082=>"101010001",
  28083=>"000001011",
  28084=>"011000010",
  28085=>"001101101",
  28086=>"011110101",
  28087=>"100110110",
  28088=>"101110100",
  28089=>"101010001",
  28090=>"110011000",
  28091=>"100010110",
  28092=>"011100011",
  28093=>"010011011",
  28094=>"000100001",
  28095=>"101100110",
  28096=>"111001000",
  28097=>"011100101",
  28098=>"001010110",
  28099=>"100100010",
  28100=>"110110111",
  28101=>"111100101",
  28102=>"110001000",
  28103=>"111001101",
  28104=>"011101001",
  28105=>"101100111",
  28106=>"110010010",
  28107=>"000100001",
  28108=>"110010100",
  28109=>"100100100",
  28110=>"011000100",
  28111=>"001101000",
  28112=>"001001101",
  28113=>"000000011",
  28114=>"000100000",
  28115=>"001010000",
  28116=>"101001010",
  28117=>"101100111",
  28118=>"001100110",
  28119=>"111111100",
  28120=>"010000000",
  28121=>"101110000",
  28122=>"100111010",
  28123=>"111101100",
  28124=>"111001010",
  28125=>"110100100",
  28126=>"101111011",
  28127=>"011111110",
  28128=>"101111100",
  28129=>"010010010",
  28130=>"110110000",
  28131=>"101000001",
  28132=>"101001110",
  28133=>"100001111",
  28134=>"000110100",
  28135=>"101100100",
  28136=>"011000001",
  28137=>"111101101",
  28138=>"001111010",
  28139=>"100011010",
  28140=>"101010110",
  28141=>"010000100",
  28142=>"110110010",
  28143=>"010000100",
  28144=>"110101011",
  28145=>"101101100",
  28146=>"110001101",
  28147=>"100000001",
  28148=>"100100111",
  28149=>"000101110",
  28150=>"001011110",
  28151=>"100011010",
  28152=>"100111010",
  28153=>"111011101",
  28154=>"101111001",
  28155=>"101100101",
  28156=>"111100010",
  28157=>"010000110",
  28158=>"110101100",
  28159=>"111001010",
  28160=>"000001101",
  28161=>"000101101",
  28162=>"110001110",
  28163=>"000110000",
  28164=>"011100110",
  28165=>"111001100",
  28166=>"111100000",
  28167=>"000110100",
  28168=>"001110000",
  28169=>"011000101",
  28170=>"000001100",
  28171=>"000000001",
  28172=>"111111001",
  28173=>"111001000",
  28174=>"010000110",
  28175=>"101101101",
  28176=>"011001011",
  28177=>"000000111",
  28178=>"000001101",
  28179=>"100111010",
  28180=>"101100011",
  28181=>"011010101",
  28182=>"011110100",
  28183=>"111101100",
  28184=>"101100110",
  28185=>"000000101",
  28186=>"000111010",
  28187=>"001000000",
  28188=>"111100100",
  28189=>"001001100",
  28190=>"111000111",
  28191=>"011100111",
  28192=>"100001110",
  28193=>"110101000",
  28194=>"111001001",
  28195=>"010100100",
  28196=>"110101001",
  28197=>"010010111",
  28198=>"011100101",
  28199=>"010110111",
  28200=>"111110111",
  28201=>"010110100",
  28202=>"001000100",
  28203=>"111110001",
  28204=>"011011110",
  28205=>"101011110",
  28206=>"110111111",
  28207=>"101101101",
  28208=>"100110111",
  28209=>"111111000",
  28210=>"110010010",
  28211=>"110000110",
  28212=>"100101001",
  28213=>"001011101",
  28214=>"011001111",
  28215=>"011000100",
  28216=>"110011001",
  28217=>"100100101",
  28218=>"001111000",
  28219=>"011111001",
  28220=>"100001001",
  28221=>"000001111",
  28222=>"001101001",
  28223=>"101001101",
  28224=>"111111100",
  28225=>"110000011",
  28226=>"000110001",
  28227=>"000111001",
  28228=>"001001010",
  28229=>"110000010",
  28230=>"100100100",
  28231=>"101101110",
  28232=>"000010010",
  28233=>"100100000",
  28234=>"100110001",
  28235=>"101101111",
  28236=>"101010010",
  28237=>"101110100",
  28238=>"110111110",
  28239=>"101011001",
  28240=>"001110100",
  28241=>"111101000",
  28242=>"100000100",
  28243=>"111011000",
  28244=>"100010111",
  28245=>"010110011",
  28246=>"010111001",
  28247=>"011110110",
  28248=>"001001011",
  28249=>"001100110",
  28250=>"001000010",
  28251=>"010011011",
  28252=>"111001010",
  28253=>"110000101",
  28254=>"100100111",
  28255=>"111101000",
  28256=>"010001001",
  28257=>"100110011",
  28258=>"111100010",
  28259=>"000001110",
  28260=>"011001011",
  28261=>"100111100",
  28262=>"000000111",
  28263=>"100111010",
  28264=>"000000011",
  28265=>"111110001",
  28266=>"010001010",
  28267=>"110110100",
  28268=>"010000001",
  28269=>"001001001",
  28270=>"011110100",
  28271=>"000010010",
  28272=>"100111011",
  28273=>"001100010",
  28274=>"101010010",
  28275=>"100000011",
  28276=>"101101010",
  28277=>"000100010",
  28278=>"100111101",
  28279=>"100100010",
  28280=>"010001001",
  28281=>"110100100",
  28282=>"010111100",
  28283=>"001111000",
  28284=>"111000010",
  28285=>"010010111",
  28286=>"101100100",
  28287=>"100011111",
  28288=>"101010100",
  28289=>"101110011",
  28290=>"110100110",
  28291=>"001010000",
  28292=>"100000010",
  28293=>"000111000",
  28294=>"111101011",
  28295=>"111111010",
  28296=>"010100011",
  28297=>"010110001",
  28298=>"011111010",
  28299=>"011010000",
  28300=>"000000111",
  28301=>"101111101",
  28302=>"111101001",
  28303=>"110110111",
  28304=>"111001000",
  28305=>"000110100",
  28306=>"000100101",
  28307=>"111010100",
  28308=>"011111100",
  28309=>"010001011",
  28310=>"010000111",
  28311=>"001000110",
  28312=>"011101010",
  28313=>"100101110",
  28314=>"111010011",
  28315=>"111101111",
  28316=>"000000111",
  28317=>"100101110",
  28318=>"110011101",
  28319=>"111010100",
  28320=>"101100110",
  28321=>"001100001",
  28322=>"100100101",
  28323=>"110011011",
  28324=>"101100100",
  28325=>"000000101",
  28326=>"100110110",
  28327=>"101100101",
  28328=>"110001000",
  28329=>"110000100",
  28330=>"101000001",
  28331=>"000100100",
  28332=>"011111010",
  28333=>"100011110",
  28334=>"010010000",
  28335=>"001110001",
  28336=>"000101000",
  28337=>"100001111",
  28338=>"011100011",
  28339=>"100111100",
  28340=>"001101111",
  28341=>"000100110",
  28342=>"010001001",
  28343=>"001010100",
  28344=>"110000110",
  28345=>"111011011",
  28346=>"100001010",
  28347=>"000100110",
  28348=>"101101100",
  28349=>"000000110",
  28350=>"111100111",
  28351=>"111111110",
  28352=>"000110111",
  28353=>"001001011",
  28354=>"000100100",
  28355=>"001001100",
  28356=>"000001001",
  28357=>"110111110",
  28358=>"100111001",
  28359=>"010100110",
  28360=>"111110111",
  28361=>"000010101",
  28362=>"011011011",
  28363=>"001001010",
  28364=>"000010011",
  28365=>"110011110",
  28366=>"100000001",
  28367=>"110101100",
  28368=>"000111000",
  28369=>"101111101",
  28370=>"101000010",
  28371=>"010111111",
  28372=>"011101001",
  28373=>"110001001",
  28374=>"111100110",
  28375=>"101111101",
  28376=>"110000101",
  28377=>"000001011",
  28378=>"110111110",
  28379=>"000000001",
  28380=>"001010000",
  28381=>"100111000",
  28382=>"111001011",
  28383=>"000000011",
  28384=>"111100101",
  28385=>"011011110",
  28386=>"101111100",
  28387=>"001110100",
  28388=>"101110000",
  28389=>"011001001",
  28390=>"100000110",
  28391=>"010001110",
  28392=>"000000110",
  28393=>"101100101",
  28394=>"000001000",
  28395=>"100001100",
  28396=>"000000100",
  28397=>"010100111",
  28398=>"110011101",
  28399=>"101101100",
  28400=>"110110000",
  28401=>"100010101",
  28402=>"010000111",
  28403=>"101101001",
  28404=>"001110101",
  28405=>"011101001",
  28406=>"100011011",
  28407=>"111100100",
  28408=>"000000001",
  28409=>"100110100",
  28410=>"001001010",
  28411=>"000010110",
  28412=>"000101110",
  28413=>"110101110",
  28414=>"110100101",
  28415=>"101100010",
  28416=>"010011100",
  28417=>"101111101",
  28418=>"000110101",
  28419=>"101110101",
  28420=>"100001011",
  28421=>"110110011",
  28422=>"101001101",
  28423=>"101101000",
  28424=>"100001101",
  28425=>"100111001",
  28426=>"010010111",
  28427=>"011001111",
  28428=>"110010000",
  28429=>"110111001",
  28430=>"011000111",
  28431=>"111100001",
  28432=>"110110010",
  28433=>"110101100",
  28434=>"000111000",
  28435=>"111111111",
  28436=>"110111001",
  28437=>"110111010",
  28438=>"101100011",
  28439=>"000100101",
  28440=>"010000000",
  28441=>"001010110",
  28442=>"000011100",
  28443=>"100111001",
  28444=>"010000010",
  28445=>"101010011",
  28446=>"111000111",
  28447=>"011011000",
  28448=>"011110111",
  28449=>"001001001",
  28450=>"000111101",
  28451=>"110100011",
  28452=>"100111101",
  28453=>"111111010",
  28454=>"001111000",
  28455=>"010001110",
  28456=>"101010001",
  28457=>"100001000",
  28458=>"110111110",
  28459=>"010110100",
  28460=>"001000001",
  28461=>"100001001",
  28462=>"101100100",
  28463=>"110110101",
  28464=>"000100010",
  28465=>"000111111",
  28466=>"000011001",
  28467=>"001001111",
  28468=>"001000110",
  28469=>"011010000",
  28470=>"100111011",
  28471=>"011011011",
  28472=>"101100100",
  28473=>"010110101",
  28474=>"001101010",
  28475=>"101010110",
  28476=>"011011100",
  28477=>"100100101",
  28478=>"001000000",
  28479=>"100001011",
  28480=>"101000001",
  28481=>"111100010",
  28482=>"100101100",
  28483=>"111011100",
  28484=>"110100001",
  28485=>"010011101",
  28486=>"100111010",
  28487=>"011010100",
  28488=>"100000011",
  28489=>"010010000",
  28490=>"101001110",
  28491=>"000111100",
  28492=>"111001000",
  28493=>"100101100",
  28494=>"001111111",
  28495=>"001101111",
  28496=>"100110111",
  28497=>"011111000",
  28498=>"110101111",
  28499=>"000010011",
  28500=>"000111000",
  28501=>"001001111",
  28502=>"001100001",
  28503=>"001110011",
  28504=>"101101110",
  28505=>"011011010",
  28506=>"001010110",
  28507=>"001100110",
  28508=>"101100000",
  28509=>"011000001",
  28510=>"111110110",
  28511=>"101000100",
  28512=>"111010100",
  28513=>"111100100",
  28514=>"101000001",
  28515=>"001110000",
  28516=>"110111110",
  28517=>"111010001",
  28518=>"111010001",
  28519=>"001101111",
  28520=>"100110000",
  28521=>"101010001",
  28522=>"000011001",
  28523=>"100100100",
  28524=>"100000100",
  28525=>"000000000",
  28526=>"110101110",
  28527=>"010001001",
  28528=>"011000000",
  28529=>"011111011",
  28530=>"101010011",
  28531=>"101000101",
  28532=>"100010000",
  28533=>"111110111",
  28534=>"011100001",
  28535=>"110101101",
  28536=>"110101100",
  28537=>"110111100",
  28538=>"110111101",
  28539=>"000000011",
  28540=>"000100100",
  28541=>"110110001",
  28542=>"110101110",
  28543=>"111111101",
  28544=>"101010000",
  28545=>"101101011",
  28546=>"001000111",
  28547=>"011111101",
  28548=>"100000111",
  28549=>"000100001",
  28550=>"110000110",
  28551=>"111011100",
  28552=>"110000010",
  28553=>"100010110",
  28554=>"010001101",
  28555=>"101110101",
  28556=>"111010011",
  28557=>"111010001",
  28558=>"010011001",
  28559=>"111111100",
  28560=>"110001111",
  28561=>"001111010",
  28562=>"110110110",
  28563=>"010101110",
  28564=>"100000001",
  28565=>"001110111",
  28566=>"000110100",
  28567=>"100011000",
  28568=>"111001111",
  28569=>"110101111",
  28570=>"110000010",
  28571=>"110000111",
  28572=>"011111001",
  28573=>"011000000",
  28574=>"111111110",
  28575=>"011011101",
  28576=>"111110010",
  28577=>"000010000",
  28578=>"000011010",
  28579=>"111000011",
  28580=>"101001001",
  28581=>"010111100",
  28582=>"001011101",
  28583=>"000100111",
  28584=>"010001111",
  28585=>"001001111",
  28586=>"010111110",
  28587=>"011101111",
  28588=>"101100011",
  28589=>"011011000",
  28590=>"100101111",
  28591=>"110111110",
  28592=>"101000010",
  28593=>"111011011",
  28594=>"111111011",
  28595=>"101111000",
  28596=>"111111011",
  28597=>"000000011",
  28598=>"001011011",
  28599=>"100001101",
  28600=>"111011011",
  28601=>"011001111",
  28602=>"110001111",
  28603=>"001110001",
  28604=>"010010000",
  28605=>"101011100",
  28606=>"101010010",
  28607=>"100101110",
  28608=>"001001010",
  28609=>"011000010",
  28610=>"011000000",
  28611=>"011100110",
  28612=>"010011001",
  28613=>"100101100",
  28614=>"110000100",
  28615=>"011000100",
  28616=>"000010001",
  28617=>"100100101",
  28618=>"011001110",
  28619=>"111101010",
  28620=>"111110000",
  28621=>"101100100",
  28622=>"010011111",
  28623=>"010111001",
  28624=>"001111110",
  28625=>"001100111",
  28626=>"011111010",
  28627=>"011000110",
  28628=>"110100010",
  28629=>"100011001",
  28630=>"110100101",
  28631=>"001011011",
  28632=>"111100011",
  28633=>"110101101",
  28634=>"001100010",
  28635=>"111001011",
  28636=>"110010010",
  28637=>"010110111",
  28638=>"111101100",
  28639=>"011101101",
  28640=>"010011000",
  28641=>"000101001",
  28642=>"001001001",
  28643=>"110100100",
  28644=>"100010110",
  28645=>"110100101",
  28646=>"110101100",
  28647=>"110001001",
  28648=>"110100000",
  28649=>"011000111",
  28650=>"011100010",
  28651=>"110100101",
  28652=>"111001001",
  28653=>"101011010",
  28654=>"101111010",
  28655=>"011110000",
  28656=>"001001111",
  28657=>"111110101",
  28658=>"001011100",
  28659=>"110100001",
  28660=>"001111111",
  28661=>"000110110",
  28662=>"010000110",
  28663=>"111111011",
  28664=>"001000101",
  28665=>"011010000",
  28666=>"110001111",
  28667=>"110010110",
  28668=>"110110100",
  28669=>"010001100",
  28670=>"001011100",
  28671=>"000001111",
  28672=>"001000001",
  28673=>"010011010",
  28674=>"101011001",
  28675=>"001000101",
  28676=>"001000101",
  28677=>"010100010",
  28678=>"011001101",
  28679=>"011101010",
  28680=>"111010010",
  28681=>"111011001",
  28682=>"110001110",
  28683=>"100101000",
  28684=>"010110110",
  28685=>"110010100",
  28686=>"001110110",
  28687=>"001111010",
  28688=>"010000000",
  28689=>"000101011",
  28690=>"110100101",
  28691=>"001001110",
  28692=>"000100000",
  28693=>"100001000",
  28694=>"110010001",
  28695=>"111001100",
  28696=>"000101111",
  28697=>"011000010",
  28698=>"110111000",
  28699=>"011100110",
  28700=>"001010001",
  28701=>"111110100",
  28702=>"010100100",
  28703=>"101000111",
  28704=>"011110000",
  28705=>"111001001",
  28706=>"110000011",
  28707=>"000101110",
  28708=>"111111011",
  28709=>"101010001",
  28710=>"100000000",
  28711=>"100000000",
  28712=>"000000110",
  28713=>"100011110",
  28714=>"010011101",
  28715=>"000011100",
  28716=>"010110001",
  28717=>"101111110",
  28718=>"011010000",
  28719=>"010100100",
  28720=>"111101100",
  28721=>"001100110",
  28722=>"011111011",
  28723=>"000101110",
  28724=>"000010011",
  28725=>"001110000",
  28726=>"111000110",
  28727=>"111101010",
  28728=>"111000000",
  28729=>"011010001",
  28730=>"010110100",
  28731=>"111101100",
  28732=>"110010101",
  28733=>"110010101",
  28734=>"110101100",
  28735=>"000100100",
  28736=>"010010001",
  28737=>"000000001",
  28738=>"110100011",
  28739=>"110111001",
  28740=>"000011011",
  28741=>"111011011",
  28742=>"111011000",
  28743=>"111011110",
  28744=>"001111010",
  28745=>"001111000",
  28746=>"110011000",
  28747=>"010011001",
  28748=>"110111111",
  28749=>"001101101",
  28750=>"111110001",
  28751=>"100010110",
  28752=>"110000010",
  28753=>"101010100",
  28754=>"100100010",
  28755=>"110101111",
  28756=>"000011001",
  28757=>"110111101",
  28758=>"011000111",
  28759=>"110111100",
  28760=>"011000111",
  28761=>"010111001",
  28762=>"110011101",
  28763=>"000001111",
  28764=>"100100100",
  28765=>"011101001",
  28766=>"001010010",
  28767=>"100000011",
  28768=>"111010010",
  28769=>"111101001",
  28770=>"000001000",
  28771=>"101100000",
  28772=>"011101000",
  28773=>"110011110",
  28774=>"000101010",
  28775=>"101111010",
  28776=>"000010101",
  28777=>"111101011",
  28778=>"001011000",
  28779=>"000001111",
  28780=>"000110010",
  28781=>"010100010",
  28782=>"001001000",
  28783=>"001110000",
  28784=>"010000100",
  28785=>"010000000",
  28786=>"111000011",
  28787=>"111110011",
  28788=>"000110111",
  28789=>"111011001",
  28790=>"100111101",
  28791=>"010111010",
  28792=>"100000100",
  28793=>"010000011",
  28794=>"010000110",
  28795=>"101111010",
  28796=>"010001000",
  28797=>"111001111",
  28798=>"000011110",
  28799=>"100111000",
  28800=>"001000011",
  28801=>"110111000",
  28802=>"111010011",
  28803=>"001001111",
  28804=>"000101011",
  28805=>"111111111",
  28806=>"110101101",
  28807=>"001101001",
  28808=>"100000011",
  28809=>"101001111",
  28810=>"000000100",
  28811=>"100001111",
  28812=>"011010110",
  28813=>"000110111",
  28814=>"110000110",
  28815=>"100101001",
  28816=>"100001001",
  28817=>"111110001",
  28818=>"100010011",
  28819=>"000100000",
  28820=>"010000010",
  28821=>"000101001",
  28822=>"000101001",
  28823=>"000011110",
  28824=>"001010100",
  28825=>"000111011",
  28826=>"111101111",
  28827=>"111111100",
  28828=>"001010110",
  28829=>"001001011",
  28830=>"010100000",
  28831=>"101101111",
  28832=>"110100101",
  28833=>"000000100",
  28834=>"101100100",
  28835=>"010111011",
  28836=>"100011110",
  28837=>"110001001",
  28838=>"011101100",
  28839=>"101000111",
  28840=>"000100000",
  28841=>"111110000",
  28842=>"000011000",
  28843=>"101010100",
  28844=>"111000110",
  28845=>"011101011",
  28846=>"110000001",
  28847=>"000111101",
  28848=>"110110010",
  28849=>"111011111",
  28850=>"110101010",
  28851=>"100110000",
  28852=>"101100011",
  28853=>"010100000",
  28854=>"111001100",
  28855=>"001010000",
  28856=>"110011110",
  28857=>"100100011",
  28858=>"001110110",
  28859=>"101010110",
  28860=>"000110110",
  28861=>"101000001",
  28862=>"111111010",
  28863=>"110100100",
  28864=>"011101110",
  28865=>"000100100",
  28866=>"000001000",
  28867=>"101111000",
  28868=>"001000000",
  28869=>"011110111",
  28870=>"100111110",
  28871=>"001001000",
  28872=>"110100111",
  28873=>"011110010",
  28874=>"101001110",
  28875=>"110110100",
  28876=>"000000101",
  28877=>"000010010",
  28878=>"000000011",
  28879=>"110110000",
  28880=>"011101100",
  28881=>"010111010",
  28882=>"000101001",
  28883=>"001101011",
  28884=>"010001100",
  28885=>"100101100",
  28886=>"110010011",
  28887=>"001000001",
  28888=>"011111000",
  28889=>"001110100",
  28890=>"010111010",
  28891=>"100110001",
  28892=>"011100001",
  28893=>"100010001",
  28894=>"111010001",
  28895=>"011101111",
  28896=>"000001000",
  28897=>"010010011",
  28898=>"011101101",
  28899=>"110101100",
  28900=>"000010101",
  28901=>"101111111",
  28902=>"001111001",
  28903=>"010011000",
  28904=>"010111011",
  28905=>"101000010",
  28906=>"000100101",
  28907=>"110000111",
  28908=>"000110001",
  28909=>"101111000",
  28910=>"011010001",
  28911=>"000011100",
  28912=>"010010101",
  28913=>"100101011",
  28914=>"001010100",
  28915=>"000101101",
  28916=>"001110000",
  28917=>"011101101",
  28918=>"011101110",
  28919=>"010010010",
  28920=>"011111011",
  28921=>"110110000",
  28922=>"010011111",
  28923=>"010111001",
  28924=>"010011000",
  28925=>"000100111",
  28926=>"100010000",
  28927=>"011000100",
  28928=>"000011101",
  28929=>"011101011",
  28930=>"111101011",
  28931=>"011000111",
  28932=>"001001100",
  28933=>"011111100",
  28934=>"000000010",
  28935=>"011010010",
  28936=>"101001110",
  28937=>"010001000",
  28938=>"000111010",
  28939=>"000001101",
  28940=>"001110001",
  28941=>"001110101",
  28942=>"000111110",
  28943=>"111000001",
  28944=>"000010100",
  28945=>"001011000",
  28946=>"000111100",
  28947=>"100100111",
  28948=>"001110011",
  28949=>"001010101",
  28950=>"001011010",
  28951=>"000011001",
  28952=>"010100100",
  28953=>"101111101",
  28954=>"010001010",
  28955=>"101000001",
  28956=>"100001110",
  28957=>"101011100",
  28958=>"001011000",
  28959=>"000111011",
  28960=>"001110110",
  28961=>"000010000",
  28962=>"100001100",
  28963=>"100000001",
  28964=>"011010001",
  28965=>"101100000",
  28966=>"011100100",
  28967=>"100110101",
  28968=>"110100100",
  28969=>"100001011",
  28970=>"010101000",
  28971=>"011110101",
  28972=>"011110101",
  28973=>"101110100",
  28974=>"100000000",
  28975=>"100000010",
  28976=>"010001110",
  28977=>"010000011",
  28978=>"111101010",
  28979=>"111100000",
  28980=>"100101011",
  28981=>"101011111",
  28982=>"100100110",
  28983=>"001110111",
  28984=>"010001110",
  28985=>"001100000",
  28986=>"001101101",
  28987=>"111000111",
  28988=>"010011111",
  28989=>"111100110",
  28990=>"110000101",
  28991=>"110001101",
  28992=>"000000011",
  28993=>"011000110",
  28994=>"111111101",
  28995=>"111010110",
  28996=>"010111001",
  28997=>"010010100",
  28998=>"000010111",
  28999=>"011011001",
  29000=>"010010100",
  29001=>"110010011",
  29002=>"001000010",
  29003=>"001110011",
  29004=>"011001100",
  29005=>"111110101",
  29006=>"000100001",
  29007=>"101111010",
  29008=>"001000000",
  29009=>"011001100",
  29010=>"100001010",
  29011=>"000111001",
  29012=>"110110111",
  29013=>"000010000",
  29014=>"110010011",
  29015=>"100111100",
  29016=>"101001111",
  29017=>"101010000",
  29018=>"111110101",
  29019=>"000100001",
  29020=>"001101101",
  29021=>"011010001",
  29022=>"000100000",
  29023=>"001010010",
  29024=>"101111011",
  29025=>"010010111",
  29026=>"100011101",
  29027=>"100001110",
  29028=>"000010000",
  29029=>"110110110",
  29030=>"011110011",
  29031=>"101111010",
  29032=>"110111100",
  29033=>"011010110",
  29034=>"101110111",
  29035=>"010110101",
  29036=>"110111101",
  29037=>"011111001",
  29038=>"011001010",
  29039=>"100100101",
  29040=>"000001001",
  29041=>"101001001",
  29042=>"011000000",
  29043=>"110000110",
  29044=>"010011111",
  29045=>"111100001",
  29046=>"000101000",
  29047=>"000110001",
  29048=>"011111101",
  29049=>"010011011",
  29050=>"010101100",
  29051=>"101101100",
  29052=>"100111100",
  29053=>"111011111",
  29054=>"000100110",
  29055=>"001000111",
  29056=>"000000010",
  29057=>"111000000",
  29058=>"010011001",
  29059=>"001001010",
  29060=>"100101011",
  29061=>"000101010",
  29062=>"110101110",
  29063=>"100111110",
  29064=>"101111110",
  29065=>"011111011",
  29066=>"000101011",
  29067=>"110111101",
  29068=>"010000111",
  29069=>"001010000",
  29070=>"010000101",
  29071=>"011111111",
  29072=>"000101110",
  29073=>"100001110",
  29074=>"110101011",
  29075=>"100011111",
  29076=>"000000100",
  29077=>"110110000",
  29078=>"011101010",
  29079=>"100101011",
  29080=>"111001101",
  29081=>"101111101",
  29082=>"010110111",
  29083=>"110001010",
  29084=>"011100010",
  29085=>"100110001",
  29086=>"110011100",
  29087=>"111110000",
  29088=>"010010000",
  29089=>"010100011",
  29090=>"100111111",
  29091=>"010101110",
  29092=>"111101101",
  29093=>"000111011",
  29094=>"111100110",
  29095=>"110010110",
  29096=>"001001101",
  29097=>"111001111",
  29098=>"100001001",
  29099=>"000110001",
  29100=>"110101111",
  29101=>"010111011",
  29102=>"101110111",
  29103=>"001000010",
  29104=>"101000011",
  29105=>"001111110",
  29106=>"110010001",
  29107=>"100100001",
  29108=>"011010100",
  29109=>"100011001",
  29110=>"101010010",
  29111=>"110010111",
  29112=>"010000000",
  29113=>"010110000",
  29114=>"010001110",
  29115=>"111101101",
  29116=>"110111000",
  29117=>"111111000",
  29118=>"101010001",
  29119=>"000101100",
  29120=>"101000001",
  29121=>"110010110",
  29122=>"101010110",
  29123=>"010110000",
  29124=>"000000101",
  29125=>"101011001",
  29126=>"010100110",
  29127=>"000010110",
  29128=>"001101110",
  29129=>"011101011",
  29130=>"000001010",
  29131=>"100001100",
  29132=>"101011001",
  29133=>"101010001",
  29134=>"000001010",
  29135=>"101000010",
  29136=>"111101011",
  29137=>"001000000",
  29138=>"010010000",
  29139=>"100111010",
  29140=>"000111111",
  29141=>"001100100",
  29142=>"000100110",
  29143=>"011000001",
  29144=>"111101110",
  29145=>"100011001",
  29146=>"101001011",
  29147=>"001011001",
  29148=>"101100001",
  29149=>"010110111",
  29150=>"011111101",
  29151=>"111011101",
  29152=>"010010010",
  29153=>"101101001",
  29154=>"111011110",
  29155=>"111110010",
  29156=>"000101111",
  29157=>"000110111",
  29158=>"010011100",
  29159=>"111010000",
  29160=>"110111110",
  29161=>"000110111",
  29162=>"000100101",
  29163=>"000101101",
  29164=>"001111100",
  29165=>"111011110",
  29166=>"100101101",
  29167=>"110101010",
  29168=>"011000111",
  29169=>"111110001",
  29170=>"101101111",
  29171=>"100000111",
  29172=>"101100111",
  29173=>"101110110",
  29174=>"000001101",
  29175=>"001101100",
  29176=>"110000010",
  29177=>"001101100",
  29178=>"000001100",
  29179=>"110101111",
  29180=>"010000111",
  29181=>"110100010",
  29182=>"000011011",
  29183=>"100100000",
  29184=>"100110100",
  29185=>"011110110",
  29186=>"101100111",
  29187=>"000110011",
  29188=>"010101101",
  29189=>"110111001",
  29190=>"001100000",
  29191=>"001010001",
  29192=>"011111101",
  29193=>"000011110",
  29194=>"100101111",
  29195=>"011110100",
  29196=>"001010100",
  29197=>"100110111",
  29198=>"011111110",
  29199=>"001000001",
  29200=>"000011001",
  29201=>"101110111",
  29202=>"101001110",
  29203=>"110110000",
  29204=>"110100001",
  29205=>"001011110",
  29206=>"111111101",
  29207=>"111111101",
  29208=>"101111100",
  29209=>"010011001",
  29210=>"100001010",
  29211=>"110011110",
  29212=>"100100101",
  29213=>"001001000",
  29214=>"010001011",
  29215=>"100010000",
  29216=>"101000001",
  29217=>"010111110",
  29218=>"100001000",
  29219=>"111011110",
  29220=>"011111000",
  29221=>"100010101",
  29222=>"001100100",
  29223=>"100110000",
  29224=>"110111011",
  29225=>"111110110",
  29226=>"111101110",
  29227=>"001010111",
  29228=>"001110111",
  29229=>"101000110",
  29230=>"110110010",
  29231=>"110110011",
  29232=>"001011001",
  29233=>"001110100",
  29234=>"000111111",
  29235=>"000010100",
  29236=>"101111000",
  29237=>"001000100",
  29238=>"101010011",
  29239=>"101000111",
  29240=>"001110101",
  29241=>"111100100",
  29242=>"110101011",
  29243=>"101011000",
  29244=>"010010001",
  29245=>"000100110",
  29246=>"000010011",
  29247=>"111101000",
  29248=>"111110000",
  29249=>"011101111",
  29250=>"010100001",
  29251=>"010101100",
  29252=>"100110111",
  29253=>"100001100",
  29254=>"010110111",
  29255=>"001110001",
  29256=>"000111111",
  29257=>"111111101",
  29258=>"100010011",
  29259=>"010001010",
  29260=>"110011010",
  29261=>"100001011",
  29262=>"101100010",
  29263=>"110101011",
  29264=>"110111100",
  29265=>"011011000",
  29266=>"001110011",
  29267=>"100110110",
  29268=>"100010001",
  29269=>"001011001",
  29270=>"011011111",
  29271=>"000101011",
  29272=>"001100111",
  29273=>"010000010",
  29274=>"111110000",
  29275=>"100011010",
  29276=>"001001110",
  29277=>"111000100",
  29278=>"000101011",
  29279=>"111100100",
  29280=>"111110110",
  29281=>"010011111",
  29282=>"101101001",
  29283=>"011101000",
  29284=>"110111011",
  29285=>"001001111",
  29286=>"011101110",
  29287=>"110010010",
  29288=>"011000100",
  29289=>"101001000",
  29290=>"100110011",
  29291=>"101100101",
  29292=>"001001010",
  29293=>"010010111",
  29294=>"111101010",
  29295=>"000110101",
  29296=>"000000110",
  29297=>"100100010",
  29298=>"001001000",
  29299=>"111100011",
  29300=>"111110101",
  29301=>"100010111",
  29302=>"100001110",
  29303=>"000110101",
  29304=>"110001010",
  29305=>"010111010",
  29306=>"011011000",
  29307=>"111101110",
  29308=>"000101000",
  29309=>"110110111",
  29310=>"100000011",
  29311=>"110011010",
  29312=>"011110111",
  29313=>"011001110",
  29314=>"011010100",
  29315=>"100000101",
  29316=>"001001010",
  29317=>"011001111",
  29318=>"000101100",
  29319=>"001001011",
  29320=>"000000101",
  29321=>"000101011",
  29322=>"110000111",
  29323=>"001011111",
  29324=>"100000011",
  29325=>"000010010",
  29326=>"010010011",
  29327=>"000100110",
  29328=>"000100100",
  29329=>"101011110",
  29330=>"100101001",
  29331=>"001111101",
  29332=>"110111111",
  29333=>"001111100",
  29334=>"101111000",
  29335=>"001001000",
  29336=>"100111000",
  29337=>"001010000",
  29338=>"111000000",
  29339=>"011101100",
  29340=>"111110100",
  29341=>"001100000",
  29342=>"110000011",
  29343=>"010001001",
  29344=>"010010101",
  29345=>"011111011",
  29346=>"111110101",
  29347=>"111101111",
  29348=>"010111110",
  29349=>"011101110",
  29350=>"010011100",
  29351=>"101010100",
  29352=>"011010110",
  29353=>"000010111",
  29354=>"101100010",
  29355=>"100100011",
  29356=>"111110000",
  29357=>"010001100",
  29358=>"011110000",
  29359=>"011001100",
  29360=>"000010111",
  29361=>"010101110",
  29362=>"100001000",
  29363=>"010111010",
  29364=>"111000111",
  29365=>"111001001",
  29366=>"000000111",
  29367=>"101010100",
  29368=>"010101001",
  29369=>"110011101",
  29370=>"011000011",
  29371=>"000110000",
  29372=>"101010100",
  29373=>"010001010",
  29374=>"010001100",
  29375=>"100110110",
  29376=>"000010000",
  29377=>"010111100",
  29378=>"100101110",
  29379=>"010010100",
  29380=>"111010010",
  29381=>"110111111",
  29382=>"001100110",
  29383=>"000100111",
  29384=>"000000100",
  29385=>"101111110",
  29386=>"110011110",
  29387=>"000111010",
  29388=>"111111010",
  29389=>"001000100",
  29390=>"101011010",
  29391=>"010001110",
  29392=>"001101111",
  29393=>"000010000",
  29394=>"101001010",
  29395=>"001000110",
  29396=>"111110011",
  29397=>"010000111",
  29398=>"000101110",
  29399=>"001100100",
  29400=>"100101110",
  29401=>"011101000",
  29402=>"101110100",
  29403=>"011001000",
  29404=>"001100000",
  29405=>"101011110",
  29406=>"001111110",
  29407=>"101101010",
  29408=>"110110010",
  29409=>"011111000",
  29410=>"101010110",
  29411=>"010001100",
  29412=>"110100011",
  29413=>"000110110",
  29414=>"111001010",
  29415=>"100100100",
  29416=>"000000010",
  29417=>"100001101",
  29418=>"111101011",
  29419=>"110111111",
  29420=>"001010010",
  29421=>"110101000",
  29422=>"110101001",
  29423=>"100100100",
  29424=>"111100011",
  29425=>"000110111",
  29426=>"010011110",
  29427=>"000001110",
  29428=>"011010000",
  29429=>"001111101",
  29430=>"110111110",
  29431=>"111100101",
  29432=>"010000000",
  29433=>"110010101",
  29434=>"001111101",
  29435=>"110011100",
  29436=>"010001101",
  29437=>"110110110",
  29438=>"000010001",
  29439=>"011011001",
  29440=>"011010000",
  29441=>"001000111",
  29442=>"000110111",
  29443=>"000110111",
  29444=>"000011000",
  29445=>"001000101",
  29446=>"111101111",
  29447=>"111111101",
  29448=>"011000010",
  29449=>"100010100",
  29450=>"110011000",
  29451=>"010100100",
  29452=>"101001011",
  29453=>"101111100",
  29454=>"001101001",
  29455=>"010110011",
  29456=>"001101111",
  29457=>"111110111",
  29458=>"011101010",
  29459=>"100111001",
  29460=>"001000101",
  29461=>"010111110",
  29462=>"001111010",
  29463=>"101100001",
  29464=>"010110010",
  29465=>"011000110",
  29466=>"001111000",
  29467=>"101101100",
  29468=>"111000001",
  29469=>"001000010",
  29470=>"000000010",
  29471=>"011010010",
  29472=>"111100000",
  29473=>"110100110",
  29474=>"110110001",
  29475=>"111110100",
  29476=>"111001011",
  29477=>"111001000",
  29478=>"000001100",
  29479=>"111010011",
  29480=>"000010111",
  29481=>"001100100",
  29482=>"101001010",
  29483=>"110010111",
  29484=>"011111110",
  29485=>"010110001",
  29486=>"101101100",
  29487=>"000000111",
  29488=>"111010000",
  29489=>"110111101",
  29490=>"100001111",
  29491=>"100100100",
  29492=>"011100101",
  29493=>"101110101",
  29494=>"000111100",
  29495=>"010100011",
  29496=>"110000010",
  29497=>"111000100",
  29498=>"111111011",
  29499=>"110110110",
  29500=>"000010001",
  29501=>"011110000",
  29502=>"011110010",
  29503=>"001110001",
  29504=>"000100001",
  29505=>"100101101",
  29506=>"100111100",
  29507=>"010111010",
  29508=>"001101000",
  29509=>"001100001",
  29510=>"100001101",
  29511=>"101000010",
  29512=>"110011000",
  29513=>"000000111",
  29514=>"111111001",
  29515=>"001101110",
  29516=>"010011100",
  29517=>"111111110",
  29518=>"000000101",
  29519=>"000011101",
  29520=>"111100101",
  29521=>"011101001",
  29522=>"111111100",
  29523=>"100010101",
  29524=>"000010000",
  29525=>"110111001",
  29526=>"010100010",
  29527=>"111001000",
  29528=>"110111111",
  29529=>"101111111",
  29530=>"100110100",
  29531=>"101010001",
  29532=>"111101111",
  29533=>"111100011",
  29534=>"010000100",
  29535=>"000110011",
  29536=>"101111111",
  29537=>"111010100",
  29538=>"010010110",
  29539=>"101001011",
  29540=>"100010000",
  29541=>"100000110",
  29542=>"111100000",
  29543=>"101000100",
  29544=>"111000001",
  29545=>"010011011",
  29546=>"010101000",
  29547=>"100100001",
  29548=>"110000011",
  29549=>"010100110",
  29550=>"100110111",
  29551=>"010100110",
  29552=>"111101111",
  29553=>"011001101",
  29554=>"011101001",
  29555=>"011011011",
  29556=>"110110001",
  29557=>"110010110",
  29558=>"110000000",
  29559=>"011000111",
  29560=>"001011111",
  29561=>"010000111",
  29562=>"111100011",
  29563=>"110010010",
  29564=>"000110101",
  29565=>"011001010",
  29566=>"100111000",
  29567=>"010111110",
  29568=>"000011010",
  29569=>"101010001",
  29570=>"100011011",
  29571=>"000000111",
  29572=>"001001011",
  29573=>"010001000",
  29574=>"010110101",
  29575=>"010001010",
  29576=>"111100101",
  29577=>"010100100",
  29578=>"001100010",
  29579=>"010110011",
  29580=>"110100110",
  29581=>"010101010",
  29582=>"101001111",
  29583=>"110001111",
  29584=>"111101011",
  29585=>"101111101",
  29586=>"010000110",
  29587=>"000011000",
  29588=>"011000001",
  29589=>"011111011",
  29590=>"011000011",
  29591=>"000010001",
  29592=>"001101100",
  29593=>"000001000",
  29594=>"011010000",
  29595=>"000011111",
  29596=>"110111111",
  29597=>"101100100",
  29598=>"011010111",
  29599=>"011010010",
  29600=>"000000110",
  29601=>"011010001",
  29602=>"001000010",
  29603=>"111010010",
  29604=>"110110001",
  29605=>"100110001",
  29606=>"000100111",
  29607=>"101011110",
  29608=>"000011001",
  29609=>"011001100",
  29610=>"100101101",
  29611=>"010010100",
  29612=>"100000001",
  29613=>"001100111",
  29614=>"101000010",
  29615=>"100001110",
  29616=>"010000111",
  29617=>"111001100",
  29618=>"111100011",
  29619=>"010010101",
  29620=>"110110010",
  29621=>"111011001",
  29622=>"110010110",
  29623=>"010111100",
  29624=>"010110111",
  29625=>"000011100",
  29626=>"111011001",
  29627=>"100001001",
  29628=>"111000110",
  29629=>"000111111",
  29630=>"001110000",
  29631=>"001111010",
  29632=>"011110111",
  29633=>"000000110",
  29634=>"100100011",
  29635=>"110000110",
  29636=>"100000100",
  29637=>"110110110",
  29638=>"111111110",
  29639=>"000111011",
  29640=>"111101101",
  29641=>"100001100",
  29642=>"100101110",
  29643=>"001010001",
  29644=>"001101000",
  29645=>"001110011",
  29646=>"010000000",
  29647=>"111010000",
  29648=>"011011001",
  29649=>"011110110",
  29650=>"001011010",
  29651=>"000100011",
  29652=>"000011101",
  29653=>"011101000",
  29654=>"111110111",
  29655=>"101001111",
  29656=>"001001111",
  29657=>"000001001",
  29658=>"010001110",
  29659=>"101000010",
  29660=>"100101111",
  29661=>"110101010",
  29662=>"101000101",
  29663=>"011101000",
  29664=>"100101110",
  29665=>"110111111",
  29666=>"110111010",
  29667=>"101001001",
  29668=>"010010110",
  29669=>"000000111",
  29670=>"100011100",
  29671=>"110010001",
  29672=>"100011000",
  29673=>"010010110",
  29674=>"110100100",
  29675=>"100000101",
  29676=>"110000011",
  29677=>"101101010",
  29678=>"010001101",
  29679=>"100111001",
  29680=>"000111101",
  29681=>"111110001",
  29682=>"000101111",
  29683=>"111011111",
  29684=>"000010110",
  29685=>"110010111",
  29686=>"110001110",
  29687=>"101000000",
  29688=>"111011111",
  29689=>"110000000",
  29690=>"001011010",
  29691=>"101111100",
  29692=>"110100111",
  29693=>"010010000",
  29694=>"000000000",
  29695=>"110011001",
  29696=>"101011111",
  29697=>"101100010",
  29698=>"001101100",
  29699=>"101111010",
  29700=>"000010011",
  29701=>"010001011",
  29702=>"011010000",
  29703=>"100000010",
  29704=>"000111110",
  29705=>"000100010",
  29706=>"111010001",
  29707=>"101111110",
  29708=>"100001010",
  29709=>"001001001",
  29710=>"000011100",
  29711=>"100100001",
  29712=>"110101001",
  29713=>"011110001",
  29714=>"010110010",
  29715=>"000100010",
  29716=>"101110000",
  29717=>"100110001",
  29718=>"001010111",
  29719=>"000111000",
  29720=>"111000001",
  29721=>"100001001",
  29722=>"000110000",
  29723=>"101011111",
  29724=>"001111001",
  29725=>"101010101",
  29726=>"000010010",
  29727=>"010110010",
  29728=>"110001110",
  29729=>"000100010",
  29730=>"000011000",
  29731=>"111100101",
  29732=>"100101000",
  29733=>"000101100",
  29734=>"010101011",
  29735=>"010000011",
  29736=>"011001110",
  29737=>"011001111",
  29738=>"101010110",
  29739=>"100010010",
  29740=>"010011111",
  29741=>"100010001",
  29742=>"111010000",
  29743=>"000010011",
  29744=>"111101100",
  29745=>"011010011",
  29746=>"011110001",
  29747=>"001000101",
  29748=>"011101111",
  29749=>"110110001",
  29750=>"100111010",
  29751=>"000110100",
  29752=>"001100000",
  29753=>"000001011",
  29754=>"111100001",
  29755=>"010000111",
  29756=>"101100011",
  29757=>"001111111",
  29758=>"110000000",
  29759=>"100101011",
  29760=>"100001101",
  29761=>"000000111",
  29762=>"000100111",
  29763=>"100011001",
  29764=>"001110001",
  29765=>"110001011",
  29766=>"110001101",
  29767=>"001000011",
  29768=>"000011011",
  29769=>"111101111",
  29770=>"000100111",
  29771=>"110111000",
  29772=>"000001101",
  29773=>"011011110",
  29774=>"111110100",
  29775=>"111111000",
  29776=>"100001010",
  29777=>"100101110",
  29778=>"000011111",
  29779=>"101111010",
  29780=>"100010101",
  29781=>"000000100",
  29782=>"110011000",
  29783=>"001100101",
  29784=>"110000010",
  29785=>"110011111",
  29786=>"001100111",
  29787=>"111011010",
  29788=>"101101010",
  29789=>"100000010",
  29790=>"111001101",
  29791=>"110111101",
  29792=>"100100111",
  29793=>"111110100",
  29794=>"001000101",
  29795=>"001010010",
  29796=>"111000100",
  29797=>"101111100",
  29798=>"010000101",
  29799=>"001000001",
  29800=>"111101001",
  29801=>"001111111",
  29802=>"010001010",
  29803=>"000000111",
  29804=>"100010001",
  29805=>"100111111",
  29806=>"101011111",
  29807=>"111000111",
  29808=>"110110000",
  29809=>"000100001",
  29810=>"011100111",
  29811=>"101000110",
  29812=>"010001111",
  29813=>"100101000",
  29814=>"110011101",
  29815=>"001001111",
  29816=>"000101111",
  29817=>"110001010",
  29818=>"011101110",
  29819=>"001100000",
  29820=>"101111100",
  29821=>"111010100",
  29822=>"111000111",
  29823=>"000000010",
  29824=>"010001100",
  29825=>"001001001",
  29826=>"101101010",
  29827=>"111000011",
  29828=>"011001010",
  29829=>"100000001",
  29830=>"000000100",
  29831=>"010111101",
  29832=>"001100111",
  29833=>"000111010",
  29834=>"110010010",
  29835=>"100111111",
  29836=>"010011111",
  29837=>"110111001",
  29838=>"011111100",
  29839=>"001101010",
  29840=>"111001001",
  29841=>"111101010",
  29842=>"101111110",
  29843=>"111110101",
  29844=>"000000000",
  29845=>"001000001",
  29846=>"010000110",
  29847=>"010101010",
  29848=>"101000010",
  29849=>"001000101",
  29850=>"101110111",
  29851=>"110111010",
  29852=>"111001110",
  29853=>"010101011",
  29854=>"000001010",
  29855=>"000000010",
  29856=>"100101001",
  29857=>"100111110",
  29858=>"101001000",
  29859=>"100000101",
  29860=>"101100110",
  29861=>"101100101",
  29862=>"011110111",
  29863=>"001010110",
  29864=>"010001001",
  29865=>"000110110",
  29866=>"101011011",
  29867=>"010111110",
  29868=>"100101100",
  29869=>"111100111",
  29870=>"111100001",
  29871=>"101011110",
  29872=>"000011000",
  29873=>"000011110",
  29874=>"111111111",
  29875=>"000100110",
  29876=>"110000011",
  29877=>"001000001",
  29878=>"110001011",
  29879=>"011011000",
  29880=>"001000011",
  29881=>"001011000",
  29882=>"110110001",
  29883=>"011000111",
  29884=>"110101110",
  29885=>"011000000",
  29886=>"011010010",
  29887=>"000101011",
  29888=>"101010110",
  29889=>"010101111",
  29890=>"101010000",
  29891=>"010110111",
  29892=>"111001011",
  29893=>"000111100",
  29894=>"011111111",
  29895=>"000010110",
  29896=>"001110101",
  29897=>"100101110",
  29898=>"001011010",
  29899=>"000101010",
  29900=>"010000000",
  29901=>"011000001",
  29902=>"111001010",
  29903=>"101101010",
  29904=>"100011000",
  29905=>"001011101",
  29906=>"111001001",
  29907=>"001011010",
  29908=>"010001001",
  29909=>"000110111",
  29910=>"001000111",
  29911=>"111001110",
  29912=>"101101100",
  29913=>"110111010",
  29914=>"011001011",
  29915=>"101111001",
  29916=>"011111000",
  29917=>"110000011",
  29918=>"100101000",
  29919=>"011100110",
  29920=>"000000100",
  29921=>"101001101",
  29922=>"010110010",
  29923=>"100100010",
  29924=>"001100000",
  29925=>"001111000",
  29926=>"101010100",
  29927=>"000111001",
  29928=>"110001110",
  29929=>"001111101",
  29930=>"000011011",
  29931=>"001111100",
  29932=>"001000000",
  29933=>"110101101",
  29934=>"110001000",
  29935=>"001011000",
  29936=>"000101110",
  29937=>"111110111",
  29938=>"111000101",
  29939=>"000010001",
  29940=>"001010101",
  29941=>"001111001",
  29942=>"010010100",
  29943=>"010010100",
  29944=>"001110100",
  29945=>"010001001",
  29946=>"001100000",
  29947=>"110000111",
  29948=>"010000000",
  29949=>"001111110",
  29950=>"010110110",
  29951=>"111110110",
  29952=>"110001011",
  29953=>"010010111",
  29954=>"000111100",
  29955=>"100100000",
  29956=>"010111001",
  29957=>"011101001",
  29958=>"110011111",
  29959=>"111011110",
  29960=>"010000111",
  29961=>"110111100",
  29962=>"011111111",
  29963=>"011110100",
  29964=>"110101101",
  29965=>"000001101",
  29966=>"011011001",
  29967=>"111110111",
  29968=>"100100101",
  29969=>"110001101",
  29970=>"110100100",
  29971=>"101100110",
  29972=>"100100111",
  29973=>"101100111",
  29974=>"011001110",
  29975=>"011000100",
  29976=>"111010100",
  29977=>"101101000",
  29978=>"001010001",
  29979=>"001101100",
  29980=>"111011010",
  29981=>"111100000",
  29982=>"000000001",
  29983=>"110001001",
  29984=>"010010000",
  29985=>"101101101",
  29986=>"111111111",
  29987=>"000000011",
  29988=>"100101110",
  29989=>"011000011",
  29990=>"000001000",
  29991=>"111000100",
  29992=>"010001100",
  29993=>"011101010",
  29994=>"010000011",
  29995=>"001001011",
  29996=>"010011000",
  29997=>"111111011",
  29998=>"001000110",
  29999=>"000011111",
  30000=>"001010000",
  30001=>"010000000",
  30002=>"110111010",
  30003=>"100010101",
  30004=>"010111100",
  30005=>"100001100",
  30006=>"010001110",
  30007=>"101110000",
  30008=>"101100111",
  30009=>"000001110",
  30010=>"111111100",
  30011=>"010101000",
  30012=>"010000101",
  30013=>"111000001",
  30014=>"010100110",
  30015=>"101111000",
  30016=>"101110010",
  30017=>"111000100",
  30018=>"110010100",
  30019=>"101101011",
  30020=>"101011100",
  30021=>"110000001",
  30022=>"100010101",
  30023=>"101011111",
  30024=>"001100001",
  30025=>"010001001",
  30026=>"101101001",
  30027=>"111001111",
  30028=>"011001101",
  30029=>"010011101",
  30030=>"010101001",
  30031=>"101000000",
  30032=>"111100001",
  30033=>"110110010",
  30034=>"011001100",
  30035=>"010101001",
  30036=>"000001001",
  30037=>"011110001",
  30038=>"011010101",
  30039=>"011111101",
  30040=>"100100010",
  30041=>"000000110",
  30042=>"001110000",
  30043=>"000100111",
  30044=>"101100011",
  30045=>"000110011",
  30046=>"110110011",
  30047=>"010001001",
  30048=>"010110111",
  30049=>"011110000",
  30050=>"000011000",
  30051=>"000110010",
  30052=>"111001110",
  30053=>"101011011",
  30054=>"000101001",
  30055=>"011110000",
  30056=>"110110011",
  30057=>"011100011",
  30058=>"111000000",
  30059=>"010110001",
  30060=>"100000001",
  30061=>"111011011",
  30062=>"001011110",
  30063=>"110111001",
  30064=>"101010101",
  30065=>"001010100",
  30066=>"011011100",
  30067=>"111010010",
  30068=>"010101011",
  30069=>"101001111",
  30070=>"000000100",
  30071=>"000010111",
  30072=>"000001001",
  30073=>"010111011",
  30074=>"000101010",
  30075=>"100111101",
  30076=>"101001111",
  30077=>"101100101",
  30078=>"100101011",
  30079=>"111111010",
  30080=>"011010010",
  30081=>"111100011",
  30082=>"100111000",
  30083=>"001111001",
  30084=>"010101101",
  30085=>"111001011",
  30086=>"011000111",
  30087=>"110010010",
  30088=>"001000001",
  30089=>"010000100",
  30090=>"100011001",
  30091=>"011000010",
  30092=>"111011111",
  30093=>"000000100",
  30094=>"100110111",
  30095=>"011100101",
  30096=>"011010011",
  30097=>"101100011",
  30098=>"000100000",
  30099=>"110000100",
  30100=>"001010100",
  30101=>"000110011",
  30102=>"000010100",
  30103=>"001000001",
  30104=>"111010011",
  30105=>"000001111",
  30106=>"111111000",
  30107=>"111101000",
  30108=>"010001110",
  30109=>"110101001",
  30110=>"011011101",
  30111=>"100110010",
  30112=>"010010101",
  30113=>"011110100",
  30114=>"010101000",
  30115=>"000000100",
  30116=>"110001010",
  30117=>"011010111",
  30118=>"111100111",
  30119=>"011101111",
  30120=>"111010101",
  30121=>"110000001",
  30122=>"000111101",
  30123=>"100000011",
  30124=>"000000110",
  30125=>"011111110",
  30126=>"011101010",
  30127=>"001010111",
  30128=>"010111111",
  30129=>"100000100",
  30130=>"111101010",
  30131=>"100111011",
  30132=>"001111000",
  30133=>"011100010",
  30134=>"101001010",
  30135=>"101110110",
  30136=>"100011100",
  30137=>"111110110",
  30138=>"111110010",
  30139=>"001101100",
  30140=>"101100101",
  30141=>"101011111",
  30142=>"010001001",
  30143=>"011111011",
  30144=>"110110001",
  30145=>"001011010",
  30146=>"100100111",
  30147=>"011010011",
  30148=>"010000101",
  30149=>"001011001",
  30150=>"001000000",
  30151=>"011011011",
  30152=>"110110000",
  30153=>"011000110",
  30154=>"011000000",
  30155=>"000101011",
  30156=>"010011110",
  30157=>"101011001",
  30158=>"110001011",
  30159=>"001010010",
  30160=>"010011111",
  30161=>"001011001",
  30162=>"001011101",
  30163=>"011111111",
  30164=>"010110100",
  30165=>"100101101",
  30166=>"001000000",
  30167=>"000001101",
  30168=>"101010011",
  30169=>"101110000",
  30170=>"000010001",
  30171=>"010000000",
  30172=>"010111100",
  30173=>"111110001",
  30174=>"001010000",
  30175=>"000110001",
  30176=>"010011011",
  30177=>"001000000",
  30178=>"110110011",
  30179=>"010000011",
  30180=>"100011111",
  30181=>"010011101",
  30182=>"000000011",
  30183=>"001001000",
  30184=>"000010100",
  30185=>"010001101",
  30186=>"001101110",
  30187=>"001100101",
  30188=>"110001110",
  30189=>"100000101",
  30190=>"110000110",
  30191=>"001001010",
  30192=>"001011000",
  30193=>"000000000",
  30194=>"010100001",
  30195=>"100110010",
  30196=>"011101011",
  30197=>"011101101",
  30198=>"010110011",
  30199=>"100110101",
  30200=>"011000010",
  30201=>"011001001",
  30202=>"001011111",
  30203=>"000010010",
  30204=>"110101101",
  30205=>"001110001",
  30206=>"011001000",
  30207=>"000000110",
  30208=>"000001001",
  30209=>"011011011",
  30210=>"100111101",
  30211=>"011000011",
  30212=>"110101110",
  30213=>"110111111",
  30214=>"011011000",
  30215=>"101001010",
  30216=>"111100111",
  30217=>"111000000",
  30218=>"010000001",
  30219=>"011010101",
  30220=>"000110100",
  30221=>"101000011",
  30222=>"100010111",
  30223=>"010111010",
  30224=>"101101100",
  30225=>"011111100",
  30226=>"001100000",
  30227=>"111000100",
  30228=>"111011000",
  30229=>"100100101",
  30230=>"011000011",
  30231=>"101101100",
  30232=>"011000001",
  30233=>"110001001",
  30234=>"101001011",
  30235=>"001100010",
  30236=>"101011001",
  30237=>"000010111",
  30238=>"010001010",
  30239=>"101011101",
  30240=>"011011011",
  30241=>"100110100",
  30242=>"101100100",
  30243=>"100010001",
  30244=>"011000011",
  30245=>"011100101",
  30246=>"110110000",
  30247=>"001110010",
  30248=>"000001001",
  30249=>"110000001",
  30250=>"111011110",
  30251=>"111001010",
  30252=>"110101110",
  30253=>"100000010",
  30254=>"000000100",
  30255=>"111001100",
  30256=>"011111100",
  30257=>"100001000",
  30258=>"001100100",
  30259=>"010000011",
  30260=>"010100000",
  30261=>"011011101",
  30262=>"110011000",
  30263=>"100110111",
  30264=>"011110011",
  30265=>"100011011",
  30266=>"110100011",
  30267=>"010110001",
  30268=>"100110110",
  30269=>"110001101",
  30270=>"100111111",
  30271=>"001100010",
  30272=>"001101110",
  30273=>"100001111",
  30274=>"111011011",
  30275=>"011101000",
  30276=>"001011100",
  30277=>"011001101",
  30278=>"110100111",
  30279=>"001000001",
  30280=>"111100101",
  30281=>"000111011",
  30282=>"011001001",
  30283=>"010011001",
  30284=>"101111111",
  30285=>"010010111",
  30286=>"010001111",
  30287=>"010111100",
  30288=>"101011110",
  30289=>"011101011",
  30290=>"110011010",
  30291=>"111101100",
  30292=>"010100000",
  30293=>"001111001",
  30294=>"110000000",
  30295=>"101011111",
  30296=>"101011101",
  30297=>"100101010",
  30298=>"101011101",
  30299=>"000000000",
  30300=>"001100010",
  30301=>"100010100",
  30302=>"000010100",
  30303=>"000011111",
  30304=>"111001000",
  30305=>"001111001",
  30306=>"011000101",
  30307=>"100101010",
  30308=>"110111001",
  30309=>"101011101",
  30310=>"101110000",
  30311=>"000001110",
  30312=>"101011100",
  30313=>"010110110",
  30314=>"010111100",
  30315=>"110010010",
  30316=>"000010110",
  30317=>"111101000",
  30318=>"001000101",
  30319=>"011010101",
  30320=>"110001000",
  30321=>"111111101",
  30322=>"100001011",
  30323=>"000100110",
  30324=>"111000101",
  30325=>"010000011",
  30326=>"000101010",
  30327=>"011110011",
  30328=>"010000001",
  30329=>"000010111",
  30330=>"101101100",
  30331=>"010000100",
  30332=>"111000010",
  30333=>"110100011",
  30334=>"011100001",
  30335=>"010110000",
  30336=>"100101001",
  30337=>"011111111",
  30338=>"011001011",
  30339=>"001111111",
  30340=>"010001011",
  30341=>"000000100",
  30342=>"110001010",
  30343=>"110000110",
  30344=>"110101101",
  30345=>"101010100",
  30346=>"110111100",
  30347=>"011110101",
  30348=>"101111001",
  30349=>"010101111",
  30350=>"011111011",
  30351=>"101011011",
  30352=>"010000010",
  30353=>"100111111",
  30354=>"010110100",
  30355=>"101111111",
  30356=>"101000010",
  30357=>"001101000",
  30358=>"100101111",
  30359=>"010110010",
  30360=>"100100001",
  30361=>"100110000",
  30362=>"110101010",
  30363=>"001110100",
  30364=>"011101101",
  30365=>"010110100",
  30366=>"000100100",
  30367=>"111111010",
  30368=>"011111000",
  30369=>"000010001",
  30370=>"101111111",
  30371=>"001100000",
  30372=>"001001111",
  30373=>"100110110",
  30374=>"111111010",
  30375=>"000011110",
  30376=>"100000000",
  30377=>"111000110",
  30378=>"010100111",
  30379=>"100111011",
  30380=>"000101111",
  30381=>"110000010",
  30382=>"010000000",
  30383=>"011011001",
  30384=>"001101101",
  30385=>"001111100",
  30386=>"010010111",
  30387=>"110111111",
  30388=>"000001101",
  30389=>"001000011",
  30390=>"010010000",
  30391=>"011111000",
  30392=>"001111000",
  30393=>"101111010",
  30394=>"010111110",
  30395=>"010110110",
  30396=>"000110101",
  30397=>"000001100",
  30398=>"010100011",
  30399=>"101101011",
  30400=>"010000010",
  30401=>"001110100",
  30402=>"100101101",
  30403=>"001010000",
  30404=>"111110111",
  30405=>"101100101",
  30406=>"101010001",
  30407=>"100001000",
  30408=>"011111110",
  30409=>"010101101",
  30410=>"111100100",
  30411=>"010110011",
  30412=>"000000101",
  30413=>"101010011",
  30414=>"111111011",
  30415=>"010111100",
  30416=>"101111011",
  30417=>"000111101",
  30418=>"110100000",
  30419=>"110100011",
  30420=>"101001000",
  30421=>"001111010",
  30422=>"010000101",
  30423=>"001001100",
  30424=>"011101100",
  30425=>"110110001",
  30426=>"111000000",
  30427=>"111000101",
  30428=>"100110011",
  30429=>"100110000",
  30430=>"000000110",
  30431=>"111110100",
  30432=>"111100001",
  30433=>"000001100",
  30434=>"111011100",
  30435=>"100110110",
  30436=>"111110000",
  30437=>"010010010",
  30438=>"110000100",
  30439=>"100101101",
  30440=>"001001110",
  30441=>"101100001",
  30442=>"110111111",
  30443=>"101010111",
  30444=>"101111111",
  30445=>"110000001",
  30446=>"100011010",
  30447=>"011110001",
  30448=>"111111010",
  30449=>"001001010",
  30450=>"010010011",
  30451=>"011011100",
  30452=>"100110011",
  30453=>"100100000",
  30454=>"011111010",
  30455=>"011011001",
  30456=>"100101001",
  30457=>"001000000",
  30458=>"100011100",
  30459=>"111010110",
  30460=>"000001111",
  30461=>"010011000",
  30462=>"110001000",
  30463=>"000010111",
  30464=>"011011010",
  30465=>"110010100",
  30466=>"101101010",
  30467=>"101101100",
  30468=>"011101010",
  30469=>"011100100",
  30470=>"000010000",
  30471=>"101111100",
  30472=>"010001111",
  30473=>"100011000",
  30474=>"101001001",
  30475=>"100111010",
  30476=>"111110101",
  30477=>"011000010",
  30478=>"001101001",
  30479=>"001000110",
  30480=>"111101010",
  30481=>"010100100",
  30482=>"001000110",
  30483=>"001000101",
  30484=>"100110010",
  30485=>"101011110",
  30486=>"110111100",
  30487=>"010100000",
  30488=>"000000011",
  30489=>"000100100",
  30490=>"010001100",
  30491=>"101010101",
  30492=>"101110010",
  30493=>"100110101",
  30494=>"011111010",
  30495=>"010011001",
  30496=>"000001100",
  30497=>"101110010",
  30498=>"101011110",
  30499=>"110001111",
  30500=>"000101011",
  30501=>"110110100",
  30502=>"010000010",
  30503=>"010001010",
  30504=>"001101011",
  30505=>"101010011",
  30506=>"011110110",
  30507=>"001011001",
  30508=>"000100001",
  30509=>"111100011",
  30510=>"110111100",
  30511=>"100001000",
  30512=>"001000110",
  30513=>"000101011",
  30514=>"011000101",
  30515=>"111010111",
  30516=>"010111011",
  30517=>"101101011",
  30518=>"010000101",
  30519=>"001110100",
  30520=>"110010001",
  30521=>"001110010",
  30522=>"001010001",
  30523=>"100010101",
  30524=>"111110011",
  30525=>"010100011",
  30526=>"010001000",
  30527=>"101011011",
  30528=>"010000111",
  30529=>"010000100",
  30530=>"011111111",
  30531=>"001010011",
  30532=>"111111001",
  30533=>"010110101",
  30534=>"111101000",
  30535=>"011110110",
  30536=>"110101011",
  30537=>"011111100",
  30538=>"111010110",
  30539=>"001000111",
  30540=>"111010011",
  30541=>"100111011",
  30542=>"110110111",
  30543=>"110100010",
  30544=>"011010111",
  30545=>"101010111",
  30546=>"101101010",
  30547=>"111111011",
  30548=>"000010100",
  30549=>"011000000",
  30550=>"100110100",
  30551=>"000111010",
  30552=>"011100100",
  30553=>"101000011",
  30554=>"111111011",
  30555=>"110100010",
  30556=>"100001101",
  30557=>"110100000",
  30558=>"001111011",
  30559=>"001010010",
  30560=>"010110010",
  30561=>"000000000",
  30562=>"000010110",
  30563=>"100101010",
  30564=>"100100011",
  30565=>"100011001",
  30566=>"101111111",
  30567=>"111101010",
  30568=>"000010011",
  30569=>"100110010",
  30570=>"010001101",
  30571=>"101111110",
  30572=>"100111110",
  30573=>"000001100",
  30574=>"010100000",
  30575=>"011110010",
  30576=>"001001010",
  30577=>"010010111",
  30578=>"011011000",
  30579=>"011000101",
  30580=>"100100010",
  30581=>"000101101",
  30582=>"001101011",
  30583=>"011101000",
  30584=>"101110110",
  30585=>"100010001",
  30586=>"000101000",
  30587=>"010001000",
  30588=>"000110010",
  30589=>"110000101",
  30590=>"110010110",
  30591=>"101011010",
  30592=>"110111110",
  30593=>"010101010",
  30594=>"010100001",
  30595=>"101111101",
  30596=>"111101100",
  30597=>"100111101",
  30598=>"001001110",
  30599=>"011101100",
  30600=>"000110110",
  30601=>"010011011",
  30602=>"001101100",
  30603=>"100110100",
  30604=>"010001110",
  30605=>"100001000",
  30606=>"001011011",
  30607=>"011001001",
  30608=>"000111000",
  30609=>"110010111",
  30610=>"100001010",
  30611=>"100101000",
  30612=>"100001001",
  30613=>"100011001",
  30614=>"000011100",
  30615=>"110111010",
  30616=>"010111000",
  30617=>"110000110",
  30618=>"011000011",
  30619=>"000000100",
  30620=>"000111001",
  30621=>"010100000",
  30622=>"000000100",
  30623=>"011011011",
  30624=>"011000000",
  30625=>"001110100",
  30626=>"010111011",
  30627=>"010111000",
  30628=>"101011011",
  30629=>"001010101",
  30630=>"011100011",
  30631=>"101111011",
  30632=>"100001111",
  30633=>"000001011",
  30634=>"101101111",
  30635=>"100001001",
  30636=>"011100110",
  30637=>"101111101",
  30638=>"010110101",
  30639=>"010011110",
  30640=>"110000100",
  30641=>"010100111",
  30642=>"011011010",
  30643=>"000001000",
  30644=>"100101101",
  30645=>"111110110",
  30646=>"101000000",
  30647=>"001011110",
  30648=>"010010001",
  30649=>"111110100",
  30650=>"101111100",
  30651=>"110101000",
  30652=>"011010011",
  30653=>"000100001",
  30654=>"111001101",
  30655=>"010110011",
  30656=>"001100010",
  30657=>"010010011",
  30658=>"101010010",
  30659=>"000000011",
  30660=>"010101101",
  30661=>"000111101",
  30662=>"001111101",
  30663=>"001110100",
  30664=>"101101101",
  30665=>"111100011",
  30666=>"001010101",
  30667=>"001101010",
  30668=>"010110110",
  30669=>"111110111",
  30670=>"110011100",
  30671=>"100011001",
  30672=>"011011001",
  30673=>"010011110",
  30674=>"011100100",
  30675=>"111000010",
  30676=>"011010101",
  30677=>"111010101",
  30678=>"010001010",
  30679=>"000100110",
  30680=>"000110011",
  30681=>"111001011",
  30682=>"011001101",
  30683=>"111111011",
  30684=>"100000000",
  30685=>"010100000",
  30686=>"000000101",
  30687=>"110001101",
  30688=>"110100110",
  30689=>"111000100",
  30690=>"011110010",
  30691=>"101100010",
  30692=>"001001001",
  30693=>"010010001",
  30694=>"000001000",
  30695=>"001110100",
  30696=>"100001100",
  30697=>"010111110",
  30698=>"011000010",
  30699=>"010000101",
  30700=>"110001100",
  30701=>"011111001",
  30702=>"100100011",
  30703=>"011101011",
  30704=>"101011011",
  30705=>"111111010",
  30706=>"111001001",
  30707=>"100110101",
  30708=>"000110111",
  30709=>"101010000",
  30710=>"010110010",
  30711=>"100111100",
  30712=>"100010100",
  30713=>"111010010",
  30714=>"101111100",
  30715=>"111001010",
  30716=>"011111011",
  30717=>"100111010",
  30718=>"011100011",
  30719=>"011100110",
  30720=>"001011101",
  30721=>"011110000",
  30722=>"011111110",
  30723=>"010000110",
  30724=>"111100011",
  30725=>"110001000",
  30726=>"110110110",
  30727=>"001001111",
  30728=>"110100100",
  30729=>"101100101",
  30730=>"000100111",
  30731=>"011101010",
  30732=>"010111001",
  30733=>"010000111",
  30734=>"001001010",
  30735=>"111101000",
  30736=>"101101010",
  30737=>"111111001",
  30738=>"001001000",
  30739=>"110000001",
  30740=>"111100100",
  30741=>"001000001",
  30742=>"100101111",
  30743=>"001000100",
  30744=>"000110111",
  30745=>"000010011",
  30746=>"010100100",
  30747=>"011001010",
  30748=>"000100100",
  30749=>"010011000",
  30750=>"000011110",
  30751=>"101001000",
  30752=>"101010011",
  30753=>"100100101",
  30754=>"111000010",
  30755=>"001000101",
  30756=>"011000010",
  30757=>"111000010",
  30758=>"001101110",
  30759=>"110011010",
  30760=>"001100111",
  30761=>"000000001",
  30762=>"000000111",
  30763=>"111101010",
  30764=>"111011100",
  30765=>"100101111",
  30766=>"100110010",
  30767=>"101100100",
  30768=>"100110011",
  30769=>"100101010",
  30770=>"000110010",
  30771=>"011101101",
  30772=>"000000011",
  30773=>"001111111",
  30774=>"100010100",
  30775=>"001010011",
  30776=>"010000100",
  30777=>"000110010",
  30778=>"000111100",
  30779=>"101011011",
  30780=>"000010000",
  30781=>"010011111",
  30782=>"101100101",
  30783=>"111110110",
  30784=>"000001111",
  30785=>"011110100",
  30786=>"100010000",
  30787=>"111110001",
  30788=>"000110111",
  30789=>"100101010",
  30790=>"011010001",
  30791=>"001100000",
  30792=>"111010100",
  30793=>"011111011",
  30794=>"011001100",
  30795=>"001011000",
  30796=>"011000010",
  30797=>"101010111",
  30798=>"101010100",
  30799=>"101101011",
  30800=>"011011010",
  30801=>"011010011",
  30802=>"011100001",
  30803=>"000110101",
  30804=>"100110101",
  30805=>"001000001",
  30806=>"001000001",
  30807=>"110111111",
  30808=>"101011000",
  30809=>"101011110",
  30810=>"000000001",
  30811=>"010000011",
  30812=>"111000000",
  30813=>"001011010",
  30814=>"001000011",
  30815=>"011111110",
  30816=>"111100101",
  30817=>"000110001",
  30818=>"100100001",
  30819=>"011011111",
  30820=>"001010000",
  30821=>"010101100",
  30822=>"100111010",
  30823=>"010110100",
  30824=>"101100101",
  30825=>"101100111",
  30826=>"001101011",
  30827=>"100011111",
  30828=>"000100111",
  30829=>"010001111",
  30830=>"011111011",
  30831=>"000100000",
  30832=>"010111011",
  30833=>"111110010",
  30834=>"011010101",
  30835=>"110010011",
  30836=>"111110000",
  30837=>"111110011",
  30838=>"111000001",
  30839=>"110010001",
  30840=>"010001101",
  30841=>"100100000",
  30842=>"011000010",
  30843=>"111010101",
  30844=>"001110111",
  30845=>"101000001",
  30846=>"110101011",
  30847=>"100000110",
  30848=>"010110000",
  30849=>"101011110",
  30850=>"001001100",
  30851=>"100011001",
  30852=>"001100110",
  30853=>"011001111",
  30854=>"100010011",
  30855=>"011101000",
  30856=>"100111110",
  30857=>"011110111",
  30858=>"000100100",
  30859=>"110111101",
  30860=>"111110000",
  30861=>"100010011",
  30862=>"111101011",
  30863=>"010001100",
  30864=>"001100100",
  30865=>"011000000",
  30866=>"100111110",
  30867=>"010111111",
  30868=>"001011001",
  30869=>"000101111",
  30870=>"101010010",
  30871=>"101100010",
  30872=>"010000011",
  30873=>"110111011",
  30874=>"110110101",
  30875=>"110010010",
  30876=>"110010101",
  30877=>"111101100",
  30878=>"011110011",
  30879=>"010110111",
  30880=>"010101100",
  30881=>"000001100",
  30882=>"010100111",
  30883=>"111110010",
  30884=>"101001011",
  30885=>"010111111",
  30886=>"000100001",
  30887=>"000101000",
  30888=>"110111101",
  30889=>"001001100",
  30890=>"111110001",
  30891=>"110001001",
  30892=>"010100111",
  30893=>"011110100",
  30894=>"101011101",
  30895=>"000101100",
  30896=>"011011110",
  30897=>"000110100",
  30898=>"010001101",
  30899=>"000101111",
  30900=>"000001001",
  30901=>"010100010",
  30902=>"100111010",
  30903=>"001000100",
  30904=>"111011011",
  30905=>"110111100",
  30906=>"100010100",
  30907=>"001010110",
  30908=>"001010010",
  30909=>"011111110",
  30910=>"110011101",
  30911=>"000001110",
  30912=>"000001101",
  30913=>"010011010",
  30914=>"000000000",
  30915=>"000111100",
  30916=>"110000110",
  30917=>"111110011",
  30918=>"100110110",
  30919=>"000010101",
  30920=>"011001001",
  30921=>"110111001",
  30922=>"010100010",
  30923=>"001000111",
  30924=>"101010000",
  30925=>"001101111",
  30926=>"110001111",
  30927=>"000101000",
  30928=>"001110000",
  30929=>"110010010",
  30930=>"101110000",
  30931=>"100011100",
  30932=>"100100001",
  30933=>"011000011",
  30934=>"011000111",
  30935=>"100101001",
  30936=>"100101000",
  30937=>"110001010",
  30938=>"010001001",
  30939=>"111001011",
  30940=>"001110011",
  30941=>"100101010",
  30942=>"111010000",
  30943=>"010010111",
  30944=>"110000000",
  30945=>"101101010",
  30946=>"100000001",
  30947=>"110010100",
  30948=>"111100001",
  30949=>"010000111",
  30950=>"001010000",
  30951=>"000111100",
  30952=>"111111100",
  30953=>"000100000",
  30954=>"110111010",
  30955=>"101000110",
  30956=>"101111101",
  30957=>"110001001",
  30958=>"100001100",
  30959=>"001110100",
  30960=>"101100101",
  30961=>"110110001",
  30962=>"011011001",
  30963=>"001111111",
  30964=>"010101110",
  30965=>"001001100",
  30966=>"111010111",
  30967=>"000111011",
  30968=>"111001001",
  30969=>"101110110",
  30970=>"101011110",
  30971=>"111110010",
  30972=>"011001111",
  30973=>"010010001",
  30974=>"101110110",
  30975=>"101001110",
  30976=>"100000001",
  30977=>"011101111",
  30978=>"100100001",
  30979=>"000011101",
  30980=>"101101100",
  30981=>"010010100",
  30982=>"011101000",
  30983=>"101100010",
  30984=>"001011000",
  30985=>"110110010",
  30986=>"001010010",
  30987=>"110110100",
  30988=>"000010010",
  30989=>"000110100",
  30990=>"011101101",
  30991=>"000001111",
  30992=>"001011010",
  30993=>"101111111",
  30994=>"001000000",
  30995=>"000000100",
  30996=>"011100100",
  30997=>"001010011",
  30998=>"100000010",
  30999=>"101001101",
  31000=>"010000000",
  31001=>"001000101",
  31002=>"100001000",
  31003=>"000000111",
  31004=>"011010001",
  31005=>"010101010",
  31006=>"110100011",
  31007=>"010111101",
  31008=>"000101000",
  31009=>"111001000",
  31010=>"101011011",
  31011=>"011110101",
  31012=>"110111100",
  31013=>"110101100",
  31014=>"101000000",
  31015=>"001011010",
  31016=>"111100010",
  31017=>"101101110",
  31018=>"011101101",
  31019=>"110001100",
  31020=>"001001100",
  31021=>"001101011",
  31022=>"010111000",
  31023=>"100100111",
  31024=>"111101110",
  31025=>"001001010",
  31026=>"011010010",
  31027=>"011101110",
  31028=>"101010100",
  31029=>"010100000",
  31030=>"011111011",
  31031=>"011000001",
  31032=>"000010100",
  31033=>"111111101",
  31034=>"000000111",
  31035=>"010101010",
  31036=>"001000100",
  31037=>"110101000",
  31038=>"000110110",
  31039=>"011100110",
  31040=>"111111111",
  31041=>"000001000",
  31042=>"100011000",
  31043=>"011110011",
  31044=>"101011110",
  31045=>"001111100",
  31046=>"101101101",
  31047=>"110101000",
  31048=>"000000000",
  31049=>"110000000",
  31050=>"010111010",
  31051=>"111011110",
  31052=>"110000011",
  31053=>"101101001",
  31054=>"010011101",
  31055=>"111101010",
  31056=>"010111110",
  31057=>"010010001",
  31058=>"011010101",
  31059=>"000111100",
  31060=>"010001101",
  31061=>"001111110",
  31062=>"111011000",
  31063=>"101111101",
  31064=>"110001010",
  31065=>"100000110",
  31066=>"101111101",
  31067=>"101010100",
  31068=>"100101101",
  31069=>"111101000",
  31070=>"011000011",
  31071=>"100010001",
  31072=>"011000111",
  31073=>"111011001",
  31074=>"000101001",
  31075=>"001010010",
  31076=>"111001011",
  31077=>"100111011",
  31078=>"100101011",
  31079=>"010111110",
  31080=>"011010001",
  31081=>"000100111",
  31082=>"011100011",
  31083=>"011000100",
  31084=>"100110011",
  31085=>"010101010",
  31086=>"001100111",
  31087=>"101100011",
  31088=>"001100100",
  31089=>"110110011",
  31090=>"100000110",
  31091=>"110000001",
  31092=>"110011101",
  31093=>"010001011",
  31094=>"111001110",
  31095=>"000001001",
  31096=>"011100101",
  31097=>"010000010",
  31098=>"100001001",
  31099=>"011111000",
  31100=>"110101000",
  31101=>"001100001",
  31102=>"110111101",
  31103=>"010110100",
  31104=>"111000000",
  31105=>"000101011",
  31106=>"010111001",
  31107=>"100111110",
  31108=>"110100001",
  31109=>"000100101",
  31110=>"110100110",
  31111=>"110100110",
  31112=>"000101000",
  31113=>"110011101",
  31114=>"101010001",
  31115=>"010110010",
  31116=>"011101100",
  31117=>"000001001",
  31118=>"101011100",
  31119=>"010110010",
  31120=>"100110000",
  31121=>"000101101",
  31122=>"000101111",
  31123=>"000101101",
  31124=>"111000011",
  31125=>"000110010",
  31126=>"100100000",
  31127=>"011100000",
  31128=>"101000101",
  31129=>"000101110",
  31130=>"000000011",
  31131=>"100000000",
  31132=>"011101011",
  31133=>"111111000",
  31134=>"000100000",
  31135=>"111011111",
  31136=>"111010010",
  31137=>"111001000",
  31138=>"111011100",
  31139=>"010100011",
  31140=>"110110010",
  31141=>"000111111",
  31142=>"110010000",
  31143=>"111110101",
  31144=>"110011100",
  31145=>"010010111",
  31146=>"001101110",
  31147=>"100011111",
  31148=>"000100011",
  31149=>"011010110",
  31150=>"100110011",
  31151=>"011001000",
  31152=>"001010100",
  31153=>"011000001",
  31154=>"111110101",
  31155=>"111100000",
  31156=>"100100011",
  31157=>"000001001",
  31158=>"111000011",
  31159=>"101110000",
  31160=>"111111110",
  31161=>"001010001",
  31162=>"101001000",
  31163=>"001110010",
  31164=>"000011001",
  31165=>"110110011",
  31166=>"011111001",
  31167=>"010011101",
  31168=>"101010101",
  31169=>"011101010",
  31170=>"000111101",
  31171=>"000111111",
  31172=>"000010110",
  31173=>"100101010",
  31174=>"010100110",
  31175=>"011010000",
  31176=>"101011111",
  31177=>"011010100",
  31178=>"000010010",
  31179=>"010110011",
  31180=>"100100111",
  31181=>"010111010",
  31182=>"001001110",
  31183=>"101000101",
  31184=>"010011111",
  31185=>"011001000",
  31186=>"010000010",
  31187=>"010010010",
  31188=>"101011111",
  31189=>"001001000",
  31190=>"110101011",
  31191=>"000001010",
  31192=>"101011010",
  31193=>"000000001",
  31194=>"010100001",
  31195=>"101100001",
  31196=>"111111001",
  31197=>"100111100",
  31198=>"000010101",
  31199=>"000110011",
  31200=>"010111100",
  31201=>"100101011",
  31202=>"111011101",
  31203=>"110100111",
  31204=>"011001100",
  31205=>"101000001",
  31206=>"001001011",
  31207=>"000000010",
  31208=>"011010010",
  31209=>"000001011",
  31210=>"101111110",
  31211=>"001100010",
  31212=>"000011110",
  31213=>"111011001",
  31214=>"100001111",
  31215=>"010011101",
  31216=>"001111111",
  31217=>"111011111",
  31218=>"010110000",
  31219=>"010100010",
  31220=>"000110011",
  31221=>"001111000",
  31222=>"001011101",
  31223=>"101010011",
  31224=>"001000001",
  31225=>"101000010",
  31226=>"110000000",
  31227=>"011011101",
  31228=>"001100111",
  31229=>"011010110",
  31230=>"001001101",
  31231=>"111110001",
  31232=>"110010101",
  31233=>"011111001",
  31234=>"000011000",
  31235=>"010000110",
  31236=>"110101011",
  31237=>"001101101",
  31238=>"111011100",
  31239=>"110110000",
  31240=>"010100111",
  31241=>"110001011",
  31242=>"101001101",
  31243=>"101101101",
  31244=>"010110010",
  31245=>"101100100",
  31246=>"000101111",
  31247=>"000001100",
  31248=>"100001101",
  31249=>"110001101",
  31250=>"010011010",
  31251=>"100000100",
  31252=>"000010000",
  31253=>"011011011",
  31254=>"111111001",
  31255=>"000010000",
  31256=>"110111011",
  31257=>"100100010",
  31258=>"011001011",
  31259=>"011000101",
  31260=>"110111101",
  31261=>"011101101",
  31262=>"000010101",
  31263=>"111100011",
  31264=>"010000000",
  31265=>"010001100",
  31266=>"001100011",
  31267=>"101110100",
  31268=>"100101010",
  31269=>"111001000",
  31270=>"111011001",
  31271=>"001111010",
  31272=>"010011100",
  31273=>"101111000",
  31274=>"111010100",
  31275=>"000100101",
  31276=>"100110000",
  31277=>"111000101",
  31278=>"010100101",
  31279=>"110111100",
  31280=>"010111010",
  31281=>"000111100",
  31282=>"000110011",
  31283=>"101100011",
  31284=>"011100111",
  31285=>"011110111",
  31286=>"011111001",
  31287=>"110110000",
  31288=>"000111111",
  31289=>"111110101",
  31290=>"110101001",
  31291=>"101110111",
  31292=>"110111110",
  31293=>"000011000",
  31294=>"010101000",
  31295=>"000011100",
  31296=>"001011111",
  31297=>"100111100",
  31298=>"010100110",
  31299=>"101100111",
  31300=>"101010010",
  31301=>"011101110",
  31302=>"010000001",
  31303=>"010001001",
  31304=>"011100110",
  31305=>"010100100",
  31306=>"000110000",
  31307=>"011011100",
  31308=>"101011100",
  31309=>"100001100",
  31310=>"011110101",
  31311=>"010110101",
  31312=>"000001111",
  31313=>"001001011",
  31314=>"001011000",
  31315=>"011011001",
  31316=>"010101100",
  31317=>"100010010",
  31318=>"111000100",
  31319=>"011001001",
  31320=>"010011010",
  31321=>"100011000",
  31322=>"111000011",
  31323=>"111010011",
  31324=>"001001001",
  31325=>"001101000",
  31326=>"110001110",
  31327=>"000001101",
  31328=>"111010110",
  31329=>"111100100",
  31330=>"001101011",
  31331=>"100001001",
  31332=>"000110000",
  31333=>"001110010",
  31334=>"010011001",
  31335=>"010101010",
  31336=>"011100010",
  31337=>"101001010",
  31338=>"101100101",
  31339=>"100110111",
  31340=>"100111110",
  31341=>"101101110",
  31342=>"010001001",
  31343=>"110010110",
  31344=>"000111001",
  31345=>"000000111",
  31346=>"000000111",
  31347=>"001110111",
  31348=>"011000110",
  31349=>"001000010",
  31350=>"100000110",
  31351=>"010010110",
  31352=>"011001110",
  31353=>"011001000",
  31354=>"010111110",
  31355=>"110110010",
  31356=>"011011000",
  31357=>"011111010",
  31358=>"000110011",
  31359=>"001010000",
  31360=>"000100011",
  31361=>"010101110",
  31362=>"110101110",
  31363=>"110011011",
  31364=>"000110100",
  31365=>"010110001",
  31366=>"110010111",
  31367=>"010011101",
  31368=>"101111000",
  31369=>"001001001",
  31370=>"111101001",
  31371=>"111010001",
  31372=>"111111101",
  31373=>"001011100",
  31374=>"110010011",
  31375=>"010101101",
  31376=>"101100111",
  31377=>"010101100",
  31378=>"111100011",
  31379=>"000000011",
  31380=>"010011100",
  31381=>"101010110",
  31382=>"110111110",
  31383=>"110101100",
  31384=>"101011101",
  31385=>"011100101",
  31386=>"011011001",
  31387=>"000111111",
  31388=>"001011000",
  31389=>"010000111",
  31390=>"100100010",
  31391=>"101111100",
  31392=>"000111101",
  31393=>"001111001",
  31394=>"000001011",
  31395=>"000010100",
  31396=>"100100000",
  31397=>"100110011",
  31398=>"010011001",
  31399=>"100110001",
  31400=>"110111000",
  31401=>"000110000",
  31402=>"101111010",
  31403=>"100001010",
  31404=>"111100000",
  31405=>"100001001",
  31406=>"001111101",
  31407=>"111101110",
  31408=>"010000011",
  31409=>"101001000",
  31410=>"100100110",
  31411=>"000100011",
  31412=>"101011000",
  31413=>"100001101",
  31414=>"111001100",
  31415=>"100110000",
  31416=>"101011100",
  31417=>"010010101",
  31418=>"101111001",
  31419=>"001100011",
  31420=>"000111111",
  31421=>"101010111",
  31422=>"110001010",
  31423=>"001000000",
  31424=>"000011010",
  31425=>"010000110",
  31426=>"010100101",
  31427=>"111101100",
  31428=>"100001101",
  31429=>"010001101",
  31430=>"110111000",
  31431=>"000110111",
  31432=>"000000000",
  31433=>"011001100",
  31434=>"001011110",
  31435=>"010001000",
  31436=>"110001010",
  31437=>"100011001",
  31438=>"101010011",
  31439=>"000010101",
  31440=>"000110000",
  31441=>"101000101",
  31442=>"011001011",
  31443=>"001110100",
  31444=>"000101010",
  31445=>"000010011",
  31446=>"001011001",
  31447=>"011010100",
  31448=>"110001100",
  31449=>"010011111",
  31450=>"000101111",
  31451=>"000000101",
  31452=>"001100000",
  31453=>"110100101",
  31454=>"111000111",
  31455=>"100100110",
  31456=>"111011101",
  31457=>"101101001",
  31458=>"011111001",
  31459=>"010110001",
  31460=>"111111001",
  31461=>"001011111",
  31462=>"000010100",
  31463=>"010111101",
  31464=>"010101110",
  31465=>"011110000",
  31466=>"011000010",
  31467=>"110000111",
  31468=>"000001011",
  31469=>"101101001",
  31470=>"101110100",
  31471=>"010101010",
  31472=>"100010000",
  31473=>"111001101",
  31474=>"001101101",
  31475=>"101011101",
  31476=>"110100100",
  31477=>"000000001",
  31478=>"111110000",
  31479=>"001010010",
  31480=>"001111010",
  31481=>"100000011",
  31482=>"101110010",
  31483=>"001100011",
  31484=>"101011001",
  31485=>"111000001",
  31486=>"011101010",
  31487=>"100010001",
  31488=>"101110001",
  31489=>"001010001",
  31490=>"010000010",
  31491=>"010111101",
  31492=>"010101111",
  31493=>"011111010",
  31494=>"111101001",
  31495=>"110000000",
  31496=>"111000000",
  31497=>"101001000",
  31498=>"100100000",
  31499=>"000000011",
  31500=>"101101000",
  31501=>"011001101",
  31502=>"100111010",
  31503=>"100010100",
  31504=>"001110000",
  31505=>"111101100",
  31506=>"100101110",
  31507=>"000100010",
  31508=>"100001110",
  31509=>"010101001",
  31510=>"110001011",
  31511=>"101111111",
  31512=>"101001101",
  31513=>"000000000",
  31514=>"011001111",
  31515=>"110111110",
  31516=>"100110111",
  31517=>"110111110",
  31518=>"110000111",
  31519=>"111110111",
  31520=>"001000010",
  31521=>"010001000",
  31522=>"001011110",
  31523=>"001100110",
  31524=>"010011111",
  31525=>"100110001",
  31526=>"011111010",
  31527=>"001100100",
  31528=>"110011000",
  31529=>"110010100",
  31530=>"010001110",
  31531=>"110101100",
  31532=>"011110010",
  31533=>"011100111",
  31534=>"000010100",
  31535=>"001001100",
  31536=>"100000100",
  31537=>"111001111",
  31538=>"100000001",
  31539=>"111011110",
  31540=>"000000010",
  31541=>"110111111",
  31542=>"101101000",
  31543=>"010111110",
  31544=>"001011110",
  31545=>"000100100",
  31546=>"001010001",
  31547=>"000000000",
  31548=>"110001001",
  31549=>"001100010",
  31550=>"010010101",
  31551=>"001101110",
  31552=>"000011000",
  31553=>"001010010",
  31554=>"111111100",
  31555=>"111111101",
  31556=>"100011011",
  31557=>"111000101",
  31558=>"101110010",
  31559=>"011111011",
  31560=>"111000101",
  31561=>"000110000",
  31562=>"111101001",
  31563=>"101000001",
  31564=>"100100110",
  31565=>"101110110",
  31566=>"001001101",
  31567=>"000111000",
  31568=>"011100001",
  31569=>"101111010",
  31570=>"000111010",
  31571=>"011001000",
  31572=>"001100111",
  31573=>"011110011",
  31574=>"101001100",
  31575=>"000000001",
  31576=>"110111111",
  31577=>"110000010",
  31578=>"100101111",
  31579=>"000001111",
  31580=>"000011000",
  31581=>"111001111",
  31582=>"010101001",
  31583=>"111001100",
  31584=>"111010110",
  31585=>"101010011",
  31586=>"010001110",
  31587=>"111001100",
  31588=>"100111101",
  31589=>"010101000",
  31590=>"100001100",
  31591=>"000101101",
  31592=>"011101101",
  31593=>"101100100",
  31594=>"010001111",
  31595=>"010001110",
  31596=>"110010100",
  31597=>"001000001",
  31598=>"111100100",
  31599=>"100110110",
  31600=>"011110001",
  31601=>"100001111",
  31602=>"010001110",
  31603=>"111001110",
  31604=>"011101111",
  31605=>"010010111",
  31606=>"010110010",
  31607=>"111010101",
  31608=>"001010100",
  31609=>"011000111",
  31610=>"111010110",
  31611=>"011001001",
  31612=>"011111011",
  31613=>"110101001",
  31614=>"100110000",
  31615=>"001110001",
  31616=>"111011011",
  31617=>"001111011",
  31618=>"101100111",
  31619=>"000011101",
  31620=>"000000100",
  31621=>"110000010",
  31622=>"010000011",
  31623=>"000010111",
  31624=>"010001101",
  31625=>"000110011",
  31626=>"011000001",
  31627=>"001011100",
  31628=>"100011110",
  31629=>"010110110",
  31630=>"110111101",
  31631=>"000110111",
  31632=>"001100101",
  31633=>"111110000",
  31634=>"000101011",
  31635=>"111100011",
  31636=>"001000001",
  31637=>"010010111",
  31638=>"011100111",
  31639=>"100001000",
  31640=>"110011110",
  31641=>"000010111",
  31642=>"000100011",
  31643=>"100111111",
  31644=>"010111000",
  31645=>"000110111",
  31646=>"011111010",
  31647=>"010101100",
  31648=>"100011000",
  31649=>"111111010",
  31650=>"101001011",
  31651=>"010000111",
  31652=>"001100000",
  31653=>"000100100",
  31654=>"111010011",
  31655=>"110001101",
  31656=>"001100001",
  31657=>"011111000",
  31658=>"010101010",
  31659=>"000110111",
  31660=>"111101010",
  31661=>"111000001",
  31662=>"000001101",
  31663=>"110110110",
  31664=>"000100000",
  31665=>"011010111",
  31666=>"111000100",
  31667=>"011111010",
  31668=>"101001100",
  31669=>"100001110",
  31670=>"110001110",
  31671=>"100010111",
  31672=>"111110101",
  31673=>"101101011",
  31674=>"101101101",
  31675=>"101010000",
  31676=>"110000000",
  31677=>"101110001",
  31678=>"101000111",
  31679=>"110101000",
  31680=>"000100000",
  31681=>"011101101",
  31682=>"110110001",
  31683=>"011000001",
  31684=>"000111111",
  31685=>"001101100",
  31686=>"001101100",
  31687=>"011001010",
  31688=>"100111101",
  31689=>"001100000",
  31690=>"011010011",
  31691=>"110010011",
  31692=>"100011010",
  31693=>"000000001",
  31694=>"101001001",
  31695=>"100101011",
  31696=>"110001110",
  31697=>"100111000",
  31698=>"011110001",
  31699=>"000000100",
  31700=>"011001001",
  31701=>"001000001",
  31702=>"001101001",
  31703=>"000001000",
  31704=>"000111110",
  31705=>"000001101",
  31706=>"110100111",
  31707=>"111000111",
  31708=>"111111110",
  31709=>"011010101",
  31710=>"101101110",
  31711=>"110100011",
  31712=>"011101100",
  31713=>"000111111",
  31714=>"101001111",
  31715=>"101110111",
  31716=>"010010010",
  31717=>"101100011",
  31718=>"000100110",
  31719=>"000111000",
  31720=>"100101111",
  31721=>"110110111",
  31722=>"110111010",
  31723=>"010101011",
  31724=>"001011010",
  31725=>"110101101",
  31726=>"000100001",
  31727=>"000111011",
  31728=>"110000100",
  31729=>"101000111",
  31730=>"001001101",
  31731=>"011110011",
  31732=>"000000100",
  31733=>"000101111",
  31734=>"111011111",
  31735=>"001110000",
  31736=>"011110010",
  31737=>"101110110",
  31738=>"110101100",
  31739=>"011111111",
  31740=>"110100100",
  31741=>"010111010",
  31742=>"101000010",
  31743=>"111001100",
  31744=>"000011111",
  31745=>"001100010",
  31746=>"000011100",
  31747=>"010011100",
  31748=>"100001000",
  31749=>"010110110",
  31750=>"110110010",
  31751=>"110100011",
  31752=>"010001111",
  31753=>"110000001",
  31754=>"000000100",
  31755=>"011011001",
  31756=>"011110011",
  31757=>"010001110",
  31758=>"110111100",
  31759=>"110110001",
  31760=>"101110110",
  31761=>"100111111",
  31762=>"111100011",
  31763=>"110000101",
  31764=>"111101111",
  31765=>"010000101",
  31766=>"011001010",
  31767=>"100100011",
  31768=>"100101100",
  31769=>"000010110",
  31770=>"000110111",
  31771=>"110000101",
  31772=>"100101011",
  31773=>"011101111",
  31774=>"010101010",
  31775=>"110000110",
  31776=>"000011110",
  31777=>"110001011",
  31778=>"011000100",
  31779=>"000010010",
  31780=>"001000011",
  31781=>"101010111",
  31782=>"110010011",
  31783=>"100101110",
  31784=>"010100011",
  31785=>"101101101",
  31786=>"110110010",
  31787=>"101011010",
  31788=>"111010111",
  31789=>"111100101",
  31790=>"001100100",
  31791=>"011110111",
  31792=>"011000011",
  31793=>"001011001",
  31794=>"110101010",
  31795=>"100100100",
  31796=>"000111000",
  31797=>"111001001",
  31798=>"011110001",
  31799=>"000000000",
  31800=>"000011000",
  31801=>"110101110",
  31802=>"001000000",
  31803=>"110101101",
  31804=>"001101111",
  31805=>"100011111",
  31806=>"010110110",
  31807=>"011101101",
  31808=>"001110101",
  31809=>"100100111",
  31810=>"111001101",
  31811=>"010000100",
  31812=>"110100010",
  31813=>"011001111",
  31814=>"001001001",
  31815=>"111111001",
  31816=>"101111010",
  31817=>"000111111",
  31818=>"100010011",
  31819=>"110100001",
  31820=>"010011110",
  31821=>"110000110",
  31822=>"100001010",
  31823=>"110111100",
  31824=>"111000011",
  31825=>"000100110",
  31826=>"100110110",
  31827=>"100100101",
  31828=>"100011111",
  31829=>"110001000",
  31830=>"001010100",
  31831=>"000101000",
  31832=>"101010111",
  31833=>"101000101",
  31834=>"010010001",
  31835=>"110100110",
  31836=>"000100101",
  31837=>"101001101",
  31838=>"010111000",
  31839=>"011011111",
  31840=>"000110100",
  31841=>"101001100",
  31842=>"000010000",
  31843=>"111110110",
  31844=>"000100001",
  31845=>"011111101",
  31846=>"001110001",
  31847=>"100111001",
  31848=>"110101011",
  31849=>"001100011",
  31850=>"001100111",
  31851=>"111111101",
  31852=>"100001000",
  31853=>"100011001",
  31854=>"101011010",
  31855=>"000001110",
  31856=>"110111001",
  31857=>"010100011",
  31858=>"000001001",
  31859=>"000010111",
  31860=>"010001010",
  31861=>"100000111",
  31862=>"101101101",
  31863=>"000010110",
  31864=>"000110111",
  31865=>"011001111",
  31866=>"010100111",
  31867=>"010001010",
  31868=>"110101000",
  31869=>"101101101",
  31870=>"000100010",
  31871=>"011010100",
  31872=>"111101000",
  31873=>"111101110",
  31874=>"001101110",
  31875=>"001010000",
  31876=>"110000100",
  31877=>"100001010",
  31878=>"101000110",
  31879=>"111010101",
  31880=>"101001010",
  31881=>"101000111",
  31882=>"000000100",
  31883=>"010101111",
  31884=>"010111010",
  31885=>"010100011",
  31886=>"111110111",
  31887=>"010100010",
  31888=>"000100100",
  31889=>"010100001",
  31890=>"000010110",
  31891=>"110000011",
  31892=>"011111001",
  31893=>"001010111",
  31894=>"100000001",
  31895=>"000110111",
  31896=>"100011110",
  31897=>"000101001",
  31898=>"000111101",
  31899=>"101101100",
  31900=>"100001111",
  31901=>"010010100",
  31902=>"000100001",
  31903=>"001011111",
  31904=>"101000111",
  31905=>"000001100",
  31906=>"000000111",
  31907=>"011101110",
  31908=>"010110001",
  31909=>"111110101",
  31910=>"010100111",
  31911=>"111110010",
  31912=>"111000000",
  31913=>"010111010",
  31914=>"111000100",
  31915=>"000111100",
  31916=>"000010010",
  31917=>"100111111",
  31918=>"010001111",
  31919=>"011010000",
  31920=>"010100101",
  31921=>"011111000",
  31922=>"111111100",
  31923=>"001010000",
  31924=>"110110000",
  31925=>"010111001",
  31926=>"111010000",
  31927=>"110110101",
  31928=>"010100101",
  31929=>"111000011",
  31930=>"010111100",
  31931=>"110101011",
  31932=>"011100001",
  31933=>"101110001",
  31934=>"111011011",
  31935=>"000001101",
  31936=>"100110011",
  31937=>"011010010",
  31938=>"111001100",
  31939=>"101111111",
  31940=>"110000000",
  31941=>"101100101",
  31942=>"100010010",
  31943=>"100100000",
  31944=>"111101001",
  31945=>"110111110",
  31946=>"111110000",
  31947=>"011100001",
  31948=>"001000110",
  31949=>"011101101",
  31950=>"110010000",
  31951=>"010001110",
  31952=>"010011001",
  31953=>"001101010",
  31954=>"000100001",
  31955=>"010001110",
  31956=>"111000010",
  31957=>"101000110",
  31958=>"101000100",
  31959=>"000111101",
  31960=>"001101100",
  31961=>"110010100",
  31962=>"011100100",
  31963=>"010000000",
  31964=>"011010000",
  31965=>"010100110",
  31966=>"111101011",
  31967=>"001101111",
  31968=>"010001101",
  31969=>"110010010",
  31970=>"111001100",
  31971=>"011001100",
  31972=>"000000100",
  31973=>"010100001",
  31974=>"100110110",
  31975=>"011000100",
  31976=>"011100011",
  31977=>"100010000",
  31978=>"110101010",
  31979=>"110110010",
  31980=>"000000010",
  31981=>"100100110",
  31982=>"101110010",
  31983=>"011000001",
  31984=>"111111011",
  31985=>"011000100",
  31986=>"101100110",
  31987=>"100011101",
  31988=>"010011000",
  31989=>"010010011",
  31990=>"011111000",
  31991=>"010000110",
  31992=>"010100110",
  31993=>"101101110",
  31994=>"000100001",
  31995=>"010000111",
  31996=>"010000011",
  31997=>"101010001",
  31998=>"011011010",
  31999=>"100011001",
  32000=>"111110111",
  32001=>"100011010",
  32002=>"000001000",
  32003=>"011011100",
  32004=>"010010111",
  32005=>"001101011",
  32006=>"110111110",
  32007=>"010011101",
  32008=>"110001101",
  32009=>"101110000",
  32010=>"101000011",
  32011=>"001110101",
  32012=>"001111111",
  32013=>"010000000",
  32014=>"010110011",
  32015=>"001011111",
  32016=>"111000010",
  32017=>"100101111",
  32018=>"110111010",
  32019=>"110000100",
  32020=>"111010010",
  32021=>"111111101",
  32022=>"011100000",
  32023=>"101110100",
  32024=>"101100111",
  32025=>"010011110",
  32026=>"101011101",
  32027=>"111101000",
  32028=>"101111110",
  32029=>"110100001",
  32030=>"100111011",
  32031=>"100100110",
  32032=>"010101100",
  32033=>"101001011",
  32034=>"010101101",
  32035=>"001100110",
  32036=>"111101000",
  32037=>"011111011",
  32038=>"110110001",
  32039=>"000110001",
  32040=>"001010100",
  32041=>"010010101",
  32042=>"000110001",
  32043=>"010101100",
  32044=>"000010011",
  32045=>"110110100",
  32046=>"011101001",
  32047=>"110100001",
  32048=>"111110100",
  32049=>"101000000",
  32050=>"100111110",
  32051=>"001011101",
  32052=>"011011101",
  32053=>"100110110",
  32054=>"111010010",
  32055=>"110010010",
  32056=>"011101111",
  32057=>"000001111",
  32058=>"111100001",
  32059=>"101001000",
  32060=>"001111100",
  32061=>"101100010",
  32062=>"010110110",
  32063=>"001000101",
  32064=>"101100111",
  32065=>"010010011",
  32066=>"100011000",
  32067=>"101001001",
  32068=>"111110001",
  32069=>"011000110",
  32070=>"101010100",
  32071=>"101010110",
  32072=>"111100000",
  32073=>"000110011",
  32074=>"011101011",
  32075=>"010110010",
  32076=>"011111100",
  32077=>"110100011",
  32078=>"011001100",
  32079=>"111101110",
  32080=>"011010100",
  32081=>"100100010",
  32082=>"101010010",
  32083=>"101010000",
  32084=>"011111011",
  32085=>"011110010",
  32086=>"110000110",
  32087=>"010101001",
  32088=>"100001011",
  32089=>"011111110",
  32090=>"011011001",
  32091=>"001100100",
  32092=>"111001010",
  32093=>"110111111",
  32094=>"101001000",
  32095=>"000010011",
  32096=>"001011011",
  32097=>"010111111",
  32098=>"110010111",
  32099=>"001001101",
  32100=>"010100110",
  32101=>"000100111",
  32102=>"010101101",
  32103=>"110100101",
  32104=>"010111110",
  32105=>"001001001",
  32106=>"001010001",
  32107=>"101100101",
  32108=>"110101101",
  32109=>"010010000",
  32110=>"100010001",
  32111=>"101011110",
  32112=>"000001101",
  32113=>"110000001",
  32114=>"110101001",
  32115=>"010000111",
  32116=>"100101000",
  32117=>"011011100",
  32118=>"110010110",
  32119=>"100100001",
  32120=>"100111101",
  32121=>"011100111",
  32122=>"110011011",
  32123=>"111010010",
  32124=>"101010001",
  32125=>"010010001",
  32126=>"000110001",
  32127=>"110101000",
  32128=>"000010000",
  32129=>"000010100",
  32130=>"010100001",
  32131=>"111100011",
  32132=>"110100100",
  32133=>"000100001",
  32134=>"101010010",
  32135=>"101111100",
  32136=>"100100001",
  32137=>"011111101",
  32138=>"101011011",
  32139=>"101010101",
  32140=>"100011101",
  32141=>"110000110",
  32142=>"111010011",
  32143=>"001101111",
  32144=>"001000101",
  32145=>"011000001",
  32146=>"001010110",
  32147=>"101110110",
  32148=>"101101000",
  32149=>"000000110",
  32150=>"101010010",
  32151=>"001011000",
  32152=>"010001101",
  32153=>"100101101",
  32154=>"001101001",
  32155=>"000001111",
  32156=>"000000100",
  32157=>"000101010",
  32158=>"100000001",
  32159=>"111010011",
  32160=>"001000100",
  32161=>"110100011",
  32162=>"100110010",
  32163=>"111011001",
  32164=>"001110011",
  32165=>"011101000",
  32166=>"001001000",
  32167=>"111010011",
  32168=>"011001100",
  32169=>"101001111",
  32170=>"100011111",
  32171=>"111100110",
  32172=>"011000101",
  32173=>"000111010",
  32174=>"110111010",
  32175=>"101110001",
  32176=>"100110111",
  32177=>"110011001",
  32178=>"011100100",
  32179=>"110101100",
  32180=>"101101000",
  32181=>"011100111",
  32182=>"100101010",
  32183=>"100010011",
  32184=>"110100000",
  32185=>"010001001",
  32186=>"000000100",
  32187=>"001111001",
  32188=>"001011110",
  32189=>"000101111",
  32190=>"101111100",
  32191=>"111111101",
  32192=>"011011100",
  32193=>"001100001",
  32194=>"111110101",
  32195=>"110001111",
  32196=>"000000000",
  32197=>"111101100",
  32198=>"010010011",
  32199=>"111001110",
  32200=>"101110010",
  32201=>"111011100",
  32202=>"000110110",
  32203=>"100010001",
  32204=>"101011101",
  32205=>"101000001",
  32206=>"001111001",
  32207=>"000001101",
  32208=>"001001100",
  32209=>"110101001",
  32210=>"001010000",
  32211=>"011110110",
  32212=>"001000111",
  32213=>"001010000",
  32214=>"110000011",
  32215=>"000110101",
  32216=>"111001000",
  32217=>"001110101",
  32218=>"000111111",
  32219=>"001111000",
  32220=>"000100010",
  32221=>"111010100",
  32222=>"101111111",
  32223=>"011000110",
  32224=>"010111000",
  32225=>"101100010",
  32226=>"001111111",
  32227=>"111001010",
  32228=>"000111111",
  32229=>"100010100",
  32230=>"001000100",
  32231=>"011111001",
  32232=>"010011111",
  32233=>"110110100",
  32234=>"001110000",
  32235=>"010111111",
  32236=>"110001011",
  32237=>"111101110",
  32238=>"001000001",
  32239=>"101010101",
  32240=>"100001101",
  32241=>"111010101",
  32242=>"101111111",
  32243=>"101000110",
  32244=>"011000000",
  32245=>"010111011",
  32246=>"001000110",
  32247=>"001110010",
  32248=>"111101011",
  32249=>"101111010",
  32250=>"111110111",
  32251=>"100010110",
  32252=>"110011110",
  32253=>"010111111",
  32254=>"100010100",
  32255=>"010101011",
  32256=>"101011001",
  32257=>"110100110",
  32258=>"010010111",
  32259=>"000011011",
  32260=>"001110101",
  32261=>"110100000",
  32262=>"001101111",
  32263=>"011011001",
  32264=>"100110010",
  32265=>"000001100",
  32266=>"101100010",
  32267=>"100000000",
  32268=>"000110010",
  32269=>"110011100",
  32270=>"010001110",
  32271=>"001000100",
  32272=>"001101000",
  32273=>"101110101",
  32274=>"101000000",
  32275=>"101101010",
  32276=>"001010110",
  32277=>"001111001",
  32278=>"011111001",
  32279=>"011111101",
  32280=>"100001010",
  32281=>"101010111",
  32282=>"100101001",
  32283=>"111111010",
  32284=>"001110101",
  32285=>"100110101",
  32286=>"111001000",
  32287=>"100100100",
  32288=>"111101110",
  32289=>"011110101",
  32290=>"001100101",
  32291=>"011010111",
  32292=>"000110000",
  32293=>"010001011",
  32294=>"001011011",
  32295=>"110110001",
  32296=>"010101101",
  32297=>"111010001",
  32298=>"100001001",
  32299=>"000110000",
  32300=>"101100000",
  32301=>"100001001",
  32302=>"010011111",
  32303=>"110011011",
  32304=>"111100000",
  32305=>"111101011",
  32306=>"001101111",
  32307=>"010000101",
  32308=>"110100100",
  32309=>"101111010",
  32310=>"011100101",
  32311=>"101110101",
  32312=>"101011100",
  32313=>"110111010",
  32314=>"000101100",
  32315=>"111001001",
  32316=>"001001000",
  32317=>"000010111",
  32318=>"101101110",
  32319=>"001101100",
  32320=>"011101111",
  32321=>"010001000",
  32322=>"111101100",
  32323=>"011100011",
  32324=>"100111010",
  32325=>"011010000",
  32326=>"101000000",
  32327=>"000101010",
  32328=>"001101101",
  32329=>"001101000",
  32330=>"111000010",
  32331=>"100010000",
  32332=>"100001010",
  32333=>"000110010",
  32334=>"010111111",
  32335=>"010110000",
  32336=>"000000110",
  32337=>"101101001",
  32338=>"101101110",
  32339=>"101101000",
  32340=>"101110110",
  32341=>"101111001",
  32342=>"101001000",
  32343=>"111101101",
  32344=>"101000111",
  32345=>"101011000",
  32346=>"001000001",
  32347=>"001011101",
  32348=>"101111101",
  32349=>"110111001",
  32350=>"100011100",
  32351=>"111111101",
  32352=>"000100001",
  32353=>"100100100",
  32354=>"001000110",
  32355=>"110110111",
  32356=>"010111001",
  32357=>"010100000",
  32358=>"100111101",
  32359=>"111001111",
  32360=>"001111000",
  32361=>"111111011",
  32362=>"010100011",
  32363=>"100101101",
  32364=>"100101000",
  32365=>"101001000",
  32366=>"111101111",
  32367=>"101010000",
  32368=>"100101101",
  32369=>"101110101",
  32370=>"000000010",
  32371=>"111110110",
  32372=>"100111010",
  32373=>"001111010",
  32374=>"010101101",
  32375=>"101101010",
  32376=>"100001001",
  32377=>"101011110",
  32378=>"010111010",
  32379=>"111111000",
  32380=>"001100110",
  32381=>"101111000",
  32382=>"011011001",
  32383=>"001110111",
  32384=>"110001110",
  32385=>"001101000",
  32386=>"011111111",
  32387=>"100100000",
  32388=>"110000110",
  32389=>"101100000",
  32390=>"011110000",
  32391=>"111101001",
  32392=>"100101001",
  32393=>"110111011",
  32394=>"111110000",
  32395=>"111001010",
  32396=>"110100110",
  32397=>"111001010",
  32398=>"101010011",
  32399=>"100100000",
  32400=>"010111000",
  32401=>"011110010",
  32402=>"110010111",
  32403=>"111001011",
  32404=>"001011001",
  32405=>"011001100",
  32406=>"011101001",
  32407=>"011110100",
  32408=>"100100101",
  32409=>"110111101",
  32410=>"010010010",
  32411=>"000001100",
  32412=>"010101010",
  32413=>"101100000",
  32414=>"110100000",
  32415=>"111101101",
  32416=>"001101000",
  32417=>"110001001",
  32418=>"100010111",
  32419=>"001111000",
  32420=>"000101100",
  32421=>"000000100",
  32422=>"101111111",
  32423=>"100001100",
  32424=>"110101100",
  32425=>"000000000",
  32426=>"000101000",
  32427=>"010000111",
  32428=>"010000111",
  32429=>"111110000",
  32430=>"000001100",
  32431=>"000111101",
  32432=>"010101001",
  32433=>"110110101",
  32434=>"100100110",
  32435=>"000010000",
  32436=>"101010101",
  32437=>"101111110",
  32438=>"011000010",
  32439=>"111001100",
  32440=>"010111101",
  32441=>"111100100",
  32442=>"010001011",
  32443=>"110111110",
  32444=>"000110011",
  32445=>"000111010",
  32446=>"100011010",
  32447=>"001100101",
  32448=>"000111110",
  32449=>"010000010",
  32450=>"101001110",
  32451=>"010001111",
  32452=>"001101000",
  32453=>"110100101",
  32454=>"001111001",
  32455=>"010001100",
  32456=>"000011110",
  32457=>"000111001",
  32458=>"000100011",
  32459=>"101110000",
  32460=>"111001110",
  32461=>"000001100",
  32462=>"001110111",
  32463=>"100001100",
  32464=>"111000100",
  32465=>"011101011",
  32466=>"100000111",
  32467=>"011000001",
  32468=>"101011111",
  32469=>"001010011",
  32470=>"100010100",
  32471=>"001100101",
  32472=>"110111011",
  32473=>"011011101",
  32474=>"101000000",
  32475=>"000010001",
  32476=>"100010001",
  32477=>"010110011",
  32478=>"100100101",
  32479=>"010001011",
  32480=>"011011000",
  32481=>"110000011",
  32482=>"110101100",
  32483=>"001101111",
  32484=>"000111000",
  32485=>"100011000",
  32486=>"010011000",
  32487=>"000101101",
  32488=>"101110011",
  32489=>"101000010",
  32490=>"101101100",
  32491=>"110011011",
  32492=>"010011111",
  32493=>"010010100",
  32494=>"101011000",
  32495=>"101101000",
  32496=>"001111101",
  32497=>"011010011",
  32498=>"110010001",
  32499=>"110111111",
  32500=>"110010000",
  32501=>"101000101",
  32502=>"100010111",
  32503=>"011101100",
  32504=>"011001011",
  32505=>"001010111",
  32506=>"101100010",
  32507=>"011101000",
  32508=>"100110110",
  32509=>"101111000",
  32510=>"110110100",
  32511=>"100101010",
  32512=>"001101011",
  32513=>"000011100",
  32514=>"100111011",
  32515=>"010001110",
  32516=>"111101110",
  32517=>"001001100",
  32518=>"110101011",
  32519=>"011111001",
  32520=>"010101000",
  32521=>"100001100",
  32522=>"010000101",
  32523=>"110101111",
  32524=>"110111000",
  32525=>"010010110",
  32526=>"111100110",
  32527=>"111100100",
  32528=>"000000010",
  32529=>"110110100",
  32530=>"000111001",
  32531=>"001010100",
  32532=>"100001100",
  32533=>"110001010",
  32534=>"010100101",
  32535=>"101011111",
  32536=>"101101111",
  32537=>"100101000",
  32538=>"010010001",
  32539=>"010010111",
  32540=>"010000001",
  32541=>"011100010",
  32542=>"110111001",
  32543=>"101101111",
  32544=>"000111001",
  32545=>"101100101",
  32546=>"000010100",
  32547=>"101001100",
  32548=>"101010010",
  32549=>"000000000",
  32550=>"000000001",
  32551=>"000010101",
  32552=>"000001011",
  32553=>"111100011",
  32554=>"100110111",
  32555=>"010011110",
  32556=>"001010000",
  32557=>"010000010",
  32558=>"001010100",
  32559=>"011000100",
  32560=>"001110110",
  32561=>"010001000",
  32562=>"001000111",
  32563=>"111011010",
  32564=>"011110100",
  32565=>"101010101",
  32566=>"010110000",
  32567=>"101001100",
  32568=>"100010000",
  32569=>"001101001",
  32570=>"001101000",
  32571=>"110111100",
  32572=>"111111001",
  32573=>"110000110",
  32574=>"111101000",
  32575=>"100111010",
  32576=>"111100111",
  32577=>"010100001",
  32578=>"010101010",
  32579=>"101000111",
  32580=>"011110011",
  32581=>"110011111",
  32582=>"001111110",
  32583=>"111111111",
  32584=>"110000001",
  32585=>"001001111",
  32586=>"111110110",
  32587=>"001011001",
  32588=>"010000001",
  32589=>"011110000",
  32590=>"101100110",
  32591=>"100111101",
  32592=>"100001100",
  32593=>"011001001",
  32594=>"000010001",
  32595=>"001000111",
  32596=>"111110010",
  32597=>"001111111",
  32598=>"111101110",
  32599=>"101001000",
  32600=>"010111100",
  32601=>"101010110",
  32602=>"001100101",
  32603=>"010001001",
  32604=>"010000000",
  32605=>"101011000",
  32606=>"000100010",
  32607=>"001001010",
  32608=>"001100001",
  32609=>"000111010",
  32610=>"011011111",
  32611=>"101010000",
  32612=>"001010001",
  32613=>"110011001",
  32614=>"111111110",
  32615=>"110000000",
  32616=>"111101001",
  32617=>"001101101",
  32618=>"011111101",
  32619=>"001001101",
  32620=>"100110111",
  32621=>"001111101",
  32622=>"101110111",
  32623=>"000011000",
  32624=>"010100101",
  32625=>"110101011",
  32626=>"001101111",
  32627=>"101001101",
  32628=>"111100110",
  32629=>"001001100",
  32630=>"000010110",
  32631=>"000110111",
  32632=>"101110101",
  32633=>"111001000",
  32634=>"000100000",
  32635=>"000000000",
  32636=>"000110110",
  32637=>"011001010",
  32638=>"011001000",
  32639=>"011011101",
  32640=>"111001101",
  32641=>"100100110",
  32642=>"011111011",
  32643=>"010000110",
  32644=>"101011110",
  32645=>"000011100",
  32646=>"110011101",
  32647=>"100111001",
  32648=>"001100101",
  32649=>"110011101",
  32650=>"011001011",
  32651=>"111111110",
  32652=>"101100100",
  32653=>"010000100",
  32654=>"110100000",
  32655=>"011101010",
  32656=>"111110001",
  32657=>"111011001",
  32658=>"000111100",
  32659=>"110000101",
  32660=>"011101000",
  32661=>"000010001",
  32662=>"010011110",
  32663=>"001000101",
  32664=>"001110010",
  32665=>"010110001",
  32666=>"011010001",
  32667=>"101100111",
  32668=>"100100001",
  32669=>"000001111",
  32670=>"001101000",
  32671=>"100000001",
  32672=>"001001100",
  32673=>"010010001",
  32674=>"110001111",
  32675=>"111000111",
  32676=>"100111010",
  32677=>"110011110",
  32678=>"101011011",
  32679=>"010000100",
  32680=>"101011001",
  32681=>"001001011",
  32682=>"111000000",
  32683=>"100101111",
  32684=>"010000111",
  32685=>"011100001",
  32686=>"110110001",
  32687=>"100110110",
  32688=>"001110001",
  32689=>"111011000",
  32690=>"001001010",
  32691=>"110111110",
  32692=>"001110100",
  32693=>"001111010",
  32694=>"000111111",
  32695=>"001101011",
  32696=>"000011100",
  32697=>"111101110",
  32698=>"011000010",
  32699=>"010101010",
  32700=>"101111101",
  32701=>"111011111",
  32702=>"000000000",
  32703=>"100010111",
  32704=>"100110010",
  32705=>"110101011",
  32706=>"110011010",
  32707=>"110110100",
  32708=>"111011100",
  32709=>"111101111",
  32710=>"001110101",
  32711=>"110111110",
  32712=>"011100111",
  32713=>"001111000",
  32714=>"111111110",
  32715=>"100111111",
  32716=>"001011110",
  32717=>"110110101",
  32718=>"011001101",
  32719=>"011101000",
  32720=>"011001101",
  32721=>"101111101",
  32722=>"111111111",
  32723=>"010100100",
  32724=>"100011000",
  32725=>"100100101",
  32726=>"010000101",
  32727=>"111110110",
  32728=>"101011100",
  32729=>"000110000",
  32730=>"110000011",
  32731=>"011011111",
  32732=>"110100011",
  32733=>"100111011",
  32734=>"001000010",
  32735=>"000101011",
  32736=>"001100101",
  32737=>"111000010",
  32738=>"110101011",
  32739=>"011011110",
  32740=>"010100110",
  32741=>"110000100",
  32742=>"001100000",
  32743=>"101000001",
  32744=>"101101010",
  32745=>"001001100",
  32746=>"011011110",
  32747=>"000111010",
  32748=>"010011100",
  32749=>"101101110",
  32750=>"110110110",
  32751=>"110111001",
  32752=>"000110011",
  32753=>"100000000",
  32754=>"111001010",
  32755=>"011011001",
  32756=>"110101001",
  32757=>"011110011",
  32758=>"110000001",
  32759=>"000011101",
  32760=>"100110101",
  32761=>"111111101",
  32762=>"101101111",
  32763=>"011011000",
  32764=>"111010000",
  32765=>"100001111",
  32766=>"101011110",
  32767=>"100010001",
  32768=>"000111100",
  32769=>"010011110",
  32770=>"010110010",
  32771=>"111111101",
  32772=>"001101110",
  32773=>"000111100",
  32774=>"010110001",
  32775=>"011001111",
  32776=>"111110110",
  32777=>"000011001",
  32778=>"110011010",
  32779=>"011100100",
  32780=>"011000101",
  32781=>"010010001",
  32782=>"011001111",
  32783=>"011000111",
  32784=>"000000011",
  32785=>"111011100",
  32786=>"000101111",
  32787=>"010010111",
  32788=>"100110111",
  32789=>"010100001",
  32790=>"010101101",
  32791=>"010100110",
  32792=>"010010000",
  32793=>"000011101",
  32794=>"001100011",
  32795=>"011110110",
  32796=>"100000011",
  32797=>"001111000",
  32798=>"101001010",
  32799=>"110110111",
  32800=>"101111001",
  32801=>"111111011",
  32802=>"101010001",
  32803=>"100100011",
  32804=>"000111110",
  32805=>"010110001",
  32806=>"110100000",
  32807=>"110111111",
  32808=>"000110001",
  32809=>"000001110",
  32810=>"011000110",
  32811=>"110001000",
  32812=>"001010111",
  32813=>"000000011",
  32814=>"101000011",
  32815=>"111001100",
  32816=>"111001110",
  32817=>"011011010",
  32818=>"011011110",
  32819=>"111000100",
  32820=>"110000001",
  32821=>"101010110",
  32822=>"111111001",
  32823=>"110011000",
  32824=>"000100000",
  32825=>"100110101",
  32826=>"111001000",
  32827=>"010011111",
  32828=>"000110101",
  32829=>"100111110",
  32830=>"101101111",
  32831=>"001001011",
  32832=>"000001011",
  32833=>"000001000",
  32834=>"011011101",
  32835=>"100010111",
  32836=>"111011110",
  32837=>"000110110",
  32838=>"101001100",
  32839=>"001010011",
  32840=>"000010001",
  32841=>"111111100",
  32842=>"111101111",
  32843=>"101001001",
  32844=>"000000000",
  32845=>"000010100",
  32846=>"010110000",
  32847=>"001000010",
  32848=>"101100111",
  32849=>"000000000",
  32850=>"110011111",
  32851=>"001110000",
  32852=>"000000010",
  32853=>"000100111",
  32854=>"011010001",
  32855=>"001101101",
  32856=>"101110011",
  32857=>"010001011",
  32858=>"010001001",
  32859=>"011101010",
  32860=>"000111010",
  32861=>"101001011",
  32862=>"111010011",
  32863=>"011001001",
  32864=>"001001010",
  32865=>"110001000",
  32866=>"100100011",
  32867=>"111000010",
  32868=>"101001000",
  32869=>"110011101",
  32870=>"101001011",
  32871=>"010011011",
  32872=>"100100011",
  32873=>"101100010",
  32874=>"100010101",
  32875=>"101110110",
  32876=>"011100100",
  32877=>"001110111",
  32878=>"100010000",
  32879=>"000001000",
  32880=>"000111011",
  32881=>"000100110",
  32882=>"101010001",
  32883=>"000111010",
  32884=>"100001111",
  32885=>"101101000",
  32886=>"111000101",
  32887=>"000110100",
  32888=>"010010001",
  32889=>"010000011",
  32890=>"001011101",
  32891=>"100000011",
  32892=>"111111100",
  32893=>"010111011",
  32894=>"010010000",
  32895=>"000110100",
  32896=>"100101011",
  32897=>"101000101",
  32898=>"101011110",
  32899=>"000100001",
  32900=>"001101100",
  32901=>"000111001",
  32902=>"110011111",
  32903=>"100110001",
  32904=>"110000000",
  32905=>"000110010",
  32906=>"111101110",
  32907=>"010110111",
  32908=>"101000101",
  32909=>"100001100",
  32910=>"101001101",
  32911=>"011010111",
  32912=>"101100101",
  32913=>"100100101",
  32914=>"001010010",
  32915=>"000101111",
  32916=>"111100100",
  32917=>"101011011",
  32918=>"110111001",
  32919=>"010011001",
  32920=>"110110001",
  32921=>"001111011",
  32922=>"010100011",
  32923=>"111101001",
  32924=>"001010110",
  32925=>"111001100",
  32926=>"001001000",
  32927=>"010111101",
  32928=>"111111010",
  32929=>"000011100",
  32930=>"001100000",
  32931=>"000110111",
  32932=>"111100111",
  32933=>"100010011",
  32934=>"101000100",
  32935=>"101101111",
  32936=>"111110110",
  32937=>"010110000",
  32938=>"101110010",
  32939=>"000000111",
  32940=>"011011010",
  32941=>"101111111",
  32942=>"000110011",
  32943=>"011010000",
  32944=>"111111111",
  32945=>"000001101",
  32946=>"011101110",
  32947=>"111100000",
  32948=>"010000101",
  32949=>"110111111",
  32950=>"000101011",
  32951=>"011111101",
  32952=>"010100001",
  32953=>"101010011",
  32954=>"010101011",
  32955=>"011001010",
  32956=>"010011010",
  32957=>"001101101",
  32958=>"001011011",
  32959=>"101101111",
  32960=>"111001010",
  32961=>"110101010",
  32962=>"010010000",
  32963=>"100010000",
  32964=>"100001010",
  32965=>"000110101",
  32966=>"101001110",
  32967=>"010111010",
  32968=>"001101111",
  32969=>"101100011",
  32970=>"111000100",
  32971=>"100100100",
  32972=>"100111101",
  32973=>"001110000",
  32974=>"010111111",
  32975=>"011101100",
  32976=>"110110010",
  32977=>"000100010",
  32978=>"101110000",
  32979=>"101111000",
  32980=>"100011111",
  32981=>"011010011",
  32982=>"111000111",
  32983=>"011110010",
  32984=>"111111001",
  32985=>"000000000",
  32986=>"000000101",
  32987=>"000000011",
  32988=>"100111101",
  32989=>"001011010",
  32990=>"111010101",
  32991=>"101101110",
  32992=>"011111001",
  32993=>"000010011",
  32994=>"000100011",
  32995=>"100100011",
  32996=>"001100111",
  32997=>"111110100",
  32998=>"001110010",
  32999=>"000100111",
  33000=>"100100000",
  33001=>"100111111",
  33002=>"110110001",
  33003=>"000110011",
  33004=>"000010100",
  33005=>"010101000",
  33006=>"101011001",
  33007=>"110010000",
  33008=>"110100001",
  33009=>"101111111",
  33010=>"010101010",
  33011=>"100100000",
  33012=>"010010111",
  33013=>"100010111",
  33014=>"011110110",
  33015=>"010100110",
  33016=>"001000010",
  33017=>"000001001",
  33018=>"000001100",
  33019=>"101000111",
  33020=>"110000010",
  33021=>"011110011",
  33022=>"001010001",
  33023=>"110010001",
  33024=>"110101101",
  33025=>"101001011",
  33026=>"100111011",
  33027=>"101001101",
  33028=>"101010000",
  33029=>"011011111",
  33030=>"111101000",
  33031=>"010000100",
  33032=>"000010010",
  33033=>"000000010",
  33034=>"101101000",
  33035=>"001100010",
  33036=>"110000111",
  33037=>"010110111",
  33038=>"010101010",
  33039=>"101001101",
  33040=>"001100100",
  33041=>"011000110",
  33042=>"000100100",
  33043=>"000001101",
  33044=>"010100000",
  33045=>"000010000",
  33046=>"101001110",
  33047=>"100010100",
  33048=>"101000001",
  33049=>"010100011",
  33050=>"000111100",
  33051=>"011000001",
  33052=>"101010000",
  33053=>"110001110",
  33054=>"111010000",
  33055=>"011110000",
  33056=>"111001001",
  33057=>"100010101",
  33058=>"101000000",
  33059=>"100101001",
  33060=>"000101101",
  33061=>"101001011",
  33062=>"010011111",
  33063=>"001000101",
  33064=>"011101011",
  33065=>"110110000",
  33066=>"110010011",
  33067=>"000011100",
  33068=>"110111111",
  33069=>"111100000",
  33070=>"101101100",
  33071=>"101111110",
  33072=>"110011101",
  33073=>"011000000",
  33074=>"010000110",
  33075=>"100111110",
  33076=>"111010100",
  33077=>"100001110",
  33078=>"110101110",
  33079=>"110101000",
  33080=>"101011000",
  33081=>"011000001",
  33082=>"100011000",
  33083=>"111001111",
  33084=>"010101010",
  33085=>"010111000",
  33086=>"010001111",
  33087=>"110010100",
  33088=>"111011111",
  33089=>"011111111",
  33090=>"100110110",
  33091=>"111000010",
  33092=>"101110000",
  33093=>"000010101",
  33094=>"110010111",
  33095=>"010011100",
  33096=>"111010100",
  33097=>"110010011",
  33098=>"010110010",
  33099=>"100010100",
  33100=>"110100111",
  33101=>"001100001",
  33102=>"001001101",
  33103=>"111010001",
  33104=>"011001100",
  33105=>"100111000",
  33106=>"001101000",
  33107=>"111100101",
  33108=>"111110010",
  33109=>"010011111",
  33110=>"110011110",
  33111=>"110100101",
  33112=>"110111000",
  33113=>"111101011",
  33114=>"101000011",
  33115=>"110101111",
  33116=>"001100110",
  33117=>"111111011",
  33118=>"001011001",
  33119=>"001111100",
  33120=>"001111001",
  33121=>"111111011",
  33122=>"001010101",
  33123=>"100001111",
  33124=>"100101010",
  33125=>"010101101",
  33126=>"000000101",
  33127=>"001010010",
  33128=>"010101011",
  33129=>"000010100",
  33130=>"011001101",
  33131=>"100101001",
  33132=>"001001011",
  33133=>"101100010",
  33134=>"110010000",
  33135=>"010001001",
  33136=>"000001000",
  33137=>"000100010",
  33138=>"101100010",
  33139=>"011111001",
  33140=>"001010001",
  33141=>"011100001",
  33142=>"001101101",
  33143=>"011101000",
  33144=>"111101011",
  33145=>"001000111",
  33146=>"010111000",
  33147=>"011111000",
  33148=>"101110111",
  33149=>"111111111",
  33150=>"111111000",
  33151=>"000101100",
  33152=>"100111100",
  33153=>"111000011",
  33154=>"011000100",
  33155=>"111011101",
  33156=>"101010100",
  33157=>"101101110",
  33158=>"110100101",
  33159=>"100010101",
  33160=>"110010001",
  33161=>"101010011",
  33162=>"010000100",
  33163=>"111111110",
  33164=>"001111111",
  33165=>"101100110",
  33166=>"000000000",
  33167=>"110010110",
  33168=>"110110101",
  33169=>"010111000",
  33170=>"111010010",
  33171=>"100111100",
  33172=>"000010100",
  33173=>"010110010",
  33174=>"101110110",
  33175=>"010111000",
  33176=>"111000111",
  33177=>"000011111",
  33178=>"011000110",
  33179=>"000110001",
  33180=>"110000100",
  33181=>"001101111",
  33182=>"001111011",
  33183=>"100010010",
  33184=>"010001000",
  33185=>"101101001",
  33186=>"010110111",
  33187=>"011000100",
  33188=>"100101110",
  33189=>"000101100",
  33190=>"101100001",
  33191=>"010010101",
  33192=>"000010100",
  33193=>"011111111",
  33194=>"101001000",
  33195=>"101101010",
  33196=>"111111010",
  33197=>"010000000",
  33198=>"101011110",
  33199=>"011100000",
  33200=>"101001011",
  33201=>"111101101",
  33202=>"101110101",
  33203=>"011010100",
  33204=>"111111111",
  33205=>"110100011",
  33206=>"100100011",
  33207=>"110011010",
  33208=>"100001101",
  33209=>"011001000",
  33210=>"111101011",
  33211=>"110011101",
  33212=>"000001100",
  33213=>"110011110",
  33214=>"111001100",
  33215=>"011000001",
  33216=>"001011010",
  33217=>"010010000",
  33218=>"111001000",
  33219=>"011001001",
  33220=>"111000101",
  33221=>"111000111",
  33222=>"110101111",
  33223=>"001100000",
  33224=>"100001000",
  33225=>"000100010",
  33226=>"110000110",
  33227=>"000011001",
  33228=>"110011110",
  33229=>"111101100",
  33230=>"111001001",
  33231=>"101100001",
  33232=>"000010101",
  33233=>"101010110",
  33234=>"100010011",
  33235=>"101100101",
  33236=>"100110000",
  33237=>"010000000",
  33238=>"000011000",
  33239=>"001100010",
  33240=>"111100010",
  33241=>"111111101",
  33242=>"100000100",
  33243=>"000100100",
  33244=>"001011101",
  33245=>"001011000",
  33246=>"011100011",
  33247=>"011110110",
  33248=>"100011001",
  33249=>"101010001",
  33250=>"111101110",
  33251=>"000001001",
  33252=>"011110011",
  33253=>"100100010",
  33254=>"100011110",
  33255=>"000000001",
  33256=>"011010100",
  33257=>"011111111",
  33258=>"000110001",
  33259=>"100011100",
  33260=>"011000110",
  33261=>"111100010",
  33262=>"001010010",
  33263=>"110111001",
  33264=>"110110100",
  33265=>"000110111",
  33266=>"111100100",
  33267=>"110110011",
  33268=>"000010000",
  33269=>"111010001",
  33270=>"110110001",
  33271=>"010011000",
  33272=>"101111100",
  33273=>"111010011",
  33274=>"110001101",
  33275=>"001101100",
  33276=>"011010100",
  33277=>"011001010",
  33278=>"001011110",
  33279=>"000000011",
  33280=>"011010011",
  33281=>"101100111",
  33282=>"101100010",
  33283=>"010110101",
  33284=>"100101000",
  33285=>"011000100",
  33286=>"110100010",
  33287=>"000100001",
  33288=>"000011111",
  33289=>"110010100",
  33290=>"111110001",
  33291=>"001000001",
  33292=>"001001000",
  33293=>"001110110",
  33294=>"000001011",
  33295=>"010010100",
  33296=>"111001011",
  33297=>"010111010",
  33298=>"000101100",
  33299=>"001010110",
  33300=>"011001000",
  33301=>"000100101",
  33302=>"001100001",
  33303=>"111101100",
  33304=>"010110011",
  33305=>"000010011",
  33306=>"000001001",
  33307=>"110101001",
  33308=>"100001100",
  33309=>"110011001",
  33310=>"101111111",
  33311=>"001011000",
  33312=>"111000010",
  33313=>"100010100",
  33314=>"000100110",
  33315=>"010011011",
  33316=>"000100110",
  33317=>"011111110",
  33318=>"001000110",
  33319=>"010100011",
  33320=>"001010000",
  33321=>"100010111",
  33322=>"000110110",
  33323=>"100101011",
  33324=>"110011110",
  33325=>"000100000",
  33326=>"010000101",
  33327=>"111111010",
  33328=>"111110111",
  33329=>"111011101",
  33330=>"101110011",
  33331=>"111100110",
  33332=>"011001001",
  33333=>"110010111",
  33334=>"010000110",
  33335=>"001011111",
  33336=>"010001011",
  33337=>"111010011",
  33338=>"110110001",
  33339=>"000011011",
  33340=>"100010000",
  33341=>"000001011",
  33342=>"110000101",
  33343=>"111000010",
  33344=>"100010010",
  33345=>"110110101",
  33346=>"000001110",
  33347=>"010010001",
  33348=>"111001110",
  33349=>"011111111",
  33350=>"010111111",
  33351=>"101111011",
  33352=>"011110100",
  33353=>"000111001",
  33354=>"101111010",
  33355=>"101100001",
  33356=>"100011001",
  33357=>"100100010",
  33358=>"101110111",
  33359=>"101011000",
  33360=>"001110010",
  33361=>"000110000",
  33362=>"001110111",
  33363=>"100011111",
  33364=>"110001010",
  33365=>"000000110",
  33366=>"110101000",
  33367=>"101101101",
  33368=>"111000100",
  33369=>"000101100",
  33370=>"101001111",
  33371=>"001000011",
  33372=>"001010000",
  33373=>"001010111",
  33374=>"001010001",
  33375=>"100001011",
  33376=>"110010101",
  33377=>"111001110",
  33378=>"001110001",
  33379=>"010011111",
  33380=>"101101010",
  33381=>"111010011",
  33382=>"010100101",
  33383=>"111101100",
  33384=>"000000010",
  33385=>"011011111",
  33386=>"110111000",
  33387=>"000111100",
  33388=>"001000110",
  33389=>"100001000",
  33390=>"000001010",
  33391=>"011101101",
  33392=>"000111101",
  33393=>"111110000",
  33394=>"110100010",
  33395=>"101001111",
  33396=>"010000101",
  33397=>"100001110",
  33398=>"111011001",
  33399=>"111010111",
  33400=>"011011000",
  33401=>"001111111",
  33402=>"000011101",
  33403=>"101011001",
  33404=>"111001000",
  33405=>"100101100",
  33406=>"100101100",
  33407=>"011111110",
  33408=>"111111000",
  33409=>"001101111",
  33410=>"000100101",
  33411=>"110100001",
  33412=>"100010001",
  33413=>"001010111",
  33414=>"110000101",
  33415=>"101000100",
  33416=>"010100001",
  33417=>"111000000",
  33418=>"100011000",
  33419=>"110110010",
  33420=>"101111011",
  33421=>"001100001",
  33422=>"010000000",
  33423=>"111011001",
  33424=>"111011110",
  33425=>"001001000",
  33426=>"111110111",
  33427=>"010011100",
  33428=>"100100001",
  33429=>"011000101",
  33430=>"010000010",
  33431=>"100000010",
  33432=>"101000101",
  33433=>"001010111",
  33434=>"111000010",
  33435=>"110010111",
  33436=>"111010101",
  33437=>"010101000",
  33438=>"010011011",
  33439=>"000101111",
  33440=>"111110101",
  33441=>"110011111",
  33442=>"010101100",
  33443=>"100001011",
  33444=>"010100111",
  33445=>"111111101",
  33446=>"011001010",
  33447=>"001100001",
  33448=>"001101000",
  33449=>"010110101",
  33450=>"101101100",
  33451=>"100001010",
  33452=>"010000000",
  33453=>"000010111",
  33454=>"101010100",
  33455=>"111111111",
  33456=>"011111100",
  33457=>"001111101",
  33458=>"011010110",
  33459=>"010001001",
  33460=>"111011111",
  33461=>"011011010",
  33462=>"110100111",
  33463=>"101110110",
  33464=>"011000100",
  33465=>"111001001",
  33466=>"100000110",
  33467=>"000010011",
  33468=>"111111111",
  33469=>"100010111",
  33470=>"000000110",
  33471=>"100011110",
  33472=>"000000000",
  33473=>"100001101",
  33474=>"001001001",
  33475=>"001100100",
  33476=>"011011011",
  33477=>"111101011",
  33478=>"101111100",
  33479=>"101010110",
  33480=>"001000001",
  33481=>"110011001",
  33482=>"000000100",
  33483=>"011001000",
  33484=>"001010000",
  33485=>"110111101",
  33486=>"011001010",
  33487=>"000111010",
  33488=>"100111011",
  33489=>"000010101",
  33490=>"111111011",
  33491=>"100110110",
  33492=>"101111010",
  33493=>"101110111",
  33494=>"011111000",
  33495=>"001111010",
  33496=>"101000111",
  33497=>"100011111",
  33498=>"000110111",
  33499=>"111000000",
  33500=>"101010001",
  33501=>"000101011",
  33502=>"100101111",
  33503=>"101011111",
  33504=>"001001101",
  33505=>"011000100",
  33506=>"101111111",
  33507=>"111100110",
  33508=>"011110111",
  33509=>"000100010",
  33510=>"110000011",
  33511=>"001001001",
  33512=>"010001001",
  33513=>"011000111",
  33514=>"100011000",
  33515=>"011010100",
  33516=>"001011011",
  33517=>"100011100",
  33518=>"000001111",
  33519=>"110000010",
  33520=>"001011001",
  33521=>"111111000",
  33522=>"011111010",
  33523=>"111101111",
  33524=>"111000001",
  33525=>"011010101",
  33526=>"000000000",
  33527=>"010111100",
  33528=>"101101101",
  33529=>"010111000",
  33530=>"000100100",
  33531=>"100010010",
  33532=>"001001100",
  33533=>"101110011",
  33534=>"110101110",
  33535=>"011110011",
  33536=>"111000000",
  33537=>"010010011",
  33538=>"111110101",
  33539=>"011110111",
  33540=>"010100001",
  33541=>"111000101",
  33542=>"000101100",
  33543=>"111101000",
  33544=>"000010000",
  33545=>"010011111",
  33546=>"001101100",
  33547=>"101100000",
  33548=>"000011001",
  33549=>"110001010",
  33550=>"100010001",
  33551=>"010111111",
  33552=>"101011100",
  33553=>"001100110",
  33554=>"011100100",
  33555=>"011000010",
  33556=>"100011100",
  33557=>"000000101",
  33558=>"011001101",
  33559=>"000001001",
  33560=>"000000100",
  33561=>"000101111",
  33562=>"011010110",
  33563=>"100111110",
  33564=>"111011010",
  33565=>"010101110",
  33566=>"010100000",
  33567=>"111111010",
  33568=>"111100101",
  33569=>"100001000",
  33570=>"110101100",
  33571=>"000000010",
  33572=>"110000111",
  33573=>"000000001",
  33574=>"011100100",
  33575=>"010010100",
  33576=>"011111011",
  33577=>"000101110",
  33578=>"000110000",
  33579=>"000101101",
  33580=>"001011010",
  33581=>"111111111",
  33582=>"010000111",
  33583=>"110111111",
  33584=>"000011011",
  33585=>"100010101",
  33586=>"011010110",
  33587=>"111001001",
  33588=>"111111111",
  33589=>"011011100",
  33590=>"011011111",
  33591=>"100100001",
  33592=>"000101001",
  33593=>"100101111",
  33594=>"000000111",
  33595=>"100000111",
  33596=>"101100101",
  33597=>"100011001",
  33598=>"111001110",
  33599=>"010111011",
  33600=>"100110100",
  33601=>"010001100",
  33602=>"101100011",
  33603=>"101111101",
  33604=>"010001101",
  33605=>"100010111",
  33606=>"100110000",
  33607=>"111011101",
  33608=>"010010000",
  33609=>"100010010",
  33610=>"010011011",
  33611=>"100000011",
  33612=>"110110110",
  33613=>"001001111",
  33614=>"010011010",
  33615=>"000110001",
  33616=>"101000001",
  33617=>"100010101",
  33618=>"001001100",
  33619=>"011000101",
  33620=>"001100000",
  33621=>"010010000",
  33622=>"101000000",
  33623=>"001100100",
  33624=>"100010100",
  33625=>"000000111",
  33626=>"111110111",
  33627=>"001100000",
  33628=>"111110011",
  33629=>"101010010",
  33630=>"100111111",
  33631=>"101111110",
  33632=>"101110010",
  33633=>"111111101",
  33634=>"111101101",
  33635=>"011111101",
  33636=>"101111101",
  33637=>"101010000",
  33638=>"000111000",
  33639=>"111001000",
  33640=>"101111011",
  33641=>"000110111",
  33642=>"011100000",
  33643=>"011110000",
  33644=>"010110100",
  33645=>"111101100",
  33646=>"011110001",
  33647=>"100101101",
  33648=>"000000001",
  33649=>"111111000",
  33650=>"111100001",
  33651=>"111100111",
  33652=>"110001001",
  33653=>"111111000",
  33654=>"110110101",
  33655=>"011111000",
  33656=>"111011001",
  33657=>"110011000",
  33658=>"111101100",
  33659=>"001110101",
  33660=>"101100101",
  33661=>"111101001",
  33662=>"101011001",
  33663=>"011000001",
  33664=>"100011010",
  33665=>"100000001",
  33666=>"000010111",
  33667=>"011110101",
  33668=>"111110000",
  33669=>"110011110",
  33670=>"100110010",
  33671=>"111100100",
  33672=>"001011011",
  33673=>"010010101",
  33674=>"111000011",
  33675=>"111111101",
  33676=>"111011100",
  33677=>"100100010",
  33678=>"011111101",
  33679=>"001101111",
  33680=>"000001101",
  33681=>"111111011",
  33682=>"000100000",
  33683=>"011100011",
  33684=>"011000101",
  33685=>"010011000",
  33686=>"010000010",
  33687=>"111001000",
  33688=>"101110011",
  33689=>"000110000",
  33690=>"111011011",
  33691=>"110100101",
  33692=>"100110110",
  33693=>"100110100",
  33694=>"000100101",
  33695=>"001001111",
  33696=>"011101001",
  33697=>"000110001",
  33698=>"001010111",
  33699=>"000010001",
  33700=>"010111111",
  33701=>"011100001",
  33702=>"111011101",
  33703=>"100111011",
  33704=>"000010011",
  33705=>"000001100",
  33706=>"101000111",
  33707=>"010010110",
  33708=>"000100000",
  33709=>"011000010",
  33710=>"000111101",
  33711=>"000000101",
  33712=>"011100101",
  33713=>"110011001",
  33714=>"100010101",
  33715=>"000000110",
  33716=>"111000100",
  33717=>"111100100",
  33718=>"010001101",
  33719=>"111010000",
  33720=>"110110111",
  33721=>"001111001",
  33722=>"111111110",
  33723=>"010010110",
  33724=>"101010001",
  33725=>"101101010",
  33726=>"100011011",
  33727=>"000100010",
  33728=>"011000000",
  33729=>"000000001",
  33730=>"011100001",
  33731=>"110000111",
  33732=>"001000010",
  33733=>"101110010",
  33734=>"010101000",
  33735=>"001000011",
  33736=>"010100111",
  33737=>"001011000",
  33738=>"010011011",
  33739=>"011000010",
  33740=>"110110011",
  33741=>"000001110",
  33742=>"010110001",
  33743=>"011010001",
  33744=>"111011111",
  33745=>"010010101",
  33746=>"011101101",
  33747=>"100011000",
  33748=>"010000111",
  33749=>"100101100",
  33750=>"010111001",
  33751=>"101111001",
  33752=>"000010101",
  33753=>"010000101",
  33754=>"001100000",
  33755=>"011011110",
  33756=>"101111110",
  33757=>"100100000",
  33758=>"110101000",
  33759=>"011101100",
  33760=>"100101110",
  33761=>"000100100",
  33762=>"000101000",
  33763=>"111010001",
  33764=>"110111001",
  33765=>"001000100",
  33766=>"100001001",
  33767=>"010101101",
  33768=>"000001110",
  33769=>"110101101",
  33770=>"111111101",
  33771=>"100111111",
  33772=>"000011000",
  33773=>"101100100",
  33774=>"111111110",
  33775=>"111110000",
  33776=>"111010100",
  33777=>"100000010",
  33778=>"000100000",
  33779=>"101100101",
  33780=>"111110011",
  33781=>"101100001",
  33782=>"100100000",
  33783=>"010000001",
  33784=>"100001010",
  33785=>"101110110",
  33786=>"101011011",
  33787=>"000011101",
  33788=>"101001011",
  33789=>"000100101",
  33790=>"011001001",
  33791=>"010000100",
  33792=>"110011011",
  33793=>"100011000",
  33794=>"001001000",
  33795=>"101010010",
  33796=>"101100010",
  33797=>"000001110",
  33798=>"111001101",
  33799=>"011010010",
  33800=>"110010000",
  33801=>"111010110",
  33802=>"111101000",
  33803=>"011011111",
  33804=>"001111000",
  33805=>"010110110",
  33806=>"011100100",
  33807=>"001101111",
  33808=>"001101000",
  33809=>"110101110",
  33810=>"010000001",
  33811=>"111101110",
  33812=>"000110110",
  33813=>"100100000",
  33814=>"000001100",
  33815=>"110100000",
  33816=>"011000100",
  33817=>"101110011",
  33818=>"011011000",
  33819=>"110111100",
  33820=>"110011110",
  33821=>"011111000",
  33822=>"001010010",
  33823=>"100000001",
  33824=>"100101101",
  33825=>"101000010",
  33826=>"011010111",
  33827=>"000111010",
  33828=>"000101100",
  33829=>"111111110",
  33830=>"010110101",
  33831=>"011010111",
  33832=>"011111000",
  33833=>"100001010",
  33834=>"011011000",
  33835=>"010001110",
  33836=>"001111101",
  33837=>"111100110",
  33838=>"010100101",
  33839=>"000100000",
  33840=>"000011001",
  33841=>"111101111",
  33842=>"000110111",
  33843=>"101111000",
  33844=>"001111001",
  33845=>"001011001",
  33846=>"010111100",
  33847=>"011111111",
  33848=>"001000000",
  33849=>"101000001",
  33850=>"010000011",
  33851=>"000111101",
  33852=>"011101000",
  33853=>"110111010",
  33854=>"011110011",
  33855=>"110111001",
  33856=>"111000000",
  33857=>"001001011",
  33858=>"000011001",
  33859=>"010011010",
  33860=>"100100110",
  33861=>"011111001",
  33862=>"010111111",
  33863=>"101111111",
  33864=>"000100000",
  33865=>"011110101",
  33866=>"101111001",
  33867=>"101111000",
  33868=>"011000111",
  33869=>"111111000",
  33870=>"011101000",
  33871=>"010110010",
  33872=>"100001001",
  33873=>"000110010",
  33874=>"010101111",
  33875=>"100111001",
  33876=>"001100010",
  33877=>"010100111",
  33878=>"111001001",
  33879=>"111110110",
  33880=>"010010111",
  33881=>"110101001",
  33882=>"010011000",
  33883=>"010110011",
  33884=>"011010101",
  33885=>"011011000",
  33886=>"000001100",
  33887=>"000000111",
  33888=>"000111010",
  33889=>"001001000",
  33890=>"000111110",
  33891=>"111111000",
  33892=>"101011011",
  33893=>"100011110",
  33894=>"000001000",
  33895=>"000110001",
  33896=>"001000101",
  33897=>"101001010",
  33898=>"100010100",
  33899=>"110001000",
  33900=>"000110011",
  33901=>"001001000",
  33902=>"101111000",
  33903=>"000001101",
  33904=>"000010101",
  33905=>"110000101",
  33906=>"101000110",
  33907=>"000101011",
  33908=>"110100101",
  33909=>"101101100",
  33910=>"111101001",
  33911=>"110001000",
  33912=>"111101111",
  33913=>"010001000",
  33914=>"100101110",
  33915=>"110110010",
  33916=>"001101010",
  33917=>"110010001",
  33918=>"010111101",
  33919=>"111011001",
  33920=>"111111010",
  33921=>"010000111",
  33922=>"000111001",
  33923=>"100101110",
  33924=>"111000110",
  33925=>"001010110",
  33926=>"010111110",
  33927=>"101000111",
  33928=>"010101110",
  33929=>"101101101",
  33930=>"110110011",
  33931=>"101011110",
  33932=>"001001000",
  33933=>"100010110",
  33934=>"101110110",
  33935=>"110101100",
  33936=>"000000101",
  33937=>"111011011",
  33938=>"000110110",
  33939=>"000010111",
  33940=>"001101000",
  33941=>"001010100",
  33942=>"101010010",
  33943=>"000101110",
  33944=>"011110101",
  33945=>"100100111",
  33946=>"101100000",
  33947=>"111101001",
  33948=>"010011100",
  33949=>"001011110",
  33950=>"110110101",
  33951=>"010101010",
  33952=>"110100100",
  33953=>"001001100",
  33954=>"011001000",
  33955=>"000110110",
  33956=>"101100100",
  33957=>"111101101",
  33958=>"101000000",
  33959=>"001111000",
  33960=>"110000101",
  33961=>"111010010",
  33962=>"010000000",
  33963=>"110011111",
  33964=>"011101110",
  33965=>"010110111",
  33966=>"111010000",
  33967=>"110101100",
  33968=>"000001110",
  33969=>"001101110",
  33970=>"010010001",
  33971=>"011101100",
  33972=>"111100101",
  33973=>"000110111",
  33974=>"100010010",
  33975=>"001011010",
  33976=>"111101110",
  33977=>"100110000",
  33978=>"111100110",
  33979=>"101101111",
  33980=>"011111011",
  33981=>"100010000",
  33982=>"001010000",
  33983=>"110101001",
  33984=>"000100001",
  33985=>"001011010",
  33986=>"000100100",
  33987=>"111110110",
  33988=>"100111100",
  33989=>"001111111",
  33990=>"100010010",
  33991=>"010110001",
  33992=>"011100010",
  33993=>"011010111",
  33994=>"001100011",
  33995=>"000000000",
  33996=>"101111010",
  33997=>"100010111",
  33998=>"111101100",
  33999=>"110101100",
  34000=>"110101010",
  34001=>"000001110",
  34002=>"111000011",
  34003=>"011101111",
  34004=>"010101110",
  34005=>"110101111",
  34006=>"110111101",
  34007=>"001001110",
  34008=>"011100101",
  34009=>"110011111",
  34010=>"001111100",
  34011=>"010100011",
  34012=>"011011011",
  34013=>"100101001",
  34014=>"011100111",
  34015=>"011100001",
  34016=>"001001010",
  34017=>"001011100",
  34018=>"001001111",
  34019=>"111110001",
  34020=>"011111111",
  34021=>"011000101",
  34022=>"010010010",
  34023=>"010001111",
  34024=>"101000001",
  34025=>"101010111",
  34026=>"010000001",
  34027=>"000110001",
  34028=>"110010101",
  34029=>"000000100",
  34030=>"000110100",
  34031=>"010011111",
  34032=>"110100010",
  34033=>"000001110",
  34034=>"011000101",
  34035=>"111011000",
  34036=>"111111111",
  34037=>"111110100",
  34038=>"110100111",
  34039=>"000000000",
  34040=>"100111111",
  34041=>"101100101",
  34042=>"010110100",
  34043=>"010110100",
  34044=>"001010101",
  34045=>"001111000",
  34046=>"101110001",
  34047=>"100111101",
  34048=>"010101010",
  34049=>"000111110",
  34050=>"001111011",
  34051=>"111111111",
  34052=>"110101101",
  34053=>"010111110",
  34054=>"010111100",
  34055=>"111001010",
  34056=>"111000100",
  34057=>"001101100",
  34058=>"111011101",
  34059=>"101011000",
  34060=>"111101110",
  34061=>"110001110",
  34062=>"111101001",
  34063=>"011111011",
  34064=>"111100000",
  34065=>"011110000",
  34066=>"000000010",
  34067=>"111110111",
  34068=>"010010111",
  34069=>"101111011",
  34070=>"000010000",
  34071=>"110011101",
  34072=>"101101001",
  34073=>"100110101",
  34074=>"110000010",
  34075=>"010010111",
  34076=>"010010100",
  34077=>"001011101",
  34078=>"101010111",
  34079=>"110100001",
  34080=>"000110100",
  34081=>"010100111",
  34082=>"001000011",
  34083=>"110111110",
  34084=>"001000101",
  34085=>"001101000",
  34086=>"111000010",
  34087=>"111010101",
  34088=>"001101010",
  34089=>"000100011",
  34090=>"100000011",
  34091=>"000100101",
  34092=>"111111000",
  34093=>"011001000",
  34094=>"100001101",
  34095=>"110001100",
  34096=>"101110111",
  34097=>"101110000",
  34098=>"111111100",
  34099=>"010111111",
  34100=>"100001011",
  34101=>"011111111",
  34102=>"010000100",
  34103=>"011000110",
  34104=>"001111111",
  34105=>"001101010",
  34106=>"000111000",
  34107=>"011010000",
  34108=>"001101111",
  34109=>"111001011",
  34110=>"001000110",
  34111=>"001111110",
  34112=>"001001110",
  34113=>"010110100",
  34114=>"000010001",
  34115=>"100111110",
  34116=>"100010010",
  34117=>"000101010",
  34118=>"110001101",
  34119=>"110101000",
  34120=>"110101001",
  34121=>"101010001",
  34122=>"000111000",
  34123=>"111000010",
  34124=>"100101101",
  34125=>"110110000",
  34126=>"100100000",
  34127=>"010110010",
  34128=>"101100101",
  34129=>"100001101",
  34130=>"100110010",
  34131=>"010111010",
  34132=>"000001111",
  34133=>"011010110",
  34134=>"011101111",
  34135=>"000011100",
  34136=>"000000110",
  34137=>"111001111",
  34138=>"100011111",
  34139=>"110110011",
  34140=>"111011111",
  34141=>"000001110",
  34142=>"110111101",
  34143=>"000111110",
  34144=>"010001101",
  34145=>"101110011",
  34146=>"100000101",
  34147=>"100000010",
  34148=>"101101101",
  34149=>"100101111",
  34150=>"010101010",
  34151=>"011111001",
  34152=>"001100010",
  34153=>"110110010",
  34154=>"110101111",
  34155=>"011111101",
  34156=>"111000110",
  34157=>"111010010",
  34158=>"011111110",
  34159=>"001101010",
  34160=>"111111010",
  34161=>"101000000",
  34162=>"111010111",
  34163=>"101110001",
  34164=>"011011010",
  34165=>"100110110",
  34166=>"111001010",
  34167=>"001001011",
  34168=>"101001111",
  34169=>"111010101",
  34170=>"101010100",
  34171=>"100001111",
  34172=>"000101100",
  34173=>"001111101",
  34174=>"101010011",
  34175=>"101010100",
  34176=>"100001110",
  34177=>"010100101",
  34178=>"101000011",
  34179=>"101111010",
  34180=>"100100011",
  34181=>"101100100",
  34182=>"111001011",
  34183=>"010010010",
  34184=>"010010101",
  34185=>"101010000",
  34186=>"100100101",
  34187=>"011001100",
  34188=>"101001000",
  34189=>"001001010",
  34190=>"010010101",
  34191=>"001010010",
  34192=>"111000101",
  34193=>"000000000",
  34194=>"100111000",
  34195=>"001110001",
  34196=>"101100010",
  34197=>"010111111",
  34198=>"010000010",
  34199=>"101011000",
  34200=>"011111001",
  34201=>"000111000",
  34202=>"010110010",
  34203=>"101000100",
  34204=>"111001001",
  34205=>"001111100",
  34206=>"101001100",
  34207=>"101100001",
  34208=>"011111100",
  34209=>"010111011",
  34210=>"000111011",
  34211=>"100001001",
  34212=>"111101010",
  34213=>"000000110",
  34214=>"101010101",
  34215=>"111111110",
  34216=>"010100110",
  34217=>"010100001",
  34218=>"000000011",
  34219=>"000011000",
  34220=>"001111110",
  34221=>"101111000",
  34222=>"001010010",
  34223=>"001010000",
  34224=>"110011110",
  34225=>"101100101",
  34226=>"011001001",
  34227=>"110011011",
  34228=>"001110011",
  34229=>"100000110",
  34230=>"001010011",
  34231=>"000011101",
  34232=>"000101101",
  34233=>"001010111",
  34234=>"111010111",
  34235=>"011111111",
  34236=>"010010110",
  34237=>"111100110",
  34238=>"000100110",
  34239=>"101010011",
  34240=>"111110001",
  34241=>"100001001",
  34242=>"101110111",
  34243=>"111110101",
  34244=>"111011110",
  34245=>"010001110",
  34246=>"101101000",
  34247=>"001110100",
  34248=>"100011111",
  34249=>"101000111",
  34250=>"000100110",
  34251=>"000001101",
  34252=>"010011111",
  34253=>"101111100",
  34254=>"100101011",
  34255=>"101110011",
  34256=>"101001011",
  34257=>"110010101",
  34258=>"110001001",
  34259=>"110100011",
  34260=>"101000001",
  34261=>"011001011",
  34262=>"010111101",
  34263=>"101101001",
  34264=>"111000001",
  34265=>"100100111",
  34266=>"110010100",
  34267=>"011101101",
  34268=>"110001100",
  34269=>"100101100",
  34270=>"000111101",
  34271=>"010111100",
  34272=>"110110111",
  34273=>"000000110",
  34274=>"000010011",
  34275=>"011101110",
  34276=>"001111100",
  34277=>"010000101",
  34278=>"100111101",
  34279=>"011110111",
  34280=>"101111111",
  34281=>"010000101",
  34282=>"110101001",
  34283=>"011111101",
  34284=>"001111010",
  34285=>"111101010",
  34286=>"110111111",
  34287=>"101000001",
  34288=>"011100010",
  34289=>"100011011",
  34290=>"010111010",
  34291=>"111000110",
  34292=>"011011000",
  34293=>"101000110",
  34294=>"001011101",
  34295=>"111011100",
  34296=>"110001110",
  34297=>"000000010",
  34298=>"100000100",
  34299=>"001100011",
  34300=>"100000000",
  34301=>"011101110",
  34302=>"010001011",
  34303=>"101100000",
  34304=>"101001101",
  34305=>"101100010",
  34306=>"110010001",
  34307=>"011101110",
  34308=>"001001010",
  34309=>"000010110",
  34310=>"010000011",
  34311=>"110001101",
  34312=>"001101000",
  34313=>"010000100",
  34314=>"110111111",
  34315=>"000000000",
  34316=>"000010100",
  34317=>"111111111",
  34318=>"000010000",
  34319=>"100101010",
  34320=>"111000001",
  34321=>"101110110",
  34322=>"100111110",
  34323=>"100011100",
  34324=>"100100010",
  34325=>"111000101",
  34326=>"100110100",
  34327=>"110111101",
  34328=>"010010010",
  34329=>"001001111",
  34330=>"111000100",
  34331=>"010000101",
  34332=>"111011011",
  34333=>"001100111",
  34334=>"001011101",
  34335=>"100111111",
  34336=>"000111000",
  34337=>"101100110",
  34338=>"100100100",
  34339=>"111000100",
  34340=>"011110101",
  34341=>"100101011",
  34342=>"001011010",
  34343=>"000011000",
  34344=>"011111100",
  34345=>"110011000",
  34346=>"101111000",
  34347=>"111011000",
  34348=>"101010100",
  34349=>"101001101",
  34350=>"100001000",
  34351=>"100011011",
  34352=>"101101000",
  34353=>"000001000",
  34354=>"001100111",
  34355=>"011100001",
  34356=>"001010110",
  34357=>"101000111",
  34358=>"100110001",
  34359=>"111110100",
  34360=>"100001101",
  34361=>"110110010",
  34362=>"001100001",
  34363=>"110110111",
  34364=>"001101001",
  34365=>"000101000",
  34366=>"010010001",
  34367=>"100011000",
  34368=>"010110001",
  34369=>"101111010",
  34370=>"000101010",
  34371=>"011010011",
  34372=>"101000000",
  34373=>"001010000",
  34374=>"011011101",
  34375=>"011111101",
  34376=>"000010011",
  34377=>"111111111",
  34378=>"011010111",
  34379=>"100111110",
  34380=>"100111110",
  34381=>"100111001",
  34382=>"000010001",
  34383=>"111010011",
  34384=>"000000000",
  34385=>"001011101",
  34386=>"111101111",
  34387=>"000000111",
  34388=>"010101111",
  34389=>"001100111",
  34390=>"000100001",
  34391=>"100000001",
  34392=>"000110011",
  34393=>"001110110",
  34394=>"010110101",
  34395=>"011110100",
  34396=>"001010101",
  34397=>"100100010",
  34398=>"110111011",
  34399=>"100011011",
  34400=>"001101001",
  34401=>"101100110",
  34402=>"101100100",
  34403=>"101010110",
  34404=>"110100100",
  34405=>"010111111",
  34406=>"110101110",
  34407=>"101001100",
  34408=>"110011111",
  34409=>"001000100",
  34410=>"011110101",
  34411=>"011011000",
  34412=>"010000110",
  34413=>"100011011",
  34414=>"001011001",
  34415=>"011110111",
  34416=>"100000010",
  34417=>"011100010",
  34418=>"001101011",
  34419=>"110001000",
  34420=>"111111111",
  34421=>"101001101",
  34422=>"001100001",
  34423=>"111000000",
  34424=>"010010011",
  34425=>"101110000",
  34426=>"001000101",
  34427=>"111100100",
  34428=>"001100101",
  34429=>"000111111",
  34430=>"011100100",
  34431=>"001101101",
  34432=>"101110100",
  34433=>"000000101",
  34434=>"101101110",
  34435=>"001001011",
  34436=>"000110111",
  34437=>"101010010",
  34438=>"111011111",
  34439=>"111000010",
  34440=>"111011111",
  34441=>"010010011",
  34442=>"101101001",
  34443=>"111110111",
  34444=>"111011111",
  34445=>"010110010",
  34446=>"001000110",
  34447=>"001001011",
  34448=>"110010111",
  34449=>"111011100",
  34450=>"111100101",
  34451=>"100100010",
  34452=>"010111010",
  34453=>"000000001",
  34454=>"000010111",
  34455=>"011010010",
  34456=>"000101011",
  34457=>"110001000",
  34458=>"000001110",
  34459=>"000100111",
  34460=>"011000001",
  34461=>"010111111",
  34462=>"010110100",
  34463=>"001011110",
  34464=>"000100001",
  34465=>"000110010",
  34466=>"111101000",
  34467=>"010001100",
  34468=>"100111111",
  34469=>"000110011",
  34470=>"010001101",
  34471=>"011110101",
  34472=>"100111011",
  34473=>"001001001",
  34474=>"100010000",
  34475=>"100010000",
  34476=>"000110110",
  34477=>"111000111",
  34478=>"100110001",
  34479=>"100111100",
  34480=>"010110011",
  34481=>"000001010",
  34482=>"110110111",
  34483=>"001011100",
  34484=>"101010100",
  34485=>"011001101",
  34486=>"100001010",
  34487=>"110101010",
  34488=>"010101000",
  34489=>"010100001",
  34490=>"111000111",
  34491=>"001010101",
  34492=>"111101000",
  34493=>"101100000",
  34494=>"110111001",
  34495=>"100110010",
  34496=>"001010110",
  34497=>"101111101",
  34498=>"111011000",
  34499=>"110111100",
  34500=>"111111101",
  34501=>"011111110",
  34502=>"001100001",
  34503=>"011101001",
  34504=>"001101100",
  34505=>"110100101",
  34506=>"100111100",
  34507=>"011101100",
  34508=>"111011001",
  34509=>"111000011",
  34510=>"000110010",
  34511=>"010100000",
  34512=>"111101101",
  34513=>"111110000",
  34514=>"011100111",
  34515=>"101000001",
  34516=>"111100100",
  34517=>"101011100",
  34518=>"011111101",
  34519=>"001001110",
  34520=>"011110111",
  34521=>"110001101",
  34522=>"110100101",
  34523=>"101010111",
  34524=>"111000000",
  34525=>"111010001",
  34526=>"110011010",
  34527=>"100011100",
  34528=>"010101100",
  34529=>"001100110",
  34530=>"010100110",
  34531=>"011001111",
  34532=>"010111111",
  34533=>"011101110",
  34534=>"011111001",
  34535=>"010101101",
  34536=>"010000111",
  34537=>"100111101",
  34538=>"010010000",
  34539=>"101111111",
  34540=>"110101000",
  34541=>"011111101",
  34542=>"101011000",
  34543=>"000011100",
  34544=>"110111110",
  34545=>"001101010",
  34546=>"010100111",
  34547=>"000011111",
  34548=>"010111010",
  34549=>"111001111",
  34550=>"100111101",
  34551=>"100011101",
  34552=>"010011110",
  34553=>"001100000",
  34554=>"100011101",
  34555=>"010111110",
  34556=>"110100111",
  34557=>"111011000",
  34558=>"011100110",
  34559=>"110101100",
  34560=>"010010110",
  34561=>"110001010",
  34562=>"011101101",
  34563=>"101001010",
  34564=>"000001110",
  34565=>"111100111",
  34566=>"010010011",
  34567=>"100011001",
  34568=>"011010110",
  34569=>"000001010",
  34570=>"000000001",
  34571=>"001101000",
  34572=>"110100001",
  34573=>"010001001",
  34574=>"110000000",
  34575=>"111010010",
  34576=>"111011001",
  34577=>"111110101",
  34578=>"010000100",
  34579=>"011100110",
  34580=>"010110110",
  34581=>"100110010",
  34582=>"110111000",
  34583=>"110110011",
  34584=>"000111000",
  34585=>"000000011",
  34586=>"001010010",
  34587=>"110011101",
  34588=>"000101001",
  34589=>"001011101",
  34590=>"000111001",
  34591=>"001010000",
  34592=>"110100101",
  34593=>"001111001",
  34594=>"011100100",
  34595=>"011111101",
  34596=>"011101110",
  34597=>"111001001",
  34598=>"011111110",
  34599=>"000111101",
  34600=>"101011011",
  34601=>"001000100",
  34602=>"110000001",
  34603=>"010100111",
  34604=>"010000000",
  34605=>"101111001",
  34606=>"001100101",
  34607=>"110100011",
  34608=>"010100000",
  34609=>"101001100",
  34610=>"111000111",
  34611=>"010001011",
  34612=>"101010101",
  34613=>"101110010",
  34614=>"111001001",
  34615=>"000101010",
  34616=>"111111101",
  34617=>"010100111",
  34618=>"111010101",
  34619=>"000111000",
  34620=>"001110101",
  34621=>"110001011",
  34622=>"010100110",
  34623=>"100001100",
  34624=>"011010101",
  34625=>"001001101",
  34626=>"110111010",
  34627=>"000010100",
  34628=>"010010111",
  34629=>"001001110",
  34630=>"001000110",
  34631=>"100010010",
  34632=>"111000100",
  34633=>"110100100",
  34634=>"110011110",
  34635=>"001010010",
  34636=>"001111111",
  34637=>"001101100",
  34638=>"010100001",
  34639=>"001100000",
  34640=>"001111110",
  34641=>"110010000",
  34642=>"010100111",
  34643=>"100000000",
  34644=>"000011111",
  34645=>"000100010",
  34646=>"100110101",
  34647=>"011010100",
  34648=>"010001100",
  34649=>"110100001",
  34650=>"000100111",
  34651=>"010101100",
  34652=>"110010010",
  34653=>"011011010",
  34654=>"000011101",
  34655=>"000010111",
  34656=>"110000101",
  34657=>"111100011",
  34658=>"001111111",
  34659=>"011101011",
  34660=>"000000101",
  34661=>"001111110",
  34662=>"000011101",
  34663=>"110001101",
  34664=>"101000100",
  34665=>"111001000",
  34666=>"101010110",
  34667=>"001010100",
  34668=>"101100110",
  34669=>"011001111",
  34670=>"011111101",
  34671=>"111000101",
  34672=>"110011100",
  34673=>"101001100",
  34674=>"101100000",
  34675=>"111011010",
  34676=>"101110100",
  34677=>"111001101",
  34678=>"110000110",
  34679=>"011010100",
  34680=>"100101100",
  34681=>"011000111",
  34682=>"101101111",
  34683=>"110001011",
  34684=>"011011101",
  34685=>"010110110",
  34686=>"010111011",
  34687=>"101100111",
  34688=>"010110011",
  34689=>"101000000",
  34690=>"001110001",
  34691=>"010010011",
  34692=>"101110001",
  34693=>"110001000",
  34694=>"011100110",
  34695=>"001111111",
  34696=>"101100101",
  34697=>"100011100",
  34698=>"101110100",
  34699=>"111011011",
  34700=>"101010001",
  34701=>"101111100",
  34702=>"111100010",
  34703=>"011110110",
  34704=>"100010011",
  34705=>"000011110",
  34706=>"100000101",
  34707=>"011000110",
  34708=>"011111001",
  34709=>"011111111",
  34710=>"101010001",
  34711=>"111111010",
  34712=>"010101010",
  34713=>"101001010",
  34714=>"100110101",
  34715=>"001001101",
  34716=>"100011001",
  34717=>"111010111",
  34718=>"100100011",
  34719=>"010010010",
  34720=>"111101100",
  34721=>"100011010",
  34722=>"001111110",
  34723=>"011110111",
  34724=>"110000110",
  34725=>"001000100",
  34726=>"100110000",
  34727=>"111011101",
  34728=>"001000000",
  34729=>"000100011",
  34730=>"000110101",
  34731=>"011000111",
  34732=>"010001110",
  34733=>"000110000",
  34734=>"010011011",
  34735=>"000010000",
  34736=>"100000001",
  34737=>"011010000",
  34738=>"001010100",
  34739=>"101001010",
  34740=>"110101111",
  34741=>"011011011",
  34742=>"100101000",
  34743=>"011000100",
  34744=>"011001100",
  34745=>"110000101",
  34746=>"001010011",
  34747=>"011101001",
  34748=>"000001110",
  34749=>"010000111",
  34750=>"011001011",
  34751=>"000011000",
  34752=>"001010011",
  34753=>"110100100",
  34754=>"100011100",
  34755=>"111001000",
  34756=>"000100001",
  34757=>"111000011",
  34758=>"110101110",
  34759=>"001010000",
  34760=>"011100001",
  34761=>"111111100",
  34762=>"111100001",
  34763=>"111111110",
  34764=>"001111000",
  34765=>"011011000",
  34766=>"001111110",
  34767=>"111110111",
  34768=>"000101110",
  34769=>"000111001",
  34770=>"000011011",
  34771=>"101001001",
  34772=>"010001110",
  34773=>"001000011",
  34774=>"000010101",
  34775=>"100001010",
  34776=>"000110111",
  34777=>"000111011",
  34778=>"111100101",
  34779=>"110001010",
  34780=>"011010000",
  34781=>"110011011",
  34782=>"000100100",
  34783=>"010101101",
  34784=>"110110110",
  34785=>"111110011",
  34786=>"001010010",
  34787=>"001100111",
  34788=>"001011100",
  34789=>"100001000",
  34790=>"111110000",
  34791=>"101100000",
  34792=>"111011001",
  34793=>"100011110",
  34794=>"100000000",
  34795=>"001101111",
  34796=>"001110011",
  34797=>"111111010",
  34798=>"010101100",
  34799=>"011101001",
  34800=>"000011111",
  34801=>"111011011",
  34802=>"000011101",
  34803=>"110000111",
  34804=>"110011111",
  34805=>"101100101",
  34806=>"100100101",
  34807=>"110100011",
  34808=>"001001011",
  34809=>"000000110",
  34810=>"101101000",
  34811=>"001011111",
  34812=>"010001001",
  34813=>"001100010",
  34814=>"111101011",
  34815=>"000110010",
  34816=>"001101011",
  34817=>"011011110",
  34818=>"110011011",
  34819=>"100001101",
  34820=>"110000001",
  34821=>"101110010",
  34822=>"000010100",
  34823=>"111000111",
  34824=>"010010001",
  34825=>"101110000",
  34826=>"000111001",
  34827=>"100000001",
  34828=>"111100000",
  34829=>"000001000",
  34830=>"001111111",
  34831=>"000111100",
  34832=>"010001100",
  34833=>"010001100",
  34834=>"000000010",
  34835=>"011011001",
  34836=>"010000011",
  34837=>"101011101",
  34838=>"111110010",
  34839=>"100000101",
  34840=>"001101101",
  34841=>"010010001",
  34842=>"101000111",
  34843=>"111101011",
  34844=>"010000100",
  34845=>"010000001",
  34846=>"101010000",
  34847=>"111110100",
  34848=>"001010001",
  34849=>"110101011",
  34850=>"110011101",
  34851=>"101000100",
  34852=>"000100101",
  34853=>"001101110",
  34854=>"110111010",
  34855=>"111111010",
  34856=>"101000100",
  34857=>"000101001",
  34858=>"100011000",
  34859=>"011100000",
  34860=>"101111001",
  34861=>"011111000",
  34862=>"111001001",
  34863=>"011100001",
  34864=>"001000011",
  34865=>"110010000",
  34866=>"011100100",
  34867=>"010100100",
  34868=>"011001111",
  34869=>"001000101",
  34870=>"101100000",
  34871=>"011011110",
  34872=>"000110111",
  34873=>"110111011",
  34874=>"000001101",
  34875=>"000111000",
  34876=>"000011100",
  34877=>"011001001",
  34878=>"101010011",
  34879=>"010001011",
  34880=>"101000011",
  34881=>"101000101",
  34882=>"111111001",
  34883=>"101101000",
  34884=>"101111010",
  34885=>"101001001",
  34886=>"101100110",
  34887=>"010010000",
  34888=>"110101000",
  34889=>"100100000",
  34890=>"000110101",
  34891=>"010111000",
  34892=>"100101011",
  34893=>"101110100",
  34894=>"101110110",
  34895=>"110010010",
  34896=>"110101101",
  34897=>"101000100",
  34898=>"011111011",
  34899=>"000100111",
  34900=>"100010011",
  34901=>"011011000",
  34902=>"000110010",
  34903=>"001101101",
  34904=>"100001000",
  34905=>"100011011",
  34906=>"101010100",
  34907=>"011000010",
  34908=>"010110101",
  34909=>"001100100",
  34910=>"000101110",
  34911=>"010010101",
  34912=>"101111011",
  34913=>"000111010",
  34914=>"001000110",
  34915=>"111001001",
  34916=>"100011111",
  34917=>"010010100",
  34918=>"000000010",
  34919=>"011111011",
  34920=>"000110001",
  34921=>"100111111",
  34922=>"000101010",
  34923=>"100000111",
  34924=>"100101100",
  34925=>"000010100",
  34926=>"100000100",
  34927=>"100110000",
  34928=>"111101101",
  34929=>"011110111",
  34930=>"101101101",
  34931=>"100101110",
  34932=>"010101111",
  34933=>"100001011",
  34934=>"010111111",
  34935=>"101011001",
  34936=>"101011101",
  34937=>"001101011",
  34938=>"010011110",
  34939=>"001111000",
  34940=>"010011111",
  34941=>"001011010",
  34942=>"000010100",
  34943=>"011111001",
  34944=>"000010000",
  34945=>"111001100",
  34946=>"101010000",
  34947=>"000001011",
  34948=>"111011001",
  34949=>"101100011",
  34950=>"110101101",
  34951=>"110010010",
  34952=>"110101101",
  34953=>"000101010",
  34954=>"101000101",
  34955=>"111110111",
  34956=>"111010110",
  34957=>"110101000",
  34958=>"001011101",
  34959=>"011111100",
  34960=>"001011100",
  34961=>"111101010",
  34962=>"001010100",
  34963=>"000111110",
  34964=>"011111001",
  34965=>"101110111",
  34966=>"001011110",
  34967=>"000001010",
  34968=>"010101000",
  34969=>"010111000",
  34970=>"010100101",
  34971=>"111001110",
  34972=>"000100110",
  34973=>"100000000",
  34974=>"100001001",
  34975=>"110100001",
  34976=>"111101010",
  34977=>"101011000",
  34978=>"010100001",
  34979=>"101101000",
  34980=>"100000100",
  34981=>"110110110",
  34982=>"001010101",
  34983=>"101000000",
  34984=>"011010100",
  34985=>"101010011",
  34986=>"000000110",
  34987=>"111001100",
  34988=>"000001000",
  34989=>"001000101",
  34990=>"100010000",
  34991=>"110010000",
  34992=>"011000010",
  34993=>"101101000",
  34994=>"111011011",
  34995=>"111101110",
  34996=>"111001110",
  34997=>"000100010",
  34998=>"001011011",
  34999=>"100101110",
  35000=>"100110011",
  35001=>"101100111",
  35002=>"100001101",
  35003=>"110111101",
  35004=>"011000111",
  35005=>"111101111",
  35006=>"001011110",
  35007=>"001010110",
  35008=>"100001100",
  35009=>"011000111",
  35010=>"000111000",
  35011=>"011110101",
  35012=>"111101000",
  35013=>"101000110",
  35014=>"000000011",
  35015=>"010001100",
  35016=>"111101111",
  35017=>"001001100",
  35018=>"100111110",
  35019=>"111000100",
  35020=>"010110101",
  35021=>"011110111",
  35022=>"001001110",
  35023=>"100000010",
  35024=>"110000010",
  35025=>"000001010",
  35026=>"101101100",
  35027=>"000011101",
  35028=>"000000011",
  35029=>"010001001",
  35030=>"010011001",
  35031=>"111011100",
  35032=>"010110000",
  35033=>"100100000",
  35034=>"101000110",
  35035=>"101011001",
  35036=>"011100010",
  35037=>"111000111",
  35038=>"011100011",
  35039=>"000111100",
  35040=>"101000001",
  35041=>"101010000",
  35042=>"001001000",
  35043=>"101010101",
  35044=>"010001110",
  35045=>"011001000",
  35046=>"000001000",
  35047=>"001010011",
  35048=>"100010101",
  35049=>"100001110",
  35050=>"001111110",
  35051=>"101010101",
  35052=>"010110111",
  35053=>"011001011",
  35054=>"100000110",
  35055=>"001001000",
  35056=>"110001011",
  35057=>"001100001",
  35058=>"000101010",
  35059=>"111010101",
  35060=>"000010111",
  35061=>"011111000",
  35062=>"011111001",
  35063=>"100011010",
  35064=>"101011101",
  35065=>"111011010",
  35066=>"000110011",
  35067=>"000100001",
  35068=>"001000101",
  35069=>"110110000",
  35070=>"001010100",
  35071=>"111001011",
  35072=>"101011100",
  35073=>"110101101",
  35074=>"011110010",
  35075=>"101001001",
  35076=>"100101000",
  35077=>"000100011",
  35078=>"011101011",
  35079=>"011101001",
  35080=>"010000010",
  35081=>"100111010",
  35082=>"011001100",
  35083=>"001011011",
  35084=>"011100100",
  35085=>"101101111",
  35086=>"100111100",
  35087=>"110101110",
  35088=>"010001100",
  35089=>"111110110",
  35090=>"100001011",
  35091=>"001110011",
  35092=>"111101100",
  35093=>"011001010",
  35094=>"011000111",
  35095=>"111110011",
  35096=>"111111110",
  35097=>"011101001",
  35098=>"111110001",
  35099=>"101101010",
  35100=>"001011001",
  35101=>"111110010",
  35102=>"101100010",
  35103=>"000001001",
  35104=>"010000101",
  35105=>"010011110",
  35106=>"101011000",
  35107=>"111110111",
  35108=>"110000010",
  35109=>"101100101",
  35110=>"111101100",
  35111=>"110101110",
  35112=>"011010111",
  35113=>"001101101",
  35114=>"011110101",
  35115=>"100101100",
  35116=>"101000100",
  35117=>"011100111",
  35118=>"010100111",
  35119=>"101000000",
  35120=>"011110111",
  35121=>"100100000",
  35122=>"100001001",
  35123=>"001111010",
  35124=>"100000100",
  35125=>"000111101",
  35126=>"101001011",
  35127=>"110000010",
  35128=>"100111000",
  35129=>"110001010",
  35130=>"011111110",
  35131=>"010011110",
  35132=>"010000010",
  35133=>"100101100",
  35134=>"100000011",
  35135=>"110101110",
  35136=>"111000001",
  35137=>"011110111",
  35138=>"111100110",
  35139=>"010011010",
  35140=>"101001011",
  35141=>"001001111",
  35142=>"001100100",
  35143=>"101000000",
  35144=>"100010001",
  35145=>"110101001",
  35146=>"100000100",
  35147=>"001000010",
  35148=>"110000100",
  35149=>"001001001",
  35150=>"100000111",
  35151=>"000011000",
  35152=>"101001101",
  35153=>"100010011",
  35154=>"010110110",
  35155=>"101011011",
  35156=>"011100011",
  35157=>"010000011",
  35158=>"101000100",
  35159=>"100111010",
  35160=>"111001001",
  35161=>"011100001",
  35162=>"001111100",
  35163=>"010011010",
  35164=>"000010110",
  35165=>"001011001",
  35166=>"110011000",
  35167=>"010010111",
  35168=>"111011101",
  35169=>"011011010",
  35170=>"010010001",
  35171=>"101111011",
  35172=>"011101100",
  35173=>"100000010",
  35174=>"101101011",
  35175=>"111101101",
  35176=>"000001100",
  35177=>"010100010",
  35178=>"101001110",
  35179=>"100101100",
  35180=>"000110101",
  35181=>"011011010",
  35182=>"001101110",
  35183=>"101111011",
  35184=>"001001010",
  35185=>"010011110",
  35186=>"101001010",
  35187=>"111100011",
  35188=>"011000100",
  35189=>"001010010",
  35190=>"111011100",
  35191=>"111011111",
  35192=>"000000110",
  35193=>"111110001",
  35194=>"001000101",
  35195=>"001000000",
  35196=>"100011000",
  35197=>"111101100",
  35198=>"000011100",
  35199=>"011111110",
  35200=>"111001101",
  35201=>"111101001",
  35202=>"000000100",
  35203=>"001100001",
  35204=>"100100000",
  35205=>"000000011",
  35206=>"111100100",
  35207=>"111111101",
  35208=>"100100000",
  35209=>"110010101",
  35210=>"111110000",
  35211=>"000001001",
  35212=>"000111110",
  35213=>"100010101",
  35214=>"000011101",
  35215=>"101010111",
  35216=>"101110001",
  35217=>"001001011",
  35218=>"101011001",
  35219=>"111010111",
  35220=>"000110101",
  35221=>"000001101",
  35222=>"100000001",
  35223=>"100111110",
  35224=>"100011000",
  35225=>"101110000",
  35226=>"000011001",
  35227=>"111010000",
  35228=>"000100010",
  35229=>"010100101",
  35230=>"100000001",
  35231=>"011011101",
  35232=>"101011001",
  35233=>"010011101",
  35234=>"100000010",
  35235=>"111100101",
  35236=>"111101111",
  35237=>"011001011",
  35238=>"111110011",
  35239=>"111101011",
  35240=>"001100111",
  35241=>"010111101",
  35242=>"110111001",
  35243=>"110111111",
  35244=>"100001000",
  35245=>"111011011",
  35246=>"000110010",
  35247=>"000010000",
  35248=>"011101011",
  35249=>"001101111",
  35250=>"110000011",
  35251=>"000101110",
  35252=>"100010110",
  35253=>"000110101",
  35254=>"001111001",
  35255=>"001010101",
  35256=>"111000101",
  35257=>"100100010",
  35258=>"110100010",
  35259=>"000000100",
  35260=>"110111001",
  35261=>"011101011",
  35262=>"100010101",
  35263=>"111011111",
  35264=>"000001110",
  35265=>"010110010",
  35266=>"010100110",
  35267=>"010000001",
  35268=>"100101000",
  35269=>"000111000",
  35270=>"001101101",
  35271=>"100000100",
  35272=>"011000001",
  35273=>"000010101",
  35274=>"000011001",
  35275=>"100001011",
  35276=>"000110010",
  35277=>"011101101",
  35278=>"100110101",
  35279=>"110011111",
  35280=>"010100010",
  35281=>"110110100",
  35282=>"111000011",
  35283=>"011001011",
  35284=>"111111100",
  35285=>"010011000",
  35286=>"110101110",
  35287=>"011001000",
  35288=>"100100110",
  35289=>"100101110",
  35290=>"111000111",
  35291=>"010011001",
  35292=>"001110110",
  35293=>"110011110",
  35294=>"011011010",
  35295=>"111100110",
  35296=>"111001100",
  35297=>"100111111",
  35298=>"100101101",
  35299=>"011110001",
  35300=>"010000000",
  35301=>"011100100",
  35302=>"101101011",
  35303=>"000000001",
  35304=>"100100110",
  35305=>"100101011",
  35306=>"100101001",
  35307=>"100100100",
  35308=>"100001101",
  35309=>"010111111",
  35310=>"100111000",
  35311=>"101111101",
  35312=>"010011010",
  35313=>"000100011",
  35314=>"110000000",
  35315=>"011100101",
  35316=>"110011011",
  35317=>"110110110",
  35318=>"000100001",
  35319=>"010001100",
  35320=>"000100001",
  35321=>"101100011",
  35322=>"110101100",
  35323=>"100111101",
  35324=>"010101001",
  35325=>"111011101",
  35326=>"000000111",
  35327=>"110110111",
  35328=>"001010000",
  35329=>"010101011",
  35330=>"100101011",
  35331=>"000100000",
  35332=>"111111010",
  35333=>"111010100",
  35334=>"111010000",
  35335=>"011101000",
  35336=>"001001111",
  35337=>"000011010",
  35338=>"101010001",
  35339=>"111011110",
  35340=>"110100110",
  35341=>"100011110",
  35342=>"000011110",
  35343=>"010010000",
  35344=>"001010001",
  35345=>"000001011",
  35346=>"111100100",
  35347=>"100111001",
  35348=>"001001000",
  35349=>"001110101",
  35350=>"101111001",
  35351=>"010101110",
  35352=>"010100101",
  35353=>"110001100",
  35354=>"001000101",
  35355=>"101001011",
  35356=>"101111000",
  35357=>"110010011",
  35358=>"111101111",
  35359=>"111001101",
  35360=>"001011100",
  35361=>"000010001",
  35362=>"000110111",
  35363=>"110001010",
  35364=>"111011011",
  35365=>"100101000",
  35366=>"000110000",
  35367=>"000101001",
  35368=>"001000001",
  35369=>"101001001",
  35370=>"010101110",
  35371=>"100001000",
  35372=>"010100101",
  35373=>"110010100",
  35374=>"001010101",
  35375=>"100100100",
  35376=>"011001010",
  35377=>"001110111",
  35378=>"100000110",
  35379=>"110010011",
  35380=>"000000000",
  35381=>"011010011",
  35382=>"001000100",
  35383=>"100100100",
  35384=>"000011010",
  35385=>"100001101",
  35386=>"110010010",
  35387=>"100101010",
  35388=>"110010010",
  35389=>"111111010",
  35390=>"010110011",
  35391=>"010100100",
  35392=>"011000101",
  35393=>"000110000",
  35394=>"011110011",
  35395=>"110010110",
  35396=>"011011110",
  35397=>"101101101",
  35398=>"010101001",
  35399=>"001110110",
  35400=>"101010010",
  35401=>"111011110",
  35402=>"011100111",
  35403=>"100101011",
  35404=>"010111010",
  35405=>"001110010",
  35406=>"000011110",
  35407=>"000101001",
  35408=>"011111001",
  35409=>"110001010",
  35410=>"000110111",
  35411=>"100001011",
  35412=>"010101100",
  35413=>"111101101",
  35414=>"000110101",
  35415=>"010111100",
  35416=>"101010111",
  35417=>"100010101",
  35418=>"100001000",
  35419=>"011010111",
  35420=>"100010011",
  35421=>"000110000",
  35422=>"111100110",
  35423=>"001110111",
  35424=>"001111111",
  35425=>"111000001",
  35426=>"000100011",
  35427=>"101011100",
  35428=>"101001111",
  35429=>"100010010",
  35430=>"100101110",
  35431=>"001110101",
  35432=>"011011110",
  35433=>"100000101",
  35434=>"110111100",
  35435=>"001100111",
  35436=>"001100011",
  35437=>"101110110",
  35438=>"001111010",
  35439=>"110100111",
  35440=>"101110000",
  35441=>"101100100",
  35442=>"010101101",
  35443=>"111101011",
  35444=>"100100101",
  35445=>"010101111",
  35446=>"000101010",
  35447=>"010111011",
  35448=>"100000110",
  35449=>"001101011",
  35450=>"001000100",
  35451=>"001011010",
  35452=>"110110001",
  35453=>"010001111",
  35454=>"011000101",
  35455=>"110001000",
  35456=>"101011111",
  35457=>"010010110",
  35458=>"011111110",
  35459=>"000100100",
  35460=>"110101100",
  35461=>"101001010",
  35462=>"111100100",
  35463=>"001011101",
  35464=>"000000111",
  35465=>"010101010",
  35466=>"100010100",
  35467=>"000001011",
  35468=>"111110111",
  35469=>"110101101",
  35470=>"000010101",
  35471=>"100110101",
  35472=>"000110001",
  35473=>"100101110",
  35474=>"111101101",
  35475=>"110010111",
  35476=>"001000000",
  35477=>"110000001",
  35478=>"111101110",
  35479=>"010111101",
  35480=>"110101110",
  35481=>"110111001",
  35482=>"101100100",
  35483=>"000001111",
  35484=>"000000011",
  35485=>"000000101",
  35486=>"000010110",
  35487=>"101011111",
  35488=>"111011011",
  35489=>"110011011",
  35490=>"000110111",
  35491=>"100110011",
  35492=>"001010011",
  35493=>"010100101",
  35494=>"111010001",
  35495=>"001011110",
  35496=>"000111100",
  35497=>"010100011",
  35498=>"011101100",
  35499=>"100100101",
  35500=>"111011110",
  35501=>"001101001",
  35502=>"100010001",
  35503=>"100100111",
  35504=>"011111000",
  35505=>"010110010",
  35506=>"101100111",
  35507=>"000110101",
  35508=>"100101000",
  35509=>"100110101",
  35510=>"101001011",
  35511=>"000000000",
  35512=>"000111111",
  35513=>"000100010",
  35514=>"001111110",
  35515=>"110000110",
  35516=>"001110010",
  35517=>"100100001",
  35518=>"000010001",
  35519=>"110001101",
  35520=>"001000111",
  35521=>"101111011",
  35522=>"010010001",
  35523=>"001010110",
  35524=>"100000001",
  35525=>"000011100",
  35526=>"010101100",
  35527=>"010111110",
  35528=>"010100001",
  35529=>"101001001",
  35530=>"001101111",
  35531=>"000001100",
  35532=>"101111001",
  35533=>"111011000",
  35534=>"001110001",
  35535=>"110110010",
  35536=>"110111001",
  35537=>"000011011",
  35538=>"111101100",
  35539=>"000001011",
  35540=>"111110110",
  35541=>"111010101",
  35542=>"100001010",
  35543=>"000111101",
  35544=>"010001110",
  35545=>"011011110",
  35546=>"001101100",
  35547=>"101001100",
  35548=>"001100101",
  35549=>"100110011",
  35550=>"010101011",
  35551=>"101110000",
  35552=>"000011011",
  35553=>"100101010",
  35554=>"101011000",
  35555=>"000011110",
  35556=>"100100011",
  35557=>"110111110",
  35558=>"000011001",
  35559=>"001111111",
  35560=>"111011010",
  35561=>"111100101",
  35562=>"001101001",
  35563=>"000010100",
  35564=>"010000001",
  35565=>"001111000",
  35566=>"011101001",
  35567=>"000111111",
  35568=>"001000101",
  35569=>"000110000",
  35570=>"101110111",
  35571=>"011011011",
  35572=>"000011111",
  35573=>"100001011",
  35574=>"000111011",
  35575=>"100111001",
  35576=>"111011101",
  35577=>"001011000",
  35578=>"010110010",
  35579=>"000100101",
  35580=>"011000001",
  35581=>"110011100",
  35582=>"010011010",
  35583=>"100010001",
  35584=>"000001011",
  35585=>"000101100",
  35586=>"010101011",
  35587=>"000011000",
  35588=>"001000011",
  35589=>"000100101",
  35590=>"111011110",
  35591=>"001011110",
  35592=>"000101111",
  35593=>"110000011",
  35594=>"101000111",
  35595=>"001101100",
  35596=>"110111010",
  35597=>"010011010",
  35598=>"001000111",
  35599=>"111011000",
  35600=>"110000101",
  35601=>"111110110",
  35602=>"110111011",
  35603=>"011010000",
  35604=>"111000100",
  35605=>"101101110",
  35606=>"100001011",
  35607=>"111000001",
  35608=>"101110010",
  35609=>"010000010",
  35610=>"001101110",
  35611=>"011011001",
  35612=>"010000011",
  35613=>"101010111",
  35614=>"000000011",
  35615=>"110100010",
  35616=>"101010111",
  35617=>"010000010",
  35618=>"111111110",
  35619=>"111001100",
  35620=>"000101010",
  35621=>"001001100",
  35622=>"100101001",
  35623=>"001001100",
  35624=>"101100110",
  35625=>"011000010",
  35626=>"100000011",
  35627=>"011000001",
  35628=>"100011001",
  35629=>"001101110",
  35630=>"000101010",
  35631=>"000111101",
  35632=>"011100000",
  35633=>"001001010",
  35634=>"010001111",
  35635=>"111101100",
  35636=>"101111111",
  35637=>"101100011",
  35638=>"000000101",
  35639=>"101000111",
  35640=>"000100111",
  35641=>"110000001",
  35642=>"111000011",
  35643=>"000111101",
  35644=>"011111010",
  35645=>"000100111",
  35646=>"110001110",
  35647=>"011010111",
  35648=>"011000011",
  35649=>"110010111",
  35650=>"110111100",
  35651=>"111101011",
  35652=>"100010111",
  35653=>"101100001",
  35654=>"100001111",
  35655=>"001110001",
  35656=>"101111010",
  35657=>"110001100",
  35658=>"001010101",
  35659=>"000110000",
  35660=>"011101000",
  35661=>"001000011",
  35662=>"010010100",
  35663=>"010010001",
  35664=>"000000011",
  35665=>"010001101",
  35666=>"010000101",
  35667=>"110011100",
  35668=>"011111011",
  35669=>"000100100",
  35670=>"111011101",
  35671=>"100011010",
  35672=>"101100000",
  35673=>"110010110",
  35674=>"111011010",
  35675=>"110000111",
  35676=>"111100000",
  35677=>"001001000",
  35678=>"010101101",
  35679=>"100110011",
  35680=>"110101111",
  35681=>"101100111",
  35682=>"000001011",
  35683=>"000010010",
  35684=>"110011011",
  35685=>"000001011",
  35686=>"011101011",
  35687=>"011001111",
  35688=>"011000001",
  35689=>"111111110",
  35690=>"111001110",
  35691=>"111111111",
  35692=>"101001000",
  35693=>"110000010",
  35694=>"010010000",
  35695=>"100110101",
  35696=>"001000100",
  35697=>"010011010",
  35698=>"101011011",
  35699=>"001101100",
  35700=>"000000001",
  35701=>"001111111",
  35702=>"000000101",
  35703=>"100001011",
  35704=>"100101110",
  35705=>"000010101",
  35706=>"000000101",
  35707=>"010101011",
  35708=>"001010011",
  35709=>"011001001",
  35710=>"111000111",
  35711=>"000001001",
  35712=>"101010110",
  35713=>"111010100",
  35714=>"000110111",
  35715=>"001010101",
  35716=>"010000101",
  35717=>"010111010",
  35718=>"100110010",
  35719=>"110010111",
  35720=>"010000100",
  35721=>"000100111",
  35722=>"101011011",
  35723=>"001011010",
  35724=>"110010010",
  35725=>"010000011",
  35726=>"101110110",
  35727=>"010010010",
  35728=>"101010011",
  35729=>"110000010",
  35730=>"000101011",
  35731=>"011111011",
  35732=>"011101000",
  35733=>"001010001",
  35734=>"000100111",
  35735=>"010001110",
  35736=>"101111101",
  35737=>"101001010",
  35738=>"010100000",
  35739=>"010000001",
  35740=>"011010111",
  35741=>"101010000",
  35742=>"000100100",
  35743=>"000010011",
  35744=>"010111011",
  35745=>"100101000",
  35746=>"001000011",
  35747=>"010000001",
  35748=>"001101000",
  35749=>"101000001",
  35750=>"010100000",
  35751=>"000000100",
  35752=>"101000000",
  35753=>"001001000",
  35754=>"101010011",
  35755=>"111011100",
  35756=>"110011010",
  35757=>"000011101",
  35758=>"111000111",
  35759=>"101000010",
  35760=>"000001101",
  35761=>"111000101",
  35762=>"100101100",
  35763=>"110010001",
  35764=>"011111001",
  35765=>"100011101",
  35766=>"100001000",
  35767=>"110000010",
  35768=>"100100010",
  35769=>"111100100",
  35770=>"011101111",
  35771=>"010000100",
  35772=>"011001001",
  35773=>"010001000",
  35774=>"111010101",
  35775=>"000000011",
  35776=>"011001011",
  35777=>"000100010",
  35778=>"110100001",
  35779=>"010110100",
  35780=>"110111101",
  35781=>"010001011",
  35782=>"010100110",
  35783=>"100001110",
  35784=>"100011000",
  35785=>"011011001",
  35786=>"101100101",
  35787=>"010100010",
  35788=>"000000010",
  35789=>"111100100",
  35790=>"010001010",
  35791=>"111111011",
  35792=>"011001010",
  35793=>"010000100",
  35794=>"010001001",
  35795=>"001101111",
  35796=>"011010110",
  35797=>"111010001",
  35798=>"010010101",
  35799=>"011111000",
  35800=>"000110000",
  35801=>"111100101",
  35802=>"000011111",
  35803=>"110000110",
  35804=>"100110010",
  35805=>"000010010",
  35806=>"011001010",
  35807=>"101100011",
  35808=>"011100001",
  35809=>"111010110",
  35810=>"101110100",
  35811=>"111101010",
  35812=>"011010000",
  35813=>"001100100",
  35814=>"000001011",
  35815=>"000110010",
  35816=>"001011010",
  35817=>"000011011",
  35818=>"100000111",
  35819=>"011101110",
  35820=>"101100111",
  35821=>"111111110",
  35822=>"110001110",
  35823=>"001001010",
  35824=>"001101011",
  35825=>"001010001",
  35826=>"001101011",
  35827=>"011000010",
  35828=>"111111111",
  35829=>"101111000",
  35830=>"011011101",
  35831=>"111010001",
  35832=>"111010111",
  35833=>"111100101",
  35834=>"100111001",
  35835=>"001011110",
  35836=>"100000000",
  35837=>"000010100",
  35838=>"111111101",
  35839=>"000010000",
  35840=>"111101000",
  35841=>"101010010",
  35842=>"100110000",
  35843=>"001111111",
  35844=>"000111100",
  35845=>"001000100",
  35846=>"000111101",
  35847=>"010101010",
  35848=>"111110101",
  35849=>"101111101",
  35850=>"111010110",
  35851=>"010100001",
  35852=>"011111110",
  35853=>"011110000",
  35854=>"100011101",
  35855=>"101011011",
  35856=>"000000110",
  35857=>"001011011",
  35858=>"101000100",
  35859=>"111011100",
  35860=>"101101010",
  35861=>"000011101",
  35862=>"010010111",
  35863=>"111101000",
  35864=>"010100000",
  35865=>"011111111",
  35866=>"001010101",
  35867=>"111001001",
  35868=>"000100001",
  35869=>"111100001",
  35870=>"100110011",
  35871=>"011001000",
  35872=>"111100110",
  35873=>"101101011",
  35874=>"001101101",
  35875=>"110111001",
  35876=>"101101010",
  35877=>"111101000",
  35878=>"011000100",
  35879=>"110101011",
  35880=>"011011010",
  35881=>"111001100",
  35882=>"010011110",
  35883=>"000000111",
  35884=>"100011110",
  35885=>"010010101",
  35886=>"101111110",
  35887=>"001100001",
  35888=>"011100110",
  35889=>"110101110",
  35890=>"010011110",
  35891=>"100100011",
  35892=>"010111000",
  35893=>"111001011",
  35894=>"000011100",
  35895=>"111000111",
  35896=>"011011101",
  35897=>"011101111",
  35898=>"111100100",
  35899=>"010000010",
  35900=>"000101010",
  35901=>"111010100",
  35902=>"101000000",
  35903=>"110110110",
  35904=>"100010101",
  35905=>"010110001",
  35906=>"111101010",
  35907=>"010111010",
  35908=>"011011000",
  35909=>"011100100",
  35910=>"000101101",
  35911=>"100101111",
  35912=>"000101010",
  35913=>"101101100",
  35914=>"110011101",
  35915=>"100000001",
  35916=>"111111111",
  35917=>"100110001",
  35918=>"110100111",
  35919=>"111000101",
  35920=>"000000000",
  35921=>"010110100",
  35922=>"000101011",
  35923=>"100000111",
  35924=>"000001100",
  35925=>"100000011",
  35926=>"000001010",
  35927=>"110010101",
  35928=>"101111000",
  35929=>"111101010",
  35930=>"010110101",
  35931=>"100010010",
  35932=>"011011001",
  35933=>"000110101",
  35934=>"100111000",
  35935=>"011001010",
  35936=>"010010100",
  35937=>"100100000",
  35938=>"100001100",
  35939=>"100111001",
  35940=>"010111011",
  35941=>"000110001",
  35942=>"001010111",
  35943=>"101111101",
  35944=>"000011000",
  35945=>"111111101",
  35946=>"110000010",
  35947=>"011111001",
  35948=>"000101111",
  35949=>"001110001",
  35950=>"110111011",
  35951=>"000100100",
  35952=>"110010110",
  35953=>"000010110",
  35954=>"011100011",
  35955=>"011110111",
  35956=>"110011100",
  35957=>"110100100",
  35958=>"110110001",
  35959=>"111010000",
  35960=>"011101101",
  35961=>"000101110",
  35962=>"101101000",
  35963=>"110000111",
  35964=>"010001111",
  35965=>"000101001",
  35966=>"110101011",
  35967=>"111101001",
  35968=>"100001111",
  35969=>"100011111",
  35970=>"011010000",
  35971=>"101010101",
  35972=>"000011010",
  35973=>"101111010",
  35974=>"111111101",
  35975=>"000111000",
  35976=>"000001010",
  35977=>"100010011",
  35978=>"011110010",
  35979=>"001110100",
  35980=>"000101101",
  35981=>"110110010",
  35982=>"101010001",
  35983=>"001110010",
  35984=>"110001101",
  35985=>"111011000",
  35986=>"101011000",
  35987=>"001110101",
  35988=>"110011111",
  35989=>"001001010",
  35990=>"101001001",
  35991=>"111001001",
  35992=>"111101110",
  35993=>"010010111",
  35994=>"011001010",
  35995=>"000110000",
  35996=>"000100001",
  35997=>"010100101",
  35998=>"001110010",
  35999=>"001110110",
  36000=>"010100011",
  36001=>"101110001",
  36002=>"100101101",
  36003=>"101000111",
  36004=>"100001110",
  36005=>"101001100",
  36006=>"010010100",
  36007=>"010010000",
  36008=>"000101010",
  36009=>"100011001",
  36010=>"101010010",
  36011=>"101010100",
  36012=>"101100100",
  36013=>"111111011",
  36014=>"100001010",
  36015=>"010101111",
  36016=>"010000011",
  36017=>"001100101",
  36018=>"100110000",
  36019=>"100101110",
  36020=>"110110000",
  36021=>"101010111",
  36022=>"110000010",
  36023=>"001100100",
  36024=>"010101011",
  36025=>"000001000",
  36026=>"010111100",
  36027=>"000110101",
  36028=>"011000000",
  36029=>"010000001",
  36030=>"010001101",
  36031=>"000111010",
  36032=>"001101011",
  36033=>"000001001",
  36034=>"110111001",
  36035=>"010011000",
  36036=>"111110101",
  36037=>"110101000",
  36038=>"100001011",
  36039=>"110111101",
  36040=>"101000011",
  36041=>"011100110",
  36042=>"110010010",
  36043=>"000101101",
  36044=>"101001010",
  36045=>"011101111",
  36046=>"000011101",
  36047=>"000011101",
  36048=>"100101110",
  36049=>"011110000",
  36050=>"111101101",
  36051=>"100110011",
  36052=>"001010000",
  36053=>"011110110",
  36054=>"111011011",
  36055=>"100101010",
  36056=>"111001000",
  36057=>"011000110",
  36058=>"100000000",
  36059=>"011011001",
  36060=>"101011100",
  36061=>"111100110",
  36062=>"001111100",
  36063=>"001010001",
  36064=>"111101010",
  36065=>"110011101",
  36066=>"011101111",
  36067=>"101101110",
  36068=>"001100110",
  36069=>"000110111",
  36070=>"100111001",
  36071=>"011000011",
  36072=>"000100000",
  36073=>"011000010",
  36074=>"100110011",
  36075=>"101010000",
  36076=>"000111110",
  36077=>"101100001",
  36078=>"111001100",
  36079=>"011000011",
  36080=>"001000000",
  36081=>"000101100",
  36082=>"001101111",
  36083=>"101100110",
  36084=>"100001101",
  36085=>"110101000",
  36086=>"110111100",
  36087=>"111111111",
  36088=>"000011010",
  36089=>"110010111",
  36090=>"000111111",
  36091=>"010001000",
  36092=>"000001111",
  36093=>"000111000",
  36094=>"100101101",
  36095=>"010111000",
  36096=>"011110111",
  36097=>"111110001",
  36098=>"110100111",
  36099=>"101100110",
  36100=>"110001000",
  36101=>"000000111",
  36102=>"111001011",
  36103=>"100000001",
  36104=>"111010110",
  36105=>"000111000",
  36106=>"001110100",
  36107=>"111001010",
  36108=>"000110110",
  36109=>"100100100",
  36110=>"011111010",
  36111=>"010000111",
  36112=>"010101110",
  36113=>"000000001",
  36114=>"001011111",
  36115=>"111100011",
  36116=>"111010111",
  36117=>"010111101",
  36118=>"010010000",
  36119=>"001000100",
  36120=>"111110110",
  36121=>"110010001",
  36122=>"000100101",
  36123=>"000000001",
  36124=>"101111000",
  36125=>"110000011",
  36126=>"110011000",
  36127=>"000001101",
  36128=>"100010100",
  36129=>"100111000",
  36130=>"011000111",
  36131=>"001110001",
  36132=>"000100100",
  36133=>"001100111",
  36134=>"001111010",
  36135=>"001000010",
  36136=>"110011110",
  36137=>"000001101",
  36138=>"000000111",
  36139=>"101010111",
  36140=>"111000101",
  36141=>"001000000",
  36142=>"101011011",
  36143=>"011000111",
  36144=>"101001010",
  36145=>"001100011",
  36146=>"001100010",
  36147=>"011111010",
  36148=>"000100100",
  36149=>"101111111",
  36150=>"000001010",
  36151=>"111111001",
  36152=>"001100101",
  36153=>"111001001",
  36154=>"101001011",
  36155=>"100001110",
  36156=>"110101010",
  36157=>"110110001",
  36158=>"001100000",
  36159=>"010011011",
  36160=>"010010100",
  36161=>"110111010",
  36162=>"100100001",
  36163=>"000000101",
  36164=>"011010000",
  36165=>"111110000",
  36166=>"000100011",
  36167=>"010111111",
  36168=>"010010001",
  36169=>"001000101",
  36170=>"101110100",
  36171=>"000000101",
  36172=>"110110000",
  36173=>"110011001",
  36174=>"000110100",
  36175=>"011110110",
  36176=>"000010101",
  36177=>"101011011",
  36178=>"011011001",
  36179=>"100100010",
  36180=>"011111100",
  36181=>"100101101",
  36182=>"001000010",
  36183=>"100100000",
  36184=>"100001110",
  36185=>"100000000",
  36186=>"010111101",
  36187=>"000100010",
  36188=>"110100010",
  36189=>"001011000",
  36190=>"001010001",
  36191=>"101001000",
  36192=>"001110110",
  36193=>"001100101",
  36194=>"111111111",
  36195=>"001000001",
  36196=>"011100110",
  36197=>"101010001",
  36198=>"101001010",
  36199=>"010001111",
  36200=>"111001011",
  36201=>"110100011",
  36202=>"011011001",
  36203=>"001101110",
  36204=>"001001110",
  36205=>"101001101",
  36206=>"111011101",
  36207=>"110101110",
  36208=>"001000000",
  36209=>"101010111",
  36210=>"010000000",
  36211=>"011000010",
  36212=>"000111011",
  36213=>"010000110",
  36214=>"110000000",
  36215=>"110110001",
  36216=>"001101000",
  36217=>"000100101",
  36218=>"010001100",
  36219=>"101110100",
  36220=>"001111001",
  36221=>"111111100",
  36222=>"000101001",
  36223=>"101010001",
  36224=>"111111101",
  36225=>"110110000",
  36226=>"111011011",
  36227=>"110011100",
  36228=>"000001011",
  36229=>"000101010",
  36230=>"000110101",
  36231=>"100000010",
  36232=>"111011001",
  36233=>"010110110",
  36234=>"111001100",
  36235=>"011000001",
  36236=>"111110100",
  36237=>"010110001",
  36238=>"110101110",
  36239=>"010101110",
  36240=>"110000111",
  36241=>"111000110",
  36242=>"001001101",
  36243=>"011111101",
  36244=>"100010101",
  36245=>"110001110",
  36246=>"101010000",
  36247=>"101011110",
  36248=>"101001101",
  36249=>"001101001",
  36250=>"100100010",
  36251=>"101010101",
  36252=>"011000111",
  36253=>"101000010",
  36254=>"101001101",
  36255=>"001110111",
  36256=>"101100110",
  36257=>"000000000",
  36258=>"100111001",
  36259=>"000010100",
  36260=>"011100110",
  36261=>"110010101",
  36262=>"010000100",
  36263=>"101000110",
  36264=>"000000110",
  36265=>"000100100",
  36266=>"101011010",
  36267=>"111000100",
  36268=>"101101110",
  36269=>"010101111",
  36270=>"000000010",
  36271=>"001101001",
  36272=>"111110000",
  36273=>"111000100",
  36274=>"011100011",
  36275=>"011010010",
  36276=>"111111101",
  36277=>"111010000",
  36278=>"111101100",
  36279=>"011011011",
  36280=>"111100010",
  36281=>"001110111",
  36282=>"001000000",
  36283=>"001100101",
  36284=>"101011100",
  36285=>"111000000",
  36286=>"111100101",
  36287=>"111001100",
  36288=>"101001011",
  36289=>"010100001",
  36290=>"101010101",
  36291=>"100011011",
  36292=>"000101010",
  36293=>"001010100",
  36294=>"000100000",
  36295=>"110010010",
  36296=>"000110100",
  36297=>"111111011",
  36298=>"010001011",
  36299=>"101111001",
  36300=>"001101001",
  36301=>"110010001",
  36302=>"001010100",
  36303=>"111100111",
  36304=>"010011111",
  36305=>"100100111",
  36306=>"010010100",
  36307=>"010001000",
  36308=>"011101000",
  36309=>"110000000",
  36310=>"000100101",
  36311=>"111000101",
  36312=>"101010000",
  36313=>"011011111",
  36314=>"110100100",
  36315=>"100000100",
  36316=>"111011001",
  36317=>"110101111",
  36318=>"100100000",
  36319=>"011010110",
  36320=>"101101011",
  36321=>"110111111",
  36322=>"111011100",
  36323=>"000101011",
  36324=>"111010111",
  36325=>"100000011",
  36326=>"000111001",
  36327=>"101111100",
  36328=>"011000001",
  36329=>"001010101",
  36330=>"000000000",
  36331=>"100011010",
  36332=>"001110111",
  36333=>"011100100",
  36334=>"001001000",
  36335=>"011011110",
  36336=>"100101101",
  36337=>"100011011",
  36338=>"100111010",
  36339=>"010111101",
  36340=>"111101010",
  36341=>"110000100",
  36342=>"011111100",
  36343=>"100111010",
  36344=>"011001110",
  36345=>"000010000",
  36346=>"100000000",
  36347=>"010010001",
  36348=>"101111011",
  36349=>"101000001",
  36350=>"010110010",
  36351=>"011001000",
  36352=>"010000100",
  36353=>"101101000",
  36354=>"001011010",
  36355=>"001011111",
  36356=>"001101001",
  36357=>"000010000",
  36358=>"001000111",
  36359=>"001000110",
  36360=>"011011000",
  36361=>"111111110",
  36362=>"111100111",
  36363=>"100000011",
  36364=>"001010110",
  36365=>"110101100",
  36366=>"000111111",
  36367=>"010111000",
  36368=>"000011010",
  36369=>"011111111",
  36370=>"000101011",
  36371=>"101001001",
  36372=>"010000011",
  36373=>"001111010",
  36374=>"000110111",
  36375=>"101000011",
  36376=>"011010011",
  36377=>"110101110",
  36378=>"000001011",
  36379=>"010000010",
  36380=>"010000100",
  36381=>"010011101",
  36382=>"000000111",
  36383=>"010111111",
  36384=>"001010111",
  36385=>"011100000",
  36386=>"001100111",
  36387=>"111111101",
  36388=>"010110000",
  36389=>"101001000",
  36390=>"010000101",
  36391=>"100101010",
  36392=>"001000011",
  36393=>"010111100",
  36394=>"011001001",
  36395=>"101001011",
  36396=>"101010000",
  36397=>"010100000",
  36398=>"001101110",
  36399=>"011000000",
  36400=>"010100111",
  36401=>"101001101",
  36402=>"101000001",
  36403=>"101001111",
  36404=>"011010100",
  36405=>"111101011",
  36406=>"001101100",
  36407=>"000001100",
  36408=>"101010101",
  36409=>"101010100",
  36410=>"111101101",
  36411=>"101011000",
  36412=>"010011010",
  36413=>"010100000",
  36414=>"011011000",
  36415=>"001011110",
  36416=>"000010111",
  36417=>"001101101",
  36418=>"011111110",
  36419=>"001110101",
  36420=>"011111101",
  36421=>"000111000",
  36422=>"110101111",
  36423=>"001000100",
  36424=>"010000111",
  36425=>"100110011",
  36426=>"110011110",
  36427=>"001110110",
  36428=>"101010111",
  36429=>"011110101",
  36430=>"101110000",
  36431=>"001011001",
  36432=>"111000110",
  36433=>"110100000",
  36434=>"101111110",
  36435=>"010110110",
  36436=>"011011010",
  36437=>"010000101",
  36438=>"000101001",
  36439=>"001000011",
  36440=>"110110000",
  36441=>"001101000",
  36442=>"001111111",
  36443=>"010010011",
  36444=>"110000101",
  36445=>"110011100",
  36446=>"011011101",
  36447=>"111001110",
  36448=>"010011011",
  36449=>"010000001",
  36450=>"111101000",
  36451=>"001000000",
  36452=>"011110001",
  36453=>"001101111",
  36454=>"100100101",
  36455=>"010101001",
  36456=>"001100100",
  36457=>"000010010",
  36458=>"111100110",
  36459=>"110010001",
  36460=>"101101111",
  36461=>"110000110",
  36462=>"100111100",
  36463=>"001101010",
  36464=>"011111011",
  36465=>"000011101",
  36466=>"101000110",
  36467=>"010011010",
  36468=>"111001111",
  36469=>"010100101",
  36470=>"100000000",
  36471=>"101100111",
  36472=>"000111010",
  36473=>"001101000",
  36474=>"100111000",
  36475=>"010001000",
  36476=>"001000100",
  36477=>"000010100",
  36478=>"111101111",
  36479=>"011111101",
  36480=>"101010100",
  36481=>"101010111",
  36482=>"000110110",
  36483=>"000001100",
  36484=>"000110001",
  36485=>"000011110",
  36486=>"100111010",
  36487=>"111101010",
  36488=>"011111000",
  36489=>"110010010",
  36490=>"010011110",
  36491=>"001101010",
  36492=>"110010011",
  36493=>"100000000",
  36494=>"010010000",
  36495=>"110101010",
  36496=>"010110010",
  36497=>"101000010",
  36498=>"111101000",
  36499=>"101001001",
  36500=>"100100101",
  36501=>"100100101",
  36502=>"001001000",
  36503=>"110000100",
  36504=>"010111001",
  36505=>"101000110",
  36506=>"110110001",
  36507=>"110111111",
  36508=>"101010101",
  36509=>"110001100",
  36510=>"100010010",
  36511=>"001110100",
  36512=>"100001000",
  36513=>"000001111",
  36514=>"101110110",
  36515=>"000000000",
  36516=>"110101010",
  36517=>"100001100",
  36518=>"110101101",
  36519=>"100010010",
  36520=>"011100100",
  36521=>"010010100",
  36522=>"101111100",
  36523=>"010010010",
  36524=>"111101100",
  36525=>"101011001",
  36526=>"001100110",
  36527=>"101010000",
  36528=>"100000110",
  36529=>"110100101",
  36530=>"100101100",
  36531=>"011111111",
  36532=>"000111110",
  36533=>"011101001",
  36534=>"100011110",
  36535=>"000111101",
  36536=>"010101010",
  36537=>"101101100",
  36538=>"111000100",
  36539=>"000110000",
  36540=>"110111001",
  36541=>"101001011",
  36542=>"000100101",
  36543=>"100011100",
  36544=>"011111111",
  36545=>"111101111",
  36546=>"100001100",
  36547=>"011100011",
  36548=>"011001111",
  36549=>"000010000",
  36550=>"101010100",
  36551=>"011110110",
  36552=>"111011010",
  36553=>"101110001",
  36554=>"111000110",
  36555=>"110111000",
  36556=>"110100010",
  36557=>"000011111",
  36558=>"000000000",
  36559=>"110001001",
  36560=>"101011101",
  36561=>"110101101",
  36562=>"101101111",
  36563=>"011011011",
  36564=>"001001011",
  36565=>"100000001",
  36566=>"100010111",
  36567=>"101001000",
  36568=>"010011010",
  36569=>"110111110",
  36570=>"100010000",
  36571=>"011010001",
  36572=>"001001111",
  36573=>"100101011",
  36574=>"010110100",
  36575=>"111101011",
  36576=>"110001100",
  36577=>"101011010",
  36578=>"001101010",
  36579=>"011100111",
  36580=>"001100111",
  36581=>"010101111",
  36582=>"101101101",
  36583=>"010101011",
  36584=>"100000000",
  36585=>"000110010",
  36586=>"100010000",
  36587=>"010000011",
  36588=>"000000010",
  36589=>"101010100",
  36590=>"010110111",
  36591=>"000110010",
  36592=>"000100010",
  36593=>"110111000",
  36594=>"000100101",
  36595=>"001010001",
  36596=>"100001111",
  36597=>"000101100",
  36598=>"101101110",
  36599=>"010011111",
  36600=>"101111101",
  36601=>"101100001",
  36602=>"010010001",
  36603=>"101000001",
  36604=>"100011101",
  36605=>"001100100",
  36606=>"001110111",
  36607=>"101111010",
  36608=>"001010101",
  36609=>"001001001",
  36610=>"100000011",
  36611=>"111000000",
  36612=>"000101110",
  36613=>"000101011",
  36614=>"011010011",
  36615=>"010100101",
  36616=>"110001101",
  36617=>"000011100",
  36618=>"000110000",
  36619=>"000110000",
  36620=>"110001000",
  36621=>"000001100",
  36622=>"101001000",
  36623=>"101100001",
  36624=>"010100010",
  36625=>"001101001",
  36626=>"100001001",
  36627=>"111010110",
  36628=>"111111001",
  36629=>"000001101",
  36630=>"110101011",
  36631=>"000111001",
  36632=>"011011101",
  36633=>"001110011",
  36634=>"010000111",
  36635=>"100011011",
  36636=>"001101101",
  36637=>"001100011",
  36638=>"001001000",
  36639=>"010010110",
  36640=>"110111011",
  36641=>"110110001",
  36642=>"100010010",
  36643=>"010101001",
  36644=>"100000010",
  36645=>"110010000",
  36646=>"111010101",
  36647=>"001000100",
  36648=>"111101111",
  36649=>"011011011",
  36650=>"111010101",
  36651=>"111100101",
  36652=>"101111000",
  36653=>"001110110",
  36654=>"011101101",
  36655=>"100110010",
  36656=>"100101101",
  36657=>"010100111",
  36658=>"101110011",
  36659=>"000100000",
  36660=>"101111001",
  36661=>"000010010",
  36662=>"000110100",
  36663=>"011101000",
  36664=>"101011101",
  36665=>"101001011",
  36666=>"011110101",
  36667=>"111100110",
  36668=>"100100010",
  36669=>"011101000",
  36670=>"111000000",
  36671=>"110011001",
  36672=>"000111001",
  36673=>"010001110",
  36674=>"110000001",
  36675=>"111100100",
  36676=>"111110110",
  36677=>"010011111",
  36678=>"100000011",
  36679=>"011000000",
  36680=>"011101111",
  36681=>"111101101",
  36682=>"010100001",
  36683=>"101100101",
  36684=>"101110010",
  36685=>"101011100",
  36686=>"100010100",
  36687=>"100011011",
  36688=>"100111100",
  36689=>"010100101",
  36690=>"000111001",
  36691=>"100011110",
  36692=>"100001010",
  36693=>"011000110",
  36694=>"011010101",
  36695=>"111111011",
  36696=>"011010001",
  36697=>"110000101",
  36698=>"100110111",
  36699=>"110101101",
  36700=>"011111011",
  36701=>"100111100",
  36702=>"101011110",
  36703=>"100000100",
  36704=>"011001011",
  36705=>"111101011",
  36706=>"101000111",
  36707=>"101001101",
  36708=>"010001111",
  36709=>"101111001",
  36710=>"011101110",
  36711=>"001000001",
  36712=>"011011101",
  36713=>"101100001",
  36714=>"010001101",
  36715=>"010000101",
  36716=>"101111000",
  36717=>"110110000",
  36718=>"010000000",
  36719=>"001101110",
  36720=>"101101000",
  36721=>"010110001",
  36722=>"001110000",
  36723=>"001010000",
  36724=>"100111011",
  36725=>"111010111",
  36726=>"100000011",
  36727=>"010001101",
  36728=>"110001001",
  36729=>"010110101",
  36730=>"100111000",
  36731=>"011110010",
  36732=>"100100110",
  36733=>"110100000",
  36734=>"100000001",
  36735=>"001101110",
  36736=>"011001100",
  36737=>"100111000",
  36738=>"010001011",
  36739=>"011000100",
  36740=>"010011111",
  36741=>"011100100",
  36742=>"000010100",
  36743=>"000110001",
  36744=>"000110010",
  36745=>"111100001",
  36746=>"000011101",
  36747=>"110111000",
  36748=>"010101001",
  36749=>"100010010",
  36750=>"011110110",
  36751=>"011101011",
  36752=>"101010111",
  36753=>"101000100",
  36754=>"001000000",
  36755=>"010001010",
  36756=>"001000101",
  36757=>"111001100",
  36758=>"011100001",
  36759=>"100110111",
  36760=>"101101011",
  36761=>"100011110",
  36762=>"011100010",
  36763=>"100001110",
  36764=>"101010001",
  36765=>"000101100",
  36766=>"001000111",
  36767=>"000010100",
  36768=>"110111101",
  36769=>"100101111",
  36770=>"100100100",
  36771=>"111100000",
  36772=>"000111110",
  36773=>"101001011",
  36774=>"010100001",
  36775=>"110110010",
  36776=>"011000100",
  36777=>"100011000",
  36778=>"011010001",
  36779=>"001100100",
  36780=>"010001000",
  36781=>"011001100",
  36782=>"100111001",
  36783=>"110100100",
  36784=>"111100100",
  36785=>"001101101",
  36786=>"111111110",
  36787=>"111000100",
  36788=>"011100110",
  36789=>"000000001",
  36790=>"111110010",
  36791=>"110100000",
  36792=>"110101011",
  36793=>"011011001",
  36794=>"011000011",
  36795=>"101011001",
  36796=>"110000011",
  36797=>"111011111",
  36798=>"110100001",
  36799=>"000000010",
  36800=>"100111011",
  36801=>"101001011",
  36802=>"100001100",
  36803=>"111010111",
  36804=>"001011110",
  36805=>"001010100",
  36806=>"101101110",
  36807=>"100110010",
  36808=>"000001010",
  36809=>"011101100",
  36810=>"010010100",
  36811=>"011011111",
  36812=>"001011000",
  36813=>"011010101",
  36814=>"010101101",
  36815=>"110111001",
  36816=>"010111111",
  36817=>"010011001",
  36818=>"000100011",
  36819=>"100110101",
  36820=>"001000000",
  36821=>"011011101",
  36822=>"001000001",
  36823=>"010001111",
  36824=>"100001110",
  36825=>"001010001",
  36826=>"111111111",
  36827=>"010011011",
  36828=>"100010101",
  36829=>"100001011",
  36830=>"011000101",
  36831=>"000011010",
  36832=>"111100100",
  36833=>"100011111",
  36834=>"111110010",
  36835=>"000111100",
  36836=>"101011000",
  36837=>"100111110",
  36838=>"001101101",
  36839=>"000100000",
  36840=>"000110100",
  36841=>"010010000",
  36842=>"001110110",
  36843=>"101000000",
  36844=>"010111010",
  36845=>"010101101",
  36846=>"010100111",
  36847=>"011111001",
  36848=>"110101011",
  36849=>"101011010",
  36850=>"110100111",
  36851=>"010111101",
  36852=>"101100100",
  36853=>"111111001",
  36854=>"010011010",
  36855=>"000101111",
  36856=>"100101111",
  36857=>"111000000",
  36858=>"101000100",
  36859=>"001010011",
  36860=>"111100011",
  36861=>"011110101",
  36862=>"111001001",
  36863=>"001000001",
  36864=>"000100110",
  36865=>"111010010",
  36866=>"010001111",
  36867=>"011100000",
  36868=>"111000111",
  36869=>"101011111",
  36870=>"000011101",
  36871=>"111111110",
  36872=>"100110001",
  36873=>"010100101",
  36874=>"010010111",
  36875=>"001101011",
  36876=>"011001011",
  36877=>"111111001",
  36878=>"110100010",
  36879=>"011101101",
  36880=>"011110101",
  36881=>"111000111",
  36882=>"000100101",
  36883=>"010101011",
  36884=>"111010011",
  36885=>"111011101",
  36886=>"111111111",
  36887=>"101110101",
  36888=>"110101101",
  36889=>"001000010",
  36890=>"001111011",
  36891=>"101000111",
  36892=>"110000000",
  36893=>"010010010",
  36894=>"001111110",
  36895=>"001100110",
  36896=>"001111011",
  36897=>"101101110",
  36898=>"010111010",
  36899=>"000100111",
  36900=>"111111011",
  36901=>"001000001",
  36902=>"000111111",
  36903=>"010100011",
  36904=>"010100101",
  36905=>"110100011",
  36906=>"110011000",
  36907=>"111110001",
  36908=>"100111110",
  36909=>"111100011",
  36910=>"111110100",
  36911=>"000111111",
  36912=>"100011110",
  36913=>"011111110",
  36914=>"001000100",
  36915=>"101001001",
  36916=>"010010110",
  36917=>"001110000",
  36918=>"100111011",
  36919=>"111111101",
  36920=>"010111001",
  36921=>"111101010",
  36922=>"101001011",
  36923=>"101011101",
  36924=>"000101100",
  36925=>"011110000",
  36926=>"101010101",
  36927=>"011011011",
  36928=>"110111111",
  36929=>"000111101",
  36930=>"111000000",
  36931=>"100001100",
  36932=>"111111011",
  36933=>"101101011",
  36934=>"010111111",
  36935=>"001110110",
  36936=>"111011100",
  36937=>"111000000",
  36938=>"010001001",
  36939=>"110111111",
  36940=>"011000110",
  36941=>"101000101",
  36942=>"101001000",
  36943=>"010111101",
  36944=>"000001010",
  36945=>"111000000",
  36946=>"110001001",
  36947=>"110101000",
  36948=>"011100000",
  36949=>"000100101",
  36950=>"101101011",
  36951=>"100101101",
  36952=>"101000110",
  36953=>"011100100",
  36954=>"000101000",
  36955=>"110100100",
  36956=>"100001100",
  36957=>"111011100",
  36958=>"000001010",
  36959=>"011100100",
  36960=>"101011101",
  36961=>"010010011",
  36962=>"001100101",
  36963=>"100010110",
  36964=>"111010001",
  36965=>"111101010",
  36966=>"100010100",
  36967=>"110001101",
  36968=>"111101011",
  36969=>"001111011",
  36970=>"101001011",
  36971=>"000001010",
  36972=>"100100001",
  36973=>"001100100",
  36974=>"010100000",
  36975=>"110010001",
  36976=>"110000000",
  36977=>"011110111",
  36978=>"011111100",
  36979=>"110101111",
  36980=>"001111001",
  36981=>"011100100",
  36982=>"001010000",
  36983=>"010100111",
  36984=>"001001111",
  36985=>"110111010",
  36986=>"001101101",
  36987=>"010101111",
  36988=>"010001111",
  36989=>"010010101",
  36990=>"001101100",
  36991=>"001000101",
  36992=>"110010100",
  36993=>"011101100",
  36994=>"000010000",
  36995=>"000000000",
  36996=>"100100111",
  36997=>"111111111",
  36998=>"010000100",
  36999=>"101011010",
  37000=>"001000100",
  37001=>"101111100",
  37002=>"011010111",
  37003=>"111110100",
  37004=>"100011010",
  37005=>"001000010",
  37006=>"010011111",
  37007=>"111011000",
  37008=>"110011100",
  37009=>"011101000",
  37010=>"101000000",
  37011=>"110010100",
  37012=>"111100110",
  37013=>"011111000",
  37014=>"000100011",
  37015=>"111111011",
  37016=>"001111000",
  37017=>"001011111",
  37018=>"001100100",
  37019=>"111100011",
  37020=>"001101011",
  37021=>"011011110",
  37022=>"110101011",
  37023=>"000001100",
  37024=>"001011100",
  37025=>"110101101",
  37026=>"000010111",
  37027=>"011001000",
  37028=>"100010000",
  37029=>"111100000",
  37030=>"110101111",
  37031=>"010111110",
  37032=>"001100000",
  37033=>"000100110",
  37034=>"101100110",
  37035=>"011010101",
  37036=>"011011101",
  37037=>"000111001",
  37038=>"100100100",
  37039=>"111010011",
  37040=>"011101001",
  37041=>"001111010",
  37042=>"111100010",
  37043=>"111000001",
  37044=>"101001011",
  37045=>"001010011",
  37046=>"010111010",
  37047=>"110011101",
  37048=>"111001011",
  37049=>"011101010",
  37050=>"101111011",
  37051=>"111111001",
  37052=>"100101011",
  37053=>"101110110",
  37054=>"111011000",
  37055=>"100000001",
  37056=>"011001000",
  37057=>"011010010",
  37058=>"000011100",
  37059=>"110100010",
  37060=>"000100111",
  37061=>"001001111",
  37062=>"100110111",
  37063=>"000100001",
  37064=>"111101000",
  37065=>"001010010",
  37066=>"010101010",
  37067=>"000010110",
  37068=>"001001000",
  37069=>"010110110",
  37070=>"111111101",
  37071=>"110110001",
  37072=>"110111100",
  37073=>"100011101",
  37074=>"000010010",
  37075=>"101000111",
  37076=>"100000010",
  37077=>"101011101",
  37078=>"010001111",
  37079=>"011101000",
  37080=>"101101001",
  37081=>"101000111",
  37082=>"011111001",
  37083=>"011100010",
  37084=>"011111111",
  37085=>"010111110",
  37086=>"101100011",
  37087=>"110010111",
  37088=>"111011101",
  37089=>"110110101",
  37090=>"111011111",
  37091=>"001011000",
  37092=>"111000001",
  37093=>"110111101",
  37094=>"001001101",
  37095=>"101011111",
  37096=>"100111111",
  37097=>"101000110",
  37098=>"101001101",
  37099=>"011011001",
  37100=>"101011001",
  37101=>"000011111",
  37102=>"110101011",
  37103=>"001011001",
  37104=>"001100111",
  37105=>"111001000",
  37106=>"001110110",
  37107=>"100010000",
  37108=>"000000101",
  37109=>"011100111",
  37110=>"001101110",
  37111=>"000101000",
  37112=>"001011111",
  37113=>"011010100",
  37114=>"000100001",
  37115=>"000011010",
  37116=>"111011111",
  37117=>"001010001",
  37118=>"001000010",
  37119=>"110101010",
  37120=>"010111101",
  37121=>"110011011",
  37122=>"001000100",
  37123=>"000100001",
  37124=>"100000111",
  37125=>"011001001",
  37126=>"101101001",
  37127=>"111001110",
  37128=>"110000100",
  37129=>"110101101",
  37130=>"110011011",
  37131=>"101001101",
  37132=>"000111001",
  37133=>"000011111",
  37134=>"111111111",
  37135=>"011101111",
  37136=>"101110111",
  37137=>"111011001",
  37138=>"111010100",
  37139=>"110100011",
  37140=>"011000101",
  37141=>"000100001",
  37142=>"000111101",
  37143=>"011110110",
  37144=>"101011111",
  37145=>"000000100",
  37146=>"111010110",
  37147=>"010111001",
  37148=>"010010011",
  37149=>"111100010",
  37150=>"110010001",
  37151=>"101011011",
  37152=>"100111010",
  37153=>"111011011",
  37154=>"100011101",
  37155=>"110010101",
  37156=>"001100101",
  37157=>"011101101",
  37158=>"101011010",
  37159=>"101111010",
  37160=>"000001111",
  37161=>"000100101",
  37162=>"111100011",
  37163=>"000001110",
  37164=>"001010010",
  37165=>"001010110",
  37166=>"100110101",
  37167=>"111101001",
  37168=>"010101001",
  37169=>"001101010",
  37170=>"011001111",
  37171=>"100010111",
  37172=>"011001011",
  37173=>"001100011",
  37174=>"011011101",
  37175=>"010100010",
  37176=>"010000111",
  37177=>"000111011",
  37178=>"100011100",
  37179=>"100010100",
  37180=>"001100101",
  37181=>"001000110",
  37182=>"110111111",
  37183=>"111011010",
  37184=>"000011011",
  37185=>"100111000",
  37186=>"100000001",
  37187=>"001000011",
  37188=>"111111100",
  37189=>"100101011",
  37190=>"001000100",
  37191=>"110110001",
  37192=>"000011110",
  37193=>"011001100",
  37194=>"101111110",
  37195=>"001001111",
  37196=>"010000011",
  37197=>"001000010",
  37198=>"111011100",
  37199=>"111001100",
  37200=>"110011101",
  37201=>"101100101",
  37202=>"000001111",
  37203=>"000001111",
  37204=>"000111011",
  37205=>"111110100",
  37206=>"001001010",
  37207=>"101000000",
  37208=>"110101010",
  37209=>"111100111",
  37210=>"011101111",
  37211=>"100101111",
  37212=>"001111011",
  37213=>"000011100",
  37214=>"010000000",
  37215=>"111100100",
  37216=>"001110101",
  37217=>"110001010",
  37218=>"011000111",
  37219=>"101010000",
  37220=>"000001001",
  37221=>"010100111",
  37222=>"011101111",
  37223=>"011010100",
  37224=>"111011111",
  37225=>"010010111",
  37226=>"110011001",
  37227=>"000111110",
  37228=>"001011100",
  37229=>"100010101",
  37230=>"000011000",
  37231=>"010101000",
  37232=>"000101001",
  37233=>"001111010",
  37234=>"110100011",
  37235=>"100100000",
  37236=>"001101001",
  37237=>"100100000",
  37238=>"101010001",
  37239=>"111110101",
  37240=>"111000001",
  37241=>"111101111",
  37242=>"100011111",
  37243=>"010101111",
  37244=>"000111001",
  37245=>"000010000",
  37246=>"011111011",
  37247=>"101111101",
  37248=>"000000110",
  37249=>"010011011",
  37250=>"010011101",
  37251=>"000010001",
  37252=>"110101011",
  37253=>"011101000",
  37254=>"111000111",
  37255=>"111011011",
  37256=>"010000111",
  37257=>"010010101",
  37258=>"010011011",
  37259=>"000110011",
  37260=>"000100010",
  37261=>"101110111",
  37262=>"100101000",
  37263=>"011100101",
  37264=>"011001000",
  37265=>"101101010",
  37266=>"111000011",
  37267=>"011110010",
  37268=>"001111001",
  37269=>"101000000",
  37270=>"010101110",
  37271=>"101001001",
  37272=>"100111010",
  37273=>"001000001",
  37274=>"101100100",
  37275=>"111101101",
  37276=>"110100101",
  37277=>"000001101",
  37278=>"000111001",
  37279=>"100001001",
  37280=>"101011111",
  37281=>"000110111",
  37282=>"001001000",
  37283=>"111101000",
  37284=>"001101111",
  37285=>"101110001",
  37286=>"001001111",
  37287=>"110111001",
  37288=>"001100010",
  37289=>"101001011",
  37290=>"101100101",
  37291=>"000000110",
  37292=>"000110001",
  37293=>"100101111",
  37294=>"110111101",
  37295=>"101011001",
  37296=>"100100111",
  37297=>"010001011",
  37298=>"100100111",
  37299=>"000111101",
  37300=>"111000100",
  37301=>"100101110",
  37302=>"001010001",
  37303=>"100100111",
  37304=>"111001011",
  37305=>"011010011",
  37306=>"001000011",
  37307=>"001000011",
  37308=>"001000110",
  37309=>"110101111",
  37310=>"010000101",
  37311=>"001111111",
  37312=>"011111101",
  37313=>"000110111",
  37314=>"010100011",
  37315=>"011011000",
  37316=>"011110011",
  37317=>"101101101",
  37318=>"011010101",
  37319=>"111111110",
  37320=>"001010100",
  37321=>"000000110",
  37322=>"010001001",
  37323=>"111001001",
  37324=>"101111101",
  37325=>"001000111",
  37326=>"001001111",
  37327=>"000100111",
  37328=>"010010111",
  37329=>"001101000",
  37330=>"010000000",
  37331=>"010001000",
  37332=>"111111110",
  37333=>"101101101",
  37334=>"100001011",
  37335=>"101011001",
  37336=>"100000101",
  37337=>"101110101",
  37338=>"011011000",
  37339=>"110000000",
  37340=>"110000110",
  37341=>"101100001",
  37342=>"010010101",
  37343=>"111111100",
  37344=>"111001100",
  37345=>"001000011",
  37346=>"110001010",
  37347=>"010101000",
  37348=>"100001100",
  37349=>"010001001",
  37350=>"101110000",
  37351=>"011000000",
  37352=>"001101100",
  37353=>"001001001",
  37354=>"101000001",
  37355=>"000111101",
  37356=>"010001011",
  37357=>"100010001",
  37358=>"000000000",
  37359=>"110110000",
  37360=>"100101100",
  37361=>"000101100",
  37362=>"111110111",
  37363=>"111010110",
  37364=>"100011100",
  37365=>"000110011",
  37366=>"001001000",
  37367=>"001010110",
  37368=>"101011001",
  37369=>"010001001",
  37370=>"110110101",
  37371=>"011001101",
  37372=>"010000111",
  37373=>"011011010",
  37374=>"001010110",
  37375=>"111101111",
  37376=>"111001000",
  37377=>"101000001",
  37378=>"100000110",
  37379=>"100101011",
  37380=>"110011001",
  37381=>"000000100",
  37382=>"100111101",
  37383=>"111110111",
  37384=>"001100101",
  37385=>"001111100",
  37386=>"000101010",
  37387=>"100000011",
  37388=>"110110111",
  37389=>"000100100",
  37390=>"110000000",
  37391=>"010000001",
  37392=>"011101010",
  37393=>"011010111",
  37394=>"110001101",
  37395=>"111011000",
  37396=>"101010000",
  37397=>"001001000",
  37398=>"001110101",
  37399=>"001000100",
  37400=>"111111100",
  37401=>"011110011",
  37402=>"010100100",
  37403=>"101111001",
  37404=>"011111110",
  37405=>"100001000",
  37406=>"111010111",
  37407=>"101101100",
  37408=>"011111111",
  37409=>"111100000",
  37410=>"000000010",
  37411=>"101000111",
  37412=>"111000111",
  37413=>"001010111",
  37414=>"110011110",
  37415=>"011001011",
  37416=>"011101111",
  37417=>"000100100",
  37418=>"000010011",
  37419=>"011101011",
  37420=>"010110001",
  37421=>"001110100",
  37422=>"110110010",
  37423=>"110011010",
  37424=>"111001101",
  37425=>"111010101",
  37426=>"010000010",
  37427=>"001111000",
  37428=>"010110001",
  37429=>"000001110",
  37430=>"101001011",
  37431=>"101001010",
  37432=>"011001011",
  37433=>"100100101",
  37434=>"110011011",
  37435=>"100000100",
  37436=>"110110111",
  37437=>"011001000",
  37438=>"010100000",
  37439=>"000111100",
  37440=>"011000001",
  37441=>"011000101",
  37442=>"100111110",
  37443=>"010010100",
  37444=>"101001110",
  37445=>"000000111",
  37446=>"110010000",
  37447=>"100001011",
  37448=>"011010010",
  37449=>"001001001",
  37450=>"011110100",
  37451=>"000001101",
  37452=>"000011001",
  37453=>"100111001",
  37454=>"111101000",
  37455=>"100011111",
  37456=>"000101111",
  37457=>"110001000",
  37458=>"100000101",
  37459=>"110001111",
  37460=>"010100000",
  37461=>"111010110",
  37462=>"101011101",
  37463=>"010010010",
  37464=>"111010011",
  37465=>"111100000",
  37466=>"000111011",
  37467=>"100111011",
  37468=>"111101001",
  37469=>"100101000",
  37470=>"110000101",
  37471=>"111011101",
  37472=>"111101011",
  37473=>"000010001",
  37474=>"001110101",
  37475=>"000010110",
  37476=>"010010011",
  37477=>"110010010",
  37478=>"001011011",
  37479=>"110010011",
  37480=>"000010001",
  37481=>"101010111",
  37482=>"100000100",
  37483=>"111100000",
  37484=>"000011000",
  37485=>"000100101",
  37486=>"001010111",
  37487=>"101000010",
  37488=>"011100110",
  37489=>"001110010",
  37490=>"110010111",
  37491=>"001000010",
  37492=>"000001100",
  37493=>"010101100",
  37494=>"001111010",
  37495=>"111010101",
  37496=>"011100111",
  37497=>"010101101",
  37498=>"111000000",
  37499=>"011101101",
  37500=>"111111101",
  37501=>"011101100",
  37502=>"000110010",
  37503=>"001001010",
  37504=>"110010011",
  37505=>"001010100",
  37506=>"110001101",
  37507=>"001000110",
  37508=>"001100111",
  37509=>"001001101",
  37510=>"010101111",
  37511=>"110110101",
  37512=>"100001011",
  37513=>"100001101",
  37514=>"011110011",
  37515=>"000001011",
  37516=>"011110011",
  37517=>"010011111",
  37518=>"110100001",
  37519=>"110110110",
  37520=>"101000001",
  37521=>"001111110",
  37522=>"111010110",
  37523=>"100110001",
  37524=>"111011011",
  37525=>"100000110",
  37526=>"110000010",
  37527=>"001100010",
  37528=>"101001001",
  37529=>"110010010",
  37530=>"110100010",
  37531=>"100111111",
  37532=>"000101000",
  37533=>"100010010",
  37534=>"010100001",
  37535=>"111111111",
  37536=>"110001101",
  37537=>"110010011",
  37538=>"111111010",
  37539=>"001001011",
  37540=>"000101111",
  37541=>"010100010",
  37542=>"101000000",
  37543=>"011010110",
  37544=>"111011100",
  37545=>"000000011",
  37546=>"010110100",
  37547=>"101010011",
  37548=>"101100111",
  37549=>"001000000",
  37550=>"110101110",
  37551=>"110011000",
  37552=>"110110011",
  37553=>"001010111",
  37554=>"000100111",
  37555=>"001101011",
  37556=>"111011101",
  37557=>"011100011",
  37558=>"010001101",
  37559=>"100111011",
  37560=>"011111110",
  37561=>"101000101",
  37562=>"011110101",
  37563=>"111011011",
  37564=>"100100100",
  37565=>"010000111",
  37566=>"100100101",
  37567=>"000001110",
  37568=>"000010010",
  37569=>"010011111",
  37570=>"000011111",
  37571=>"100101010",
  37572=>"010001000",
  37573=>"111100111",
  37574=>"111100101",
  37575=>"001111011",
  37576=>"100000010",
  37577=>"110100101",
  37578=>"011110110",
  37579=>"000011101",
  37580=>"110000001",
  37581=>"111110110",
  37582=>"101010011",
  37583=>"011101011",
  37584=>"110011001",
  37585=>"010111001",
  37586=>"110011000",
  37587=>"001100001",
  37588=>"100111001",
  37589=>"111000111",
  37590=>"100100000",
  37591=>"101101111",
  37592=>"100111011",
  37593=>"101111110",
  37594=>"000111011",
  37595=>"011001011",
  37596=>"000010010",
  37597=>"001011101",
  37598=>"011011110",
  37599=>"110110100",
  37600=>"011010101",
  37601=>"011000001",
  37602=>"011011000",
  37603=>"101000010",
  37604=>"011101001",
  37605=>"101101110",
  37606=>"001100111",
  37607=>"100000100",
  37608=>"011011100",
  37609=>"010111101",
  37610=>"110111010",
  37611=>"011101000",
  37612=>"001010100",
  37613=>"011011010",
  37614=>"010110010",
  37615=>"001000001",
  37616=>"011001000",
  37617=>"110011001",
  37618=>"010011000",
  37619=>"000100110",
  37620=>"100000100",
  37621=>"111100000",
  37622=>"000110110",
  37623=>"000010111",
  37624=>"001001110",
  37625=>"111010111",
  37626=>"100000010",
  37627=>"001101110",
  37628=>"101101110",
  37629=>"001000001",
  37630=>"110101100",
  37631=>"111110011",
  37632=>"100111111",
  37633=>"001011011",
  37634=>"001011000",
  37635=>"001101100",
  37636=>"010100111",
  37637=>"100000100",
  37638=>"000111000",
  37639=>"111111110",
  37640=>"110100101",
  37641=>"000001010",
  37642=>"001100110",
  37643=>"000100001",
  37644=>"010010000",
  37645=>"100000101",
  37646=>"000011110",
  37647=>"010011010",
  37648=>"001110111",
  37649=>"010110010",
  37650=>"011101001",
  37651=>"000110000",
  37652=>"110011011",
  37653=>"111000011",
  37654=>"001110101",
  37655=>"001001100",
  37656=>"110110110",
  37657=>"000000101",
  37658=>"001100111",
  37659=>"001110110",
  37660=>"111111110",
  37661=>"111001011",
  37662=>"100011100",
  37663=>"011010000",
  37664=>"100111101",
  37665=>"001000100",
  37666=>"010000001",
  37667=>"010001100",
  37668=>"001010000",
  37669=>"110111011",
  37670=>"111101111",
  37671=>"101000010",
  37672=>"010001110",
  37673=>"111000011",
  37674=>"110000011",
  37675=>"101100110",
  37676=>"000011000",
  37677=>"101111101",
  37678=>"000101011",
  37679=>"000111101",
  37680=>"111111101",
  37681=>"000101101",
  37682=>"010001110",
  37683=>"111001100",
  37684=>"111010010",
  37685=>"111011101",
  37686=>"101010011",
  37687=>"100000100",
  37688=>"111000000",
  37689=>"001111111",
  37690=>"110001100",
  37691=>"000001011",
  37692=>"101100100",
  37693=>"011011000",
  37694=>"001100001",
  37695=>"010000101",
  37696=>"011000000",
  37697=>"000010011",
  37698=>"000111001",
  37699=>"110001100",
  37700=>"011111001",
  37701=>"101010001",
  37702=>"110111101",
  37703=>"110000111",
  37704=>"111000111",
  37705=>"110111101",
  37706=>"101101001",
  37707=>"010010011",
  37708=>"010101011",
  37709=>"110111001",
  37710=>"100010111",
  37711=>"010111011",
  37712=>"011111000",
  37713=>"100101100",
  37714=>"101011111",
  37715=>"000010110",
  37716=>"000001101",
  37717=>"110110100",
  37718=>"011100000",
  37719=>"101011000",
  37720=>"010100000",
  37721=>"111110010",
  37722=>"110110110",
  37723=>"100100111",
  37724=>"011000111",
  37725=>"111100000",
  37726=>"110110011",
  37727=>"010101111",
  37728=>"000000100",
  37729=>"101101111",
  37730=>"100100110",
  37731=>"001110000",
  37732=>"000100010",
  37733=>"000001111",
  37734=>"001111011",
  37735=>"111101110",
  37736=>"110001110",
  37737=>"110111001",
  37738=>"010100111",
  37739=>"000100111",
  37740=>"100110100",
  37741=>"111010011",
  37742=>"111001110",
  37743=>"111010110",
  37744=>"000000001",
  37745=>"011100111",
  37746=>"100100111",
  37747=>"010011101",
  37748=>"010010011",
  37749=>"000001011",
  37750=>"110111010",
  37751=>"101111000",
  37752=>"100101011",
  37753=>"101110111",
  37754=>"011011011",
  37755=>"101010011",
  37756=>"000110000",
  37757=>"101111000",
  37758=>"100010110",
  37759=>"001000000",
  37760=>"110101111",
  37761=>"000011010",
  37762=>"010000101",
  37763=>"001010111",
  37764=>"101011111",
  37765=>"100000010",
  37766=>"111101101",
  37767=>"000101001",
  37768=>"001011110",
  37769=>"101100000",
  37770=>"011010010",
  37771=>"001011111",
  37772=>"101001000",
  37773=>"110011011",
  37774=>"001111111",
  37775=>"110000110",
  37776=>"100111110",
  37777=>"111000000",
  37778=>"000101000",
  37779=>"011001100",
  37780=>"000100110",
  37781=>"110010110",
  37782=>"000010000",
  37783=>"000111101",
  37784=>"101100100",
  37785=>"100110000",
  37786=>"110111001",
  37787=>"100100011",
  37788=>"101001100",
  37789=>"001010110",
  37790=>"111010000",
  37791=>"010110100",
  37792=>"110001001",
  37793=>"001100000",
  37794=>"011101111",
  37795=>"001111011",
  37796=>"000000100",
  37797=>"011111011",
  37798=>"000111001",
  37799=>"010001000",
  37800=>"100011001",
  37801=>"010101001",
  37802=>"000010110",
  37803=>"101100001",
  37804=>"110011111",
  37805=>"000011111",
  37806=>"010000100",
  37807=>"101100101",
  37808=>"111101001",
  37809=>"111001000",
  37810=>"101000011",
  37811=>"111110000",
  37812=>"101000101",
  37813=>"010011101",
  37814=>"100010011",
  37815=>"011110101",
  37816=>"011001010",
  37817=>"100000010",
  37818=>"111101100",
  37819=>"110000010",
  37820=>"101111100",
  37821=>"011000000",
  37822=>"010010011",
  37823=>"000100000",
  37824=>"101110001",
  37825=>"011110101",
  37826=>"110101110",
  37827=>"000010101",
  37828=>"101100000",
  37829=>"010001001",
  37830=>"011011000",
  37831=>"100111010",
  37832=>"011001000",
  37833=>"010100000",
  37834=>"100010100",
  37835=>"101011101",
  37836=>"110110110",
  37837=>"001001001",
  37838=>"111100101",
  37839=>"001100000",
  37840=>"100000000",
  37841=>"011101100",
  37842=>"011111010",
  37843=>"101011001",
  37844=>"101101000",
  37845=>"001100010",
  37846=>"000000100",
  37847=>"110000001",
  37848=>"100110000",
  37849=>"110111011",
  37850=>"010100111",
  37851=>"111010011",
  37852=>"101110111",
  37853=>"010000011",
  37854=>"010000000",
  37855=>"010000000",
  37856=>"111000101",
  37857=>"011101111",
  37858=>"010000101",
  37859=>"000000001",
  37860=>"011111011",
  37861=>"100000110",
  37862=>"111011101",
  37863=>"110111011",
  37864=>"111010101",
  37865=>"110111001",
  37866=>"010111001",
  37867=>"100110101",
  37868=>"100010011",
  37869=>"001101000",
  37870=>"000100000",
  37871=>"000000000",
  37872=>"011011110",
  37873=>"010110110",
  37874=>"111000100",
  37875=>"101100111",
  37876=>"100110000",
  37877=>"010110110",
  37878=>"000110010",
  37879=>"000000101",
  37880=>"001110110",
  37881=>"101000001",
  37882=>"111110001",
  37883=>"010001011",
  37884=>"010100001",
  37885=>"111100000",
  37886=>"010000101",
  37887=>"000011000",
  37888=>"111101110",
  37889=>"010010110",
  37890=>"101001011",
  37891=>"000001001",
  37892=>"111011101",
  37893=>"011111001",
  37894=>"001111010",
  37895=>"001000100",
  37896=>"111001100",
  37897=>"101110011",
  37898=>"010101001",
  37899=>"000101011",
  37900=>"101000111",
  37901=>"110011111",
  37902=>"010000010",
  37903=>"000010000",
  37904=>"010001111",
  37905=>"000110000",
  37906=>"010100100",
  37907=>"000111110",
  37908=>"111010110",
  37909=>"011000111",
  37910=>"101110011",
  37911=>"010000010",
  37912=>"110110010",
  37913=>"101110011",
  37914=>"011110001",
  37915=>"100111110",
  37916=>"100101100",
  37917=>"010010111",
  37918=>"000110000",
  37919=>"110010010",
  37920=>"100011111",
  37921=>"111101110",
  37922=>"100000101",
  37923=>"111010101",
  37924=>"011100011",
  37925=>"001001101",
  37926=>"010111101",
  37927=>"111111011",
  37928=>"111101010",
  37929=>"101111110",
  37930=>"101011001",
  37931=>"110011001",
  37932=>"011010101",
  37933=>"100011100",
  37934=>"001101111",
  37935=>"111000001",
  37936=>"000110001",
  37937=>"110001101",
  37938=>"000111000",
  37939=>"101011001",
  37940=>"111001100",
  37941=>"001111101",
  37942=>"111100011",
  37943=>"000011001",
  37944=>"010000111",
  37945=>"110011011",
  37946=>"111101110",
  37947=>"010010100",
  37948=>"000001000",
  37949=>"011001111",
  37950=>"111100000",
  37951=>"011101011",
  37952=>"110000100",
  37953=>"000010111",
  37954=>"010100001",
  37955=>"000010100",
  37956=>"111111110",
  37957=>"111000111",
  37958=>"000000000",
  37959=>"010000001",
  37960=>"111011101",
  37961=>"111101001",
  37962=>"110001110",
  37963=>"111010010",
  37964=>"110001110",
  37965=>"101010001",
  37966=>"000111111",
  37967=>"011010011",
  37968=>"010000010",
  37969=>"011101110",
  37970=>"100010111",
  37971=>"100000110",
  37972=>"111001110",
  37973=>"111000110",
  37974=>"101000100",
  37975=>"100001001",
  37976=>"001000100",
  37977=>"011001011",
  37978=>"000100110",
  37979=>"101110110",
  37980=>"110010010",
  37981=>"000001101",
  37982=>"110010001",
  37983=>"010000100",
  37984=>"001101100",
  37985=>"110010010",
  37986=>"101110001",
  37987=>"001001110",
  37988=>"110001110",
  37989=>"100000011",
  37990=>"100100000",
  37991=>"000001101",
  37992=>"010010110",
  37993=>"100110100",
  37994=>"111000110",
  37995=>"010100111",
  37996=>"011001011",
  37997=>"010110110",
  37998=>"100011010",
  37999=>"111100111",
  38000=>"010011110",
  38001=>"110001111",
  38002=>"010110000",
  38003=>"111011101",
  38004=>"011110101",
  38005=>"010000100",
  38006=>"001100100",
  38007=>"110010101",
  38008=>"001111100",
  38009=>"110001010",
  38010=>"101110001",
  38011=>"000100100",
  38012=>"110110000",
  38013=>"100110110",
  38014=>"111011111",
  38015=>"110100000",
  38016=>"000110111",
  38017=>"000010110",
  38018=>"110101001",
  38019=>"000110110",
  38020=>"011100000",
  38021=>"101110110",
  38022=>"110111101",
  38023=>"111101101",
  38024=>"010000001",
  38025=>"001111000",
  38026=>"000110110",
  38027=>"011000001",
  38028=>"101000011",
  38029=>"100100100",
  38030=>"010000000",
  38031=>"110100110",
  38032=>"101001110",
  38033=>"010110100",
  38034=>"111100010",
  38035=>"011101011",
  38036=>"001010100",
  38037=>"111010101",
  38038=>"011100110",
  38039=>"011100001",
  38040=>"001000101",
  38041=>"000101011",
  38042=>"000110010",
  38043=>"001001111",
  38044=>"010010001",
  38045=>"010000001",
  38046=>"110001110",
  38047=>"111100100",
  38048=>"111001101",
  38049=>"110110011",
  38050=>"100101110",
  38051=>"001000100",
  38052=>"001101110",
  38053=>"001100010",
  38054=>"001000100",
  38055=>"101000010",
  38056=>"011000011",
  38057=>"000100111",
  38058=>"101001000",
  38059=>"010100000",
  38060=>"100100011",
  38061=>"111101101",
  38062=>"101111011",
  38063=>"000100111",
  38064=>"011000100",
  38065=>"001110110",
  38066=>"111101111",
  38067=>"111111000",
  38068=>"010010110",
  38069=>"011101111",
  38070=>"110101110",
  38071=>"000010111",
  38072=>"111010101",
  38073=>"011100100",
  38074=>"010101001",
  38075=>"001101100",
  38076=>"010001110",
  38077=>"010101010",
  38078=>"010110110",
  38079=>"111011111",
  38080=>"010010010",
  38081=>"011101111",
  38082=>"001100000",
  38083=>"110001101",
  38084=>"101111100",
  38085=>"100001001",
  38086=>"000000001",
  38087=>"010010111",
  38088=>"011100011",
  38089=>"111110100",
  38090=>"011100100",
  38091=>"111100111",
  38092=>"000111001",
  38093=>"100100000",
  38094=>"110100110",
  38095=>"110000000",
  38096=>"011000011",
  38097=>"001010100",
  38098=>"011111110",
  38099=>"001000110",
  38100=>"110000011",
  38101=>"010011000",
  38102=>"011010101",
  38103=>"011011101",
  38104=>"100001011",
  38105=>"001111001",
  38106=>"011110100",
  38107=>"010011110",
  38108=>"101010001",
  38109=>"101111011",
  38110=>"110111100",
  38111=>"110011100",
  38112=>"000001110",
  38113=>"101010111",
  38114=>"000001100",
  38115=>"001001000",
  38116=>"011000011",
  38117=>"001010001",
  38118=>"011101000",
  38119=>"010011100",
  38120=>"001000111",
  38121=>"011101011",
  38122=>"100100101",
  38123=>"100100101",
  38124=>"101101101",
  38125=>"001011011",
  38126=>"011000101",
  38127=>"111111000",
  38128=>"000011110",
  38129=>"101011111",
  38130=>"001000000",
  38131=>"011000101",
  38132=>"011101100",
  38133=>"000101110",
  38134=>"010000000",
  38135=>"010000110",
  38136=>"111011110",
  38137=>"001001101",
  38138=>"010010110",
  38139=>"110001100",
  38140=>"011001011",
  38141=>"110111001",
  38142=>"011000001",
  38143=>"101001110",
  38144=>"111111011",
  38145=>"011110101",
  38146=>"101001000",
  38147=>"101111101",
  38148=>"100010111",
  38149=>"011110100",
  38150=>"000101100",
  38151=>"010011111",
  38152=>"001011001",
  38153=>"001100011",
  38154=>"010101000",
  38155=>"111010000",
  38156=>"000100110",
  38157=>"010001011",
  38158=>"100101101",
  38159=>"111010110",
  38160=>"110010000",
  38161=>"100010110",
  38162=>"111001111",
  38163=>"010011110",
  38164=>"110110000",
  38165=>"100001000",
  38166=>"101000000",
  38167=>"101011010",
  38168=>"110001010",
  38169=>"010001101",
  38170=>"010010011",
  38171=>"100010011",
  38172=>"000100111",
  38173=>"110011001",
  38174=>"111001101",
  38175=>"010000101",
  38176=>"101111111",
  38177=>"010101011",
  38178=>"010110011",
  38179=>"101100011",
  38180=>"010001010",
  38181=>"001001100",
  38182=>"110101101",
  38183=>"101000110",
  38184=>"111110101",
  38185=>"001100100",
  38186=>"011011000",
  38187=>"011001011",
  38188=>"111010001",
  38189=>"001001110",
  38190=>"100100110",
  38191=>"110100011",
  38192=>"111111111",
  38193=>"010100101",
  38194=>"111010001",
  38195=>"110100111",
  38196=>"100011110",
  38197=>"100111101",
  38198=>"111000000",
  38199=>"110001100",
  38200=>"100101111",
  38201=>"101000000",
  38202=>"011110001",
  38203=>"001011110",
  38204=>"010011001",
  38205=>"100001101",
  38206=>"001011011",
  38207=>"000010011",
  38208=>"001010010",
  38209=>"011110101",
  38210=>"000000110",
  38211=>"110110110",
  38212=>"101010010",
  38213=>"000111010",
  38214=>"100011000",
  38215=>"100101110",
  38216=>"000001001",
  38217=>"111010101",
  38218=>"010101001",
  38219=>"000100001",
  38220=>"000110000",
  38221=>"010011010",
  38222=>"011101000",
  38223=>"000010100",
  38224=>"110100000",
  38225=>"111111010",
  38226=>"100111011",
  38227=>"101111001",
  38228=>"101110010",
  38229=>"000010110",
  38230=>"111000100",
  38231=>"011101111",
  38232=>"001100110",
  38233=>"010001000",
  38234=>"000110110",
  38235=>"110111100",
  38236=>"101011010",
  38237=>"101110101",
  38238=>"001011000",
  38239=>"110001100",
  38240=>"110110000",
  38241=>"100000110",
  38242=>"100100101",
  38243=>"000011011",
  38244=>"101010000",
  38245=>"100100001",
  38246=>"011110101",
  38247=>"101000001",
  38248=>"100010110",
  38249=>"001100100",
  38250=>"110111001",
  38251=>"110000010",
  38252=>"111101000",
  38253=>"110000011",
  38254=>"111110101",
  38255=>"101110011",
  38256=>"011010011",
  38257=>"001011101",
  38258=>"111000111",
  38259=>"100100010",
  38260=>"100000111",
  38261=>"100111001",
  38262=>"000001110",
  38263=>"011011010",
  38264=>"010011010",
  38265=>"011101010",
  38266=>"001001010",
  38267=>"110111110",
  38268=>"001111100",
  38269=>"111110111",
  38270=>"001101010",
  38271=>"100000101",
  38272=>"110101111",
  38273=>"100010010",
  38274=>"100011011",
  38275=>"111010111",
  38276=>"100011001",
  38277=>"101111111",
  38278=>"011000011",
  38279=>"110000000",
  38280=>"011110001",
  38281=>"001111010",
  38282=>"110111111",
  38283=>"111100111",
  38284=>"100101110",
  38285=>"101111001",
  38286=>"100010111",
  38287=>"101110111",
  38288=>"010001000",
  38289=>"101001001",
  38290=>"100100011",
  38291=>"101000110",
  38292=>"011111111",
  38293=>"000001011",
  38294=>"110111010",
  38295=>"011100011",
  38296=>"111111101",
  38297=>"101011000",
  38298=>"100101101",
  38299=>"101000010",
  38300=>"110101011",
  38301=>"011010111",
  38302=>"100100010",
  38303=>"110011100",
  38304=>"001111100",
  38305=>"100111101",
  38306=>"000100111",
  38307=>"101100101",
  38308=>"010110010",
  38309=>"101000000",
  38310=>"001111010",
  38311=>"100011001",
  38312=>"111010001",
  38313=>"010100001",
  38314=>"010111110",
  38315=>"001001001",
  38316=>"000011101",
  38317=>"110100011",
  38318=>"110001101",
  38319=>"001010000",
  38320=>"000010001",
  38321=>"110110011",
  38322=>"010001011",
  38323=>"100110111",
  38324=>"001100000",
  38325=>"110010010",
  38326=>"010000011",
  38327=>"001001101",
  38328=>"011110100",
  38329=>"110001000",
  38330=>"001000111",
  38331=>"111110000",
  38332=>"110010010",
  38333=>"100011100",
  38334=>"101010000",
  38335=>"011001110",
  38336=>"110100001",
  38337=>"100100110",
  38338=>"010111010",
  38339=>"001110111",
  38340=>"110100100",
  38341=>"011010000",
  38342=>"011111001",
  38343=>"000111000",
  38344=>"010010010",
  38345=>"101111111",
  38346=>"100000000",
  38347=>"001111000",
  38348=>"010111111",
  38349=>"001110001",
  38350=>"010010001",
  38351=>"110011011",
  38352=>"100101101",
  38353=>"101011010",
  38354=>"101101001",
  38355=>"110100100",
  38356=>"000111110",
  38357=>"010010111",
  38358=>"011111100",
  38359=>"110000100",
  38360=>"001001101",
  38361=>"111001010",
  38362=>"110110111",
  38363=>"010010001",
  38364=>"111011001",
  38365=>"100010111",
  38366=>"101110100",
  38367=>"010110001",
  38368=>"001100001",
  38369=>"000010101",
  38370=>"101000010",
  38371=>"100110100",
  38372=>"101100011",
  38373=>"000000100",
  38374=>"010010001",
  38375=>"001101010",
  38376=>"101100110",
  38377=>"001100111",
  38378=>"011100101",
  38379=>"011111110",
  38380=>"001010000",
  38381=>"110101010",
  38382=>"100100011",
  38383=>"011010001",
  38384=>"000100110",
  38385=>"110111001",
  38386=>"001010110",
  38387=>"010010110",
  38388=>"110100001",
  38389=>"101010111",
  38390=>"010010110",
  38391=>"101001010",
  38392=>"110000010",
  38393=>"100010111",
  38394=>"111000110",
  38395=>"100100111",
  38396=>"001110001",
  38397=>"000000101",
  38398=>"001110100",
  38399=>"000110000",
  38400=>"100001000",
  38401=>"111111100",
  38402=>"100001000",
  38403=>"000001100",
  38404=>"111010100",
  38405=>"101111001",
  38406=>"100111001",
  38407=>"101011010",
  38408=>"011110110",
  38409=>"110000111",
  38410=>"010110101",
  38411=>"000110101",
  38412=>"110100010",
  38413=>"110110111",
  38414=>"110100011",
  38415=>"011001000",
  38416=>"000111101",
  38417=>"110111101",
  38418=>"011110101",
  38419=>"001100100",
  38420=>"111011000",
  38421=>"001000101",
  38422=>"000110101",
  38423=>"001111101",
  38424=>"011110111",
  38425=>"111011101",
  38426=>"101000000",
  38427=>"000111111",
  38428=>"101010100",
  38429=>"010111100",
  38430=>"110010000",
  38431=>"010110100",
  38432=>"100110001",
  38433=>"101000000",
  38434=>"100000010",
  38435=>"100101011",
  38436=>"101001011",
  38437=>"100101000",
  38438=>"101111010",
  38439=>"101010001",
  38440=>"110101101",
  38441=>"011100100",
  38442=>"010010001",
  38443=>"100101110",
  38444=>"010000100",
  38445=>"011101110",
  38446=>"110111101",
  38447=>"100100001",
  38448=>"001110101",
  38449=>"011111001",
  38450=>"000000110",
  38451=>"101100001",
  38452=>"111001010",
  38453=>"011000100",
  38454=>"110000000",
  38455=>"111000000",
  38456=>"100101100",
  38457=>"111110000",
  38458=>"000111011",
  38459=>"011100110",
  38460=>"000010110",
  38461=>"010000110",
  38462=>"011101100",
  38463=>"111011101",
  38464=>"100100010",
  38465=>"010110000",
  38466=>"000010010",
  38467=>"010100001",
  38468=>"111100110",
  38469=>"001111101",
  38470=>"001000101",
  38471=>"111111001",
  38472=>"101100011",
  38473=>"011110101",
  38474=>"111011000",
  38475=>"101110010",
  38476=>"010101110",
  38477=>"101000000",
  38478=>"111111001",
  38479=>"010010010",
  38480=>"011000001",
  38481=>"100011000",
  38482=>"101100110",
  38483=>"100111101",
  38484=>"001101001",
  38485=>"101110000",
  38486=>"110011010",
  38487=>"110001110",
  38488=>"111111110",
  38489=>"110010111",
  38490=>"001010110",
  38491=>"111100100",
  38492=>"111111110",
  38493=>"100101010",
  38494=>"110101111",
  38495=>"010000000",
  38496=>"110010001",
  38497=>"011010110",
  38498=>"110011100",
  38499=>"100000000",
  38500=>"111101110",
  38501=>"110001101",
  38502=>"011100110",
  38503=>"011011111",
  38504=>"000101100",
  38505=>"110100010",
  38506=>"110010111",
  38507=>"010000011",
  38508=>"011011101",
  38509=>"111100111",
  38510=>"011101110",
  38511=>"010101101",
  38512=>"101001010",
  38513=>"000001000",
  38514=>"100100000",
  38515=>"110001101",
  38516=>"000000111",
  38517=>"110110111",
  38518=>"011010101",
  38519=>"011010101",
  38520=>"110001100",
  38521=>"100111010",
  38522=>"000011111",
  38523=>"001000010",
  38524=>"010101100",
  38525=>"001000010",
  38526=>"001011111",
  38527=>"011000111",
  38528=>"111111100",
  38529=>"110000101",
  38530=>"011101011",
  38531=>"101111010",
  38532=>"000000100",
  38533=>"000011100",
  38534=>"000001100",
  38535=>"010001111",
  38536=>"100100001",
  38537=>"100001011",
  38538=>"000111111",
  38539=>"111101100",
  38540=>"101101001",
  38541=>"010010000",
  38542=>"000001000",
  38543=>"000101000",
  38544=>"100010110",
  38545=>"101101111",
  38546=>"010000101",
  38547=>"101110001",
  38548=>"001011100",
  38549=>"010100011",
  38550=>"111010110",
  38551=>"000110110",
  38552=>"110110011",
  38553=>"110100101",
  38554=>"100101110",
  38555=>"111101000",
  38556=>"000100110",
  38557=>"101100101",
  38558=>"010000101",
  38559=>"101000110",
  38560=>"110011010",
  38561=>"100000111",
  38562=>"101001110",
  38563=>"000011101",
  38564=>"000010111",
  38565=>"101000001",
  38566=>"001000000",
  38567=>"010000001",
  38568=>"101100010",
  38569=>"000010000",
  38570=>"001011000",
  38571=>"101111101",
  38572=>"100100111",
  38573=>"111000000",
  38574=>"000010010",
  38575=>"010000000",
  38576=>"010010000",
  38577=>"001110011",
  38578=>"100100001",
  38579=>"100010010",
  38580=>"010101100",
  38581=>"100101110",
  38582=>"111001100",
  38583=>"111101010",
  38584=>"110011101",
  38585=>"011011100",
  38586=>"111110110",
  38587=>"010110001",
  38588=>"111101001",
  38589=>"101011110",
  38590=>"000011000",
  38591=>"011010100",
  38592=>"001011111",
  38593=>"100011001",
  38594=>"000111011",
  38595=>"111000100",
  38596=>"101111011",
  38597=>"101000100",
  38598=>"101000001",
  38599=>"101101011",
  38600=>"010001010",
  38601=>"010001001",
  38602=>"110000111",
  38603=>"110001010",
  38604=>"010000010",
  38605=>"011100110",
  38606=>"001111110",
  38607=>"010010000",
  38608=>"001100001",
  38609=>"100100100",
  38610=>"111110110",
  38611=>"101011010",
  38612=>"010011010",
  38613=>"110100001",
  38614=>"110001010",
  38615=>"011001100",
  38616=>"011001001",
  38617=>"101000101",
  38618=>"011110100",
  38619=>"001111010",
  38620=>"000101101",
  38621=>"000110100",
  38622=>"110001010",
  38623=>"101100101",
  38624=>"011010111",
  38625=>"101101001",
  38626=>"100101111",
  38627=>"011101100",
  38628=>"110011011",
  38629=>"100010110",
  38630=>"010001001",
  38631=>"111011101",
  38632=>"001010000",
  38633=>"010001101",
  38634=>"001001000",
  38635=>"100001101",
  38636=>"011111110",
  38637=>"000011011",
  38638=>"110111001",
  38639=>"100001001",
  38640=>"011001100",
  38641=>"100101111",
  38642=>"010010001",
  38643=>"110001110",
  38644=>"000111100",
  38645=>"100100111",
  38646=>"100100110",
  38647=>"111110010",
  38648=>"011111100",
  38649=>"111110011",
  38650=>"010111011",
  38651=>"110100001",
  38652=>"000001011",
  38653=>"000100011",
  38654=>"000110000",
  38655=>"111100110",
  38656=>"010100010",
  38657=>"100000001",
  38658=>"011000011",
  38659=>"000111110",
  38660=>"111110100",
  38661=>"111110000",
  38662=>"111011110",
  38663=>"001001010",
  38664=>"000111001",
  38665=>"010011011",
  38666=>"000111101",
  38667=>"011001111",
  38668=>"110010101",
  38669=>"101000111",
  38670=>"000001110",
  38671=>"000111000",
  38672=>"011011011",
  38673=>"100111111",
  38674=>"110100000",
  38675=>"100010011",
  38676=>"100101010",
  38677=>"111100100",
  38678=>"000001101",
  38679=>"110001110",
  38680=>"000111001",
  38681=>"001100000",
  38682=>"101000111",
  38683=>"010111110",
  38684=>"011001010",
  38685=>"010110001",
  38686=>"000100001",
  38687=>"111001111",
  38688=>"111101111",
  38689=>"011000100",
  38690=>"100100001",
  38691=>"101010110",
  38692=>"011111110",
  38693=>"100011101",
  38694=>"000010101",
  38695=>"110001101",
  38696=>"101111001",
  38697=>"010001001",
  38698=>"111001000",
  38699=>"100101001",
  38700=>"001011011",
  38701=>"101011001",
  38702=>"101101011",
  38703=>"101000101",
  38704=>"001001010",
  38705=>"110000100",
  38706=>"101101101",
  38707=>"111100001",
  38708=>"110000111",
  38709=>"101010100",
  38710=>"010010000",
  38711=>"101000100",
  38712=>"111000101",
  38713=>"100101110",
  38714=>"010001011",
  38715=>"000101000",
  38716=>"010010011",
  38717=>"001001111",
  38718=>"111001111",
  38719=>"000001111",
  38720=>"001000110",
  38721=>"010000110",
  38722=>"100000110",
  38723=>"110000101",
  38724=>"000111110",
  38725=>"100100111",
  38726=>"001111011",
  38727=>"110010100",
  38728=>"111110110",
  38729=>"011010101",
  38730=>"111010010",
  38731=>"110100010",
  38732=>"111000000",
  38733=>"001010001",
  38734=>"001111011",
  38735=>"000101001",
  38736=>"100101101",
  38737=>"101111101",
  38738=>"010110000",
  38739=>"111110000",
  38740=>"101011101",
  38741=>"010101011",
  38742=>"111011000",
  38743=>"001101001",
  38744=>"001111111",
  38745=>"001111100",
  38746=>"001010011",
  38747=>"011010111",
  38748=>"001000011",
  38749=>"100011011",
  38750=>"100000010",
  38751=>"000111110",
  38752=>"100110000",
  38753=>"100100111",
  38754=>"010001101",
  38755=>"101111011",
  38756=>"111110001",
  38757=>"100000101",
  38758=>"110000100",
  38759=>"101011100",
  38760=>"110110101",
  38761=>"101111101",
  38762=>"001010111",
  38763=>"010111101",
  38764=>"011111001",
  38765=>"101000001",
  38766=>"100001000",
  38767=>"010000111",
  38768=>"100101111",
  38769=>"000010100",
  38770=>"110000100",
  38771=>"001110100",
  38772=>"011011011",
  38773=>"100111011",
  38774=>"011011111",
  38775=>"000000100",
  38776=>"111100101",
  38777=>"001101100",
  38778=>"100100100",
  38779=>"010111100",
  38780=>"010011111",
  38781=>"111011001",
  38782=>"001101010",
  38783=>"001010110",
  38784=>"001001100",
  38785=>"111001010",
  38786=>"101000111",
  38787=>"001011010",
  38788=>"101010101",
  38789=>"110000011",
  38790=>"010111000",
  38791=>"001100010",
  38792=>"111110011",
  38793=>"111101011",
  38794=>"111011000",
  38795=>"000100000",
  38796=>"100000010",
  38797=>"110010110",
  38798=>"110100011",
  38799=>"001110000",
  38800=>"011001000",
  38801=>"101011001",
  38802=>"111001111",
  38803=>"000001110",
  38804=>"001101101",
  38805=>"110001101",
  38806=>"101101110",
  38807=>"101111110",
  38808=>"100011011",
  38809=>"000001110",
  38810=>"000101001",
  38811=>"010000101",
  38812=>"000010100",
  38813=>"000010100",
  38814=>"110000000",
  38815=>"100110010",
  38816=>"110010101",
  38817=>"100011101",
  38818=>"110110000",
  38819=>"010011001",
  38820=>"111110110",
  38821=>"110000101",
  38822=>"001011100",
  38823=>"010010011",
  38824=>"001010011",
  38825=>"110111000",
  38826=>"101111011",
  38827=>"011011011",
  38828=>"000010001",
  38829=>"110000101",
  38830=>"111000011",
  38831=>"001111011",
  38832=>"010010011",
  38833=>"111111111",
  38834=>"000001101",
  38835=>"101001110",
  38836=>"101001000",
  38837=>"011000100",
  38838=>"111001010",
  38839=>"110100110",
  38840=>"000100100",
  38841=>"111000011",
  38842=>"010100100",
  38843=>"000110011",
  38844=>"011010111",
  38845=>"010111100",
  38846=>"100101111",
  38847=>"010011000",
  38848=>"101101010",
  38849=>"011010100",
  38850=>"000001111",
  38851=>"001100110",
  38852=>"000101101",
  38853=>"100010010",
  38854=>"001110101",
  38855=>"110010010",
  38856=>"000000000",
  38857=>"011000001",
  38858=>"100001001",
  38859=>"001110010",
  38860=>"111100110",
  38861=>"100111110",
  38862=>"101110101",
  38863=>"111011111",
  38864=>"000001100",
  38865=>"000001110",
  38866=>"111000100",
  38867=>"001000111",
  38868=>"001110110",
  38869=>"000111101",
  38870=>"111001100",
  38871=>"011100111",
  38872=>"110100101",
  38873=>"011001100",
  38874=>"000010100",
  38875=>"110001101",
  38876=>"101100100",
  38877=>"101010111",
  38878=>"010111100",
  38879=>"101101010",
  38880=>"011001111",
  38881=>"111100110",
  38882=>"110000111",
  38883=>"101100010",
  38884=>"100001101",
  38885=>"010010010",
  38886=>"110000001",
  38887=>"000111110",
  38888=>"010010110",
  38889=>"000101010",
  38890=>"010100010",
  38891=>"101000110",
  38892=>"000001101",
  38893=>"000110000",
  38894=>"101100110",
  38895=>"001110101",
  38896=>"011101011",
  38897=>"001000100",
  38898=>"111100111",
  38899=>"001111001",
  38900=>"000101101",
  38901=>"001011011",
  38902=>"011010001",
  38903=>"010000111",
  38904=>"010001011",
  38905=>"010001101",
  38906=>"101101101",
  38907=>"001011001",
  38908=>"011110110",
  38909=>"101000000",
  38910=>"101100011",
  38911=>"110111011",
  38912=>"000001000",
  38913=>"111101100",
  38914=>"101100100",
  38915=>"100001111",
  38916=>"000101100",
  38917=>"010101001",
  38918=>"001110101",
  38919=>"111101101",
  38920=>"111000011",
  38921=>"101100111",
  38922=>"010101010",
  38923=>"110110110",
  38924=>"011111111",
  38925=>"110110110",
  38926=>"111010101",
  38927=>"010010110",
  38928=>"010100100",
  38929=>"001101000",
  38930=>"000001111",
  38931=>"000110101",
  38932=>"000000110",
  38933=>"000100111",
  38934=>"000111010",
  38935=>"011001010",
  38936=>"110100011",
  38937=>"111011101",
  38938=>"000111110",
  38939=>"000111001",
  38940=>"101000101",
  38941=>"111010101",
  38942=>"011101111",
  38943=>"001011000",
  38944=>"010100101",
  38945=>"001101101",
  38946=>"110100100",
  38947=>"111010111",
  38948=>"001101100",
  38949=>"000010110",
  38950=>"001110001",
  38951=>"001110001",
  38952=>"001000111",
  38953=>"101011111",
  38954=>"000000110",
  38955=>"100000001",
  38956=>"000001100",
  38957=>"101100100",
  38958=>"100110100",
  38959=>"001000110",
  38960=>"000000000",
  38961=>"001011101",
  38962=>"101001110",
  38963=>"000001000",
  38964=>"110001110",
  38965=>"101111010",
  38966=>"111010000",
  38967=>"110000110",
  38968=>"111000111",
  38969=>"101101101",
  38970=>"101001001",
  38971=>"111110101",
  38972=>"111001001",
  38973=>"001101101",
  38974=>"010000110",
  38975=>"000100011",
  38976=>"100010000",
  38977=>"001011100",
  38978=>"010111101",
  38979=>"011000111",
  38980=>"010001010",
  38981=>"110100110",
  38982=>"011010101",
  38983=>"100100110",
  38984=>"111101001",
  38985=>"100111111",
  38986=>"110110101",
  38987=>"100011010",
  38988=>"100011111",
  38989=>"100100110",
  38990=>"011111011",
  38991=>"111011100",
  38992=>"011110000",
  38993=>"001000011",
  38994=>"111111010",
  38995=>"110100110",
  38996=>"110000110",
  38997=>"011011100",
  38998=>"010101001",
  38999=>"001111110",
  39000=>"011111010",
  39001=>"111100110",
  39002=>"011000010",
  39003=>"100110101",
  39004=>"011001011",
  39005=>"000101000",
  39006=>"111010001",
  39007=>"100111101",
  39008=>"001110000",
  39009=>"011001100",
  39010=>"011001010",
  39011=>"000011000",
  39012=>"011011011",
  39013=>"111111101",
  39014=>"011100010",
  39015=>"110010001",
  39016=>"001000110",
  39017=>"100000000",
  39018=>"100101001",
  39019=>"100101000",
  39020=>"101110001",
  39021=>"010100101",
  39022=>"000000111",
  39023=>"000010010",
  39024=>"110000011",
  39025=>"100110000",
  39026=>"110000000",
  39027=>"001000101",
  39028=>"111001111",
  39029=>"001111111",
  39030=>"000011001",
  39031=>"100111000",
  39032=>"101101111",
  39033=>"010011000",
  39034=>"111101110",
  39035=>"111111100",
  39036=>"101010110",
  39037=>"101110010",
  39038=>"110100101",
  39039=>"110101110",
  39040=>"010010100",
  39041=>"111000001",
  39042=>"011001100",
  39043=>"000100111",
  39044=>"100000110",
  39045=>"000101110",
  39046=>"101010100",
  39047=>"101101100",
  39048=>"101000001",
  39049=>"001110110",
  39050=>"100111111",
  39051=>"001001010",
  39052=>"011111100",
  39053=>"100111111",
  39054=>"100001010",
  39055=>"001100000",
  39056=>"111011110",
  39057=>"101110011",
  39058=>"111001110",
  39059=>"000010100",
  39060=>"011110100",
  39061=>"001011111",
  39062=>"111111001",
  39063=>"001111110",
  39064=>"001010011",
  39065=>"111100110",
  39066=>"001001101",
  39067=>"111100110",
  39068=>"001101011",
  39069=>"111101000",
  39070=>"000010010",
  39071=>"110110110",
  39072=>"100010010",
  39073=>"000011110",
  39074=>"100001001",
  39075=>"100011101",
  39076=>"101110011",
  39077=>"111000100",
  39078=>"111001111",
  39079=>"001100011",
  39080=>"001000101",
  39081=>"000110010",
  39082=>"000100101",
  39083=>"001111011",
  39084=>"110110001",
  39085=>"001100101",
  39086=>"000001101",
  39087=>"110111111",
  39088=>"011010111",
  39089=>"110100101",
  39090=>"101110010",
  39091=>"000000000",
  39092=>"001000011",
  39093=>"110010000",
  39094=>"111110011",
  39095=>"010110000",
  39096=>"101000001",
  39097=>"110011101",
  39098=>"001110110",
  39099=>"000111111",
  39100=>"000011011",
  39101=>"010010010",
  39102=>"100100111",
  39103=>"011110011",
  39104=>"101001011",
  39105=>"110001001",
  39106=>"111010000",
  39107=>"111000011",
  39108=>"100000110",
  39109=>"011101110",
  39110=>"111110100",
  39111=>"101100011",
  39112=>"001010111",
  39113=>"010111101",
  39114=>"101100010",
  39115=>"111100000",
  39116=>"100010001",
  39117=>"000010000",
  39118=>"000011111",
  39119=>"111001011",
  39120=>"101011111",
  39121=>"110010010",
  39122=>"111111000",
  39123=>"011000011",
  39124=>"111000001",
  39125=>"001001001",
  39126=>"101100100",
  39127=>"111010110",
  39128=>"100111001",
  39129=>"001100001",
  39130=>"100110100",
  39131=>"011011100",
  39132=>"010011000",
  39133=>"000000000",
  39134=>"101001100",
  39135=>"100110001",
  39136=>"001010111",
  39137=>"001011101",
  39138=>"100111010",
  39139=>"001001000",
  39140=>"001101011",
  39141=>"111101111",
  39142=>"000111011",
  39143=>"111101110",
  39144=>"101100100",
  39145=>"110001100",
  39146=>"110100001",
  39147=>"000011100",
  39148=>"000110111",
  39149=>"001100001",
  39150=>"001001001",
  39151=>"100100000",
  39152=>"010101011",
  39153=>"111000011",
  39154=>"011100110",
  39155=>"010011101",
  39156=>"111001011",
  39157=>"010110111",
  39158=>"101010011",
  39159=>"110011000",
  39160=>"101111011",
  39161=>"000001100",
  39162=>"010111101",
  39163=>"111000000",
  39164=>"101010101",
  39165=>"000101100",
  39166=>"001010001",
  39167=>"101101010",
  39168=>"111001010",
  39169=>"000100000",
  39170=>"010000001",
  39171=>"111000010",
  39172=>"001010000",
  39173=>"001100111",
  39174=>"011000111",
  39175=>"110111100",
  39176=>"000111001",
  39177=>"101010010",
  39178=>"011001101",
  39179=>"001100000",
  39180=>"011000101",
  39181=>"011010011",
  39182=>"010100111",
  39183=>"011110110",
  39184=>"101100110",
  39185=>"011111010",
  39186=>"010011110",
  39187=>"001111010",
  39188=>"101000000",
  39189=>"001010110",
  39190=>"011011101",
  39191=>"111100101",
  39192=>"010101111",
  39193=>"110100111",
  39194=>"100100111",
  39195=>"111011010",
  39196=>"100011110",
  39197=>"110101101",
  39198=>"011000111",
  39199=>"111110001",
  39200=>"011010001",
  39201=>"000011010",
  39202=>"001000000",
  39203=>"001011000",
  39204=>"101011010",
  39205=>"011110011",
  39206=>"101010000",
  39207=>"100011100",
  39208=>"110100111",
  39209=>"010011001",
  39210=>"001011101",
  39211=>"011100101",
  39212=>"100110010",
  39213=>"010110100",
  39214=>"111000010",
  39215=>"111111100",
  39216=>"000011001",
  39217=>"101001111",
  39218=>"011010001",
  39219=>"001100111",
  39220=>"000100011",
  39221=>"011011100",
  39222=>"111110001",
  39223=>"101101000",
  39224=>"111110010",
  39225=>"100001010",
  39226=>"001111000",
  39227=>"010101011",
  39228=>"101110000",
  39229=>"110010110",
  39230=>"101100000",
  39231=>"100000100",
  39232=>"101000000",
  39233=>"001111010",
  39234=>"011111000",
  39235=>"010111001",
  39236=>"001001001",
  39237=>"011111110",
  39238=>"110100010",
  39239=>"010001111",
  39240=>"100100110",
  39241=>"011001101",
  39242=>"101011011",
  39243=>"011011110",
  39244=>"111010101",
  39245=>"011011111",
  39246=>"111011001",
  39247=>"000001100",
  39248=>"101110000",
  39249=>"000011111",
  39250=>"100001101",
  39251=>"011111001",
  39252=>"111001000",
  39253=>"000010000",
  39254=>"111101110",
  39255=>"101001110",
  39256=>"101111011",
  39257=>"000100110",
  39258=>"100001101",
  39259=>"001111010",
  39260=>"110110011",
  39261=>"101010100",
  39262=>"010001110",
  39263=>"010010101",
  39264=>"010110110",
  39265=>"110010110",
  39266=>"111110010",
  39267=>"001000000",
  39268=>"011100001",
  39269=>"111000000",
  39270=>"101111010",
  39271=>"100110111",
  39272=>"111111110",
  39273=>"000011000",
  39274=>"100111110",
  39275=>"100110110",
  39276=>"000010100",
  39277=>"011111001",
  39278=>"000101011",
  39279=>"000111100",
  39280=>"011101100",
  39281=>"110000111",
  39282=>"011001101",
  39283=>"001111001",
  39284=>"100011101",
  39285=>"110010100",
  39286=>"101010100",
  39287=>"110100110",
  39288=>"000010100",
  39289=>"101011010",
  39290=>"110101111",
  39291=>"010100110",
  39292=>"000010100",
  39293=>"100111000",
  39294=>"000111100",
  39295=>"001001001",
  39296=>"001001011",
  39297=>"000110100",
  39298=>"100101100",
  39299=>"001000101",
  39300=>"110001010",
  39301=>"010010011",
  39302=>"100010010",
  39303=>"001111000",
  39304=>"110100011",
  39305=>"110010011",
  39306=>"110001000",
  39307=>"011000000",
  39308=>"000000110",
  39309=>"100111010",
  39310=>"011111000",
  39311=>"110000010",
  39312=>"101001001",
  39313=>"001010110",
  39314=>"100001100",
  39315=>"110010111",
  39316=>"111010001",
  39317=>"101110100",
  39318=>"110010011",
  39319=>"110101011",
  39320=>"001011001",
  39321=>"000101101",
  39322=>"011100011",
  39323=>"110100110",
  39324=>"111001011",
  39325=>"011001111",
  39326=>"010110110",
  39327=>"000010100",
  39328=>"010001101",
  39329=>"001000010",
  39330=>"011101011",
  39331=>"001100001",
  39332=>"111010110",
  39333=>"101101001",
  39334=>"000100101",
  39335=>"110111111",
  39336=>"001101101",
  39337=>"011111010",
  39338=>"001001011",
  39339=>"001011110",
  39340=>"101010110",
  39341=>"111010110",
  39342=>"000110000",
  39343=>"010101000",
  39344=>"001110010",
  39345=>"011010000",
  39346=>"100011000",
  39347=>"111101111",
  39348=>"111100110",
  39349=>"101000111",
  39350=>"001101101",
  39351=>"110010000",
  39352=>"010011000",
  39353=>"000101101",
  39354=>"011011000",
  39355=>"000100110",
  39356=>"101111011",
  39357=>"100011011",
  39358=>"001001010",
  39359=>"011000001",
  39360=>"100000010",
  39361=>"110001101",
  39362=>"101111101",
  39363=>"100000111",
  39364=>"111001111",
  39365=>"010000011",
  39366=>"011100110",
  39367=>"001000101",
  39368=>"100101110",
  39369=>"110011010",
  39370=>"011000000",
  39371=>"101010100",
  39372=>"011001101",
  39373=>"001010000",
  39374=>"001001111",
  39375=>"001011000",
  39376=>"111111001",
  39377=>"001100001",
  39378=>"100011000",
  39379=>"001000110",
  39380=>"110000001",
  39381=>"110111110",
  39382=>"110011101",
  39383=>"001001011",
  39384=>"110001010",
  39385=>"011011111",
  39386=>"001100010",
  39387=>"001111100",
  39388=>"100101100",
  39389=>"011110111",
  39390=>"000000000",
  39391=>"101101011",
  39392=>"101011000",
  39393=>"000100001",
  39394=>"010000101",
  39395=>"000101110",
  39396=>"011101101",
  39397=>"111011010",
  39398=>"100101000",
  39399=>"111111001",
  39400=>"000011110",
  39401=>"010110001",
  39402=>"011000100",
  39403=>"010111110",
  39404=>"000110111",
  39405=>"000011011",
  39406=>"110110000",
  39407=>"110000000",
  39408=>"001100111",
  39409=>"110101101",
  39410=>"000100101",
  39411=>"001011010",
  39412=>"110000111",
  39413=>"001001001",
  39414=>"110001011",
  39415=>"000000100",
  39416=>"110000101",
  39417=>"111100101",
  39418=>"000100011",
  39419=>"010100100",
  39420=>"000010000",
  39421=>"101011110",
  39422=>"100010001",
  39423=>"100110010",
  39424=>"101101000",
  39425=>"010100110",
  39426=>"001110011",
  39427=>"101011001",
  39428=>"100101011",
  39429=>"111011000",
  39430=>"010011111",
  39431=>"100000101",
  39432=>"111010101",
  39433=>"110110000",
  39434=>"111000010",
  39435=>"000011000",
  39436=>"001010100",
  39437=>"010010110",
  39438=>"011001001",
  39439=>"110111110",
  39440=>"011111010",
  39441=>"111111101",
  39442=>"110000101",
  39443=>"101001101",
  39444=>"100110001",
  39445=>"101111001",
  39446=>"111011110",
  39447=>"110101110",
  39448=>"101001001",
  39449=>"111001010",
  39450=>"111111000",
  39451=>"010010011",
  39452=>"010111101",
  39453=>"101100001",
  39454=>"101101011",
  39455=>"000000011",
  39456=>"111101001",
  39457=>"000001100",
  39458=>"000010010",
  39459=>"100000111",
  39460=>"001001001",
  39461=>"101110011",
  39462=>"001111101",
  39463=>"101001110",
  39464=>"011001001",
  39465=>"000111101",
  39466=>"001010101",
  39467=>"010001100",
  39468=>"000101000",
  39469=>"111001000",
  39470=>"010110101",
  39471=>"111010101",
  39472=>"000101101",
  39473=>"011111011",
  39474=>"011101000",
  39475=>"000001001",
  39476=>"000001011",
  39477=>"110001000",
  39478=>"111101011",
  39479=>"011100000",
  39480=>"100010110",
  39481=>"101111111",
  39482=>"100100100",
  39483=>"100000010",
  39484=>"000110010",
  39485=>"101010110",
  39486=>"011110011",
  39487=>"001100100",
  39488=>"011000011",
  39489=>"010100111",
  39490=>"011101100",
  39491=>"110101100",
  39492=>"101011100",
  39493=>"111011011",
  39494=>"101011001",
  39495=>"000010011",
  39496=>"110100111",
  39497=>"001010000",
  39498=>"101101111",
  39499=>"010011010",
  39500=>"001011001",
  39501=>"001000001",
  39502=>"000100110",
  39503=>"011100010",
  39504=>"010001000",
  39505=>"010010001",
  39506=>"010101010",
  39507=>"101011111",
  39508=>"000010010",
  39509=>"000000011",
  39510=>"000001000",
  39511=>"111111000",
  39512=>"110101011",
  39513=>"011111001",
  39514=>"001001010",
  39515=>"100000010",
  39516=>"011011111",
  39517=>"001001000",
  39518=>"000000100",
  39519=>"010101001",
  39520=>"101011101",
  39521=>"110111101",
  39522=>"000000110",
  39523=>"001011101",
  39524=>"111011110",
  39525=>"000101100",
  39526=>"011001111",
  39527=>"111101010",
  39528=>"101000101",
  39529=>"101100001",
  39530=>"001100011",
  39531=>"000000001",
  39532=>"100010001",
  39533=>"110111101",
  39534=>"010111011",
  39535=>"111111111",
  39536=>"101011100",
  39537=>"001101010",
  39538=>"111111010",
  39539=>"010001010",
  39540=>"100011101",
  39541=>"010110101",
  39542=>"111011111",
  39543=>"001110111",
  39544=>"010110111",
  39545=>"111100111",
  39546=>"001101101",
  39547=>"100001101",
  39548=>"110011001",
  39549=>"000001001",
  39550=>"100100011",
  39551=>"111101011",
  39552=>"110110000",
  39553=>"100100111",
  39554=>"011011011",
  39555=>"110001101",
  39556=>"001101010",
  39557=>"001011010",
  39558=>"000110001",
  39559=>"011110100",
  39560=>"100100000",
  39561=>"111010011",
  39562=>"110000101",
  39563=>"110011000",
  39564=>"111110110",
  39565=>"101001001",
  39566=>"101001100",
  39567=>"111101011",
  39568=>"110101011",
  39569=>"001111011",
  39570=>"000001110",
  39571=>"100101010",
  39572=>"000100111",
  39573=>"100011011",
  39574=>"111000000",
  39575=>"100110100",
  39576=>"100010111",
  39577=>"101100001",
  39578=>"101000001",
  39579=>"010110100",
  39580=>"011001111",
  39581=>"001100000",
  39582=>"110100111",
  39583=>"000001010",
  39584=>"100000000",
  39585=>"011010100",
  39586=>"100001110",
  39587=>"101100111",
  39588=>"011011000",
  39589=>"010001000",
  39590=>"110001000",
  39591=>"001001111",
  39592=>"010101100",
  39593=>"111100101",
  39594=>"011001000",
  39595=>"001110110",
  39596=>"110000100",
  39597=>"000111101",
  39598=>"111111010",
  39599=>"111000101",
  39600=>"111000001",
  39601=>"101011110",
  39602=>"101110010",
  39603=>"001000001",
  39604=>"001001011",
  39605=>"101011010",
  39606=>"000011101",
  39607=>"010101001",
  39608=>"010101001",
  39609=>"100111001",
  39610=>"110110111",
  39611=>"000101011",
  39612=>"010111000",
  39613=>"011111001",
  39614=>"111101100",
  39615=>"000011100",
  39616=>"111111001",
  39617=>"011110101",
  39618=>"000100111",
  39619=>"100011011",
  39620=>"010001100",
  39621=>"010010101",
  39622=>"101101101",
  39623=>"100011010",
  39624=>"011100101",
  39625=>"100100010",
  39626=>"101000101",
  39627=>"111101011",
  39628=>"010010101",
  39629=>"000101011",
  39630=>"011000100",
  39631=>"010001001",
  39632=>"101000011",
  39633=>"101110011",
  39634=>"111110100",
  39635=>"101011010",
  39636=>"101110011",
  39637=>"111000010",
  39638=>"010111001",
  39639=>"011001011",
  39640=>"001000011",
  39641=>"110100110",
  39642=>"000001110",
  39643=>"110001111",
  39644=>"010101100",
  39645=>"011000101",
  39646=>"110001010",
  39647=>"101111101",
  39648=>"000000010",
  39649=>"000000001",
  39650=>"010000011",
  39651=>"110100111",
  39652=>"010011111",
  39653=>"110111001",
  39654=>"001000010",
  39655=>"000100010",
  39656=>"100001011",
  39657=>"000000110",
  39658=>"010101100",
  39659=>"000101111",
  39660=>"001011010",
  39661=>"110011010",
  39662=>"110010101",
  39663=>"000101110",
  39664=>"101010000",
  39665=>"001001011",
  39666=>"111111110",
  39667=>"010100010",
  39668=>"010111110",
  39669=>"101101111",
  39670=>"111000111",
  39671=>"010101011",
  39672=>"000011110",
  39673=>"111001011",
  39674=>"110010110",
  39675=>"000010110",
  39676=>"110111110",
  39677=>"010011110",
  39678=>"101100111",
  39679=>"011111000",
  39680=>"000100101",
  39681=>"010100011",
  39682=>"100111001",
  39683=>"010000101",
  39684=>"100111111",
  39685=>"000011111",
  39686=>"101100011",
  39687=>"000010001",
  39688=>"011100011",
  39689=>"010111101",
  39690=>"110110100",
  39691=>"111110001",
  39692=>"110000101",
  39693=>"110111101",
  39694=>"010011110",
  39695=>"011111011",
  39696=>"011000111",
  39697=>"001001110",
  39698=>"011111000",
  39699=>"110000111",
  39700=>"000010111",
  39701=>"100111101",
  39702=>"000011000",
  39703=>"000101001",
  39704=>"111011111",
  39705=>"100011011",
  39706=>"001011110",
  39707=>"111100010",
  39708=>"100110000",
  39709=>"111010101",
  39710=>"101000010",
  39711=>"110111000",
  39712=>"000100000",
  39713=>"100101111",
  39714=>"111101100",
  39715=>"011111011",
  39716=>"001000010",
  39717=>"101100111",
  39718=>"100110110",
  39719=>"101000000",
  39720=>"001100000",
  39721=>"110101101",
  39722=>"010011001",
  39723=>"010100111",
  39724=>"101001010",
  39725=>"000101011",
  39726=>"011001010",
  39727=>"100001011",
  39728=>"000101111",
  39729=>"101000101",
  39730=>"010101000",
  39731=>"110010101",
  39732=>"111111011",
  39733=>"111011110",
  39734=>"011110110",
  39735=>"000000011",
  39736=>"010001001",
  39737=>"101111000",
  39738=>"101101000",
  39739=>"111111000",
  39740=>"100111111",
  39741=>"100010101",
  39742=>"100100111",
  39743=>"011110111",
  39744=>"100000000",
  39745=>"010011111",
  39746=>"101010000",
  39747=>"111001000",
  39748=>"100110011",
  39749=>"101111111",
  39750=>"011001011",
  39751=>"001010001",
  39752=>"011000100",
  39753=>"011011100",
  39754=>"100110011",
  39755=>"110101001",
  39756=>"010100010",
  39757=>"110101010",
  39758=>"010000000",
  39759=>"100110001",
  39760=>"010000100",
  39761=>"110000000",
  39762=>"101110110",
  39763=>"011110000",
  39764=>"101010000",
  39765=>"011101111",
  39766=>"110100011",
  39767=>"100100000",
  39768=>"111010111",
  39769=>"101010000",
  39770=>"110001101",
  39771=>"010001010",
  39772=>"111001011",
  39773=>"010110111",
  39774=>"011011000",
  39775=>"001000010",
  39776=>"010100001",
  39777=>"011110110",
  39778=>"000000000",
  39779=>"110000101",
  39780=>"101000100",
  39781=>"000011111",
  39782=>"100111100",
  39783=>"010110101",
  39784=>"111001010",
  39785=>"100100011",
  39786=>"110101010",
  39787=>"001011111",
  39788=>"100111111",
  39789=>"111110111",
  39790=>"110001010",
  39791=>"110010110",
  39792=>"100101011",
  39793=>"110010000",
  39794=>"000011101",
  39795=>"111111000",
  39796=>"010101000",
  39797=>"100001010",
  39798=>"000001110",
  39799=>"101100111",
  39800=>"100010111",
  39801=>"000110110",
  39802=>"110000010",
  39803=>"000000001",
  39804=>"011001000",
  39805=>"011001010",
  39806=>"010101101",
  39807=>"010011100",
  39808=>"101011110",
  39809=>"111101001",
  39810=>"100100100",
  39811=>"101110001",
  39812=>"110110110",
  39813=>"111111101",
  39814=>"010000000",
  39815=>"000000100",
  39816=>"101011000",
  39817=>"100110111",
  39818=>"000010101",
  39819=>"100110100",
  39820=>"100111111",
  39821=>"011111110",
  39822=>"101001101",
  39823=>"111000010",
  39824=>"011010001",
  39825=>"101100110",
  39826=>"001000000",
  39827=>"010000001",
  39828=>"101111010",
  39829=>"001110011",
  39830=>"001101111",
  39831=>"101110101",
  39832=>"111111000",
  39833=>"011110011",
  39834=>"100110000",
  39835=>"100110000",
  39836=>"111001101",
  39837=>"010111000",
  39838=>"101110111",
  39839=>"010110100",
  39840=>"001100011",
  39841=>"001010011",
  39842=>"101010101",
  39843=>"100000100",
  39844=>"110010000",
  39845=>"011000101",
  39846=>"100101000",
  39847=>"011011110",
  39848=>"101100100",
  39849=>"001001111",
  39850=>"000000011",
  39851=>"111001100",
  39852=>"011011001",
  39853=>"101111100",
  39854=>"000101010",
  39855=>"010010100",
  39856=>"100101000",
  39857=>"000001010",
  39858=>"001000100",
  39859=>"111101010",
  39860=>"100000000",
  39861=>"110101011",
  39862=>"100000000",
  39863=>"000010101",
  39864=>"000110000",
  39865=>"111110100",
  39866=>"100000000",
  39867=>"100011001",
  39868=>"110111101",
  39869=>"010001111",
  39870=>"100001000",
  39871=>"011010011",
  39872=>"011111100",
  39873=>"010010100",
  39874=>"001010100",
  39875=>"111011100",
  39876=>"010100111",
  39877=>"001000110",
  39878=>"000011110",
  39879=>"011010011",
  39880=>"000001001",
  39881=>"010111010",
  39882=>"001110010",
  39883=>"100110101",
  39884=>"100111011",
  39885=>"010001010",
  39886=>"010101111",
  39887=>"010100100",
  39888=>"101011001",
  39889=>"011100011",
  39890=>"001000001",
  39891=>"110110111",
  39892=>"110110110",
  39893=>"011100101",
  39894=>"010000000",
  39895=>"100011000",
  39896=>"001001100",
  39897=>"110001100",
  39898=>"000010010",
  39899=>"010111001",
  39900=>"010010100",
  39901=>"010101100",
  39902=>"011111000",
  39903=>"111010100",
  39904=>"000110000",
  39905=>"101011100",
  39906=>"011100110",
  39907=>"011101010",
  39908=>"011000001",
  39909=>"001001010",
  39910=>"010101111",
  39911=>"011100001",
  39912=>"000010101",
  39913=>"000110111",
  39914=>"101011000",
  39915=>"010111010",
  39916=>"010001110",
  39917=>"000011100",
  39918=>"111111110",
  39919=>"010111001",
  39920=>"110001101",
  39921=>"111110011",
  39922=>"100001011",
  39923=>"111011101",
  39924=>"011011010",
  39925=>"000001101",
  39926=>"101010000",
  39927=>"010010000",
  39928=>"011101110",
  39929=>"100011110",
  39930=>"000100010",
  39931=>"101101111",
  39932=>"001010101",
  39933=>"010100010",
  39934=>"100100111",
  39935=>"010101111",
  39936=>"011111001",
  39937=>"110101111",
  39938=>"001100010",
  39939=>"110100110",
  39940=>"011101001",
  39941=>"000101011",
  39942=>"111000010",
  39943=>"111101010",
  39944=>"100110000",
  39945=>"010001010",
  39946=>"100110110",
  39947=>"110100111",
  39948=>"110010001",
  39949=>"011001111",
  39950=>"101111001",
  39951=>"111011111",
  39952=>"101001010",
  39953=>"101011011",
  39954=>"101111000",
  39955=>"010000000",
  39956=>"001110101",
  39957=>"001101111",
  39958=>"001100111",
  39959=>"001000001",
  39960=>"111010010",
  39961=>"101010110",
  39962=>"001001110",
  39963=>"000111101",
  39964=>"001100110",
  39965=>"111100001",
  39966=>"000000100",
  39967=>"101001010",
  39968=>"100011001",
  39969=>"110100010",
  39970=>"110000111",
  39971=>"000101101",
  39972=>"110100100",
  39973=>"100000101",
  39974=>"111101010",
  39975=>"111100001",
  39976=>"011000010",
  39977=>"011010101",
  39978=>"111110001",
  39979=>"101111011",
  39980=>"100010110",
  39981=>"010001000",
  39982=>"011011001",
  39983=>"101101000",
  39984=>"010010010",
  39985=>"110000110",
  39986=>"110111110",
  39987=>"110000000",
  39988=>"101100101",
  39989=>"100111011",
  39990=>"000011010",
  39991=>"100101101",
  39992=>"000000000",
  39993=>"001000111",
  39994=>"010110011",
  39995=>"011011001",
  39996=>"110110001",
  39997=>"100010101",
  39998=>"000100100",
  39999=>"111000010",
  40000=>"011000101",
  40001=>"000001000",
  40002=>"100110100",
  40003=>"010101110",
  40004=>"110011010",
  40005=>"001000101",
  40006=>"010000110",
  40007=>"100101111",
  40008=>"011101011",
  40009=>"111111100",
  40010=>"011001010",
  40011=>"111011000",
  40012=>"110001011",
  40013=>"000011011",
  40014=>"101010000",
  40015=>"001000100",
  40016=>"111110101",
  40017=>"000011001",
  40018=>"001000110",
  40019=>"111000010",
  40020=>"000110010",
  40021=>"100000001",
  40022=>"001101011",
  40023=>"011111111",
  40024=>"110111001",
  40025=>"100101000",
  40026=>"101011010",
  40027=>"010101101",
  40028=>"111111000",
  40029=>"110011100",
  40030=>"000011111",
  40031=>"110011000",
  40032=>"101101111",
  40033=>"001100100",
  40034=>"010011111",
  40035=>"010010001",
  40036=>"100010001",
  40037=>"000011000",
  40038=>"010010001",
  40039=>"100000010",
  40040=>"001011101",
  40041=>"000110111",
  40042=>"110101000",
  40043=>"100001100",
  40044=>"110001010",
  40045=>"111111111",
  40046=>"100111111",
  40047=>"000001000",
  40048=>"011111110",
  40049=>"000100111",
  40050=>"101000000",
  40051=>"011001110",
  40052=>"011100111",
  40053=>"110100000",
  40054=>"111011011",
  40055=>"110100110",
  40056=>"011101100",
  40057=>"110000111",
  40058=>"011111111",
  40059=>"000010011",
  40060=>"111111110",
  40061=>"000010110",
  40062=>"111010011",
  40063=>"111111010",
  40064=>"101111100",
  40065=>"010001000",
  40066=>"000010111",
  40067=>"000011011",
  40068=>"111001011",
  40069=>"100001000",
  40070=>"100111010",
  40071=>"100011000",
  40072=>"000110111",
  40073=>"001011100",
  40074=>"000100010",
  40075=>"100111111",
  40076=>"110000111",
  40077=>"101011010",
  40078=>"101000011",
  40079=>"111101011",
  40080=>"100010100",
  40081=>"110101110",
  40082=>"011111101",
  40083=>"010100110",
  40084=>"001001100",
  40085=>"111111110",
  40086=>"101110000",
  40087=>"101010000",
  40088=>"010110111",
  40089=>"000101011",
  40090=>"110101100",
  40091=>"110000101",
  40092=>"000111001",
  40093=>"011101000",
  40094=>"111011100",
  40095=>"110100010",
  40096=>"001000101",
  40097=>"101100100",
  40098=>"010010100",
  40099=>"000100101",
  40100=>"011111111",
  40101=>"110001001",
  40102=>"000000011",
  40103=>"011101010",
  40104=>"001000001",
  40105=>"001101110",
  40106=>"001111011",
  40107=>"000001110",
  40108=>"000111100",
  40109=>"000110100",
  40110=>"011111110",
  40111=>"011111111",
  40112=>"010000011",
  40113=>"000101000",
  40114=>"010001111",
  40115=>"100000011",
  40116=>"010001110",
  40117=>"001100011",
  40118=>"011101000",
  40119=>"011100011",
  40120=>"101111001",
  40121=>"000111000",
  40122=>"010101001",
  40123=>"001011111",
  40124=>"010011001",
  40125=>"110100010",
  40126=>"000011111",
  40127=>"100110011",
  40128=>"011111010",
  40129=>"001110011",
  40130=>"011110011",
  40131=>"100000000",
  40132=>"000011010",
  40133=>"001101101",
  40134=>"101001101",
  40135=>"010111011",
  40136=>"110011010",
  40137=>"101110000",
  40138=>"100100001",
  40139=>"100000100",
  40140=>"101110100",
  40141=>"111011110",
  40142=>"110001111",
  40143=>"001011111",
  40144=>"000011110",
  40145=>"011000110",
  40146=>"111010001",
  40147=>"010100100",
  40148=>"000101001",
  40149=>"111001111",
  40150=>"010110101",
  40151=>"001010101",
  40152=>"011001111",
  40153=>"010111001",
  40154=>"001000111",
  40155=>"100000011",
  40156=>"111110111",
  40157=>"100010010",
  40158=>"010111001",
  40159=>"111111111",
  40160=>"011111101",
  40161=>"000100101",
  40162=>"010001011",
  40163=>"111111110",
  40164=>"101011110",
  40165=>"011110000",
  40166=>"100111101",
  40167=>"000011100",
  40168=>"011110010",
  40169=>"110010010",
  40170=>"100010011",
  40171=>"101001011",
  40172=>"101011100",
  40173=>"101100101",
  40174=>"011010000",
  40175=>"100000100",
  40176=>"110111111",
  40177=>"111111111",
  40178=>"010110101",
  40179=>"001111111",
  40180=>"010111101",
  40181=>"010100010",
  40182=>"000111100",
  40183=>"010000100",
  40184=>"000010110",
  40185=>"100101010",
  40186=>"100000101",
  40187=>"010000000",
  40188=>"101110010",
  40189=>"100101111",
  40190=>"000010001",
  40191=>"110100110",
  40192=>"100010001",
  40193=>"111100001",
  40194=>"010001001",
  40195=>"001011110",
  40196=>"001101111",
  40197=>"000001100",
  40198=>"000011100",
  40199=>"100000010",
  40200=>"100010001",
  40201=>"000101011",
  40202=>"100000110",
  40203=>"110000110",
  40204=>"001001010",
  40205=>"001100010",
  40206=>"011010001",
  40207=>"101101000",
  40208=>"000010011",
  40209=>"010100011",
  40210=>"000000101",
  40211=>"111110100",
  40212=>"001111101",
  40213=>"110100010",
  40214=>"000010011",
  40215=>"100110100",
  40216=>"100000101",
  40217=>"110001111",
  40218=>"010011110",
  40219=>"111101010",
  40220=>"011100000",
  40221=>"100001010",
  40222=>"001011111",
  40223=>"111000100",
  40224=>"001000111",
  40225=>"001001001",
  40226=>"000000000",
  40227=>"001000010",
  40228=>"110100100",
  40229=>"001111001",
  40230=>"000000100",
  40231=>"100000010",
  40232=>"001110001",
  40233=>"110001001",
  40234=>"111010100",
  40235=>"100110101",
  40236=>"100111111",
  40237=>"010111100",
  40238=>"001110111",
  40239=>"100111111",
  40240=>"101111100",
  40241=>"101000011",
  40242=>"000001000",
  40243=>"000010011",
  40244=>"111101100",
  40245=>"110010100",
  40246=>"010111101",
  40247=>"000011001",
  40248=>"010000001",
  40249=>"001001111",
  40250=>"001110111",
  40251=>"011011000",
  40252=>"101001001",
  40253=>"010110111",
  40254=>"011110000",
  40255=>"001001010",
  40256=>"110110110",
  40257=>"101110100",
  40258=>"100010101",
  40259=>"100101011",
  40260=>"000011000",
  40261=>"110111111",
  40262=>"110000000",
  40263=>"110001000",
  40264=>"111010001",
  40265=>"000000001",
  40266=>"000011000",
  40267=>"000001101",
  40268=>"010010110",
  40269=>"111100110",
  40270=>"110111001",
  40271=>"000101001",
  40272=>"111110101",
  40273=>"010000000",
  40274=>"000110000",
  40275=>"111101100",
  40276=>"010011000",
  40277=>"110111110",
  40278=>"011111111",
  40279=>"001001001",
  40280=>"010001000",
  40281=>"000000000",
  40282=>"011010011",
  40283=>"100100101",
  40284=>"111000010",
  40285=>"101100110",
  40286=>"111001000",
  40287=>"001011011",
  40288=>"001111010",
  40289=>"100101101",
  40290=>"110000110",
  40291=>"001000111",
  40292=>"111011111",
  40293=>"110000001",
  40294=>"110101100",
  40295=>"100100010",
  40296=>"001000011",
  40297=>"111101000",
  40298=>"011010101",
  40299=>"010110110",
  40300=>"101111111",
  40301=>"011011000",
  40302=>"011000011",
  40303=>"001100011",
  40304=>"000110110",
  40305=>"100100101",
  40306=>"110111100",
  40307=>"100001110",
  40308=>"111100000",
  40309=>"111011101",
  40310=>"010110110",
  40311=>"010101101",
  40312=>"010101010",
  40313=>"101011000",
  40314=>"000011011",
  40315=>"000111101",
  40316=>"101110011",
  40317=>"100100100",
  40318=>"010011110",
  40319=>"110100100",
  40320=>"100100100",
  40321=>"011001000",
  40322=>"100100001",
  40323=>"111111010",
  40324=>"000110110",
  40325=>"110100011",
  40326=>"101111110",
  40327=>"011000001",
  40328=>"110001000",
  40329=>"110110010",
  40330=>"001111100",
  40331=>"110110110",
  40332=>"100101111",
  40333=>"001010010",
  40334=>"100000110",
  40335=>"111100000",
  40336=>"011111001",
  40337=>"000111000",
  40338=>"000001000",
  40339=>"010010000",
  40340=>"000100100",
  40341=>"000011000",
  40342=>"010101111",
  40343=>"101101001",
  40344=>"011000101",
  40345=>"000110010",
  40346=>"010100101",
  40347=>"000010000",
  40348=>"001010011",
  40349=>"011110011",
  40350=>"100011111",
  40351=>"010000100",
  40352=>"011101010",
  40353=>"101011001",
  40354=>"111100001",
  40355=>"000100010",
  40356=>"100100010",
  40357=>"010010100",
  40358=>"111101001",
  40359=>"101111111",
  40360=>"001101000",
  40361=>"101000110",
  40362=>"001011111",
  40363=>"001011001",
  40364=>"110000111",
  40365=>"000001010",
  40366=>"101000111",
  40367=>"110101110",
  40368=>"001001110",
  40369=>"111011010",
  40370=>"011101110",
  40371=>"110101000",
  40372=>"100111101",
  40373=>"001000001",
  40374=>"101110011",
  40375=>"000100110",
  40376=>"110010001",
  40377=>"101001111",
  40378=>"001111111",
  40379=>"001010010",
  40380=>"100001101",
  40381=>"111110000",
  40382=>"100111000",
  40383=>"010001111",
  40384=>"001000000",
  40385=>"000001110",
  40386=>"010110100",
  40387=>"001010101",
  40388=>"001000000",
  40389=>"111000000",
  40390=>"100011011",
  40391=>"111011100",
  40392=>"000000001",
  40393=>"011000111",
  40394=>"001000000",
  40395=>"001100110",
  40396=>"010100111",
  40397=>"110100011",
  40398=>"101110011",
  40399=>"000001111",
  40400=>"011001101",
  40401=>"111010011",
  40402=>"001001010",
  40403=>"011011110",
  40404=>"010011010",
  40405=>"000010010",
  40406=>"011010010",
  40407=>"110110101",
  40408=>"101101000",
  40409=>"001100101",
  40410=>"011000000",
  40411=>"110000001",
  40412=>"101100101",
  40413=>"010010001",
  40414=>"111101010",
  40415=>"010101000",
  40416=>"110000110",
  40417=>"001011001",
  40418=>"111011110",
  40419=>"000100010",
  40420=>"110000001",
  40421=>"000001101",
  40422=>"110100000",
  40423=>"001101101",
  40424=>"011110000",
  40425=>"101011001",
  40426=>"111100010",
  40427=>"011110010",
  40428=>"110100011",
  40429=>"000001101",
  40430=>"111011110",
  40431=>"001011010",
  40432=>"011001011",
  40433=>"101101010",
  40434=>"110010110",
  40435=>"011100000",
  40436=>"010111001",
  40437=>"100000001",
  40438=>"100110000",
  40439=>"111001010",
  40440=>"000111100",
  40441=>"111001100",
  40442=>"111000010",
  40443=>"100100000",
  40444=>"110100011",
  40445=>"101010100",
  40446=>"100000010",
  40447=>"010111010",
  40448=>"011111111",
  40449=>"101100110",
  40450=>"111101010",
  40451=>"010000111",
  40452=>"110001000",
  40453=>"111101001",
  40454=>"011011000",
  40455=>"000111000",
  40456=>"110011000",
  40457=>"001010010",
  40458=>"010000010",
  40459=>"100001001",
  40460=>"110001101",
  40461=>"000000110",
  40462=>"000000000",
  40463=>"011111001",
  40464=>"101000101",
  40465=>"110001101",
  40466=>"110010010",
  40467=>"010010001",
  40468=>"011111111",
  40469=>"100101011",
  40470=>"011000000",
  40471=>"101110010",
  40472=>"011110001",
  40473=>"000111010",
  40474=>"011000110",
  40475=>"001000001",
  40476=>"100010001",
  40477=>"101100011",
  40478=>"000111001",
  40479=>"101100100",
  40480=>"011101111",
  40481=>"100001100",
  40482=>"010111101",
  40483=>"010010100",
  40484=>"101001100",
  40485=>"001111110",
  40486=>"100011110",
  40487=>"000100110",
  40488=>"101000011",
  40489=>"111100011",
  40490=>"100000001",
  40491=>"101111101",
  40492=>"111101100",
  40493=>"001000001",
  40494=>"110101001",
  40495=>"110110101",
  40496=>"011000010",
  40497=>"011010010",
  40498=>"010010011",
  40499=>"100100111",
  40500=>"010110000",
  40501=>"011011000",
  40502=>"100010100",
  40503=>"000101011",
  40504=>"001101100",
  40505=>"111011001",
  40506=>"100001001",
  40507=>"001011000",
  40508=>"100010101",
  40509=>"110110111",
  40510=>"010001100",
  40511=>"101100001",
  40512=>"000001010",
  40513=>"011101100",
  40514=>"000111110",
  40515=>"111101100",
  40516=>"100101100",
  40517=>"111111000",
  40518=>"101101011",
  40519=>"010001001",
  40520=>"001100100",
  40521=>"001110110",
  40522=>"110010100",
  40523=>"000010001",
  40524=>"101000000",
  40525=>"001110100",
  40526=>"100101110",
  40527=>"001101100",
  40528=>"001111001",
  40529=>"101001010",
  40530=>"000101001",
  40531=>"100000111",
  40532=>"000100110",
  40533=>"110001010",
  40534=>"011011000",
  40535=>"000010100",
  40536=>"101101101",
  40537=>"001111110",
  40538=>"001011101",
  40539=>"110010000",
  40540=>"011000100",
  40541=>"010000110",
  40542=>"100111111",
  40543=>"000000000",
  40544=>"101101100",
  40545=>"001010001",
  40546=>"111110101",
  40547=>"100000010",
  40548=>"111110110",
  40549=>"001011000",
  40550=>"010010010",
  40551=>"001001000",
  40552=>"110101011",
  40553=>"110100001",
  40554=>"011111101",
  40555=>"000010100",
  40556=>"110011000",
  40557=>"101110001",
  40558=>"100110000",
  40559=>"011011011",
  40560=>"010100111",
  40561=>"111110111",
  40562=>"011011110",
  40563=>"000011000",
  40564=>"010000001",
  40565=>"110111101",
  40566=>"000001100",
  40567=>"111101110",
  40568=>"100011101",
  40569=>"100010101",
  40570=>"100011110",
  40571=>"101110100",
  40572=>"101101100",
  40573=>"000101000",
  40574=>"000010000",
  40575=>"000001001",
  40576=>"101001011",
  40577=>"100000011",
  40578=>"100111010",
  40579=>"110111011",
  40580=>"100110111",
  40581=>"101111010",
  40582=>"100000010",
  40583=>"111110011",
  40584=>"111111101",
  40585=>"000111101",
  40586=>"010010100",
  40587=>"010011100",
  40588=>"101001101",
  40589=>"110010011",
  40590=>"111000100",
  40591=>"101011110",
  40592=>"010000101",
  40593=>"111010101",
  40594=>"010100001",
  40595=>"101010011",
  40596=>"101010101",
  40597=>"101111100",
  40598=>"000101100",
  40599=>"010101001",
  40600=>"100010000",
  40601=>"100101000",
  40602=>"010000100",
  40603=>"110011001",
  40604=>"110000001",
  40605=>"001111111",
  40606=>"010000110",
  40607=>"001000001",
  40608=>"111000010",
  40609=>"000000111",
  40610=>"000011100",
  40611=>"001101011",
  40612=>"110101000",
  40613=>"011101011",
  40614=>"001000100",
  40615=>"001011010",
  40616=>"000010010",
  40617=>"111101000",
  40618=>"000001001",
  40619=>"010001101",
  40620=>"010100000",
  40621=>"011100010",
  40622=>"000110100",
  40623=>"101011100",
  40624=>"010101010",
  40625=>"001100011",
  40626=>"010001010",
  40627=>"101110001",
  40628=>"010010110",
  40629=>"010111000",
  40630=>"001100001",
  40631=>"111011101",
  40632=>"000100100",
  40633=>"100001110",
  40634=>"000011000",
  40635=>"101001010",
  40636=>"010011110",
  40637=>"010110100",
  40638=>"011101001",
  40639=>"110010100",
  40640=>"001110100",
  40641=>"011001100",
  40642=>"000111001",
  40643=>"111100000",
  40644=>"111000001",
  40645=>"001001001",
  40646=>"100001000",
  40647=>"000000110",
  40648=>"001101101",
  40649=>"001000010",
  40650=>"000001010",
  40651=>"111111000",
  40652=>"001110101",
  40653=>"110010000",
  40654=>"111010111",
  40655=>"000000100",
  40656=>"010011101",
  40657=>"010001111",
  40658=>"110111101",
  40659=>"010110111",
  40660=>"101101000",
  40661=>"101111101",
  40662=>"010010000",
  40663=>"011001000",
  40664=>"100000010",
  40665=>"111001100",
  40666=>"111001101",
  40667=>"001101101",
  40668=>"101110000",
  40669=>"001101000",
  40670=>"100111011",
  40671=>"000011101",
  40672=>"101010100",
  40673=>"111010101",
  40674=>"010011110",
  40675=>"011010110",
  40676=>"011110111",
  40677=>"010011110",
  40678=>"110001000",
  40679=>"000101011",
  40680=>"100111111",
  40681=>"001101000",
  40682=>"101001001",
  40683=>"111101010",
  40684=>"010001101",
  40685=>"000101010",
  40686=>"000001111",
  40687=>"111011010",
  40688=>"000101011",
  40689=>"100101010",
  40690=>"111100100",
  40691=>"111110010",
  40692=>"110111111",
  40693=>"111110010",
  40694=>"000100110",
  40695=>"011101110",
  40696=>"010001111",
  40697=>"110100010",
  40698=>"110110000",
  40699=>"010100000",
  40700=>"010110001",
  40701=>"110000111",
  40702=>"000011111",
  40703=>"111000101",
  40704=>"100100001",
  40705=>"001010011",
  40706=>"000010000",
  40707=>"011010001",
  40708=>"100010111",
  40709=>"101101001",
  40710=>"110010100",
  40711=>"001100101",
  40712=>"001111100",
  40713=>"010100100",
  40714=>"000011111",
  40715=>"110110010",
  40716=>"010101010",
  40717=>"011110111",
  40718=>"100100101",
  40719=>"011010110",
  40720=>"011110011",
  40721=>"001110011",
  40722=>"011011111",
  40723=>"110101111",
  40724=>"101100000",
  40725=>"011000001",
  40726=>"010010011",
  40727=>"000110101",
  40728=>"000101101",
  40729=>"101111101",
  40730=>"110110010",
  40731=>"101000000",
  40732=>"011111111",
  40733=>"011011010",
  40734=>"010001010",
  40735=>"110110010",
  40736=>"101010110",
  40737=>"011001010",
  40738=>"001010111",
  40739=>"010100110",
  40740=>"011001000",
  40741=>"010010101",
  40742=>"001111100",
  40743=>"011110101",
  40744=>"111111010",
  40745=>"101010111",
  40746=>"101111100",
  40747=>"001111110",
  40748=>"111100111",
  40749=>"111100011",
  40750=>"110000101",
  40751=>"111100100",
  40752=>"111000000",
  40753=>"010010010",
  40754=>"100110000",
  40755=>"001000001",
  40756=>"110111000",
  40757=>"011000111",
  40758=>"110110000",
  40759=>"100111111",
  40760=>"011010000",
  40761=>"000001000",
  40762=>"011100110",
  40763=>"001110100",
  40764=>"111111100",
  40765=>"100010011",
  40766=>"000010011",
  40767=>"100101101",
  40768=>"101011100",
  40769=>"010111110",
  40770=>"111010000",
  40771=>"010110010",
  40772=>"110001001",
  40773=>"110100111",
  40774=>"110011100",
  40775=>"110010110",
  40776=>"010000010",
  40777=>"000000010",
  40778=>"001100011",
  40779=>"000111010",
  40780=>"011000110",
  40781=>"001110101",
  40782=>"000100001",
  40783=>"000000010",
  40784=>"001111011",
  40785=>"100000101",
  40786=>"000000110",
  40787=>"010001010",
  40788=>"000000011",
  40789=>"100101000",
  40790=>"101001001",
  40791=>"111000011",
  40792=>"010100011",
  40793=>"010000010",
  40794=>"111010010",
  40795=>"001010001",
  40796=>"111010011",
  40797=>"001001010",
  40798=>"000000000",
  40799=>"010010011",
  40800=>"000110111",
  40801=>"010001010",
  40802=>"010010111",
  40803=>"110010111",
  40804=>"111111011",
  40805=>"001000110",
  40806=>"101011110",
  40807=>"000000010",
  40808=>"100100101",
  40809=>"010011110",
  40810=>"011100100",
  40811=>"000000111",
  40812=>"101100011",
  40813=>"110100010",
  40814=>"010111001",
  40815=>"011101000",
  40816=>"100011101",
  40817=>"111100101",
  40818=>"000011111",
  40819=>"101110000",
  40820=>"111100101",
  40821=>"100011111",
  40822=>"010101001",
  40823=>"101101010",
  40824=>"110100110",
  40825=>"011111101",
  40826=>"110001011",
  40827=>"101010000",
  40828=>"011011000",
  40829=>"011000011",
  40830=>"111011010",
  40831=>"001110100",
  40832=>"011110000",
  40833=>"000100010",
  40834=>"110000101",
  40835=>"000001001",
  40836=>"000001001",
  40837=>"111001101",
  40838=>"010100100",
  40839=>"100110101",
  40840=>"001010111",
  40841=>"100110000",
  40842=>"111101001",
  40843=>"010100110",
  40844=>"011101111",
  40845=>"000001100",
  40846=>"110110101",
  40847=>"100001101",
  40848=>"100001111",
  40849=>"000110101",
  40850=>"010111101",
  40851=>"011001010",
  40852=>"001101010",
  40853=>"011011100",
  40854=>"001000111",
  40855=>"100000001",
  40856=>"011010001",
  40857=>"010000101",
  40858=>"001001100",
  40859=>"110101011",
  40860=>"001001100",
  40861=>"100001101",
  40862=>"000010110",
  40863=>"000010100",
  40864=>"101101010",
  40865=>"011011001",
  40866=>"000011010",
  40867=>"010001010",
  40868=>"111101001",
  40869=>"101011001",
  40870=>"100010100",
  40871=>"101111011",
  40872=>"111010111",
  40873=>"110011001",
  40874=>"111111011",
  40875=>"100111001",
  40876=>"101010000",
  40877=>"000110000",
  40878=>"111100011",
  40879=>"001110000",
  40880=>"111001011",
  40881=>"100001111",
  40882=>"111110001",
  40883=>"110111010",
  40884=>"000000010",
  40885=>"101101100",
  40886=>"110101101",
  40887=>"111011010",
  40888=>"001000001",
  40889=>"010110111",
  40890=>"111010110",
  40891=>"110000011",
  40892=>"001101101",
  40893=>"110010001",
  40894=>"001101001",
  40895=>"100000101",
  40896=>"011000100",
  40897=>"101101111",
  40898=>"100010101",
  40899=>"000010101",
  40900=>"001010110",
  40901=>"110000100",
  40902=>"000010110",
  40903=>"100111101",
  40904=>"111000010",
  40905=>"111011010",
  40906=>"111100110",
  40907=>"000000000",
  40908=>"010000101",
  40909=>"111100101",
  40910=>"000011100",
  40911=>"100010111",
  40912=>"010001101",
  40913=>"011101001",
  40914=>"000001110",
  40915=>"111010011",
  40916=>"011111111",
  40917=>"000010001",
  40918=>"111010111",
  40919=>"000011001",
  40920=>"111111101",
  40921=>"001000100",
  40922=>"111010011",
  40923=>"011110000",
  40924=>"010001100",
  40925=>"011001000",
  40926=>"010110111",
  40927=>"101011111",
  40928=>"101011111",
  40929=>"010111011",
  40930=>"100101000",
  40931=>"001110111",
  40932=>"110110010",
  40933=>"001111000",
  40934=>"110010010",
  40935=>"110001111",
  40936=>"001010110",
  40937=>"101000000",
  40938=>"010101100",
  40939=>"100101101",
  40940=>"000000111",
  40941=>"011010000",
  40942=>"000101001",
  40943=>"110010001",
  40944=>"100100110",
  40945=>"010001100",
  40946=>"100010100",
  40947=>"010010111",
  40948=>"110010000",
  40949=>"000010100",
  40950=>"101110001",
  40951=>"011010010",
  40952=>"000001110",
  40953=>"001100111",
  40954=>"001111011",
  40955=>"101111000",
  40956=>"100111101",
  40957=>"100000000",
  40958=>"100000000",
  40959=>"110011010",
  40960=>"100011001",
  40961=>"101100111",
  40962=>"010011110",
  40963=>"010011010",
  40964=>"100101010",
  40965=>"110100101",
  40966=>"100000110",
  40967=>"011110000",
  40968=>"010000100",
  40969=>"101001100",
  40970=>"001001010",
  40971=>"001001010",
  40972=>"001101000",
  40973=>"101111111",
  40974=>"111011000",
  40975=>"000011111",
  40976=>"110111100",
  40977=>"001001001",
  40978=>"001110101",
  40979=>"010101000",
  40980=>"101010111",
  40981=>"110011101",
  40982=>"111101011",
  40983=>"100010011",
  40984=>"110010111",
  40985=>"110000000",
  40986=>"010110110",
  40987=>"101001000",
  40988=>"010001110",
  40989=>"001101110",
  40990=>"101100100",
  40991=>"110100111",
  40992=>"101111010",
  40993=>"011000000",
  40994=>"001000111",
  40995=>"100101000",
  40996=>"010011000",
  40997=>"100010101",
  40998=>"010011000",
  40999=>"000001111",
  41000=>"001010110",
  41001=>"010010000",
  41002=>"010010100",
  41003=>"011000001",
  41004=>"001101000",
  41005=>"110100000",
  41006=>"001100110",
  41007=>"111101000",
  41008=>"111010100",
  41009=>"011111110",
  41010=>"001111111",
  41011=>"010111001",
  41012=>"011110101",
  41013=>"000110000",
  41014=>"111101001",
  41015=>"001111011",
  41016=>"100000101",
  41017=>"000111100",
  41018=>"000001100",
  41019=>"100001001",
  41020=>"100111100",
  41021=>"100011010",
  41022=>"111000010",
  41023=>"011010000",
  41024=>"101100000",
  41025=>"001110011",
  41026=>"011000011",
  41027=>"110100100",
  41028=>"110011100",
  41029=>"000111000",
  41030=>"001001000",
  41031=>"010101011",
  41032=>"110111010",
  41033=>"110101100",
  41034=>"000001000",
  41035=>"000011011",
  41036=>"110011000",
  41037=>"000000111",
  41038=>"001111101",
  41039=>"101100101",
  41040=>"100110011",
  41041=>"000010110",
  41042=>"110101000",
  41043=>"011011110",
  41044=>"010101101",
  41045=>"100001110",
  41046=>"110100110",
  41047=>"101011010",
  41048=>"011111011",
  41049=>"110000000",
  41050=>"110101100",
  41051=>"011111010",
  41052=>"110110010",
  41053=>"000101110",
  41054=>"011000000",
  41055=>"100000110",
  41056=>"111100110",
  41057=>"100010110",
  41058=>"100011101",
  41059=>"001001000",
  41060=>"011110011",
  41061=>"001100001",
  41062=>"100101110",
  41063=>"100110111",
  41064=>"101100010",
  41065=>"010111110",
  41066=>"110100110",
  41067=>"100100010",
  41068=>"000111011",
  41069=>"100011011",
  41070=>"001100110",
  41071=>"101010000",
  41072=>"001110010",
  41073=>"011010100",
  41074=>"100001010",
  41075=>"000111110",
  41076=>"101101110",
  41077=>"101100000",
  41078=>"001000000",
  41079=>"101001000",
  41080=>"011001000",
  41081=>"000111110",
  41082=>"000000010",
  41083=>"011010101",
  41084=>"111100101",
  41085=>"111000001",
  41086=>"010111000",
  41087=>"110011001",
  41088=>"000010110",
  41089=>"110100101",
  41090=>"000001001",
  41091=>"000011011",
  41092=>"111101001",
  41093=>"111010101",
  41094=>"111111100",
  41095=>"110001110",
  41096=>"000000010",
  41097=>"100011001",
  41098=>"100011000",
  41099=>"000110111",
  41100=>"000001101",
  41101=>"010000000",
  41102=>"010010001",
  41103=>"000010100",
  41104=>"110000000",
  41105=>"111101101",
  41106=>"111100111",
  41107=>"001000110",
  41108=>"100011111",
  41109=>"000101000",
  41110=>"101010000",
  41111=>"101001011",
  41112=>"000000111",
  41113=>"001110001",
  41114=>"110101111",
  41115=>"010100100",
  41116=>"010101111",
  41117=>"111110111",
  41118=>"001101001",
  41119=>"001110010",
  41120=>"100011010",
  41121=>"011110111",
  41122=>"111000111",
  41123=>"100010111",
  41124=>"011110010",
  41125=>"000011001",
  41126=>"001000001",
  41127=>"000110000",
  41128=>"011000011",
  41129=>"010000001",
  41130=>"001011000",
  41131=>"111010001",
  41132=>"010011101",
  41133=>"101111011",
  41134=>"101011101",
  41135=>"001111100",
  41136=>"111010011",
  41137=>"000100100",
  41138=>"000101100",
  41139=>"000111001",
  41140=>"001101011",
  41141=>"110110011",
  41142=>"100001001",
  41143=>"101000100",
  41144=>"101011011",
  41145=>"111011111",
  41146=>"001101100",
  41147=>"110001101",
  41148=>"100110011",
  41149=>"001010000",
  41150=>"000000110",
  41151=>"100011010",
  41152=>"111011100",
  41153=>"101000010",
  41154=>"001100100",
  41155=>"111100101",
  41156=>"011110001",
  41157=>"101010011",
  41158=>"011100111",
  41159=>"111001001",
  41160=>"111000100",
  41161=>"001110000",
  41162=>"010000110",
  41163=>"111010110",
  41164=>"011011101",
  41165=>"111000001",
  41166=>"001111000",
  41167=>"001000101",
  41168=>"110011011",
  41169=>"100000110",
  41170=>"110100011",
  41171=>"001001000",
  41172=>"010100111",
  41173=>"000010101",
  41174=>"001110100",
  41175=>"000000000",
  41176=>"011100001",
  41177=>"100011101",
  41178=>"001010100",
  41179=>"110100000",
  41180=>"101101100",
  41181=>"001101110",
  41182=>"101001101",
  41183=>"110111001",
  41184=>"011101010",
  41185=>"111000110",
  41186=>"101100111",
  41187=>"100101000",
  41188=>"100101101",
  41189=>"101011111",
  41190=>"000010011",
  41191=>"001000000",
  41192=>"010110010",
  41193=>"000001100",
  41194=>"110111101",
  41195=>"111111110",
  41196=>"011011100",
  41197=>"011111101",
  41198=>"101010011",
  41199=>"101110011",
  41200=>"001001001",
  41201=>"101110101",
  41202=>"000011110",
  41203=>"111111100",
  41204=>"011110111",
  41205=>"100110110",
  41206=>"101000011",
  41207=>"110011000",
  41208=>"010100101",
  41209=>"001011100",
  41210=>"001000001",
  41211=>"110100101",
  41212=>"001101011",
  41213=>"101011111",
  41214=>"010000000",
  41215=>"110011101",
  41216=>"001100001",
  41217=>"000100111",
  41218=>"000111010",
  41219=>"111011100",
  41220=>"110110110",
  41221=>"101110111",
  41222=>"011100001",
  41223=>"100000010",
  41224=>"111110101",
  41225=>"110001010",
  41226=>"010111001",
  41227=>"101100100",
  41228=>"110010100",
  41229=>"000000000",
  41230=>"100100011",
  41231=>"101001011",
  41232=>"111010011",
  41233=>"001000110",
  41234=>"100010000",
  41235=>"111000010",
  41236=>"010000100",
  41237=>"011110010",
  41238=>"000101000",
  41239=>"111000000",
  41240=>"101001001",
  41241=>"001011001",
  41242=>"010001001",
  41243=>"100010011",
  41244=>"010101000",
  41245=>"001001111",
  41246=>"111111110",
  41247=>"000110100",
  41248=>"000110101",
  41249=>"111111000",
  41250=>"101101000",
  41251=>"001110101",
  41252=>"001001110",
  41253=>"111001000",
  41254=>"100100111",
  41255=>"110111011",
  41256=>"010111001",
  41257=>"011010001",
  41258=>"100111101",
  41259=>"111010101",
  41260=>"010000011",
  41261=>"101010001",
  41262=>"010011001",
  41263=>"100110100",
  41264=>"001101101",
  41265=>"110001101",
  41266=>"110100110",
  41267=>"110011111",
  41268=>"101001111",
  41269=>"011011111",
  41270=>"000000100",
  41271=>"001010000",
  41272=>"110001000",
  41273=>"010011101",
  41274=>"100100100",
  41275=>"100010000",
  41276=>"000111101",
  41277=>"011010010",
  41278=>"100101101",
  41279=>"000010000",
  41280=>"011100110",
  41281=>"010101011",
  41282=>"110111111",
  41283=>"100010100",
  41284=>"001000011",
  41285=>"110110000",
  41286=>"011010011",
  41287=>"010111000",
  41288=>"011101000",
  41289=>"110110111",
  41290=>"101101000",
  41291=>"110111110",
  41292=>"001110000",
  41293=>"000001011",
  41294=>"000111011",
  41295=>"010000010",
  41296=>"110100001",
  41297=>"110100110",
  41298=>"100101110",
  41299=>"011001101",
  41300=>"010100001",
  41301=>"111001111",
  41302=>"111110000",
  41303=>"110101100",
  41304=>"000001000",
  41305=>"000011001",
  41306=>"101001011",
  41307=>"001010011",
  41308=>"011111110",
  41309=>"000011111",
  41310=>"110011011",
  41311=>"111100001",
  41312=>"011001101",
  41313=>"000111010",
  41314=>"000110000",
  41315=>"011011111",
  41316=>"110100101",
  41317=>"100001000",
  41318=>"110001111",
  41319=>"010000000",
  41320=>"010111110",
  41321=>"001011010",
  41322=>"111110111",
  41323=>"101001000",
  41324=>"010110000",
  41325=>"110101111",
  41326=>"011001000",
  41327=>"010100111",
  41328=>"110010011",
  41329=>"001110100",
  41330=>"001011110",
  41331=>"111001111",
  41332=>"010010111",
  41333=>"101000100",
  41334=>"010001010",
  41335=>"011111011",
  41336=>"000010011",
  41337=>"001100011",
  41338=>"100000101",
  41339=>"101010111",
  41340=>"110001111",
  41341=>"111011111",
  41342=>"011000001",
  41343=>"111111001",
  41344=>"101111111",
  41345=>"000011100",
  41346=>"000101110",
  41347=>"111100011",
  41348=>"111000101",
  41349=>"011000110",
  41350=>"101101111",
  41351=>"101100000",
  41352=>"100111100",
  41353=>"110011011",
  41354=>"101100101",
  41355=>"111111011",
  41356=>"110010000",
  41357=>"001000000",
  41358=>"111010001",
  41359=>"011001101",
  41360=>"101100110",
  41361=>"100011111",
  41362=>"010111101",
  41363=>"110010011",
  41364=>"001101110",
  41365=>"010011111",
  41366=>"001011000",
  41367=>"000101000",
  41368=>"111010011",
  41369=>"100100000",
  41370=>"000100001",
  41371=>"101001100",
  41372=>"001101100",
  41373=>"011010001",
  41374=>"100001000",
  41375=>"111001100",
  41376=>"110101100",
  41377=>"011101001",
  41378=>"011101110",
  41379=>"100110010",
  41380=>"011110000",
  41381=>"101110011",
  41382=>"011001001",
  41383=>"010110100",
  41384=>"110011111",
  41385=>"001000111",
  41386=>"010111011",
  41387=>"110111111",
  41388=>"111011101",
  41389=>"010000011",
  41390=>"000110101",
  41391=>"100001101",
  41392=>"100111110",
  41393=>"110100111",
  41394=>"110100110",
  41395=>"111110101",
  41396=>"110110111",
  41397=>"000000000",
  41398=>"110111101",
  41399=>"100110011",
  41400=>"010110101",
  41401=>"000110000",
  41402=>"101110100",
  41403=>"101110110",
  41404=>"100111110",
  41405=>"111011101",
  41406=>"001010100",
  41407=>"111000101",
  41408=>"010011010",
  41409=>"011011011",
  41410=>"000100010",
  41411=>"111011010",
  41412=>"010101000",
  41413=>"111000011",
  41414=>"101111111",
  41415=>"110000000",
  41416=>"010101001",
  41417=>"010001101",
  41418=>"000000011",
  41419=>"101000011",
  41420=>"001011011",
  41421=>"101100011",
  41422=>"101111101",
  41423=>"000111110",
  41424=>"001001110",
  41425=>"001001010",
  41426=>"001010000",
  41427=>"111100101",
  41428=>"110100101",
  41429=>"101010010",
  41430=>"111111010",
  41431=>"100110000",
  41432=>"101010100",
  41433=>"100011101",
  41434=>"010111110",
  41435=>"011100001",
  41436=>"110011001",
  41437=>"010000011",
  41438=>"010100001",
  41439=>"000001000",
  41440=>"010110010",
  41441=>"000110000",
  41442=>"011111110",
  41443=>"000111011",
  41444=>"011110111",
  41445=>"011011100",
  41446=>"100111001",
  41447=>"000011111",
  41448=>"100000110",
  41449=>"111011111",
  41450=>"011111010",
  41451=>"111100110",
  41452=>"100000100",
  41453=>"101010000",
  41454=>"100001111",
  41455=>"100001101",
  41456=>"011001110",
  41457=>"010010010",
  41458=>"010001111",
  41459=>"010001100",
  41460=>"001011110",
  41461=>"101010011",
  41462=>"100111000",
  41463=>"111000011",
  41464=>"100001100",
  41465=>"101011011",
  41466=>"001001011",
  41467=>"010111011",
  41468=>"011010110",
  41469=>"111110011",
  41470=>"110000111",
  41471=>"000100010",
  41472=>"010111011",
  41473=>"010111011",
  41474=>"111010101",
  41475=>"010000111",
  41476=>"011101100",
  41477=>"110111100",
  41478=>"111000011",
  41479=>"001011111",
  41480=>"111100100",
  41481=>"000010110",
  41482=>"000011101",
  41483=>"010001100",
  41484=>"010001010",
  41485=>"111111001",
  41486=>"111000000",
  41487=>"100101011",
  41488=>"110001001",
  41489=>"011101101",
  41490=>"000000001",
  41491=>"100101000",
  41492=>"101000001",
  41493=>"011000100",
  41494=>"011101101",
  41495=>"101000011",
  41496=>"110000010",
  41497=>"001001100",
  41498=>"101010010",
  41499=>"001010011",
  41500=>"010110101",
  41501=>"111010101",
  41502=>"101111111",
  41503=>"000110000",
  41504=>"101000000",
  41505=>"011001100",
  41506=>"110010010",
  41507=>"001110000",
  41508=>"110011110",
  41509=>"010110100",
  41510=>"111110000",
  41511=>"010111111",
  41512=>"000010100",
  41513=>"101110100",
  41514=>"010010101",
  41515=>"111001111",
  41516=>"001101111",
  41517=>"101101010",
  41518=>"110101010",
  41519=>"011100110",
  41520=>"011111110",
  41521=>"110111001",
  41522=>"000000100",
  41523=>"010001000",
  41524=>"011101100",
  41525=>"010010000",
  41526=>"000100100",
  41527=>"100110011",
  41528=>"011110101",
  41529=>"111110000",
  41530=>"110101001",
  41531=>"010001111",
  41532=>"010001100",
  41533=>"000011000",
  41534=>"010100010",
  41535=>"001110010",
  41536=>"111111111",
  41537=>"100001110",
  41538=>"111110011",
  41539=>"110011000",
  41540=>"000000111",
  41541=>"010000000",
  41542=>"000001000",
  41543=>"011000001",
  41544=>"011101011",
  41545=>"001111111",
  41546=>"100001000",
  41547=>"100110110",
  41548=>"100000011",
  41549=>"100101101",
  41550=>"110110111",
  41551=>"110011001",
  41552=>"000001010",
  41553=>"000001011",
  41554=>"001011110",
  41555=>"101100000",
  41556=>"010001111",
  41557=>"100011001",
  41558=>"010010001",
  41559=>"011010001",
  41560=>"010010000",
  41561=>"000110000",
  41562=>"101000100",
  41563=>"100000101",
  41564=>"111100000",
  41565=>"110100011",
  41566=>"010000110",
  41567=>"011000111",
  41568=>"010001101",
  41569=>"100001000",
  41570=>"011101010",
  41571=>"111111100",
  41572=>"010011101",
  41573=>"010100011",
  41574=>"000011011",
  41575=>"100011111",
  41576=>"001110000",
  41577=>"110010110",
  41578=>"111010001",
  41579=>"011010010",
  41580=>"111010101",
  41581=>"010010010",
  41582=>"000010100",
  41583=>"000110000",
  41584=>"010010100",
  41585=>"100111010",
  41586=>"011001011",
  41587=>"110101111",
  41588=>"111110011",
  41589=>"110000001",
  41590=>"111110101",
  41591=>"100001011",
  41592=>"010010000",
  41593=>"101001010",
  41594=>"010000001",
  41595=>"010110011",
  41596=>"010001001",
  41597=>"111010110",
  41598=>"000100000",
  41599=>"010010001",
  41600=>"010000001",
  41601=>"101101111",
  41602=>"011101001",
  41603=>"100101010",
  41604=>"001001111",
  41605=>"111001111",
  41606=>"111110100",
  41607=>"101110100",
  41608=>"001011100",
  41609=>"001011100",
  41610=>"011001101",
  41611=>"011101101",
  41612=>"101100111",
  41613=>"001000111",
  41614=>"101010000",
  41615=>"011001000",
  41616=>"001001000",
  41617=>"101010001",
  41618=>"111001111",
  41619=>"111101101",
  41620=>"110111100",
  41621=>"001111101",
  41622=>"101110110",
  41623=>"001011011",
  41624=>"111010110",
  41625=>"000100101",
  41626=>"011100000",
  41627=>"011001010",
  41628=>"001010010",
  41629=>"000110010",
  41630=>"000011000",
  41631=>"100001001",
  41632=>"010101011",
  41633=>"001001111",
  41634=>"111111110",
  41635=>"000110100",
  41636=>"010010101",
  41637=>"111110101",
  41638=>"011010101",
  41639=>"000111111",
  41640=>"011110011",
  41641=>"010000011",
  41642=>"000011000",
  41643=>"000001101",
  41644=>"011010000",
  41645=>"011000101",
  41646=>"010100100",
  41647=>"111011011",
  41648=>"001100010",
  41649=>"100000000",
  41650=>"100010010",
  41651=>"010100011",
  41652=>"101111000",
  41653=>"011001110",
  41654=>"110100000",
  41655=>"010001101",
  41656=>"101001110",
  41657=>"100101000",
  41658=>"001110101",
  41659=>"001111100",
  41660=>"000011011",
  41661=>"010101011",
  41662=>"001010000",
  41663=>"000101110",
  41664=>"000011000",
  41665=>"011100100",
  41666=>"111101000",
  41667=>"111010011",
  41668=>"000001010",
  41669=>"100100101",
  41670=>"010111111",
  41671=>"100111001",
  41672=>"001000111",
  41673=>"010100011",
  41674=>"111100101",
  41675=>"001010000",
  41676=>"010011110",
  41677=>"111011001",
  41678=>"010101110",
  41679=>"110000010",
  41680=>"001011000",
  41681=>"100100101",
  41682=>"110101010",
  41683=>"001111001",
  41684=>"111011001",
  41685=>"001001010",
  41686=>"000011000",
  41687=>"110000011",
  41688=>"100111100",
  41689=>"100110000",
  41690=>"101100011",
  41691=>"001011010",
  41692=>"010101101",
  41693=>"010001011",
  41694=>"101011101",
  41695=>"001110001",
  41696=>"010110100",
  41697=>"000001100",
  41698=>"000011001",
  41699=>"011010010",
  41700=>"110010100",
  41701=>"010110010",
  41702=>"011100000",
  41703=>"011010010",
  41704=>"010100011",
  41705=>"101111110",
  41706=>"101101000",
  41707=>"110001001",
  41708=>"100100110",
  41709=>"111110100",
  41710=>"111110110",
  41711=>"100001000",
  41712=>"101011011",
  41713=>"001101011",
  41714=>"111001110",
  41715=>"011111100",
  41716=>"110011011",
  41717=>"001110001",
  41718=>"011111000",
  41719=>"110010111",
  41720=>"000101111",
  41721=>"111011000",
  41722=>"000110001",
  41723=>"011010110",
  41724=>"000101011",
  41725=>"011011001",
  41726=>"110011101",
  41727=>"010101111",
  41728=>"101011011",
  41729=>"001110010",
  41730=>"010110110",
  41731=>"000000110",
  41732=>"101101001",
  41733=>"000101101",
  41734=>"010001000",
  41735=>"000000110",
  41736=>"111000111",
  41737=>"001100011",
  41738=>"100001111",
  41739=>"100001001",
  41740=>"010001000",
  41741=>"110000111",
  41742=>"000100101",
  41743=>"110110000",
  41744=>"111111111",
  41745=>"101000010",
  41746=>"111000101",
  41747=>"100101100",
  41748=>"111101111",
  41749=>"101110000",
  41750=>"010011101",
  41751=>"100101000",
  41752=>"111111001",
  41753=>"101001110",
  41754=>"000101100",
  41755=>"010000001",
  41756=>"010011011",
  41757=>"100001100",
  41758=>"100110001",
  41759=>"011001001",
  41760=>"000001100",
  41761=>"110100000",
  41762=>"100010011",
  41763=>"001110110",
  41764=>"110100001",
  41765=>"001001101",
  41766=>"010111001",
  41767=>"001110100",
  41768=>"011111101",
  41769=>"100001100",
  41770=>"000011100",
  41771=>"101010110",
  41772=>"101011100",
  41773=>"010001101",
  41774=>"001000001",
  41775=>"000011101",
  41776=>"010100110",
  41777=>"001110100",
  41778=>"000100000",
  41779=>"110010100",
  41780=>"111100101",
  41781=>"101100010",
  41782=>"100100000",
  41783=>"000001001",
  41784=>"000110110",
  41785=>"000000010",
  41786=>"111000111",
  41787=>"010010010",
  41788=>"010011111",
  41789=>"100010110",
  41790=>"011010100",
  41791=>"101100111",
  41792=>"001110001",
  41793=>"001101011",
  41794=>"111101110",
  41795=>"111111001",
  41796=>"001011001",
  41797=>"111010111",
  41798=>"110111100",
  41799=>"111001111",
  41800=>"111001110",
  41801=>"111011100",
  41802=>"011101111",
  41803=>"101001110",
  41804=>"110110001",
  41805=>"111001110",
  41806=>"001001100",
  41807=>"101110100",
  41808=>"110010010",
  41809=>"011000011",
  41810=>"101010100",
  41811=>"000001100",
  41812=>"110110100",
  41813=>"011101111",
  41814=>"010111101",
  41815=>"110111011",
  41816=>"000010011",
  41817=>"010011000",
  41818=>"001110100",
  41819=>"111000001",
  41820=>"111100001",
  41821=>"110010101",
  41822=>"000011110",
  41823=>"000100110",
  41824=>"100110101",
  41825=>"000100011",
  41826=>"101110010",
  41827=>"100111010",
  41828=>"000111111",
  41829=>"010111100",
  41830=>"111101011",
  41831=>"100101001",
  41832=>"100000101",
  41833=>"010101100",
  41834=>"001011000",
  41835=>"010100011",
  41836=>"000000101",
  41837=>"100101101",
  41838=>"000011101",
  41839=>"010100011",
  41840=>"001000110",
  41841=>"011100011",
  41842=>"110110110",
  41843=>"101010011",
  41844=>"100101001",
  41845=>"111000110",
  41846=>"100000001",
  41847=>"011101000",
  41848=>"011100110",
  41849=>"100100101",
  41850=>"000110110",
  41851=>"011010100",
  41852=>"000011011",
  41853=>"110010111",
  41854=>"000110011",
  41855=>"110010100",
  41856=>"010011111",
  41857=>"111111101",
  41858=>"001100010",
  41859=>"101011000",
  41860=>"100101010",
  41861=>"110110011",
  41862=>"111111011",
  41863=>"011111101",
  41864=>"001111101",
  41865=>"000110010",
  41866=>"001000010",
  41867=>"101110111",
  41868=>"001110000",
  41869=>"100110111",
  41870=>"001011100",
  41871=>"111110111",
  41872=>"100000001",
  41873=>"111011011",
  41874=>"000100110",
  41875=>"001100000",
  41876=>"001010101",
  41877=>"100010110",
  41878=>"110110111",
  41879=>"111000100",
  41880=>"100011101",
  41881=>"110000000",
  41882=>"010110110",
  41883=>"000001101",
  41884=>"100010101",
  41885=>"001011001",
  41886=>"011111011",
  41887=>"000110110",
  41888=>"110111111",
  41889=>"101001000",
  41890=>"011010001",
  41891=>"111110010",
  41892=>"100010011",
  41893=>"101100111",
  41894=>"100101001",
  41895=>"000001100",
  41896=>"000000100",
  41897=>"010001101",
  41898=>"000111111",
  41899=>"010011110",
  41900=>"010001110",
  41901=>"001010010",
  41902=>"111110100",
  41903=>"110100100",
  41904=>"111000111",
  41905=>"010010000",
  41906=>"101111111",
  41907=>"010010010",
  41908=>"111011100",
  41909=>"000111011",
  41910=>"110110111",
  41911=>"101010100",
  41912=>"010010000",
  41913=>"110101111",
  41914=>"111001111",
  41915=>"001010100",
  41916=>"001110001",
  41917=>"101000011",
  41918=>"110011001",
  41919=>"011111111",
  41920=>"110111001",
  41921=>"101100010",
  41922=>"011100010",
  41923=>"001001010",
  41924=>"101101111",
  41925=>"101011101",
  41926=>"111101101",
  41927=>"000001101",
  41928=>"011001010",
  41929=>"111101011",
  41930=>"001000111",
  41931=>"010111000",
  41932=>"010100110",
  41933=>"000101110",
  41934=>"001100000",
  41935=>"111000010",
  41936=>"010110011",
  41937=>"100110111",
  41938=>"011010010",
  41939=>"010001101",
  41940=>"100101110",
  41941=>"010111000",
  41942=>"001101110",
  41943=>"100000101",
  41944=>"111001011",
  41945=>"011101110",
  41946=>"111100100",
  41947=>"010100010",
  41948=>"011101000",
  41949=>"011000011",
  41950=>"011101001",
  41951=>"111111111",
  41952=>"101111111",
  41953=>"001111111",
  41954=>"010001101",
  41955=>"000101111",
  41956=>"011110001",
  41957=>"011001101",
  41958=>"010111011",
  41959=>"101100100",
  41960=>"111111001",
  41961=>"101101010",
  41962=>"111110100",
  41963=>"010010010",
  41964=>"000000010",
  41965=>"101010011",
  41966=>"000000011",
  41967=>"001001011",
  41968=>"111111011",
  41969=>"100001101",
  41970=>"001100101",
  41971=>"010000010",
  41972=>"111110101",
  41973=>"111011001",
  41974=>"011011001",
  41975=>"100100111",
  41976=>"111001101",
  41977=>"000101101",
  41978=>"010101011",
  41979=>"000001011",
  41980=>"000011111",
  41981=>"111010111",
  41982=>"010001100",
  41983=>"001010001",
  41984=>"001101101",
  41985=>"001101111",
  41986=>"100110110",
  41987=>"000001101",
  41988=>"011001010",
  41989=>"111000100",
  41990=>"110010110",
  41991=>"100110010",
  41992=>"000001100",
  41993=>"000010011",
  41994=>"111101001",
  41995=>"110001010",
  41996=>"111011101",
  41997=>"011010110",
  41998=>"101010101",
  41999=>"101100100",
  42000=>"010110000",
  42001=>"110000110",
  42002=>"010111000",
  42003=>"010000110",
  42004=>"100001000",
  42005=>"000101110",
  42006=>"101110010",
  42007=>"000001111",
  42008=>"100100110",
  42009=>"110000101",
  42010=>"000111101",
  42011=>"100100101",
  42012=>"100000001",
  42013=>"111110010",
  42014=>"100110100",
  42015=>"100011101",
  42016=>"100011011",
  42017=>"100111000",
  42018=>"001011101",
  42019=>"111110100",
  42020=>"101111111",
  42021=>"010100000",
  42022=>"000000111",
  42023=>"000010000",
  42024=>"001000001",
  42025=>"100011110",
  42026=>"111100111",
  42027=>"011100000",
  42028=>"100100000",
  42029=>"010010010",
  42030=>"011110101",
  42031=>"111010100",
  42032=>"011111110",
  42033=>"110011111",
  42034=>"010111010",
  42035=>"111110001",
  42036=>"100000010",
  42037=>"001011010",
  42038=>"100011101",
  42039=>"110010110",
  42040=>"101110110",
  42041=>"010110110",
  42042=>"111000111",
  42043=>"101101101",
  42044=>"001101100",
  42045=>"000001110",
  42046=>"100101001",
  42047=>"011100001",
  42048=>"100000010",
  42049=>"100000001",
  42050=>"101001001",
  42051=>"100000101",
  42052=>"000100101",
  42053=>"011000011",
  42054=>"111111000",
  42055=>"010011100",
  42056=>"101101110",
  42057=>"101110010",
  42058=>"010000101",
  42059=>"110100111",
  42060=>"000000010",
  42061=>"001101000",
  42062=>"000001011",
  42063=>"111000111",
  42064=>"100110101",
  42065=>"110100000",
  42066=>"110101010",
  42067=>"101010011",
  42068=>"010000000",
  42069=>"101000111",
  42070=>"000011111",
  42071=>"100101000",
  42072=>"110110010",
  42073=>"100101110",
  42074=>"000100001",
  42075=>"111101100",
  42076=>"011101110",
  42077=>"001000101",
  42078=>"100110111",
  42079=>"001100011",
  42080=>"010001111",
  42081=>"001000000",
  42082=>"111011001",
  42083=>"101001111",
  42084=>"010001001",
  42085=>"011001010",
  42086=>"010100111",
  42087=>"000011111",
  42088=>"011000011",
  42089=>"110011110",
  42090=>"110001000",
  42091=>"111101000",
  42092=>"101001011",
  42093=>"011000101",
  42094=>"101101010",
  42095=>"001010011",
  42096=>"000101110",
  42097=>"010101101",
  42098=>"111101111",
  42099=>"111001011",
  42100=>"000110101",
  42101=>"010011011",
  42102=>"011110010",
  42103=>"001100011",
  42104=>"011001000",
  42105=>"011011010",
  42106=>"111101111",
  42107=>"100011100",
  42108=>"110000100",
  42109=>"010000000",
  42110=>"000100100",
  42111=>"100100000",
  42112=>"110000000",
  42113=>"011010111",
  42114=>"111100000",
  42115=>"010110011",
  42116=>"100001011",
  42117=>"100000001",
  42118=>"000110011",
  42119=>"111111110",
  42120=>"010001001",
  42121=>"010011011",
  42122=>"110100000",
  42123=>"000111110",
  42124=>"000000000",
  42125=>"001111000",
  42126=>"101110111",
  42127=>"111100000",
  42128=>"111101100",
  42129=>"001100010",
  42130=>"111000000",
  42131=>"111101011",
  42132=>"101110010",
  42133=>"000011100",
  42134=>"100011101",
  42135=>"000101011",
  42136=>"100101000",
  42137=>"101100100",
  42138=>"111110001",
  42139=>"111111111",
  42140=>"110000000",
  42141=>"101100000",
  42142=>"011100000",
  42143=>"001010011",
  42144=>"101010101",
  42145=>"000001101",
  42146=>"001000001",
  42147=>"001001000",
  42148=>"010010000",
  42149=>"000100111",
  42150=>"110101001",
  42151=>"001100000",
  42152=>"100101000",
  42153=>"011111101",
  42154=>"010100100",
  42155=>"001111010",
  42156=>"100100100",
  42157=>"110000101",
  42158=>"001101111",
  42159=>"001100110",
  42160=>"011001111",
  42161=>"000110001",
  42162=>"001011100",
  42163=>"010101001",
  42164=>"101101111",
  42165=>"001010111",
  42166=>"111111100",
  42167=>"001011000",
  42168=>"101010011",
  42169=>"000000101",
  42170=>"101110101",
  42171=>"000000010",
  42172=>"011000101",
  42173=>"110010011",
  42174=>"000000001",
  42175=>"111110111",
  42176=>"111100100",
  42177=>"101111011",
  42178=>"100111001",
  42179=>"101100010",
  42180=>"101100010",
  42181=>"000010100",
  42182=>"100011011",
  42183=>"110101001",
  42184=>"111011001",
  42185=>"011100010",
  42186=>"101111100",
  42187=>"110110010",
  42188=>"000101110",
  42189=>"010100001",
  42190=>"011001101",
  42191=>"101111111",
  42192=>"101000000",
  42193=>"010110101",
  42194=>"100001101",
  42195=>"000101100",
  42196=>"111000000",
  42197=>"011110011",
  42198=>"110010011",
  42199=>"100001000",
  42200=>"100000101",
  42201=>"010100101",
  42202=>"000101011",
  42203=>"010001011",
  42204=>"010111010",
  42205=>"111111111",
  42206=>"001000111",
  42207=>"001001000",
  42208=>"101100001",
  42209=>"100100010",
  42210=>"001010000",
  42211=>"100000000",
  42212=>"010001101",
  42213=>"000011001",
  42214=>"001000100",
  42215=>"011000001",
  42216=>"001010010",
  42217=>"000101011",
  42218=>"011100011",
  42219=>"100101110",
  42220=>"100100100",
  42221=>"100011001",
  42222=>"000001011",
  42223=>"100000111",
  42224=>"111010000",
  42225=>"100100011",
  42226=>"000000001",
  42227=>"101100100",
  42228=>"010011000",
  42229=>"011101001",
  42230=>"110111111",
  42231=>"000101100",
  42232=>"000000110",
  42233=>"101000011",
  42234=>"000011000",
  42235=>"111001101",
  42236=>"101011001",
  42237=>"000011110",
  42238=>"101101111",
  42239=>"011010111",
  42240=>"101010111",
  42241=>"111001101",
  42242=>"111001000",
  42243=>"010100111",
  42244=>"001001100",
  42245=>"100011001",
  42246=>"010101100",
  42247=>"010000100",
  42248=>"001011000",
  42249=>"001011111",
  42250=>"011101001",
  42251=>"010100010",
  42252=>"000011001",
  42253=>"011101101",
  42254=>"100010110",
  42255=>"011000011",
  42256=>"111100001",
  42257=>"111000111",
  42258=>"100101110",
  42259=>"111111000",
  42260=>"010110001",
  42261=>"000001001",
  42262=>"000011111",
  42263=>"001101010",
  42264=>"111011100",
  42265=>"001101011",
  42266=>"000110011",
  42267=>"010111001",
  42268=>"011100001",
  42269=>"000101001",
  42270=>"110000111",
  42271=>"011001001",
  42272=>"010010011",
  42273=>"100010110",
  42274=>"101011000",
  42275=>"001011011",
  42276=>"111000100",
  42277=>"110001001",
  42278=>"011010101",
  42279=>"101000110",
  42280=>"011101110",
  42281=>"110011001",
  42282=>"101010010",
  42283=>"011110011",
  42284=>"100010001",
  42285=>"000000011",
  42286=>"011100100",
  42287=>"011110010",
  42288=>"111000000",
  42289=>"000011110",
  42290=>"111011110",
  42291=>"111001001",
  42292=>"010100100",
  42293=>"101010000",
  42294=>"011011010",
  42295=>"101110111",
  42296=>"000000000",
  42297=>"110110100",
  42298=>"100101110",
  42299=>"101010010",
  42300=>"100011000",
  42301=>"101101110",
  42302=>"001100001",
  42303=>"111111010",
  42304=>"001000000",
  42305=>"000001011",
  42306=>"001101011",
  42307=>"100111100",
  42308=>"111001110",
  42309=>"010011011",
  42310=>"110000001",
  42311=>"101110000",
  42312=>"000101011",
  42313=>"100100011",
  42314=>"010000101",
  42315=>"110001010",
  42316=>"001111111",
  42317=>"111101011",
  42318=>"001100101",
  42319=>"011011101",
  42320=>"100000010",
  42321=>"100110001",
  42322=>"111110000",
  42323=>"101000110",
  42324=>"111011000",
  42325=>"111010100",
  42326=>"000100011",
  42327=>"001111100",
  42328=>"001100001",
  42329=>"010100011",
  42330=>"000001001",
  42331=>"011010110",
  42332=>"010010010",
  42333=>"011011101",
  42334=>"011011000",
  42335=>"000100001",
  42336=>"010100001",
  42337=>"011100100",
  42338=>"010000011",
  42339=>"010001001",
  42340=>"101111001",
  42341=>"101100000",
  42342=>"111111011",
  42343=>"111110101",
  42344=>"100100001",
  42345=>"001110011",
  42346=>"010010110",
  42347=>"001101010",
  42348=>"000011110",
  42349=>"010111111",
  42350=>"000100011",
  42351=>"010001111",
  42352=>"000001001",
  42353=>"011100100",
  42354=>"001110001",
  42355=>"010111001",
  42356=>"110101110",
  42357=>"100011011",
  42358=>"111110010",
  42359=>"111110101",
  42360=>"011110000",
  42361=>"000111101",
  42362=>"001000110",
  42363=>"001011100",
  42364=>"010011010",
  42365=>"111111111",
  42366=>"011101011",
  42367=>"101000100",
  42368=>"010000101",
  42369=>"001010101",
  42370=>"101010101",
  42371=>"010010010",
  42372=>"110100000",
  42373=>"100010100",
  42374=>"000101011",
  42375=>"011010000",
  42376=>"001000001",
  42377=>"000100001",
  42378=>"000100011",
  42379=>"101001101",
  42380=>"101011111",
  42381=>"010110111",
  42382=>"100101111",
  42383=>"001110000",
  42384=>"111010000",
  42385=>"000000111",
  42386=>"001001110",
  42387=>"000110001",
  42388=>"111011100",
  42389=>"100001100",
  42390=>"101110001",
  42391=>"000001111",
  42392=>"111111000",
  42393=>"111100100",
  42394=>"101110110",
  42395=>"001000100",
  42396=>"100010111",
  42397=>"110100010",
  42398=>"110111011",
  42399=>"111010011",
  42400=>"101100111",
  42401=>"000000000",
  42402=>"110010001",
  42403=>"010000100",
  42404=>"010010100",
  42405=>"000000110",
  42406=>"000101110",
  42407=>"011110101",
  42408=>"011000111",
  42409=>"011011101",
  42410=>"000100010",
  42411=>"000010000",
  42412=>"110010000",
  42413=>"010100101",
  42414=>"010000001",
  42415=>"111101111",
  42416=>"011100100",
  42417=>"011110001",
  42418=>"011010001",
  42419=>"110000110",
  42420=>"110011011",
  42421=>"001011110",
  42422=>"010110010",
  42423=>"111011001",
  42424=>"001011011",
  42425=>"111110011",
  42426=>"001000100",
  42427=>"111001111",
  42428=>"010000100",
  42429=>"010011101",
  42430=>"100111110",
  42431=>"001111010",
  42432=>"000111101",
  42433=>"000000010",
  42434=>"100100010",
  42435=>"001010101",
  42436=>"000001000",
  42437=>"110000000",
  42438=>"011111100",
  42439=>"000110011",
  42440=>"000001010",
  42441=>"110000100",
  42442=>"000000100",
  42443=>"100111101",
  42444=>"000000111",
  42445=>"100100011",
  42446=>"101000001",
  42447=>"111100011",
  42448=>"100100111",
  42449=>"001111110",
  42450=>"101111111",
  42451=>"010110100",
  42452=>"001111111",
  42453=>"000100000",
  42454=>"011001000",
  42455=>"111001111",
  42456=>"000010101",
  42457=>"101010110",
  42458=>"101010110",
  42459=>"111001000",
  42460=>"110001101",
  42461=>"100011100",
  42462=>"010111000",
  42463=>"000000101",
  42464=>"010011100",
  42465=>"010100000",
  42466=>"100001111",
  42467=>"101010000",
  42468=>"110001010",
  42469=>"110111110",
  42470=>"010010110",
  42471=>"001000000",
  42472=>"001001110",
  42473=>"000100101",
  42474=>"010000000",
  42475=>"010001111",
  42476=>"001110001",
  42477=>"011101111",
  42478=>"110111001",
  42479=>"111111000",
  42480=>"100010110",
  42481=>"010001011",
  42482=>"011010000",
  42483=>"001000010",
  42484=>"111000000",
  42485=>"000110010",
  42486=>"001010001",
  42487=>"000000011",
  42488=>"111001010",
  42489=>"111010010",
  42490=>"110101110",
  42491=>"111001000",
  42492=>"010111100",
  42493=>"010010000",
  42494=>"010111000",
  42495=>"111001101",
  42496=>"111011001",
  42497=>"110100011",
  42498=>"000111001",
  42499=>"001011001",
  42500=>"101100110",
  42501=>"000100010",
  42502=>"111100000",
  42503=>"010110001",
  42504=>"010101001",
  42505=>"000101011",
  42506=>"000101100",
  42507=>"000110010",
  42508=>"110101000",
  42509=>"000010000",
  42510=>"101101001",
  42511=>"101100011",
  42512=>"111010010",
  42513=>"111111000",
  42514=>"000111111",
  42515=>"101111000",
  42516=>"111100110",
  42517=>"010011111",
  42518=>"000100010",
  42519=>"100011111",
  42520=>"000110000",
  42521=>"011100010",
  42522=>"100000000",
  42523=>"011000011",
  42524=>"000100100",
  42525=>"101000010",
  42526=>"000001010",
  42527=>"000000001",
  42528=>"011010010",
  42529=>"011100110",
  42530=>"101100010",
  42531=>"100001110",
  42532=>"100011000",
  42533=>"000110010",
  42534=>"111100001",
  42535=>"010011010",
  42536=>"000101011",
  42537=>"100100100",
  42538=>"101001100",
  42539=>"101111101",
  42540=>"010101101",
  42541=>"000001011",
  42542=>"100001100",
  42543=>"011110000",
  42544=>"101001010",
  42545=>"101101001",
  42546=>"101001101",
  42547=>"111010101",
  42548=>"110000100",
  42549=>"111000001",
  42550=>"110011111",
  42551=>"010000111",
  42552=>"001110101",
  42553=>"101011000",
  42554=>"000000011",
  42555=>"100111000",
  42556=>"000011000",
  42557=>"011111011",
  42558=>"010110101",
  42559=>"010000110",
  42560=>"100000110",
  42561=>"010000000",
  42562=>"000100101",
  42563=>"011011111",
  42564=>"001111001",
  42565=>"100101000",
  42566=>"000000010",
  42567=>"011011111",
  42568=>"011000000",
  42569=>"101011001",
  42570=>"010111111",
  42571=>"010010110",
  42572=>"100000000",
  42573=>"000110101",
  42574=>"101111111",
  42575=>"000011011",
  42576=>"100101010",
  42577=>"001001010",
  42578=>"011100001",
  42579=>"001111110",
  42580=>"011000000",
  42581=>"000000000",
  42582=>"000011000",
  42583=>"000010000",
  42584=>"010111000",
  42585=>"000100011",
  42586=>"100101100",
  42587=>"101001111",
  42588=>"101100001",
  42589=>"000101111",
  42590=>"000111101",
  42591=>"111001010",
  42592=>"110001010",
  42593=>"010001000",
  42594=>"100110000",
  42595=>"010000100",
  42596=>"100111100",
  42597=>"111101110",
  42598=>"100001011",
  42599=>"000110101",
  42600=>"011100010",
  42601=>"000100001",
  42602=>"111101111",
  42603=>"101111111",
  42604=>"000100101",
  42605=>"011001111",
  42606=>"110010000",
  42607=>"111101000",
  42608=>"001100010",
  42609=>"000001100",
  42610=>"010001010",
  42611=>"000000011",
  42612=>"001100101",
  42613=>"100000010",
  42614=>"100110001",
  42615=>"111111000",
  42616=>"101001101",
  42617=>"101010110",
  42618=>"111010100",
  42619=>"010111001",
  42620=>"100110000",
  42621=>"011100111",
  42622=>"100100001",
  42623=>"100010100",
  42624=>"011010111",
  42625=>"110100111",
  42626=>"101100111",
  42627=>"110001011",
  42628=>"100001101",
  42629=>"111001010",
  42630=>"001000001",
  42631=>"010111101",
  42632=>"000011111",
  42633=>"100010111",
  42634=>"101101111",
  42635=>"111000101",
  42636=>"001101101",
  42637=>"001011000",
  42638=>"100111000",
  42639=>"111011010",
  42640=>"111101000",
  42641=>"001000010",
  42642=>"000000100",
  42643=>"111111011",
  42644=>"000100101",
  42645=>"010001001",
  42646=>"100111110",
  42647=>"111000100",
  42648=>"001101001",
  42649=>"011110010",
  42650=>"101101111",
  42651=>"100100101",
  42652=>"010110011",
  42653=>"110111111",
  42654=>"100101111",
  42655=>"001010000",
  42656=>"111001101",
  42657=>"010010100",
  42658=>"100001110",
  42659=>"000000011",
  42660=>"111101100",
  42661=>"001111110",
  42662=>"110000111",
  42663=>"101000000",
  42664=>"011111011",
  42665=>"101000000",
  42666=>"100001010",
  42667=>"101100010",
  42668=>"001110000",
  42669=>"000000001",
  42670=>"010100011",
  42671=>"101110111",
  42672=>"100111111",
  42673=>"011101011",
  42674=>"000001011",
  42675=>"110000110",
  42676=>"010100100",
  42677=>"000111001",
  42678=>"011100011",
  42679=>"100000010",
  42680=>"010111000",
  42681=>"010110110",
  42682=>"101101100",
  42683=>"001011101",
  42684=>"010001101",
  42685=>"101001110",
  42686=>"001110101",
  42687=>"000001010",
  42688=>"010000100",
  42689=>"100011011",
  42690=>"010000001",
  42691=>"011100001",
  42692=>"000111111",
  42693=>"000000000",
  42694=>"111100101",
  42695=>"001011000",
  42696=>"110000001",
  42697=>"111010100",
  42698=>"101010101",
  42699=>"011100011",
  42700=>"110101011",
  42701=>"000011110",
  42702=>"001111010",
  42703=>"000111110",
  42704=>"111000111",
  42705=>"000100100",
  42706=>"111110100",
  42707=>"001000001",
  42708=>"000011010",
  42709=>"100000011",
  42710=>"011001011",
  42711=>"110111001",
  42712=>"100010110",
  42713=>"010001101",
  42714=>"000000010",
  42715=>"010111010",
  42716=>"000100110",
  42717=>"001111011",
  42718=>"010010000",
  42719=>"110001011",
  42720=>"110111000",
  42721=>"011001101",
  42722=>"000001000",
  42723=>"011100000",
  42724=>"101001101",
  42725=>"100000001",
  42726=>"010111000",
  42727=>"100000001",
  42728=>"100110101",
  42729=>"011110001",
  42730=>"010001111",
  42731=>"001001111",
  42732=>"011100100",
  42733=>"011110000",
  42734=>"110010100",
  42735=>"010001010",
  42736=>"110011110",
  42737=>"010100110",
  42738=>"000100100",
  42739=>"100011010",
  42740=>"110111000",
  42741=>"001000111",
  42742=>"101110111",
  42743=>"111110100",
  42744=>"111111101",
  42745=>"111010011",
  42746=>"001111110",
  42747=>"011000010",
  42748=>"100001001",
  42749=>"001010100",
  42750=>"001100011",
  42751=>"111111001",
  42752=>"010111100",
  42753=>"111111110",
  42754=>"000100101",
  42755=>"000001101",
  42756=>"011101001",
  42757=>"000101111",
  42758=>"001111010",
  42759=>"010101110",
  42760=>"100110111",
  42761=>"011010111",
  42762=>"111100110",
  42763=>"110011101",
  42764=>"000100111",
  42765=>"000010110",
  42766=>"110000101",
  42767=>"010010011",
  42768=>"000011110",
  42769=>"101000011",
  42770=>"100110111",
  42771=>"001101010",
  42772=>"101010001",
  42773=>"110011000",
  42774=>"110110011",
  42775=>"010000010",
  42776=>"111000100",
  42777=>"011000001",
  42778=>"000010101",
  42779=>"111100110",
  42780=>"100000101",
  42781=>"000111111",
  42782=>"101111111",
  42783=>"010001101",
  42784=>"101100101",
  42785=>"011010110",
  42786=>"000101010",
  42787=>"101001010",
  42788=>"001011011",
  42789=>"010001000",
  42790=>"001010101",
  42791=>"100110101",
  42792=>"001111001",
  42793=>"101000110",
  42794=>"010101101",
  42795=>"110101100",
  42796=>"000101101",
  42797=>"000000010",
  42798=>"001000000",
  42799=>"110101000",
  42800=>"010111011",
  42801=>"101110011",
  42802=>"010110000",
  42803=>"100000010",
  42804=>"100110101",
  42805=>"100100101",
  42806=>"101000100",
  42807=>"010110101",
  42808=>"010110011",
  42809=>"100011001",
  42810=>"010011101",
  42811=>"111110110",
  42812=>"001111001",
  42813=>"000001011",
  42814=>"001000010",
  42815=>"110010100",
  42816=>"100100111",
  42817=>"110001011",
  42818=>"111011010",
  42819=>"111100111",
  42820=>"001101001",
  42821=>"000010001",
  42822=>"001100000",
  42823=>"111101011",
  42824=>"010100010",
  42825=>"111101100",
  42826=>"110010110",
  42827=>"111101100",
  42828=>"011100011",
  42829=>"000001000",
  42830=>"111111101",
  42831=>"100111001",
  42832=>"101001100",
  42833=>"111111110",
  42834=>"000001010",
  42835=>"101010111",
  42836=>"101010000",
  42837=>"101010000",
  42838=>"011001101",
  42839=>"100001000",
  42840=>"100001100",
  42841=>"111011101",
  42842=>"110110000",
  42843=>"100001110",
  42844=>"001001100",
  42845=>"000010011",
  42846=>"101100101",
  42847=>"111100100",
  42848=>"000000110",
  42849=>"010000110",
  42850=>"000110110",
  42851=>"101101010",
  42852=>"001001001",
  42853=>"101110010",
  42854=>"001101000",
  42855=>"011111000",
  42856=>"011100001",
  42857=>"110101111",
  42858=>"001010001",
  42859=>"100001000",
  42860=>"011111011",
  42861=>"101110100",
  42862=>"100101000",
  42863=>"111011000",
  42864=>"110100000",
  42865=>"110111001",
  42866=>"001100111",
  42867=>"010010111",
  42868=>"100010000",
  42869=>"011010100",
  42870=>"111010100",
  42871=>"010110011",
  42872=>"000110110",
  42873=>"111000111",
  42874=>"110010011",
  42875=>"000000001",
  42876=>"011110011",
  42877=>"010000100",
  42878=>"101011011",
  42879=>"110011100",
  42880=>"010101000",
  42881=>"100011100",
  42882=>"110001000",
  42883=>"100010110",
  42884=>"010001100",
  42885=>"001100001",
  42886=>"111000001",
  42887=>"111100011",
  42888=>"010101001",
  42889=>"100000001",
  42890=>"000010010",
  42891=>"100100010",
  42892=>"101100011",
  42893=>"011000001",
  42894=>"110100001",
  42895=>"000100001",
  42896=>"000110110",
  42897=>"110101101",
  42898=>"000101010",
  42899=>"000000110",
  42900=>"111101111",
  42901=>"111010111",
  42902=>"100100101",
  42903=>"000000010",
  42904=>"100101001",
  42905=>"100100001",
  42906=>"000011101",
  42907=>"100001011",
  42908=>"000010011",
  42909=>"000011100",
  42910=>"110001000",
  42911=>"011000000",
  42912=>"010000000",
  42913=>"010010100",
  42914=>"110110111",
  42915=>"100111110",
  42916=>"000000101",
  42917=>"001001011",
  42918=>"111101100",
  42919=>"101101001",
  42920=>"100011011",
  42921=>"110010100",
  42922=>"010111011",
  42923=>"111101100",
  42924=>"000111001",
  42925=>"011101111",
  42926=>"000011101",
  42927=>"100000000",
  42928=>"000111111",
  42929=>"111011111",
  42930=>"010000000",
  42931=>"010110011",
  42932=>"011000101",
  42933=>"111110111",
  42934=>"100011111",
  42935=>"101100000",
  42936=>"101011101",
  42937=>"001111100",
  42938=>"101101000",
  42939=>"110001111",
  42940=>"101000101",
  42941=>"110110100",
  42942=>"111100011",
  42943=>"100010001",
  42944=>"000111101",
  42945=>"100110011",
  42946=>"101010000",
  42947=>"110110011",
  42948=>"100111110",
  42949=>"000100100",
  42950=>"000001111",
  42951=>"101111100",
  42952=>"000100001",
  42953=>"011000001",
  42954=>"011111111",
  42955=>"001011011",
  42956=>"011101010",
  42957=>"111000111",
  42958=>"100001011",
  42959=>"000100110",
  42960=>"100100000",
  42961=>"001010000",
  42962=>"011110010",
  42963=>"010110100",
  42964=>"101110100",
  42965=>"110010011",
  42966=>"011110101",
  42967=>"110101101",
  42968=>"001001010",
  42969=>"101011100",
  42970=>"101100001",
  42971=>"100111111",
  42972=>"111000011",
  42973=>"110010111",
  42974=>"110110101",
  42975=>"100001011",
  42976=>"001011100",
  42977=>"011011100",
  42978=>"100111101",
  42979=>"100010100",
  42980=>"000000001",
  42981=>"010110000",
  42982=>"000111000",
  42983=>"001100011",
  42984=>"000010000",
  42985=>"011111001",
  42986=>"000111011",
  42987=>"101011110",
  42988=>"100011111",
  42989=>"111110000",
  42990=>"001010001",
  42991=>"111011111",
  42992=>"010101100",
  42993=>"001010000",
  42994=>"000100101",
  42995=>"001111100",
  42996=>"010110001",
  42997=>"000110010",
  42998=>"011000011",
  42999=>"101111011",
  43000=>"011100101",
  43001=>"010100000",
  43002=>"000001110",
  43003=>"111000011",
  43004=>"110101011",
  43005=>"100111111",
  43006=>"110010100",
  43007=>"010001000",
  43008=>"011000001",
  43009=>"101111010",
  43010=>"010101100",
  43011=>"110110111",
  43012=>"101101011",
  43013=>"111011011",
  43014=>"001110010",
  43015=>"100011001",
  43016=>"010111111",
  43017=>"000101100",
  43018=>"010101000",
  43019=>"001100101",
  43020=>"110011110",
  43021=>"000011111",
  43022=>"110000111",
  43023=>"011010110",
  43024=>"010001110",
  43025=>"111111111",
  43026=>"111100001",
  43027=>"001000111",
  43028=>"111100111",
  43029=>"111001111",
  43030=>"010100001",
  43031=>"000011110",
  43032=>"110101100",
  43033=>"001001011",
  43034=>"001110111",
  43035=>"111110100",
  43036=>"011110010",
  43037=>"110000010",
  43038=>"010011010",
  43039=>"000110011",
  43040=>"010011111",
  43041=>"101110111",
  43042=>"111100110",
  43043=>"111111111",
  43044=>"110000011",
  43045=>"001010010",
  43046=>"110101111",
  43047=>"111111000",
  43048=>"111010000",
  43049=>"110000001",
  43050=>"111100100",
  43051=>"101110100",
  43052=>"011000111",
  43053=>"011110110",
  43054=>"111101011",
  43055=>"011000111",
  43056=>"111011111",
  43057=>"000101010",
  43058=>"100111111",
  43059=>"000100000",
  43060=>"001100000",
  43061=>"000000101",
  43062=>"111111111",
  43063=>"101100101",
  43064=>"011110101",
  43065=>"011000111",
  43066=>"000101100",
  43067=>"010100111",
  43068=>"010001000",
  43069=>"011000010",
  43070=>"010111111",
  43071=>"111111101",
  43072=>"111111110",
  43073=>"011111000",
  43074=>"100101010",
  43075=>"111000001",
  43076=>"001001010",
  43077=>"110001001",
  43078=>"000010000",
  43079=>"000001001",
  43080=>"110101001",
  43081=>"011101011",
  43082=>"010110000",
  43083=>"101010110",
  43084=>"000100011",
  43085=>"000000010",
  43086=>"010100010",
  43087=>"001011000",
  43088=>"111011100",
  43089=>"111111011",
  43090=>"100011100",
  43091=>"100101101",
  43092=>"111010010",
  43093=>"011101100",
  43094=>"000110110",
  43095=>"101001000",
  43096=>"001001010",
  43097=>"011100011",
  43098=>"010001101",
  43099=>"111110000",
  43100=>"010010101",
  43101=>"000001010",
  43102=>"101100110",
  43103=>"100100011",
  43104=>"001101000",
  43105=>"001000110",
  43106=>"100110010",
  43107=>"001000101",
  43108=>"101000110",
  43109=>"100000000",
  43110=>"110100101",
  43111=>"000111010",
  43112=>"110010001",
  43113=>"100111000",
  43114=>"000100001",
  43115=>"111110110",
  43116=>"010001100",
  43117=>"111110010",
  43118=>"111011100",
  43119=>"000111001",
  43120=>"110001101",
  43121=>"101001010",
  43122=>"111110110",
  43123=>"110110111",
  43124=>"101000111",
  43125=>"110101100",
  43126=>"101101010",
  43127=>"111010001",
  43128=>"100010111",
  43129=>"010110110",
  43130=>"010001100",
  43131=>"111000001",
  43132=>"111000011",
  43133=>"100010110",
  43134=>"011110010",
  43135=>"011000001",
  43136=>"000000100",
  43137=>"100101011",
  43138=>"010110001",
  43139=>"101110001",
  43140=>"000110111",
  43141=>"101010100",
  43142=>"100011011",
  43143=>"111011011",
  43144=>"110101100",
  43145=>"111001111",
  43146=>"010000001",
  43147=>"011010100",
  43148=>"001101100",
  43149=>"101011100",
  43150=>"111001011",
  43151=>"001000110",
  43152=>"110100000",
  43153=>"000010111",
  43154=>"110010001",
  43155=>"011000111",
  43156=>"010010000",
  43157=>"000110111",
  43158=>"001111011",
  43159=>"101011000",
  43160=>"000001000",
  43161=>"010100111",
  43162=>"000010111",
  43163=>"001100010",
  43164=>"011101011",
  43165=>"010010000",
  43166=>"101101100",
  43167=>"110010110",
  43168=>"110001101",
  43169=>"001001000",
  43170=>"010111111",
  43171=>"011000100",
  43172=>"011110000",
  43173=>"100100111",
  43174=>"111110000",
  43175=>"001111001",
  43176=>"000101011",
  43177=>"011111000",
  43178=>"010111000",
  43179=>"000111001",
  43180=>"101111111",
  43181=>"101001000",
  43182=>"001110100",
  43183=>"011001100",
  43184=>"010010110",
  43185=>"000101000",
  43186=>"101111011",
  43187=>"000010111",
  43188=>"111001000",
  43189=>"011101101",
  43190=>"000000000",
  43191=>"111110001",
  43192=>"001000101",
  43193=>"010011100",
  43194=>"000000011",
  43195=>"110010101",
  43196=>"001010100",
  43197=>"111110010",
  43198=>"101011001",
  43199=>"100101010",
  43200=>"000100001",
  43201=>"001011001",
  43202=>"011011100",
  43203=>"001111110",
  43204=>"011001111",
  43205=>"000010000",
  43206=>"111001111",
  43207=>"110011100",
  43208=>"101100101",
  43209=>"000101111",
  43210=>"000010001",
  43211=>"010000110",
  43212=>"111100111",
  43213=>"110111100",
  43214=>"001000101",
  43215=>"100010010",
  43216=>"011010110",
  43217=>"110000111",
  43218=>"001011001",
  43219=>"110100111",
  43220=>"101101000",
  43221=>"010111011",
  43222=>"001111011",
  43223=>"001101101",
  43224=>"000000101",
  43225=>"010011011",
  43226=>"100101001",
  43227=>"011100011",
  43228=>"001010100",
  43229=>"001010001",
  43230=>"011011011",
  43231=>"010101001",
  43232=>"111101111",
  43233=>"111110100",
  43234=>"001001011",
  43235=>"100011010",
  43236=>"100100110",
  43237=>"000010111",
  43238=>"101001101",
  43239=>"110101101",
  43240=>"011000000",
  43241=>"101010110",
  43242=>"101010101",
  43243=>"100101001",
  43244=>"001000011",
  43245=>"000000100",
  43246=>"010101011",
  43247=>"000000101",
  43248=>"011111001",
  43249=>"100101100",
  43250=>"010000000",
  43251=>"001001000",
  43252=>"011001011",
  43253=>"010011000",
  43254=>"011000001",
  43255=>"111000100",
  43256=>"011010010",
  43257=>"000110001",
  43258=>"001111011",
  43259=>"010001001",
  43260=>"000111101",
  43261=>"111111001",
  43262=>"100110000",
  43263=>"111101001",
  43264=>"011010101",
  43265=>"110111100",
  43266=>"101001100",
  43267=>"100000000",
  43268=>"101100000",
  43269=>"111011110",
  43270=>"111111100",
  43271=>"011110000",
  43272=>"100100000",
  43273=>"010110111",
  43274=>"111101110",
  43275=>"100111111",
  43276=>"000110001",
  43277=>"000010100",
  43278=>"000100000",
  43279=>"101100101",
  43280=>"101011110",
  43281=>"111000010",
  43282=>"110111110",
  43283=>"100101111",
  43284=>"000001011",
  43285=>"001011101",
  43286=>"110111111",
  43287=>"010101110",
  43288=>"110000011",
  43289=>"110000011",
  43290=>"111111001",
  43291=>"000100101",
  43292=>"100000100",
  43293=>"110011011",
  43294=>"011011101",
  43295=>"110001010",
  43296=>"100000110",
  43297=>"110011001",
  43298=>"010101010",
  43299=>"000001111",
  43300=>"100100110",
  43301=>"010011010",
  43302=>"000101111",
  43303=>"000011111",
  43304=>"010000110",
  43305=>"101110010",
  43306=>"101100010",
  43307=>"111111001",
  43308=>"010101100",
  43309=>"111001000",
  43310=>"000011010",
  43311=>"011110100",
  43312=>"010110010",
  43313=>"010110110",
  43314=>"000101000",
  43315=>"010110001",
  43316=>"110111001",
  43317=>"100110110",
  43318=>"101010110",
  43319=>"001011111",
  43320=>"011100001",
  43321=>"000100110",
  43322=>"111000101",
  43323=>"000110111",
  43324=>"110001001",
  43325=>"011101001",
  43326=>"100001100",
  43327=>"100100110",
  43328=>"111101011",
  43329=>"100111100",
  43330=>"011111011",
  43331=>"011110100",
  43332=>"010011111",
  43333=>"010100000",
  43334=>"001110000",
  43335=>"001101110",
  43336=>"001111001",
  43337=>"000100100",
  43338=>"010101110",
  43339=>"010110001",
  43340=>"010001011",
  43341=>"010001011",
  43342=>"011100110",
  43343=>"100100110",
  43344=>"011001011",
  43345=>"001100010",
  43346=>"100101000",
  43347=>"111000011",
  43348=>"010101111",
  43349=>"001100001",
  43350=>"000000111",
  43351=>"100111001",
  43352=>"000000110",
  43353=>"000100100",
  43354=>"010010101",
  43355=>"001011110",
  43356=>"100000100",
  43357=>"001110110",
  43358=>"010101100",
  43359=>"111110110",
  43360=>"001010001",
  43361=>"111000110",
  43362=>"111100000",
  43363=>"000000000",
  43364=>"100000010",
  43365=>"001000001",
  43366=>"001101100",
  43367=>"011010100",
  43368=>"100101100",
  43369=>"000001111",
  43370=>"101111010",
  43371=>"000010001",
  43372=>"000000000",
  43373=>"110111000",
  43374=>"010111011",
  43375=>"100100111",
  43376=>"100011010",
  43377=>"110111001",
  43378=>"111001011",
  43379=>"100101100",
  43380=>"101111111",
  43381=>"100011101",
  43382=>"010101011",
  43383=>"001000011",
  43384=>"101001101",
  43385=>"001001101",
  43386=>"111000101",
  43387=>"000111011",
  43388=>"000111100",
  43389=>"010101110",
  43390=>"001011111",
  43391=>"010000010",
  43392=>"000010110",
  43393=>"100101011",
  43394=>"000110111",
  43395=>"010101101",
  43396=>"000110111",
  43397=>"100000100",
  43398=>"011101011",
  43399=>"110010000",
  43400=>"111001010",
  43401=>"110010011",
  43402=>"100100111",
  43403=>"000011011",
  43404=>"001011101",
  43405=>"100010100",
  43406=>"111111000",
  43407=>"100000110",
  43408=>"000000010",
  43409=>"111100000",
  43410=>"000111101",
  43411=>"101110110",
  43412=>"001110011",
  43413=>"101011001",
  43414=>"100110011",
  43415=>"011111101",
  43416=>"010111111",
  43417=>"001001111",
  43418=>"100111101",
  43419=>"100001100",
  43420=>"110010100",
  43421=>"010010011",
  43422=>"000011001",
  43423=>"111001110",
  43424=>"101010000",
  43425=>"000000100",
  43426=>"010110111",
  43427=>"000001000",
  43428=>"001011100",
  43429=>"110000010",
  43430=>"010101111",
  43431=>"000101110",
  43432=>"100101101",
  43433=>"100010000",
  43434=>"001000010",
  43435=>"101011111",
  43436=>"110100010",
  43437=>"111011101",
  43438=>"101000100",
  43439=>"100110111",
  43440=>"001010110",
  43441=>"110111001",
  43442=>"100111010",
  43443=>"110111001",
  43444=>"010010000",
  43445=>"010111010",
  43446=>"010101110",
  43447=>"110010001",
  43448=>"000001100",
  43449=>"011010000",
  43450=>"010001101",
  43451=>"011100010",
  43452=>"000011001",
  43453=>"110000010",
  43454=>"100000000",
  43455=>"011110111",
  43456=>"101011101",
  43457=>"110001010",
  43458=>"001100011",
  43459=>"010001011",
  43460=>"111110111",
  43461=>"001001000",
  43462=>"010101000",
  43463=>"100110110",
  43464=>"110101111",
  43465=>"110110010",
  43466=>"011010001",
  43467=>"010010100",
  43468=>"010001101",
  43469=>"000000011",
  43470=>"101100101",
  43471=>"010001110",
  43472=>"010011100",
  43473=>"101001000",
  43474=>"010000111",
  43475=>"010100111",
  43476=>"001100111",
  43477=>"111001111",
  43478=>"000110000",
  43479=>"011000010",
  43480=>"001010001",
  43481=>"101101111",
  43482=>"000000000",
  43483=>"010000001",
  43484=>"110010100",
  43485=>"010010111",
  43486=>"110100110",
  43487=>"001011000",
  43488=>"010011010",
  43489=>"101011110",
  43490=>"110010111",
  43491=>"000001010",
  43492=>"100000010",
  43493=>"111011010",
  43494=>"010000011",
  43495=>"111010101",
  43496=>"000100001",
  43497=>"101001011",
  43498=>"101001101",
  43499=>"011111001",
  43500=>"100000001",
  43501=>"101101111",
  43502=>"000101000",
  43503=>"000011001",
  43504=>"110100000",
  43505=>"011011000",
  43506=>"000101010",
  43507=>"101110011",
  43508=>"000111011",
  43509=>"000000100",
  43510=>"100001110",
  43511=>"000000010",
  43512=>"011010001",
  43513=>"001011001",
  43514=>"111001000",
  43515=>"001101101",
  43516=>"111000101",
  43517=>"111111010",
  43518=>"000001001",
  43519=>"111011101",
  43520=>"101110100",
  43521=>"010111100",
  43522=>"000110111",
  43523=>"110010011",
  43524=>"000100010",
  43525=>"110010010",
  43526=>"010000001",
  43527=>"110110111",
  43528=>"011010010",
  43529=>"001011011",
  43530=>"010001110",
  43531=>"101111111",
  43532=>"011111110",
  43533=>"101101110",
  43534=>"001101000",
  43535=>"001110010",
  43536=>"000000011",
  43537=>"110011001",
  43538=>"011111010",
  43539=>"000100000",
  43540=>"001100010",
  43541=>"110101011",
  43542=>"100111111",
  43543=>"010011010",
  43544=>"111111001",
  43545=>"000100000",
  43546=>"101110100",
  43547=>"111101100",
  43548=>"100000000",
  43549=>"001100101",
  43550=>"001010010",
  43551=>"101011110",
  43552=>"111001001",
  43553=>"011111111",
  43554=>"111111111",
  43555=>"000001100",
  43556=>"110011110",
  43557=>"010000001",
  43558=>"001110011",
  43559=>"110000000",
  43560=>"101001011",
  43561=>"010010111",
  43562=>"011100110",
  43563=>"011101111",
  43564=>"011100100",
  43565=>"100000001",
  43566=>"100111100",
  43567=>"011010110",
  43568=>"011010101",
  43569=>"100100101",
  43570=>"110101101",
  43571=>"100011010",
  43572=>"100001011",
  43573=>"010001100",
  43574=>"111011100",
  43575=>"001110101",
  43576=>"000010101",
  43577=>"111110011",
  43578=>"011110000",
  43579=>"000001011",
  43580=>"110011100",
  43581=>"111111000",
  43582=>"001011000",
  43583=>"010101010",
  43584=>"101010101",
  43585=>"001100110",
  43586=>"010111110",
  43587=>"110011100",
  43588=>"110101110",
  43589=>"001000110",
  43590=>"000011001",
  43591=>"111111011",
  43592=>"011011000",
  43593=>"111101011",
  43594=>"001111110",
  43595=>"100001001",
  43596=>"001001110",
  43597=>"100100110",
  43598=>"111001010",
  43599=>"100001000",
  43600=>"001001011",
  43601=>"111100101",
  43602=>"001001111",
  43603=>"000000010",
  43604=>"000000100",
  43605=>"011100101",
  43606=>"101110110",
  43607=>"000001100",
  43608=>"100001001",
  43609=>"110000010",
  43610=>"010111000",
  43611=>"111110001",
  43612=>"101011110",
  43613=>"110101010",
  43614=>"011111110",
  43615=>"010111110",
  43616=>"000100100",
  43617=>"100111111",
  43618=>"001001110",
  43619=>"100111100",
  43620=>"110100100",
  43621=>"111111110",
  43622=>"000010100",
  43623=>"000010110",
  43624=>"011011101",
  43625=>"111100111",
  43626=>"111110100",
  43627=>"001100010",
  43628=>"000010010",
  43629=>"111100110",
  43630=>"110110011",
  43631=>"110111001",
  43632=>"110111101",
  43633=>"000010111",
  43634=>"000110000",
  43635=>"111010000",
  43636=>"000000110",
  43637=>"100100101",
  43638=>"001010101",
  43639=>"000011110",
  43640=>"001100110",
  43641=>"111111111",
  43642=>"011001110",
  43643=>"111101011",
  43644=>"001100001",
  43645=>"011101100",
  43646=>"010101110",
  43647=>"111100010",
  43648=>"100001001",
  43649=>"100111000",
  43650=>"001101011",
  43651=>"101010011",
  43652=>"100110100",
  43653=>"100111111",
  43654=>"011011111",
  43655=>"011111000",
  43656=>"000101001",
  43657=>"110100000",
  43658=>"000001000",
  43659=>"011111010",
  43660=>"010101001",
  43661=>"000111111",
  43662=>"100111000",
  43663=>"000001000",
  43664=>"000110011",
  43665=>"100010101",
  43666=>"111010110",
  43667=>"101001001",
  43668=>"101000000",
  43669=>"101100100",
  43670=>"111100010",
  43671=>"000110101",
  43672=>"111011000",
  43673=>"010111000",
  43674=>"110100010",
  43675=>"110111011",
  43676=>"000010001",
  43677=>"010010110",
  43678=>"100001010",
  43679=>"010010000",
  43680=>"010100010",
  43681=>"001000100",
  43682=>"011110110",
  43683=>"001001101",
  43684=>"001001101",
  43685=>"101000100",
  43686=>"000100000",
  43687=>"101001100",
  43688=>"111011011",
  43689=>"111011000",
  43690=>"111111101",
  43691=>"000010111",
  43692=>"100111110",
  43693=>"111101000",
  43694=>"010000001",
  43695=>"001011010",
  43696=>"110111100",
  43697=>"010100101",
  43698=>"111100000",
  43699=>"011000000",
  43700=>"011101011",
  43701=>"111111111",
  43702=>"111101111",
  43703=>"011001000",
  43704=>"100101111",
  43705=>"000100110",
  43706=>"011011101",
  43707=>"101100011",
  43708=>"111110111",
  43709=>"000100001",
  43710=>"101010011",
  43711=>"100010001",
  43712=>"000110101",
  43713=>"011110110",
  43714=>"111101111",
  43715=>"110000100",
  43716=>"011110100",
  43717=>"101101110",
  43718=>"111111001",
  43719=>"100111001",
  43720=>"000110010",
  43721=>"011001111",
  43722=>"000110001",
  43723=>"000110110",
  43724=>"001000001",
  43725=>"101111110",
  43726=>"010001011",
  43727=>"111111111",
  43728=>"000001110",
  43729=>"110100010",
  43730=>"011110111",
  43731=>"111110001",
  43732=>"110000010",
  43733=>"001001000",
  43734=>"111010000",
  43735=>"000011010",
  43736=>"101101100",
  43737=>"010111011",
  43738=>"001011101",
  43739=>"001111010",
  43740=>"000110100",
  43741=>"110111100",
  43742=>"011001111",
  43743=>"000011000",
  43744=>"000010010",
  43745=>"100010110",
  43746=>"010000111",
  43747=>"010111010",
  43748=>"110101001",
  43749=>"011101111",
  43750=>"010010000",
  43751=>"111110011",
  43752=>"011000101",
  43753=>"001100011",
  43754=>"100001000",
  43755=>"100111000",
  43756=>"100110011",
  43757=>"100011101",
  43758=>"011110101",
  43759=>"000100001",
  43760=>"110001110",
  43761=>"010101111",
  43762=>"110001000",
  43763=>"010001111",
  43764=>"100100110",
  43765=>"110001101",
  43766=>"100110100",
  43767=>"101011111",
  43768=>"111010011",
  43769=>"010110111",
  43770=>"011110110",
  43771=>"011000011",
  43772=>"111011011",
  43773=>"110000010",
  43774=>"001010001",
  43775=>"101010001",
  43776=>"110101111",
  43777=>"001010110",
  43778=>"110010100",
  43779=>"000000011",
  43780=>"101100100",
  43781=>"001001011",
  43782=>"000011100",
  43783=>"100100000",
  43784=>"011001100",
  43785=>"101101011",
  43786=>"111001010",
  43787=>"110100010",
  43788=>"010001101",
  43789=>"101001001",
  43790=>"011011011",
  43791=>"000000110",
  43792=>"101100010",
  43793=>"111110000",
  43794=>"010010000",
  43795=>"111000100",
  43796=>"100001101",
  43797=>"011110100",
  43798=>"110000001",
  43799=>"101010001",
  43800=>"011111111",
  43801=>"011000111",
  43802=>"111101011",
  43803=>"111001001",
  43804=>"111000111",
  43805=>"101010010",
  43806=>"111001001",
  43807=>"010100100",
  43808=>"100010000",
  43809=>"101100011",
  43810=>"000001000",
  43811=>"011011001",
  43812=>"011101000",
  43813=>"111000011",
  43814=>"000001011",
  43815=>"110100001",
  43816=>"001000101",
  43817=>"000010000",
  43818=>"001101000",
  43819=>"000001110",
  43820=>"100110100",
  43821=>"000001011",
  43822=>"110111100",
  43823=>"101101000",
  43824=>"011001111",
  43825=>"000100011",
  43826=>"000010011",
  43827=>"111010110",
  43828=>"110110110",
  43829=>"010100000",
  43830=>"101000110",
  43831=>"011100110",
  43832=>"111010011",
  43833=>"111100101",
  43834=>"000000000",
  43835=>"110111111",
  43836=>"110111101",
  43837=>"100100001",
  43838=>"011101111",
  43839=>"101000111",
  43840=>"110110100",
  43841=>"001110000",
  43842=>"110000001",
  43843=>"111100101",
  43844=>"010011110",
  43845=>"110011111",
  43846=>"010110111",
  43847=>"101111111",
  43848=>"110110100",
  43849=>"000001101",
  43850=>"000011110",
  43851=>"010010011",
  43852=>"001000000",
  43853=>"101101101",
  43854=>"100010111",
  43855=>"110101111",
  43856=>"001000100",
  43857=>"101011100",
  43858=>"110010001",
  43859=>"001001111",
  43860=>"010101111",
  43861=>"111001100",
  43862=>"110011000",
  43863=>"111100001",
  43864=>"000111101",
  43865=>"011011100",
  43866=>"001001000",
  43867=>"110111101",
  43868=>"110011100",
  43869=>"110101100",
  43870=>"010101111",
  43871=>"010001001",
  43872=>"001111011",
  43873=>"010001011",
  43874=>"001001111",
  43875=>"111010010",
  43876=>"110011111",
  43877=>"000111100",
  43878=>"011101111",
  43879=>"110000001",
  43880=>"111000101",
  43881=>"110111000",
  43882=>"010011110",
  43883=>"010000010",
  43884=>"011000001",
  43885=>"010100101",
  43886=>"111111111",
  43887=>"011100001",
  43888=>"111110100",
  43889=>"000110010",
  43890=>"101101111",
  43891=>"101010000",
  43892=>"001111001",
  43893=>"011010000",
  43894=>"101100000",
  43895=>"101110001",
  43896=>"110010001",
  43897=>"010011001",
  43898=>"010101001",
  43899=>"011101011",
  43900=>"011010001",
  43901=>"000111000",
  43902=>"100001000",
  43903=>"101011000",
  43904=>"010011110",
  43905=>"011000011",
  43906=>"000100010",
  43907=>"110000111",
  43908=>"001110001",
  43909=>"111101110",
  43910=>"001100001",
  43911=>"000010111",
  43912=>"011101101",
  43913=>"110110011",
  43914=>"110111100",
  43915=>"110110011",
  43916=>"001111011",
  43917=>"110101101",
  43918=>"001000010",
  43919=>"001001001",
  43920=>"110111111",
  43921=>"111010000",
  43922=>"101111110",
  43923=>"110011001",
  43924=>"001110101",
  43925=>"010000101",
  43926=>"111010000",
  43927=>"110100010",
  43928=>"010010000",
  43929=>"101110101",
  43930=>"110111101",
  43931=>"001111001",
  43932=>"011001111",
  43933=>"011010001",
  43934=>"001100010",
  43935=>"010010100",
  43936=>"101100110",
  43937=>"110110011",
  43938=>"100011011",
  43939=>"110100100",
  43940=>"001011111",
  43941=>"110111010",
  43942=>"110110011",
  43943=>"100010000",
  43944=>"111001111",
  43945=>"111110000",
  43946=>"110011010",
  43947=>"010010000",
  43948=>"011011010",
  43949=>"010100101",
  43950=>"010110100",
  43951=>"111110111",
  43952=>"010100011",
  43953=>"111010011",
  43954=>"101010011",
  43955=>"011100001",
  43956=>"100011110",
  43957=>"000101111",
  43958=>"011010110",
  43959=>"001110000",
  43960=>"001100011",
  43961=>"010110111",
  43962=>"001101101",
  43963=>"111011001",
  43964=>"111010101",
  43965=>"101001000",
  43966=>"011110101",
  43967=>"100001110",
  43968=>"001110001",
  43969=>"001101001",
  43970=>"110100111",
  43971=>"000110010",
  43972=>"100001000",
  43973=>"010000011",
  43974=>"000010000",
  43975=>"001001100",
  43976=>"010100101",
  43977=>"110100101",
  43978=>"100110110",
  43979=>"000010100",
  43980=>"011111111",
  43981=>"110111111",
  43982=>"100111010",
  43983=>"110100101",
  43984=>"010000001",
  43985=>"001100101",
  43986=>"011000000",
  43987=>"111110110",
  43988=>"000000101",
  43989=>"101000110",
  43990=>"000110000",
  43991=>"111000011",
  43992=>"001101010",
  43993=>"110110110",
  43994=>"111011111",
  43995=>"111000010",
  43996=>"000110110",
  43997=>"010000101",
  43998=>"010101001",
  43999=>"111010010",
  44000=>"001010011",
  44001=>"001111010",
  44002=>"100111001",
  44003=>"100111111",
  44004=>"100011000",
  44005=>"000100100",
  44006=>"111000000",
  44007=>"010110011",
  44008=>"100000001",
  44009=>"110001000",
  44010=>"110001000",
  44011=>"101000001",
  44012=>"111110111",
  44013=>"010100101",
  44014=>"111100100",
  44015=>"001000010",
  44016=>"000000111",
  44017=>"001110101",
  44018=>"101000100",
  44019=>"000001111",
  44020=>"011010010",
  44021=>"000001100",
  44022=>"000100010",
  44023=>"111111010",
  44024=>"110111010",
  44025=>"111001110",
  44026=>"001011010",
  44027=>"000010100",
  44028=>"100001011",
  44029=>"101011101",
  44030=>"011111100",
  44031=>"011011000",
  44032=>"001110000",
  44033=>"000011111",
  44034=>"011101010",
  44035=>"100111100",
  44036=>"101111011",
  44037=>"011110100",
  44038=>"001101001",
  44039=>"101000100",
  44040=>"101110010",
  44041=>"011110111",
  44042=>"110010110",
  44043=>"000001111",
  44044=>"010111000",
  44045=>"010101100",
  44046=>"111000100",
  44047=>"001100111",
  44048=>"111010011",
  44049=>"001001011",
  44050=>"111001011",
  44051=>"111111111",
  44052=>"001000000",
  44053=>"111001100",
  44054=>"111111010",
  44055=>"101101111",
  44056=>"010001011",
  44057=>"000010001",
  44058=>"110000101",
  44059=>"110110100",
  44060=>"110101101",
  44061=>"101101111",
  44062=>"001110000",
  44063=>"001101111",
  44064=>"001100101",
  44065=>"011100000",
  44066=>"111010010",
  44067=>"100011111",
  44068=>"111101110",
  44069=>"101110101",
  44070=>"100011011",
  44071=>"100110100",
  44072=>"011110110",
  44073=>"100100000",
  44074=>"111101001",
  44075=>"010010001",
  44076=>"010110100",
  44077=>"001010001",
  44078=>"001001010",
  44079=>"001101010",
  44080=>"011110111",
  44081=>"101111000",
  44082=>"011100000",
  44083=>"001110111",
  44084=>"001111011",
  44085=>"001011001",
  44086=>"011111000",
  44087=>"101000010",
  44088=>"001001110",
  44089=>"011100100",
  44090=>"110001011",
  44091=>"011011100",
  44092=>"110011111",
  44093=>"110101110",
  44094=>"000111101",
  44095=>"010011111",
  44096=>"011010001",
  44097=>"100101011",
  44098=>"101101100",
  44099=>"000011111",
  44100=>"010000000",
  44101=>"000010111",
  44102=>"101101110",
  44103=>"110111101",
  44104=>"001111111",
  44105=>"011101100",
  44106=>"111111000",
  44107=>"001110101",
  44108=>"111101010",
  44109=>"100010011",
  44110=>"100001101",
  44111=>"111111111",
  44112=>"111111111",
  44113=>"111101001",
  44114=>"001111010",
  44115=>"011100111",
  44116=>"010000101",
  44117=>"100110110",
  44118=>"001101001",
  44119=>"111000111",
  44120=>"100001110",
  44121=>"101110101",
  44122=>"001010100",
  44123=>"011110000",
  44124=>"011000001",
  44125=>"011000100",
  44126=>"010000011",
  44127=>"010111110",
  44128=>"110010010",
  44129=>"001011100",
  44130=>"011001010",
  44131=>"111101010",
  44132=>"001010001",
  44133=>"001000001",
  44134=>"011010100",
  44135=>"010110011",
  44136=>"010011100",
  44137=>"111110000",
  44138=>"000000110",
  44139=>"110100110",
  44140=>"000110000",
  44141=>"110100011",
  44142=>"111111001",
  44143=>"010000110",
  44144=>"101000010",
  44145=>"000011111",
  44146=>"010110100",
  44147=>"110110110",
  44148=>"010100110",
  44149=>"101111100",
  44150=>"100100001",
  44151=>"111111010",
  44152=>"001100111",
  44153=>"000111011",
  44154=>"111111101",
  44155=>"100110011",
  44156=>"000010001",
  44157=>"001011000",
  44158=>"000000000",
  44159=>"100101001",
  44160=>"011010000",
  44161=>"110001100",
  44162=>"110001011",
  44163=>"000011000",
  44164=>"101001101",
  44165=>"010011111",
  44166=>"011100111",
  44167=>"101000110",
  44168=>"000010011",
  44169=>"000100100",
  44170=>"100100000",
  44171=>"111101010",
  44172=>"100100101",
  44173=>"010110100",
  44174=>"001011000",
  44175=>"010000111",
  44176=>"111111110",
  44177=>"011110101",
  44178=>"011010100",
  44179=>"010011101",
  44180=>"001101101",
  44181=>"110011111",
  44182=>"111001000",
  44183=>"001101000",
  44184=>"110101111",
  44185=>"011111111",
  44186=>"011110011",
  44187=>"011011101",
  44188=>"011100011",
  44189=>"000011011",
  44190=>"001100111",
  44191=>"000001000",
  44192=>"000101001",
  44193=>"010110111",
  44194=>"000001111",
  44195=>"000111110",
  44196=>"011110110",
  44197=>"000001110",
  44198=>"001010010",
  44199=>"101001001",
  44200=>"100011011",
  44201=>"101111111",
  44202=>"010001010",
  44203=>"100111010",
  44204=>"111101100",
  44205=>"110010111",
  44206=>"001101010",
  44207=>"110111010",
  44208=>"001100111",
  44209=>"111001101",
  44210=>"110100101",
  44211=>"100011000",
  44212=>"000001111",
  44213=>"000000100",
  44214=>"011011101",
  44215=>"000110111",
  44216=>"110101011",
  44217=>"011111000",
  44218=>"111111100",
  44219=>"001111100",
  44220=>"111011000",
  44221=>"101000111",
  44222=>"111111110",
  44223=>"001010001",
  44224=>"100000101",
  44225=>"000101001",
  44226=>"010111001",
  44227=>"100110100",
  44228=>"101101000",
  44229=>"000110000",
  44230=>"010000000",
  44231=>"010011011",
  44232=>"111010111",
  44233=>"000101101",
  44234=>"000101001",
  44235=>"001100100",
  44236=>"001001010",
  44237=>"000110000",
  44238=>"010111011",
  44239=>"111110000",
  44240=>"111110010",
  44241=>"101000010",
  44242=>"101110011",
  44243=>"001010000",
  44244=>"110110010",
  44245=>"000100110",
  44246=>"010111101",
  44247=>"100111100",
  44248=>"100010011",
  44249=>"101001011",
  44250=>"101110011",
  44251=>"110010010",
  44252=>"100010000",
  44253=>"100111011",
  44254=>"010010001",
  44255=>"111001001",
  44256=>"001000011",
  44257=>"101011110",
  44258=>"110101000",
  44259=>"111110001",
  44260=>"001001001",
  44261=>"110010000",
  44262=>"011000000",
  44263=>"011000100",
  44264=>"100001000",
  44265=>"011111101",
  44266=>"000000010",
  44267=>"000001110",
  44268=>"010101010",
  44269=>"011011000",
  44270=>"000111010",
  44271=>"001000001",
  44272=>"101010111",
  44273=>"101010000",
  44274=>"000100000",
  44275=>"110110011",
  44276=>"011111100",
  44277=>"000101110",
  44278=>"101100111",
  44279=>"010000110",
  44280=>"110111011",
  44281=>"101101010",
  44282=>"011111011",
  44283=>"111101011",
  44284=>"110000001",
  44285=>"100110110",
  44286=>"100011111",
  44287=>"111110111",
  44288=>"011110010",
  44289=>"100010000",
  44290=>"101101010",
  44291=>"000010110",
  44292=>"001110110",
  44293=>"000001010",
  44294=>"101110001",
  44295=>"000010010",
  44296=>"010010110",
  44297=>"010011110",
  44298=>"111000110",
  44299=>"010000100",
  44300=>"101101000",
  44301=>"101111001",
  44302=>"110000010",
  44303=>"111101110",
  44304=>"100101110",
  44305=>"111001111",
  44306=>"100001101",
  44307=>"101100010",
  44308=>"110001100",
  44309=>"000110001",
  44310=>"110100100",
  44311=>"000000000",
  44312=>"010000110",
  44313=>"100100111",
  44314=>"111010100",
  44315=>"101010011",
  44316=>"111111001",
  44317=>"011111000",
  44318=>"111010101",
  44319=>"001001010",
  44320=>"010100011",
  44321=>"001101101",
  44322=>"101110001",
  44323=>"010010001",
  44324=>"000001011",
  44325=>"001100101",
  44326=>"010111000",
  44327=>"101011000",
  44328=>"001100101",
  44329=>"110011101",
  44330=>"001100100",
  44331=>"010010001",
  44332=>"011100110",
  44333=>"100111101",
  44334=>"111101110",
  44335=>"011110010",
  44336=>"110110011",
  44337=>"100110111",
  44338=>"010011101",
  44339=>"111001000",
  44340=>"101110101",
  44341=>"011110100",
  44342=>"111000011",
  44343=>"101011001",
  44344=>"000000010",
  44345=>"000111000",
  44346=>"111111111",
  44347=>"100000111",
  44348=>"110101111",
  44349=>"100111110",
  44350=>"110100111",
  44351=>"111110110",
  44352=>"100110110",
  44353=>"111011100",
  44354=>"100000110",
  44355=>"111010000",
  44356=>"100101110",
  44357=>"000111101",
  44358=>"100000001",
  44359=>"000101010",
  44360=>"111011000",
  44361=>"111010000",
  44362=>"101111010",
  44363=>"111110000",
  44364=>"110000000",
  44365=>"010010100",
  44366=>"100101111",
  44367=>"101000011",
  44368=>"001111100",
  44369=>"011011001",
  44370=>"001101100",
  44371=>"101110110",
  44372=>"000001110",
  44373=>"101111011",
  44374=>"000000110",
  44375=>"001010011",
  44376=>"010110011",
  44377=>"000000000",
  44378=>"100000001",
  44379=>"001101110",
  44380=>"001110010",
  44381=>"001100100",
  44382=>"011111110",
  44383=>"100111100",
  44384=>"110001111",
  44385=>"110111011",
  44386=>"000101100",
  44387=>"001101001",
  44388=>"110010100",
  44389=>"101000110",
  44390=>"000110111",
  44391=>"011101100",
  44392=>"110110101",
  44393=>"110111111",
  44394=>"110011010",
  44395=>"000101100",
  44396=>"111010011",
  44397=>"011111101",
  44398=>"111000100",
  44399=>"010110101",
  44400=>"010110000",
  44401=>"001100111",
  44402=>"101111000",
  44403=>"101010101",
  44404=>"000000001",
  44405=>"001010111",
  44406=>"000111110",
  44407=>"110111100",
  44408=>"101111011",
  44409=>"011011010",
  44410=>"100110001",
  44411=>"100011100",
  44412=>"101100000",
  44413=>"000100000",
  44414=>"010010010",
  44415=>"110100101",
  44416=>"001011110",
  44417=>"111100001",
  44418=>"001110111",
  44419=>"101000010",
  44420=>"101001101",
  44421=>"001110100",
  44422=>"111011001",
  44423=>"111111011",
  44424=>"001100101",
  44425=>"010010111",
  44426=>"100111110",
  44427=>"001000000",
  44428=>"101111110",
  44429=>"000110011",
  44430=>"010001011",
  44431=>"000011001",
  44432=>"111101111",
  44433=>"000010010",
  44434=>"011000001",
  44435=>"101101010",
  44436=>"011100011",
  44437=>"001101001",
  44438=>"110111011",
  44439=>"111010110",
  44440=>"011000111",
  44441=>"101011110",
  44442=>"001000100",
  44443=>"100000010",
  44444=>"011101111",
  44445=>"100011111",
  44446=>"001101000",
  44447=>"001010000",
  44448=>"011110011",
  44449=>"110001000",
  44450=>"000011001",
  44451=>"011111110",
  44452=>"110111000",
  44453=>"011010101",
  44454=>"100111100",
  44455=>"001101010",
  44456=>"101101101",
  44457=>"111111111",
  44458=>"010100000",
  44459=>"110000101",
  44460=>"110010101",
  44461=>"111001011",
  44462=>"000100001",
  44463=>"111001011",
  44464=>"000100100",
  44465=>"001011011",
  44466=>"000110101",
  44467=>"000010110",
  44468=>"100000000",
  44469=>"001110011",
  44470=>"000101111",
  44471=>"000100011",
  44472=>"110111110",
  44473=>"110101110",
  44474=>"111000011",
  44475=>"110111010",
  44476=>"111101011",
  44477=>"111000110",
  44478=>"010011001",
  44479=>"000010001",
  44480=>"111010010",
  44481=>"011101000",
  44482=>"000000010",
  44483=>"101101010",
  44484=>"110101001",
  44485=>"000001100",
  44486=>"110011111",
  44487=>"000010001",
  44488=>"011000000",
  44489=>"111010011",
  44490=>"101001101",
  44491=>"010110100",
  44492=>"101000101",
  44493=>"001110111",
  44494=>"000001001",
  44495=>"111110011",
  44496=>"010110000",
  44497=>"100111110",
  44498=>"101111000",
  44499=>"101000001",
  44500=>"100100011",
  44501=>"010101000",
  44502=>"111101111",
  44503=>"000111111",
  44504=>"011010101",
  44505=>"111100101",
  44506=>"111101000",
  44507=>"000110111",
  44508=>"101110000",
  44509=>"100110000",
  44510=>"100101000",
  44511=>"011110101",
  44512=>"110110110",
  44513=>"001001111",
  44514=>"001011000",
  44515=>"001111100",
  44516=>"010011101",
  44517=>"111011000",
  44518=>"001100101",
  44519=>"001100011",
  44520=>"111101010",
  44521=>"010110111",
  44522=>"111110011",
  44523=>"010001010",
  44524=>"001100000",
  44525=>"100010010",
  44526=>"011111011",
  44527=>"111001100",
  44528=>"000101110",
  44529=>"100111100",
  44530=>"001100011",
  44531=>"110111001",
  44532=>"101001010",
  44533=>"111000101",
  44534=>"110011100",
  44535=>"001011110",
  44536=>"110011100",
  44537=>"000100010",
  44538=>"111111111",
  44539=>"011010110",
  44540=>"111111110",
  44541=>"010111010",
  44542=>"100100011",
  44543=>"101010110",
  44544=>"011001010",
  44545=>"111001100",
  44546=>"101110000",
  44547=>"111111101",
  44548=>"010101010",
  44549=>"100001010",
  44550=>"001100000",
  44551=>"010101010",
  44552=>"111010010",
  44553=>"110000001",
  44554=>"111111111",
  44555=>"110110111",
  44556=>"101101000",
  44557=>"010010000",
  44558=>"101011100",
  44559=>"010011111",
  44560=>"111101010",
  44561=>"011101011",
  44562=>"100001111",
  44563=>"000001010",
  44564=>"101011111",
  44565=>"101000011",
  44566=>"000111101",
  44567=>"101111100",
  44568=>"010100100",
  44569=>"110101010",
  44570=>"111101100",
  44571=>"010110111",
  44572=>"110111111",
  44573=>"011110001",
  44574=>"111101111",
  44575=>"100001011",
  44576=>"001001111",
  44577=>"011101101",
  44578=>"010001110",
  44579=>"011000000",
  44580=>"100000101",
  44581=>"010000111",
  44582=>"100110101",
  44583=>"111000111",
  44584=>"101111101",
  44585=>"000011111",
  44586=>"010101010",
  44587=>"011111001",
  44588=>"110100100",
  44589=>"110111111",
  44590=>"010000001",
  44591=>"100001000",
  44592=>"100010011",
  44593=>"110100000",
  44594=>"001011000",
  44595=>"011001101",
  44596=>"111100000",
  44597=>"000011111",
  44598=>"101010001",
  44599=>"100111011",
  44600=>"011010101",
  44601=>"111010101",
  44602=>"001000011",
  44603=>"111101110",
  44604=>"101010000",
  44605=>"010001100",
  44606=>"110100100",
  44607=>"010111001",
  44608=>"101111011",
  44609=>"111010110",
  44610=>"100010001",
  44611=>"101000011",
  44612=>"000110101",
  44613=>"000101100",
  44614=>"000001101",
  44615=>"001011001",
  44616=>"101000100",
  44617=>"111100011",
  44618=>"011010011",
  44619=>"010000110",
  44620=>"010101100",
  44621=>"100110000",
  44622=>"100101011",
  44623=>"001100000",
  44624=>"101000000",
  44625=>"000011010",
  44626=>"011010110",
  44627=>"011110000",
  44628=>"110000000",
  44629=>"100010010",
  44630=>"010111111",
  44631=>"001011011",
  44632=>"110111011",
  44633=>"111100100",
  44634=>"011010000",
  44635=>"011010001",
  44636=>"010100010",
  44637=>"000000011",
  44638=>"000100001",
  44639=>"110011101",
  44640=>"100011000",
  44641=>"000010100",
  44642=>"011101010",
  44643=>"000101001",
  44644=>"111001001",
  44645=>"000100100",
  44646=>"000000001",
  44647=>"010111011",
  44648=>"010000000",
  44649=>"111100111",
  44650=>"101001010",
  44651=>"000100000",
  44652=>"111000111",
  44653=>"111001011",
  44654=>"101001010",
  44655=>"001110010",
  44656=>"000001111",
  44657=>"110010010",
  44658=>"100010101",
  44659=>"100111101",
  44660=>"110100110",
  44661=>"010010111",
  44662=>"100111101",
  44663=>"010000001",
  44664=>"101001010",
  44665=>"000010000",
  44666=>"100010111",
  44667=>"001001000",
  44668=>"101010100",
  44669=>"011011110",
  44670=>"110000111",
  44671=>"111010000",
  44672=>"010111001",
  44673=>"111000001",
  44674=>"101001100",
  44675=>"000000010",
  44676=>"110110101",
  44677=>"001010110",
  44678=>"011001100",
  44679=>"110010101",
  44680=>"101010010",
  44681=>"000001010",
  44682=>"011110110",
  44683=>"100001100",
  44684=>"111011010",
  44685=>"001001110",
  44686=>"001010110",
  44687=>"101000000",
  44688=>"101111111",
  44689=>"000010010",
  44690=>"011001001",
  44691=>"000000111",
  44692=>"000110000",
  44693=>"100101010",
  44694=>"001010110",
  44695=>"100001101",
  44696=>"111100100",
  44697=>"010100000",
  44698=>"011111100",
  44699=>"101010001",
  44700=>"000110100",
  44701=>"001010100",
  44702=>"111000111",
  44703=>"010110001",
  44704=>"000100000",
  44705=>"000000011",
  44706=>"000011001",
  44707=>"011010010",
  44708=>"101000110",
  44709=>"100111101",
  44710=>"101011011",
  44711=>"000100000",
  44712=>"110011101",
  44713=>"001000010",
  44714=>"100011011",
  44715=>"101111001",
  44716=>"010011001",
  44717=>"001101100",
  44718=>"001111011",
  44719=>"011100000",
  44720=>"100111001",
  44721=>"111001110",
  44722=>"101000001",
  44723=>"111110001",
  44724=>"110010110",
  44725=>"111101010",
  44726=>"110001000",
  44727=>"101010001",
  44728=>"011000011",
  44729=>"001011110",
  44730=>"010001111",
  44731=>"001010101",
  44732=>"101101111",
  44733=>"100010010",
  44734=>"000010110",
  44735=>"000000010",
  44736=>"011011010",
  44737=>"000111110",
  44738=>"010001000",
  44739=>"011001000",
  44740=>"110011010",
  44741=>"000000110",
  44742=>"000001010",
  44743=>"110001111",
  44744=>"000101110",
  44745=>"111110011",
  44746=>"010011100",
  44747=>"000010101",
  44748=>"001100000",
  44749=>"000100001",
  44750=>"101011010",
  44751=>"001111001",
  44752=>"010000101",
  44753=>"000001001",
  44754=>"101100001",
  44755=>"010100010",
  44756=>"011011111",
  44757=>"010010101",
  44758=>"011011011",
  44759=>"111100110",
  44760=>"010010011",
  44761=>"010111100",
  44762=>"110100010",
  44763=>"101000011",
  44764=>"011100010",
  44765=>"100001111",
  44766=>"001111111",
  44767=>"000000101",
  44768=>"001000000",
  44769=>"011100101",
  44770=>"011100001",
  44771=>"011101100",
  44772=>"011010011",
  44773=>"011011001",
  44774=>"010100010",
  44775=>"010010110",
  44776=>"001100001",
  44777=>"011010000",
  44778=>"000001110",
  44779=>"100000001",
  44780=>"110011011",
  44781=>"101100001",
  44782=>"111010101",
  44783=>"010111011",
  44784=>"011101100",
  44785=>"100110101",
  44786=>"000000000",
  44787=>"000010100",
  44788=>"010001101",
  44789=>"011011100",
  44790=>"010001000",
  44791=>"110100011",
  44792=>"110100011",
  44793=>"111111001",
  44794=>"111000101",
  44795=>"111011001",
  44796=>"011011010",
  44797=>"111011111",
  44798=>"010001101",
  44799=>"111100000",
  44800=>"001111000",
  44801=>"100101111",
  44802=>"110101111",
  44803=>"101000010",
  44804=>"100010111",
  44805=>"000010000",
  44806=>"010101111",
  44807=>"011001111",
  44808=>"101110011",
  44809=>"101000101",
  44810=>"000001110",
  44811=>"110111001",
  44812=>"111011100",
  44813=>"000000010",
  44814=>"011111110",
  44815=>"011000101",
  44816=>"100111010",
  44817=>"001101000",
  44818=>"011111011",
  44819=>"111001101",
  44820=>"000010001",
  44821=>"000010000",
  44822=>"000101100",
  44823=>"100000001",
  44824=>"110110001",
  44825=>"111110110",
  44826=>"110110010",
  44827=>"000010011",
  44828=>"100011011",
  44829=>"011001000",
  44830=>"000011110",
  44831=>"100110000",
  44832=>"101110010",
  44833=>"011001101",
  44834=>"001100011",
  44835=>"110111010",
  44836=>"100011010",
  44837=>"010100010",
  44838=>"010000110",
  44839=>"100110101",
  44840=>"111100010",
  44841=>"100010111",
  44842=>"100011011",
  44843=>"110010111",
  44844=>"101011011",
  44845=>"000001111",
  44846=>"010000010",
  44847=>"000000100",
  44848=>"111000001",
  44849=>"010101000",
  44850=>"000010010",
  44851=>"111100101",
  44852=>"010100110",
  44853=>"110101010",
  44854=>"110010011",
  44855=>"001111111",
  44856=>"101100001",
  44857=>"101001110",
  44858=>"111000011",
  44859=>"110111011",
  44860=>"111010000",
  44861=>"101101010",
  44862=>"011100000",
  44863=>"001000110",
  44864=>"111001000",
  44865=>"000010111",
  44866=>"011000101",
  44867=>"000100011",
  44868=>"011010100",
  44869=>"100100011",
  44870=>"011110011",
  44871=>"010101011",
  44872=>"100000010",
  44873=>"011100100",
  44874=>"111000000",
  44875=>"010010011",
  44876=>"101100101",
  44877=>"111000011",
  44878=>"101101000",
  44879=>"110100010",
  44880=>"000010011",
  44881=>"000100111",
  44882=>"010110110",
  44883=>"110011111",
  44884=>"110000101",
  44885=>"011011001",
  44886=>"001111101",
  44887=>"111011001",
  44888=>"101001010",
  44889=>"011001111",
  44890=>"011001110",
  44891=>"100000000",
  44892=>"111001011",
  44893=>"001010011",
  44894=>"101011110",
  44895=>"000001100",
  44896=>"011111100",
  44897=>"101110010",
  44898=>"111110001",
  44899=>"101100000",
  44900=>"010110110",
  44901=>"100001010",
  44902=>"001011111",
  44903=>"010100011",
  44904=>"000111110",
  44905=>"010110011",
  44906=>"010000001",
  44907=>"001001101",
  44908=>"010100111",
  44909=>"000100101",
  44910=>"111101000",
  44911=>"010000110",
  44912=>"111110011",
  44913=>"000101110",
  44914=>"101110010",
  44915=>"100011010",
  44916=>"100000010",
  44917=>"011101000",
  44918=>"011110100",
  44919=>"001111000",
  44920=>"000011100",
  44921=>"110111111",
  44922=>"001010010",
  44923=>"010011011",
  44924=>"110001000",
  44925=>"010100000",
  44926=>"001101110",
  44927=>"100101100",
  44928=>"000100000",
  44929=>"111100111",
  44930=>"011011110",
  44931=>"100111000",
  44932=>"000101011",
  44933=>"001000001",
  44934=>"111001001",
  44935=>"010001101",
  44936=>"010101100",
  44937=>"100000111",
  44938=>"010011010",
  44939=>"000111001",
  44940=>"010011111",
  44941=>"100001111",
  44942=>"110110110",
  44943=>"100000000",
  44944=>"110110000",
  44945=>"011101010",
  44946=>"010000011",
  44947=>"000110111",
  44948=>"011110001",
  44949=>"110000101",
  44950=>"000110100",
  44951=>"111101110",
  44952=>"111000101",
  44953=>"000010000",
  44954=>"000100110",
  44955=>"001111000",
  44956=>"110111111",
  44957=>"110100111",
  44958=>"100010100",
  44959=>"110100000",
  44960=>"111100111",
  44961=>"100000011",
  44962=>"110100001",
  44963=>"001011010",
  44964=>"001011000",
  44965=>"111001001",
  44966=>"101111111",
  44967=>"010100100",
  44968=>"011000111",
  44969=>"101010011",
  44970=>"100110000",
  44971=>"110010101",
  44972=>"000100010",
  44973=>"111010011",
  44974=>"001111011",
  44975=>"011011111",
  44976=>"100010010",
  44977=>"001101111",
  44978=>"001010010",
  44979=>"001101010",
  44980=>"010010011",
  44981=>"001111010",
  44982=>"001001110",
  44983=>"111000011",
  44984=>"010100010",
  44985=>"110100010",
  44986=>"010110011",
  44987=>"010010010",
  44988=>"111011000",
  44989=>"001111000",
  44990=>"001110100",
  44991=>"111011111",
  44992=>"000101100",
  44993=>"101101101",
  44994=>"100101101",
  44995=>"011011010",
  44996=>"100011110",
  44997=>"101001000",
  44998=>"010110001",
  44999=>"100100000",
  45000=>"101011101",
  45001=>"101111101",
  45002=>"101100010",
  45003=>"101011000",
  45004=>"011111110",
  45005=>"101001101",
  45006=>"101010101",
  45007=>"010110011",
  45008=>"000110101",
  45009=>"101101000",
  45010=>"011000111",
  45011=>"101001000",
  45012=>"101011111",
  45013=>"100011100",
  45014=>"100110000",
  45015=>"101001011",
  45016=>"100101100",
  45017=>"100110110",
  45018=>"000110100",
  45019=>"001001011",
  45020=>"110110100",
  45021=>"101001011",
  45022=>"011100100",
  45023=>"000010011",
  45024=>"000000101",
  45025=>"111001001",
  45026=>"001100101",
  45027=>"010110000",
  45028=>"001011000",
  45029=>"000010001",
  45030=>"000010010",
  45031=>"000110100",
  45032=>"000011101",
  45033=>"001110001",
  45034=>"000100100",
  45035=>"011011101",
  45036=>"111000000",
  45037=>"111000111",
  45038=>"101000110",
  45039=>"111101001",
  45040=>"101010101",
  45041=>"010010001",
  45042=>"110011000",
  45043=>"110111111",
  45044=>"011010000",
  45045=>"110110001",
  45046=>"000011011",
  45047=>"100000010",
  45048=>"101011111",
  45049=>"110010010",
  45050=>"010110000",
  45051=>"111011011",
  45052=>"100011101",
  45053=>"000110110",
  45054=>"000000000",
  45055=>"100100000",
  45056=>"100001101",
  45057=>"101101001",
  45058=>"010111111",
  45059=>"001001110",
  45060=>"100101001",
  45061=>"110010001",
  45062=>"111100000",
  45063=>"000011111",
  45064=>"110101101",
  45065=>"110110000",
  45066=>"000101011",
  45067=>"110001110",
  45068=>"010000110",
  45069=>"101110111",
  45070=>"111111010",
  45071=>"100110001",
  45072=>"101000111",
  45073=>"000010010",
  45074=>"011110010",
  45075=>"100000001",
  45076=>"011010100",
  45077=>"011001001",
  45078=>"101101101",
  45079=>"010110011",
  45080=>"101111100",
  45081=>"110001101",
  45082=>"110101101",
  45083=>"110101101",
  45084=>"011001010",
  45085=>"000000110",
  45086=>"000101100",
  45087=>"111101110",
  45088=>"101100111",
  45089=>"110011110",
  45090=>"000110010",
  45091=>"010000110",
  45092=>"000100010",
  45093=>"101110001",
  45094=>"011010100",
  45095=>"100111101",
  45096=>"000000101",
  45097=>"000011111",
  45098=>"010110001",
  45099=>"100000101",
  45100=>"101000011",
  45101=>"101111101",
  45102=>"000000011",
  45103=>"100011101",
  45104=>"100001010",
  45105=>"010101101",
  45106=>"000110110",
  45107=>"010011110",
  45108=>"101110110",
  45109=>"000011001",
  45110=>"100110001",
  45111=>"111101101",
  45112=>"111000001",
  45113=>"110010000",
  45114=>"110000000",
  45115=>"000100001",
  45116=>"000000000",
  45117=>"101110001",
  45118=>"011111011",
  45119=>"001011101",
  45120=>"010100100",
  45121=>"000010101",
  45122=>"000111000",
  45123=>"001111110",
  45124=>"011001101",
  45125=>"101100001",
  45126=>"001010100",
  45127=>"100010010",
  45128=>"110011011",
  45129=>"010011110",
  45130=>"001110101",
  45131=>"101000110",
  45132=>"011111011",
  45133=>"011001101",
  45134=>"010111100",
  45135=>"111000000",
  45136=>"010110011",
  45137=>"000001001",
  45138=>"011011011",
  45139=>"101100011",
  45140=>"100001111",
  45141=>"111011101",
  45142=>"000011010",
  45143=>"010101001",
  45144=>"000010011",
  45145=>"111000111",
  45146=>"100010000",
  45147=>"111000111",
  45148=>"010110110",
  45149=>"101001001",
  45150=>"110100010",
  45151=>"101001000",
  45152=>"011101001",
  45153=>"010111011",
  45154=>"000111011",
  45155=>"000010011",
  45156=>"000101001",
  45157=>"110100010",
  45158=>"001000101",
  45159=>"011101110",
  45160=>"111000100",
  45161=>"000010110",
  45162=>"001110101",
  45163=>"001100001",
  45164=>"101001001",
  45165=>"111100101",
  45166=>"010001101",
  45167=>"110000110",
  45168=>"101010111",
  45169=>"101001110",
  45170=>"000011000",
  45171=>"011000011",
  45172=>"000100011",
  45173=>"000010110",
  45174=>"101100111",
  45175=>"101100010",
  45176=>"000001010",
  45177=>"100010011",
  45178=>"000010011",
  45179=>"001010111",
  45180=>"100101001",
  45181=>"010000001",
  45182=>"010110110",
  45183=>"111000000",
  45184=>"000111011",
  45185=>"000001101",
  45186=>"011110011",
  45187=>"001101111",
  45188=>"000011110",
  45189=>"000010110",
  45190=>"111000110",
  45191=>"110100101",
  45192=>"010001010",
  45193=>"001001000",
  45194=>"000011101",
  45195=>"000110001",
  45196=>"100111111",
  45197=>"101101111",
  45198=>"111111111",
  45199=>"001100001",
  45200=>"010101000",
  45201=>"100001101",
  45202=>"111011011",
  45203=>"011100100",
  45204=>"010000101",
  45205=>"110001011",
  45206=>"001010111",
  45207=>"001111100",
  45208=>"010001001",
  45209=>"010001101",
  45210=>"000111100",
  45211=>"000000101",
  45212=>"111111111",
  45213=>"100011101",
  45214=>"010100011",
  45215=>"010111101",
  45216=>"001010001",
  45217=>"110011110",
  45218=>"010101010",
  45219=>"110000010",
  45220=>"011011001",
  45221=>"011010010",
  45222=>"000110100",
  45223=>"100101011",
  45224=>"011001010",
  45225=>"101000000",
  45226=>"000100100",
  45227=>"001110111",
  45228=>"000111011",
  45229=>"001001000",
  45230=>"110010001",
  45231=>"000101000",
  45232=>"010110001",
  45233=>"100010010",
  45234=>"110110011",
  45235=>"111011100",
  45236=>"000100100",
  45237=>"011110110",
  45238=>"010110101",
  45239=>"010000000",
  45240=>"011001110",
  45241=>"011001111",
  45242=>"011101011",
  45243=>"111101101",
  45244=>"001011001",
  45245=>"101000011",
  45246=>"001110111",
  45247=>"101000001",
  45248=>"011001111",
  45249=>"011110011",
  45250=>"011101011",
  45251=>"001111011",
  45252=>"011011011",
  45253=>"010000110",
  45254=>"100011110",
  45255=>"011010000",
  45256=>"101001110",
  45257=>"110100000",
  45258=>"001111000",
  45259=>"000011000",
  45260=>"111100100",
  45261=>"101011000",
  45262=>"100110000",
  45263=>"000010100",
  45264=>"110010100",
  45265=>"000111001",
  45266=>"110111000",
  45267=>"110111000",
  45268=>"110101000",
  45269=>"001011111",
  45270=>"001001101",
  45271=>"101011110",
  45272=>"111101101",
  45273=>"111011010",
  45274=>"010110010",
  45275=>"011101010",
  45276=>"010111001",
  45277=>"001010101",
  45278=>"111001001",
  45279=>"101100000",
  45280=>"110011000",
  45281=>"010010101",
  45282=>"101001110",
  45283=>"011010110",
  45284=>"011011110",
  45285=>"000001001",
  45286=>"000100010",
  45287=>"101110111",
  45288=>"100000100",
  45289=>"111011111",
  45290=>"011110101",
  45291=>"111111000",
  45292=>"011010111",
  45293=>"000000010",
  45294=>"001110000",
  45295=>"100000100",
  45296=>"010010111",
  45297=>"111000110",
  45298=>"011111100",
  45299=>"100000101",
  45300=>"011001011",
  45301=>"011001110",
  45302=>"110000110",
  45303=>"011010001",
  45304=>"100101011",
  45305=>"111100010",
  45306=>"111111101",
  45307=>"101100111",
  45308=>"000010011",
  45309=>"001000100",
  45310=>"110100111",
  45311=>"110000110",
  45312=>"010011100",
  45313=>"000000111",
  45314=>"001100100",
  45315=>"000110011",
  45316=>"111110000",
  45317=>"011110000",
  45318=>"100110110",
  45319=>"010111101",
  45320=>"111111010",
  45321=>"110011010",
  45322=>"000010001",
  45323=>"000101001",
  45324=>"110011001",
  45325=>"110011000",
  45326=>"000010001",
  45327=>"000001000",
  45328=>"011111111",
  45329=>"101011010",
  45330=>"000000010",
  45331=>"101100111",
  45332=>"011111111",
  45333=>"010001101",
  45334=>"100001111",
  45335=>"001011100",
  45336=>"111010100",
  45337=>"001011101",
  45338=>"011111100",
  45339=>"111101011",
  45340=>"001110011",
  45341=>"000101111",
  45342=>"111011110",
  45343=>"001000010",
  45344=>"000101000",
  45345=>"111110110",
  45346=>"001010000",
  45347=>"100100101",
  45348=>"100111011",
  45349=>"100101111",
  45350=>"100011111",
  45351=>"111101111",
  45352=>"100010001",
  45353=>"100010100",
  45354=>"011100100",
  45355=>"010010111",
  45356=>"000110000",
  45357=>"010101100",
  45358=>"011100010",
  45359=>"000010000",
  45360=>"111101001",
  45361=>"000100000",
  45362=>"010110101",
  45363=>"000111010",
  45364=>"110101110",
  45365=>"101110100",
  45366=>"110001111",
  45367=>"111111011",
  45368=>"101101111",
  45369=>"111011001",
  45370=>"001001111",
  45371=>"001110001",
  45372=>"000100100",
  45373=>"001000100",
  45374=>"000100011",
  45375=>"101111010",
  45376=>"101101110",
  45377=>"001111100",
  45378=>"110110101",
  45379=>"000010011",
  45380=>"010011000",
  45381=>"000001001",
  45382=>"100111110",
  45383=>"010111001",
  45384=>"100100010",
  45385=>"000011001",
  45386=>"100000001",
  45387=>"001110110",
  45388=>"010010100",
  45389=>"101100000",
  45390=>"001100100",
  45391=>"111010100",
  45392=>"100001111",
  45393=>"010010010",
  45394=>"010000010",
  45395=>"101000010",
  45396=>"011011011",
  45397=>"100111011",
  45398=>"110111000",
  45399=>"101100101",
  45400=>"001000110",
  45401=>"111111011",
  45402=>"001001111",
  45403=>"010011000",
  45404=>"010000001",
  45405=>"100001111",
  45406=>"111011001",
  45407=>"101011111",
  45408=>"111110011",
  45409=>"110001111",
  45410=>"011001010",
  45411=>"000110001",
  45412=>"000100001",
  45413=>"100111111",
  45414=>"100100101",
  45415=>"011101010",
  45416=>"011011000",
  45417=>"000110000",
  45418=>"000011000",
  45419=>"001011101",
  45420=>"101010011",
  45421=>"010000010",
  45422=>"100011011",
  45423=>"011100101",
  45424=>"000000001",
  45425=>"111101010",
  45426=>"100001011",
  45427=>"001011101",
  45428=>"110111100",
  45429=>"011100110",
  45430=>"101010010",
  45431=>"100001001",
  45432=>"011001010",
  45433=>"110100101",
  45434=>"100000101",
  45435=>"111110101",
  45436=>"011010001",
  45437=>"111010000",
  45438=>"101110110",
  45439=>"100111111",
  45440=>"000110111",
  45441=>"001100101",
  45442=>"100100011",
  45443=>"111011111",
  45444=>"100011000",
  45445=>"010011011",
  45446=>"111100011",
  45447=>"000101000",
  45448=>"011001010",
  45449=>"011100001",
  45450=>"000011101",
  45451=>"010110101",
  45452=>"000100111",
  45453=>"001110011",
  45454=>"000111011",
  45455=>"111010011",
  45456=>"010010101",
  45457=>"111100010",
  45458=>"001110010",
  45459=>"110011110",
  45460=>"010011101",
  45461=>"001000001",
  45462=>"111001011",
  45463=>"000101100",
  45464=>"001001010",
  45465=>"000000100",
  45466=>"010010000",
  45467=>"010100010",
  45468=>"001000110",
  45469=>"001110111",
  45470=>"000101110",
  45471=>"101101100",
  45472=>"001100001",
  45473=>"011010001",
  45474=>"111110110",
  45475=>"011001011",
  45476=>"101001100",
  45477=>"001011111",
  45478=>"001111101",
  45479=>"011000010",
  45480=>"101010010",
  45481=>"111011000",
  45482=>"111111011",
  45483=>"100010100",
  45484=>"011011101",
  45485=>"100111001",
  45486=>"001111010",
  45487=>"011000000",
  45488=>"000101110",
  45489=>"100001001",
  45490=>"001011101",
  45491=>"111110010",
  45492=>"101100010",
  45493=>"001111110",
  45494=>"011000010",
  45495=>"010001000",
  45496=>"001000111",
  45497=>"000110110",
  45498=>"110100000",
  45499=>"011110011",
  45500=>"001110000",
  45501=>"000110110",
  45502=>"000000110",
  45503=>"111110111",
  45504=>"101101111",
  45505=>"011000101",
  45506=>"001011011",
  45507=>"000001011",
  45508=>"011110001",
  45509=>"100100000",
  45510=>"101110110",
  45511=>"000100000",
  45512=>"111111101",
  45513=>"111110111",
  45514=>"010000100",
  45515=>"111000010",
  45516=>"111100101",
  45517=>"100000110",
  45518=>"101001010",
  45519=>"100011110",
  45520=>"111001110",
  45521=>"101000001",
  45522=>"110000010",
  45523=>"000011101",
  45524=>"111111001",
  45525=>"100101000",
  45526=>"111000001",
  45527=>"110100011",
  45528=>"100001110",
  45529=>"101111101",
  45530=>"101101100",
  45531=>"110100101",
  45532=>"100111111",
  45533=>"001101110",
  45534=>"101100111",
  45535=>"011111000",
  45536=>"111010110",
  45537=>"111000110",
  45538=>"010000010",
  45539=>"011111111",
  45540=>"111110110",
  45541=>"110010100",
  45542=>"101010101",
  45543=>"100110001",
  45544=>"001110100",
  45545=>"100101100",
  45546=>"110111000",
  45547=>"110111101",
  45548=>"011110111",
  45549=>"111011100",
  45550=>"001101000",
  45551=>"100010100",
  45552=>"111010011",
  45553=>"101100100",
  45554=>"111000001",
  45555=>"101101100",
  45556=>"001100100",
  45557=>"001010011",
  45558=>"000101101",
  45559=>"000101101",
  45560=>"110010101",
  45561=>"011010010",
  45562=>"001111001",
  45563=>"111101011",
  45564=>"011010110",
  45565=>"011110101",
  45566=>"010001001",
  45567=>"100111010",
  45568=>"110111110",
  45569=>"000101010",
  45570=>"110001000",
  45571=>"111000100",
  45572=>"001101100",
  45573=>"001010101",
  45574=>"110111011",
  45575=>"100010100",
  45576=>"010001011",
  45577=>"101010010",
  45578=>"001000000",
  45579=>"010000100",
  45580=>"001010010",
  45581=>"101101100",
  45582=>"000000001",
  45583=>"111011101",
  45584=>"010011100",
  45585=>"100101000",
  45586=>"100010010",
  45587=>"111111101",
  45588=>"100111111",
  45589=>"100010010",
  45590=>"110011000",
  45591=>"101111101",
  45592=>"000101000",
  45593=>"000111111",
  45594=>"011001010",
  45595=>"001111101",
  45596=>"011100001",
  45597=>"001111111",
  45598=>"111011111",
  45599=>"100101111",
  45600=>"010110111",
  45601=>"010001111",
  45602=>"000000100",
  45603=>"110111000",
  45604=>"010010001",
  45605=>"010001011",
  45606=>"010011101",
  45607=>"000110010",
  45608=>"000111110",
  45609=>"001001010",
  45610=>"101011101",
  45611=>"001011110",
  45612=>"000110101",
  45613=>"000010000",
  45614=>"000110110",
  45615=>"101010011",
  45616=>"111100110",
  45617=>"010101001",
  45618=>"010101000",
  45619=>"000011101",
  45620=>"000110010",
  45621=>"010000010",
  45622=>"010100101",
  45623=>"000111000",
  45624=>"110111010",
  45625=>"000100110",
  45626=>"101101001",
  45627=>"111000010",
  45628=>"000100101",
  45629=>"110001000",
  45630=>"111110110",
  45631=>"000110101",
  45632=>"101101110",
  45633=>"101110011",
  45634=>"001010001",
  45635=>"110001101",
  45636=>"000110100",
  45637=>"111110001",
  45638=>"110110001",
  45639=>"110000111",
  45640=>"100100111",
  45641=>"100101110",
  45642=>"011010000",
  45643=>"000000001",
  45644=>"011010101",
  45645=>"001000100",
  45646=>"000101010",
  45647=>"111000001",
  45648=>"100010110",
  45649=>"011000110",
  45650=>"010111000",
  45651=>"100111110",
  45652=>"011011001",
  45653=>"011000000",
  45654=>"111101100",
  45655=>"100000000",
  45656=>"011110101",
  45657=>"111000001",
  45658=>"111000010",
  45659=>"111100011",
  45660=>"100001100",
  45661=>"011110110",
  45662=>"111110000",
  45663=>"110000000",
  45664=>"001000001",
  45665=>"011111100",
  45666=>"101010001",
  45667=>"110000111",
  45668=>"011000100",
  45669=>"101110011",
  45670=>"100110110",
  45671=>"011101010",
  45672=>"100010000",
  45673=>"010000000",
  45674=>"001101111",
  45675=>"000101101",
  45676=>"001010010",
  45677=>"101010000",
  45678=>"110101011",
  45679=>"111000011",
  45680=>"001111101",
  45681=>"111101001",
  45682=>"001001011",
  45683=>"011100010",
  45684=>"001110011",
  45685=>"111001001",
  45686=>"001010101",
  45687=>"101001001",
  45688=>"000110101",
  45689=>"011000100",
  45690=>"001010101",
  45691=>"110110011",
  45692=>"000101010",
  45693=>"100010110",
  45694=>"011111001",
  45695=>"000010001",
  45696=>"010000110",
  45697=>"100000101",
  45698=>"100111101",
  45699=>"111001101",
  45700=>"000010100",
  45701=>"101110101",
  45702=>"110111000",
  45703=>"011111111",
  45704=>"011100011",
  45705=>"110001001",
  45706=>"011110001",
  45707=>"101000011",
  45708=>"001010000",
  45709=>"000111000",
  45710=>"001010100",
  45711=>"100000000",
  45712=>"010111101",
  45713=>"111011000",
  45714=>"011111000",
  45715=>"101001100",
  45716=>"001010100",
  45717=>"000000101",
  45718=>"001100100",
  45719=>"011101000",
  45720=>"101001110",
  45721=>"111100010",
  45722=>"010111010",
  45723=>"110100111",
  45724=>"000110100",
  45725=>"110001010",
  45726=>"001001110",
  45727=>"011001100",
  45728=>"011010010",
  45729=>"000111111",
  45730=>"010100000",
  45731=>"101111110",
  45732=>"001001111",
  45733=>"000010100",
  45734=>"101100001",
  45735=>"101111110",
  45736=>"100000100",
  45737=>"110011000",
  45738=>"001011110",
  45739=>"110111011",
  45740=>"000100011",
  45741=>"000010010",
  45742=>"001001100",
  45743=>"110010010",
  45744=>"111010000",
  45745=>"001101100",
  45746=>"000111111",
  45747=>"011101001",
  45748=>"111111101",
  45749=>"011001100",
  45750=>"010011100",
  45751=>"111001100",
  45752=>"110010101",
  45753=>"111000110",
  45754=>"011100001",
  45755=>"110011111",
  45756=>"101100001",
  45757=>"110001100",
  45758=>"000010001",
  45759=>"100110010",
  45760=>"101111000",
  45761=>"010011110",
  45762=>"101011101",
  45763=>"100000110",
  45764=>"010010100",
  45765=>"000110000",
  45766=>"010000111",
  45767=>"100000100",
  45768=>"110111011",
  45769=>"001000100",
  45770=>"010011010",
  45771=>"110101001",
  45772=>"101101111",
  45773=>"100011110",
  45774=>"100101110",
  45775=>"010010100",
  45776=>"011010010",
  45777=>"000111001",
  45778=>"110110100",
  45779=>"010101100",
  45780=>"111011000",
  45781=>"101001110",
  45782=>"110000010",
  45783=>"101000101",
  45784=>"101110010",
  45785=>"000000000",
  45786=>"010111011",
  45787=>"111000000",
  45788=>"110100101",
  45789=>"000010001",
  45790=>"101110101",
  45791=>"011000011",
  45792=>"111111001",
  45793=>"010010111",
  45794=>"000101011",
  45795=>"011011111",
  45796=>"101001001",
  45797=>"000000000",
  45798=>"010001000",
  45799=>"101111001",
  45800=>"001110100",
  45801=>"011011000",
  45802=>"111101111",
  45803=>"101000001",
  45804=>"001111111",
  45805=>"000101000",
  45806=>"001010010",
  45807=>"001010001",
  45808=>"000100011",
  45809=>"000010010",
  45810=>"001000101",
  45811=>"001101110",
  45812=>"000110100",
  45813=>"011000000",
  45814=>"001110100",
  45815=>"110100100",
  45816=>"101011011",
  45817=>"010100011",
  45818=>"001111100",
  45819=>"000000101",
  45820=>"000101101",
  45821=>"011010011",
  45822=>"110100000",
  45823=>"000000000",
  45824=>"000001111",
  45825=>"010011011",
  45826=>"110000101",
  45827=>"011111110",
  45828=>"011010010",
  45829=>"100110001",
  45830=>"001110000",
  45831=>"001011010",
  45832=>"110010010",
  45833=>"110000111",
  45834=>"000001010",
  45835=>"111011111",
  45836=>"000011011",
  45837=>"011011010",
  45838=>"111111110",
  45839=>"001101111",
  45840=>"010101101",
  45841=>"000000000",
  45842=>"101100101",
  45843=>"110010000",
  45844=>"011110001",
  45845=>"011011010",
  45846=>"100000101",
  45847=>"011111000",
  45848=>"101111000",
  45849=>"011001111",
  45850=>"110001010",
  45851=>"110011011",
  45852=>"101000110",
  45853=>"101101101",
  45854=>"000001101",
  45855=>"001101111",
  45856=>"101001100",
  45857=>"000001101",
  45858=>"110110010",
  45859=>"000101001",
  45860=>"000010100",
  45861=>"000000110",
  45862=>"000000101",
  45863=>"011010000",
  45864=>"011111000",
  45865=>"111011000",
  45866=>"011100100",
  45867=>"101011110",
  45868=>"110101010",
  45869=>"001101101",
  45870=>"111010101",
  45871=>"010010001",
  45872=>"010001000",
  45873=>"101101001",
  45874=>"101101100",
  45875=>"010010101",
  45876=>"010110000",
  45877=>"011101100",
  45878=>"100010010",
  45879=>"000010010",
  45880=>"111111011",
  45881=>"001000100",
  45882=>"011000000",
  45883=>"110011001",
  45884=>"101001100",
  45885=>"101100000",
  45886=>"101110111",
  45887=>"111100001",
  45888=>"100010101",
  45889=>"101010111",
  45890=>"100000011",
  45891=>"010011011",
  45892=>"101000010",
  45893=>"011100000",
  45894=>"101100110",
  45895=>"101110000",
  45896=>"101110010",
  45897=>"010110101",
  45898=>"001010000",
  45899=>"000100110",
  45900=>"001011000",
  45901=>"110100000",
  45902=>"010101110",
  45903=>"111110001",
  45904=>"110100110",
  45905=>"011001111",
  45906=>"010101111",
  45907=>"111011100",
  45908=>"101011011",
  45909=>"100000000",
  45910=>"001100011",
  45911=>"000001110",
  45912=>"011111110",
  45913=>"100001101",
  45914=>"000001101",
  45915=>"000001101",
  45916=>"101110000",
  45917=>"111111000",
  45918=>"100110001",
  45919=>"000110111",
  45920=>"101101110",
  45921=>"101100010",
  45922=>"100011100",
  45923=>"111111001",
  45924=>"101111011",
  45925=>"111101100",
  45926=>"001010000",
  45927=>"110111101",
  45928=>"000011001",
  45929=>"000110110",
  45930=>"011011111",
  45931=>"010000000",
  45932=>"111110101",
  45933=>"000000001",
  45934=>"110010000",
  45935=>"111001110",
  45936=>"100000111",
  45937=>"011111101",
  45938=>"010011010",
  45939=>"111111001",
  45940=>"101101110",
  45941=>"111011000",
  45942=>"001111010",
  45943=>"110100000",
  45944=>"010101011",
  45945=>"000000000",
  45946=>"100001001",
  45947=>"011101110",
  45948=>"110000110",
  45949=>"100000001",
  45950=>"101111111",
  45951=>"101000011",
  45952=>"100101111",
  45953=>"010011111",
  45954=>"111110001",
  45955=>"110111000",
  45956=>"101101000",
  45957=>"100001110",
  45958=>"111010101",
  45959=>"100110111",
  45960=>"111010100",
  45961=>"110111000",
  45962=>"000011111",
  45963=>"011001000",
  45964=>"010100110",
  45965=>"111111010",
  45966=>"101101000",
  45967=>"011000010",
  45968=>"110010101",
  45969=>"001101100",
  45970=>"000000110",
  45971=>"000000001",
  45972=>"011110101",
  45973=>"100100101",
  45974=>"100000010",
  45975=>"110011010",
  45976=>"111011010",
  45977=>"000100111",
  45978=>"000010100",
  45979=>"101001110",
  45980=>"110101001",
  45981=>"101101011",
  45982=>"100101100",
  45983=>"011111011",
  45984=>"101111110",
  45985=>"001110110",
  45986=>"110100101",
  45987=>"001101101",
  45988=>"000100010",
  45989=>"000010110",
  45990=>"000001101",
  45991=>"000101011",
  45992=>"101011111",
  45993=>"111010011",
  45994=>"011110010",
  45995=>"110110111",
  45996=>"000000000",
  45997=>"011110010",
  45998=>"111111010",
  45999=>"000111000",
  46000=>"100110110",
  46001=>"111001100",
  46002=>"101111010",
  46003=>"101111001",
  46004=>"110111100",
  46005=>"010111001",
  46006=>"011101000",
  46007=>"011101100",
  46008=>"110000111",
  46009=>"100001110",
  46010=>"011100011",
  46011=>"011111111",
  46012=>"011001110",
  46013=>"111101011",
  46014=>"011001010",
  46015=>"110110010",
  46016=>"000010010",
  46017=>"011000111",
  46018=>"101000010",
  46019=>"100010010",
  46020=>"101001101",
  46021=>"101011111",
  46022=>"001001101",
  46023=>"110011011",
  46024=>"101000100",
  46025=>"100001011",
  46026=>"100000101",
  46027=>"001000011",
  46028=>"011011111",
  46029=>"010010101",
  46030=>"110100011",
  46031=>"111100000",
  46032=>"010101011",
  46033=>"111111110",
  46034=>"011011110",
  46035=>"111010010",
  46036=>"011111000",
  46037=>"101011101",
  46038=>"110110010",
  46039=>"010111110",
  46040=>"010110011",
  46041=>"010010101",
  46042=>"010100101",
  46043=>"111110110",
  46044=>"000000011",
  46045=>"110010000",
  46046=>"000000111",
  46047=>"010000111",
  46048=>"000010010",
  46049=>"001111000",
  46050=>"000000010",
  46051=>"100110111",
  46052=>"101010110",
  46053=>"011111000",
  46054=>"000001001",
  46055=>"010011111",
  46056=>"000001111",
  46057=>"101110011",
  46058=>"111010110",
  46059=>"000101111",
  46060=>"010000001",
  46061=>"111101101",
  46062=>"010010010",
  46063=>"101101111",
  46064=>"010001101",
  46065=>"000101011",
  46066=>"100110111",
  46067=>"000101000",
  46068=>"101111100",
  46069=>"111101011",
  46070=>"100000001",
  46071=>"111001110",
  46072=>"110101100",
  46073=>"100101110",
  46074=>"001010111",
  46075=>"010000000",
  46076=>"010001001",
  46077=>"110001001",
  46078=>"111000011",
  46079=>"101101010",
  46080=>"000101001",
  46081=>"011111110",
  46082=>"101110111",
  46083=>"110011010",
  46084=>"101111100",
  46085=>"011011011",
  46086=>"000111010",
  46087=>"010010101",
  46088=>"010010000",
  46089=>"001110101",
  46090=>"001001010",
  46091=>"011101011",
  46092=>"101100101",
  46093=>"110101010",
  46094=>"000101000",
  46095=>"001001010",
  46096=>"110000101",
  46097=>"000101101",
  46098=>"110111110",
  46099=>"110101010",
  46100=>"000101000",
  46101=>"100100000",
  46102=>"101011001",
  46103=>"111011111",
  46104=>"111110000",
  46105=>"111111011",
  46106=>"111110010",
  46107=>"001110110",
  46108=>"011101010",
  46109=>"000010001",
  46110=>"100100000",
  46111=>"100000010",
  46112=>"101001111",
  46113=>"101010101",
  46114=>"010111011",
  46115=>"011111001",
  46116=>"010011001",
  46117=>"010001100",
  46118=>"000100001",
  46119=>"011111101",
  46120=>"000010011",
  46121=>"101000000",
  46122=>"011000000",
  46123=>"100010011",
  46124=>"011010011",
  46125=>"010101101",
  46126=>"000000111",
  46127=>"101100101",
  46128=>"110010010",
  46129=>"001101101",
  46130=>"010110100",
  46131=>"011010100",
  46132=>"111011110",
  46133=>"001001000",
  46134=>"011001100",
  46135=>"010011011",
  46136=>"011001000",
  46137=>"100010110",
  46138=>"011100111",
  46139=>"101110000",
  46140=>"100101000",
  46141=>"100010100",
  46142=>"101100011",
  46143=>"010110011",
  46144=>"101011010",
  46145=>"000100010",
  46146=>"111000010",
  46147=>"111000101",
  46148=>"110101111",
  46149=>"100011101",
  46150=>"000000010",
  46151=>"011000001",
  46152=>"011111100",
  46153=>"100100111",
  46154=>"011110011",
  46155=>"100001001",
  46156=>"111110001",
  46157=>"100001111",
  46158=>"011110001",
  46159=>"101010011",
  46160=>"000110000",
  46161=>"001111000",
  46162=>"111111111",
  46163=>"100111101",
  46164=>"110011100",
  46165=>"011000101",
  46166=>"011011111",
  46167=>"001001110",
  46168=>"011001100",
  46169=>"000010110",
  46170=>"111001010",
  46171=>"100001100",
  46172=>"111111010",
  46173=>"000101111",
  46174=>"000010010",
  46175=>"011000111",
  46176=>"011001000",
  46177=>"111111101",
  46178=>"000010011",
  46179=>"000000011",
  46180=>"101000110",
  46181=>"111010100",
  46182=>"000010000",
  46183=>"110110010",
  46184=>"110001110",
  46185=>"110111101",
  46186=>"100110110",
  46187=>"100000101",
  46188=>"010110010",
  46189=>"010001011",
  46190=>"000001100",
  46191=>"110010111",
  46192=>"011000001",
  46193=>"010110000",
  46194=>"010010111",
  46195=>"110110000",
  46196=>"110010010",
  46197=>"000000101",
  46198=>"001111000",
  46199=>"111100010",
  46200=>"010000001",
  46201=>"100110100",
  46202=>"010110000",
  46203=>"111001000",
  46204=>"101100111",
  46205=>"000010111",
  46206=>"100011001",
  46207=>"000001011",
  46208=>"011000010",
  46209=>"001001011",
  46210=>"101100101",
  46211=>"010000100",
  46212=>"110000110",
  46213=>"111011000",
  46214=>"100010000",
  46215=>"110110111",
  46216=>"110100010",
  46217=>"000010110",
  46218=>"100010011",
  46219=>"111101010",
  46220=>"000111010",
  46221=>"111010011",
  46222=>"101100000",
  46223=>"001000000",
  46224=>"111101100",
  46225=>"110100011",
  46226=>"011110111",
  46227=>"011000110",
  46228=>"000000110",
  46229=>"100111100",
  46230=>"011100101",
  46231=>"110001000",
  46232=>"110110101",
  46233=>"111101001",
  46234=>"110010110",
  46235=>"001001001",
  46236=>"100110111",
  46237=>"010011010",
  46238=>"101100101",
  46239=>"011001011",
  46240=>"000100011",
  46241=>"111001001",
  46242=>"011101000",
  46243=>"000110001",
  46244=>"000001110",
  46245=>"111100110",
  46246=>"001100101",
  46247=>"101110101",
  46248=>"101110011",
  46249=>"000111001",
  46250=>"110111111",
  46251=>"010011111",
  46252=>"010101000",
  46253=>"110001100",
  46254=>"000101000",
  46255=>"010000100",
  46256=>"000100111",
  46257=>"100100100",
  46258=>"101001100",
  46259=>"110100111",
  46260=>"100101011",
  46261=>"010011001",
  46262=>"111001001",
  46263=>"110011000",
  46264=>"001010010",
  46265=>"100101100",
  46266=>"001110001",
  46267=>"000110000",
  46268=>"100100100",
  46269=>"100111010",
  46270=>"111100111",
  46271=>"101110001",
  46272=>"001010010",
  46273=>"101000111",
  46274=>"111101000",
  46275=>"101100010",
  46276=>"101110100",
  46277=>"000101110",
  46278=>"101000001",
  46279=>"000001000",
  46280=>"111011111",
  46281=>"111000000",
  46282=>"110000110",
  46283=>"001111011",
  46284=>"000111101",
  46285=>"100001111",
  46286=>"110011000",
  46287=>"101011011",
  46288=>"101001100",
  46289=>"100101110",
  46290=>"111000001",
  46291=>"000101101",
  46292=>"110000011",
  46293=>"111000111",
  46294=>"011110111",
  46295=>"000000001",
  46296=>"101001000",
  46297=>"101001001",
  46298=>"010110000",
  46299=>"101100000",
  46300=>"011001010",
  46301=>"110001011",
  46302=>"111010101",
  46303=>"010101010",
  46304=>"011111111",
  46305=>"101100001",
  46306=>"000001010",
  46307=>"101111100",
  46308=>"110000110",
  46309=>"011100111",
  46310=>"101101000",
  46311=>"101110111",
  46312=>"010110111",
  46313=>"100000100",
  46314=>"111011100",
  46315=>"010111101",
  46316=>"111111111",
  46317=>"111000110",
  46318=>"011110100",
  46319=>"101010100",
  46320=>"101011100",
  46321=>"010011001",
  46322=>"101110000",
  46323=>"110000010",
  46324=>"100011001",
  46325=>"000111100",
  46326=>"111110111",
  46327=>"010110110",
  46328=>"101101010",
  46329=>"100000110",
  46330=>"111101111",
  46331=>"010111001",
  46332=>"101000101",
  46333=>"111100100",
  46334=>"010010111",
  46335=>"010011111",
  46336=>"000100011",
  46337=>"111010110",
  46338=>"111111111",
  46339=>"010011111",
  46340=>"101000100",
  46341=>"011001000",
  46342=>"111000110",
  46343=>"100110110",
  46344=>"111110100",
  46345=>"000000011",
  46346=>"001001100",
  46347=>"010100101",
  46348=>"100000010",
  46349=>"011100101",
  46350=>"001100011",
  46351=>"010010101",
  46352=>"110000010",
  46353=>"011111111",
  46354=>"110100100",
  46355=>"110111110",
  46356=>"110100010",
  46357=>"001101011",
  46358=>"000001111",
  46359=>"110111111",
  46360=>"001100000",
  46361=>"001010000",
  46362=>"000111111",
  46363=>"110100011",
  46364=>"001001001",
  46365=>"111101011",
  46366=>"010101111",
  46367=>"001101110",
  46368=>"010000100",
  46369=>"100011000",
  46370=>"001001100",
  46371=>"111101000",
  46372=>"100111100",
  46373=>"100101100",
  46374=>"100011000",
  46375=>"111001111",
  46376=>"110001101",
  46377=>"100110110",
  46378=>"101110000",
  46379=>"010011011",
  46380=>"011100010",
  46381=>"010000000",
  46382=>"000000001",
  46383=>"111010011",
  46384=>"010000010",
  46385=>"010000110",
  46386=>"101110111",
  46387=>"111101111",
  46388=>"111000101",
  46389=>"000110010",
  46390=>"001001111",
  46391=>"000101111",
  46392=>"010110000",
  46393=>"001010010",
  46394=>"110001110",
  46395=>"000000001",
  46396=>"110001011",
  46397=>"111110000",
  46398=>"000001110",
  46399=>"001100010",
  46400=>"110000111",
  46401=>"110001000",
  46402=>"100001100",
  46403=>"101101011",
  46404=>"100100101",
  46405=>"111111110",
  46406=>"000000001",
  46407=>"111111010",
  46408=>"100010010",
  46409=>"010101111",
  46410=>"000011100",
  46411=>"000101101",
  46412=>"100010010",
  46413=>"110110100",
  46414=>"010100001",
  46415=>"111010111",
  46416=>"111010000",
  46417=>"110111110",
  46418=>"011101111",
  46419=>"100000001",
  46420=>"001111000",
  46421=>"101100000",
  46422=>"110000011",
  46423=>"111111111",
  46424=>"101001110",
  46425=>"000100100",
  46426=>"000110110",
  46427=>"010101011",
  46428=>"011010100",
  46429=>"001000000",
  46430=>"011100011",
  46431=>"110101011",
  46432=>"011111010",
  46433=>"110101001",
  46434=>"101100100",
  46435=>"001011000",
  46436=>"010010000",
  46437=>"010000000",
  46438=>"011000110",
  46439=>"101000110",
  46440=>"101110011",
  46441=>"001001100",
  46442=>"010000010",
  46443=>"011100001",
  46444=>"001011010",
  46445=>"111010000",
  46446=>"110100111",
  46447=>"111111000",
  46448=>"100101101",
  46449=>"110001011",
  46450=>"010100011",
  46451=>"000110111",
  46452=>"101000111",
  46453=>"010001100",
  46454=>"110110110",
  46455=>"001110110",
  46456=>"000110000",
  46457=>"011110100",
  46458=>"000000001",
  46459=>"111001010",
  46460=>"000100011",
  46461=>"110100011",
  46462=>"010110010",
  46463=>"100011111",
  46464=>"101111111",
  46465=>"100010101",
  46466=>"001101001",
  46467=>"110010000",
  46468=>"010110011",
  46469=>"010100110",
  46470=>"111101111",
  46471=>"111111111",
  46472=>"011110011",
  46473=>"101001111",
  46474=>"111010100",
  46475=>"101001101",
  46476=>"000010011",
  46477=>"110101100",
  46478=>"101111100",
  46479=>"110011000",
  46480=>"010011001",
  46481=>"010001100",
  46482=>"000000110",
  46483=>"011100110",
  46484=>"010000011",
  46485=>"111001111",
  46486=>"000011000",
  46487=>"001001110",
  46488=>"000101001",
  46489=>"001000011",
  46490=>"010000001",
  46491=>"100011001",
  46492=>"010000100",
  46493=>"100111101",
  46494=>"000100001",
  46495=>"101010111",
  46496=>"110011000",
  46497=>"000011011",
  46498=>"111110100",
  46499=>"010010101",
  46500=>"111000100",
  46501=>"001100111",
  46502=>"010111111",
  46503=>"101100000",
  46504=>"100111010",
  46505=>"101110101",
  46506=>"111011101",
  46507=>"010001101",
  46508=>"110101101",
  46509=>"001111110",
  46510=>"000010001",
  46511=>"001110011",
  46512=>"101010000",
  46513=>"100001101",
  46514=>"110111011",
  46515=>"110011001",
  46516=>"010110100",
  46517=>"001101011",
  46518=>"001110100",
  46519=>"111001010",
  46520=>"101101101",
  46521=>"110010100",
  46522=>"010101110",
  46523=>"001010111",
  46524=>"000000000",
  46525=>"110000111",
  46526=>"000110011",
  46527=>"111011110",
  46528=>"001100100",
  46529=>"010101010",
  46530=>"000010110",
  46531=>"010101001",
  46532=>"100000001",
  46533=>"000111100",
  46534=>"110011100",
  46535=>"010000000",
  46536=>"011000000",
  46537=>"101010011",
  46538=>"000001100",
  46539=>"111110001",
  46540=>"100010110",
  46541=>"100100001",
  46542=>"110010101",
  46543=>"011101101",
  46544=>"001011011",
  46545=>"110110111",
  46546=>"100011000",
  46547=>"111111001",
  46548=>"000000011",
  46549=>"011011110",
  46550=>"011110000",
  46551=>"101110000",
  46552=>"000000111",
  46553=>"111000110",
  46554=>"000011000",
  46555=>"011110011",
  46556=>"011001000",
  46557=>"100100010",
  46558=>"111010010",
  46559=>"010000110",
  46560=>"111110000",
  46561=>"101100110",
  46562=>"011101100",
  46563=>"011001000",
  46564=>"011100100",
  46565=>"100001000",
  46566=>"000100111",
  46567=>"110101111",
  46568=>"100000001",
  46569=>"001011100",
  46570=>"011110111",
  46571=>"001100100",
  46572=>"100001000",
  46573=>"010110111",
  46574=>"101000000",
  46575=>"010101111",
  46576=>"101010101",
  46577=>"100101111",
  46578=>"101001000",
  46579=>"100111000",
  46580=>"000001000",
  46581=>"011110011",
  46582=>"001101111",
  46583=>"000110000",
  46584=>"011111010",
  46585=>"000000100",
  46586=>"000001000",
  46587=>"111011100",
  46588=>"110100001",
  46589=>"001111100",
  46590=>"000110100",
  46591=>"010100101",
  46592=>"000110000",
  46593=>"000110010",
  46594=>"100100000",
  46595=>"111011010",
  46596=>"101111100",
  46597=>"100000010",
  46598=>"110010110",
  46599=>"011100011",
  46600=>"110011111",
  46601=>"000000111",
  46602=>"100010001",
  46603=>"011010011",
  46604=>"100110001",
  46605=>"111011111",
  46606=>"001001011",
  46607=>"001000011",
  46608=>"110101001",
  46609=>"101001010",
  46610=>"011001101",
  46611=>"011000011",
  46612=>"001110000",
  46613=>"110001101",
  46614=>"111100100",
  46615=>"100100110",
  46616=>"101110100",
  46617=>"101011111",
  46618=>"001001110",
  46619=>"101011101",
  46620=>"001100110",
  46621=>"011010100",
  46622=>"110110110",
  46623=>"010001010",
  46624=>"001011010",
  46625=>"010100011",
  46626=>"101111011",
  46627=>"100000111",
  46628=>"001010111",
  46629=>"110001000",
  46630=>"110010010",
  46631=>"111000110",
  46632=>"101001110",
  46633=>"000110101",
  46634=>"000011011",
  46635=>"001100010",
  46636=>"101101001",
  46637=>"010011100",
  46638=>"101000000",
  46639=>"010000000",
  46640=>"000000010",
  46641=>"011000011",
  46642=>"000101110",
  46643=>"000110100",
  46644=>"100001110",
  46645=>"010100101",
  46646=>"101000000",
  46647=>"000000010",
  46648=>"011011010",
  46649=>"110000111",
  46650=>"001010010",
  46651=>"101100100",
  46652=>"010001100",
  46653=>"000100111",
  46654=>"011010010",
  46655=>"111111011",
  46656=>"000001000",
  46657=>"101001010",
  46658=>"100011011",
  46659=>"110010101",
  46660=>"111001010",
  46661=>"100000111",
  46662=>"010000010",
  46663=>"011111011",
  46664=>"011010101",
  46665=>"110101000",
  46666=>"100011110",
  46667=>"000010001",
  46668=>"011100010",
  46669=>"101010011",
  46670=>"111000000",
  46671=>"100010010",
  46672=>"110010011",
  46673=>"011010000",
  46674=>"000100111",
  46675=>"101011000",
  46676=>"111111011",
  46677=>"111001011",
  46678=>"011011100",
  46679=>"111100111",
  46680=>"111001011",
  46681=>"111110001",
  46682=>"011101111",
  46683=>"101100011",
  46684=>"100010110",
  46685=>"010001010",
  46686=>"101111001",
  46687=>"010100100",
  46688=>"100110110",
  46689=>"111101010",
  46690=>"111010110",
  46691=>"000100110",
  46692=>"111011110",
  46693=>"110001101",
  46694=>"010101111",
  46695=>"011001010",
  46696=>"100010011",
  46697=>"011101011",
  46698=>"101000011",
  46699=>"100000000",
  46700=>"110010000",
  46701=>"111100011",
  46702=>"011101101",
  46703=>"000101000",
  46704=>"001001011",
  46705=>"110100001",
  46706=>"001100001",
  46707=>"001000010",
  46708=>"101111000",
  46709=>"010111110",
  46710=>"010110101",
  46711=>"111010000",
  46712=>"010000110",
  46713=>"011011010",
  46714=>"101101101",
  46715=>"101110110",
  46716=>"100111111",
  46717=>"000101100",
  46718=>"110011110",
  46719=>"101010011",
  46720=>"001000111",
  46721=>"111101101",
  46722=>"111110111",
  46723=>"100011010",
  46724=>"100011001",
  46725=>"100011011",
  46726=>"001010101",
  46727=>"111001000",
  46728=>"111111110",
  46729=>"000000010",
  46730=>"011010010",
  46731=>"111010001",
  46732=>"001011101",
  46733=>"011010100",
  46734=>"000000111",
  46735=>"100000010",
  46736=>"101010100",
  46737=>"000100101",
  46738=>"110110101",
  46739=>"000101110",
  46740=>"010000110",
  46741=>"101001111",
  46742=>"111000000",
  46743=>"110011000",
  46744=>"101000101",
  46745=>"001111101",
  46746=>"101001000",
  46747=>"011001011",
  46748=>"100110110",
  46749=>"000111111",
  46750=>"100001111",
  46751=>"111110110",
  46752=>"011111111",
  46753=>"111001000",
  46754=>"001011111",
  46755=>"100111111",
  46756=>"101010110",
  46757=>"101101101",
  46758=>"110001000",
  46759=>"001000101",
  46760=>"101011110",
  46761=>"110101111",
  46762=>"010000001",
  46763=>"110011001",
  46764=>"000011100",
  46765=>"111111001",
  46766=>"111001100",
  46767=>"100010100",
  46768=>"100100100",
  46769=>"011100101",
  46770=>"001110011",
  46771=>"001110000",
  46772=>"101100000",
  46773=>"110100111",
  46774=>"101100100",
  46775=>"111101000",
  46776=>"100100110",
  46777=>"000000000",
  46778=>"011010001",
  46779=>"001010100",
  46780=>"100011110",
  46781=>"010100011",
  46782=>"001010100",
  46783=>"011010001",
  46784=>"010000111",
  46785=>"100010110",
  46786=>"110110001",
  46787=>"001001010",
  46788=>"000100010",
  46789=>"001011000",
  46790=>"010001000",
  46791=>"000100101",
  46792=>"000000001",
  46793=>"110000000",
  46794=>"011011000",
  46795=>"100000111",
  46796=>"111101001",
  46797=>"010110111",
  46798=>"010010100",
  46799=>"111010001",
  46800=>"101111000",
  46801=>"001010000",
  46802=>"010110101",
  46803=>"100000001",
  46804=>"101010110",
  46805=>"010000010",
  46806=>"110000011",
  46807=>"111111010",
  46808=>"110110001",
  46809=>"111110110",
  46810=>"001101111",
  46811=>"000010011",
  46812=>"101011110",
  46813=>"010011111",
  46814=>"100001001",
  46815=>"010000010",
  46816=>"110011000",
  46817=>"100010110",
  46818=>"001111010",
  46819=>"110010011",
  46820=>"110010011",
  46821=>"111111110",
  46822=>"111111101",
  46823=>"111111110",
  46824=>"101100000",
  46825=>"111001010",
  46826=>"011100001",
  46827=>"010011001",
  46828=>"100101001",
  46829=>"011010101",
  46830=>"001100010",
  46831=>"000110111",
  46832=>"000110010",
  46833=>"110010011",
  46834=>"100000100",
  46835=>"001010111",
  46836=>"011011000",
  46837=>"001110010",
  46838=>"000010111",
  46839=>"111111100",
  46840=>"000010000",
  46841=>"011000111",
  46842=>"101100100",
  46843=>"110101010",
  46844=>"011100010",
  46845=>"000000001",
  46846=>"010000000",
  46847=>"001011111",
  46848=>"000111010",
  46849=>"110100111",
  46850=>"101000100",
  46851=>"011001100",
  46852=>"011010101",
  46853=>"100000000",
  46854=>"000011010",
  46855=>"001001011",
  46856=>"000101001",
  46857=>"000111000",
  46858=>"100010001",
  46859=>"011101000",
  46860=>"100011100",
  46861=>"011101111",
  46862=>"111100011",
  46863=>"010011101",
  46864=>"001100111",
  46865=>"000100000",
  46866=>"110110101",
  46867=>"011101110",
  46868=>"100101100",
  46869=>"111000000",
  46870=>"010100000",
  46871=>"010111110",
  46872=>"100000100",
  46873=>"000000101",
  46874=>"110001011",
  46875=>"000001101",
  46876=>"100000101",
  46877=>"011100011",
  46878=>"100101010",
  46879=>"100011001",
  46880=>"110111010",
  46881=>"000111111",
  46882=>"100100010",
  46883=>"100010110",
  46884=>"110100011",
  46885=>"110111101",
  46886=>"010001110",
  46887=>"101111101",
  46888=>"111100111",
  46889=>"100110010",
  46890=>"010101100",
  46891=>"100101000",
  46892=>"111010101",
  46893=>"111000100",
  46894=>"010011000",
  46895=>"000110101",
  46896=>"110110000",
  46897=>"110010111",
  46898=>"100110000",
  46899=>"010000100",
  46900=>"100010000",
  46901=>"101000001",
  46902=>"100011000",
  46903=>"001000101",
  46904=>"011000010",
  46905=>"000001001",
  46906=>"011110100",
  46907=>"011000101",
  46908=>"101111010",
  46909=>"100001101",
  46910=>"101001101",
  46911=>"100010111",
  46912=>"111101000",
  46913=>"101101000",
  46914=>"101111110",
  46915=>"010111110",
  46916=>"001100100",
  46917=>"111101111",
  46918=>"110010111",
  46919=>"000000001",
  46920=>"010100001",
  46921=>"111010111",
  46922=>"100000001",
  46923=>"010011000",
  46924=>"011110011",
  46925=>"011100011",
  46926=>"011010010",
  46927=>"101111100",
  46928=>"010101111",
  46929=>"111000001",
  46930=>"100001001",
  46931=>"000101101",
  46932=>"001001010",
  46933=>"111011111",
  46934=>"010001001",
  46935=>"011000010",
  46936=>"011011010",
  46937=>"000101010",
  46938=>"000000000",
  46939=>"110110101",
  46940=>"101011011",
  46941=>"100010001",
  46942=>"010000100",
  46943=>"000011010",
  46944=>"111011110",
  46945=>"000110010",
  46946=>"111100000",
  46947=>"011101110",
  46948=>"100110101",
  46949=>"111100000",
  46950=>"011001000",
  46951=>"101010011",
  46952=>"010001100",
  46953=>"110010000",
  46954=>"000000001",
  46955=>"110010110",
  46956=>"011010010",
  46957=>"000101100",
  46958=>"010001011",
  46959=>"001100010",
  46960=>"101010100",
  46961=>"101111000",
  46962=>"010100011",
  46963=>"001011101",
  46964=>"001100111",
  46965=>"111100000",
  46966=>"010110110",
  46967=>"011110001",
  46968=>"011111000",
  46969=>"110011110",
  46970=>"110111010",
  46971=>"111000000",
  46972=>"011001001",
  46973=>"011010001",
  46974=>"011111010",
  46975=>"101001111",
  46976=>"000000110",
  46977=>"010010011",
  46978=>"011011010",
  46979=>"111001100",
  46980=>"011010100",
  46981=>"111011110",
  46982=>"100110101",
  46983=>"101101010",
  46984=>"100000011",
  46985=>"011101100",
  46986=>"011011100",
  46987=>"000101010",
  46988=>"000001110",
  46989=>"000110111",
  46990=>"101110111",
  46991=>"111101101",
  46992=>"010010101",
  46993=>"111000000",
  46994=>"001101100",
  46995=>"010010111",
  46996=>"100000010",
  46997=>"001101100",
  46998=>"110100001",
  46999=>"111001111",
  47000=>"110101101",
  47001=>"010011111",
  47002=>"110101000",
  47003=>"011011110",
  47004=>"000010001",
  47005=>"000010011",
  47006=>"111001100",
  47007=>"100110100",
  47008=>"101101101",
  47009=>"000100100",
  47010=>"010101011",
  47011=>"111100100",
  47012=>"001000000",
  47013=>"010111011",
  47014=>"110110111",
  47015=>"101010010",
  47016=>"000011011",
  47017=>"111101101",
  47018=>"011110111",
  47019=>"101101011",
  47020=>"010011000",
  47021=>"101101100",
  47022=>"100000001",
  47023=>"101011100",
  47024=>"101111110",
  47025=>"110100010",
  47026=>"010011111",
  47027=>"101111011",
  47028=>"101110010",
  47029=>"010000100",
  47030=>"100011011",
  47031=>"001010011",
  47032=>"110101010",
  47033=>"001000011",
  47034=>"101101001",
  47035=>"010000100",
  47036=>"100111011",
  47037=>"001011110",
  47038=>"101000110",
  47039=>"010001000",
  47040=>"000010110",
  47041=>"111010101",
  47042=>"101100010",
  47043=>"101101001",
  47044=>"000111110",
  47045=>"111000010",
  47046=>"010110010",
  47047=>"011101001",
  47048=>"110010101",
  47049=>"100010110",
  47050=>"111011010",
  47051=>"010111010",
  47052=>"011011101",
  47053=>"110001111",
  47054=>"001101110",
  47055=>"110001001",
  47056=>"011010110",
  47057=>"111101010",
  47058=>"111001100",
  47059=>"001111111",
  47060=>"000010000",
  47061=>"011000000",
  47062=>"001011111",
  47063=>"101111001",
  47064=>"110000110",
  47065=>"111100101",
  47066=>"100011101",
  47067=>"001001100",
  47068=>"011011001",
  47069=>"111110011",
  47070=>"100011001",
  47071=>"011011100",
  47072=>"011101100",
  47073=>"101011101",
  47074=>"000111101",
  47075=>"000110110",
  47076=>"010111000",
  47077=>"000011010",
  47078=>"101110101",
  47079=>"110001010",
  47080=>"111001101",
  47081=>"000111100",
  47082=>"110110010",
  47083=>"001101100",
  47084=>"110001100",
  47085=>"010110101",
  47086=>"001011010",
  47087=>"010010001",
  47088=>"001011000",
  47089=>"000000011",
  47090=>"011011110",
  47091=>"100010101",
  47092=>"110100000",
  47093=>"001111101",
  47094=>"111101111",
  47095=>"011000010",
  47096=>"111111111",
  47097=>"101000111",
  47098=>"110011101",
  47099=>"111010010",
  47100=>"111001111",
  47101=>"010100010",
  47102=>"100101001",
  47103=>"110100011",
  47104=>"010111010",
  47105=>"001000110",
  47106=>"101110011",
  47107=>"111000110",
  47108=>"100100110",
  47109=>"111101100",
  47110=>"111101001",
  47111=>"011101000",
  47112=>"111101001",
  47113=>"111010111",
  47114=>"101011010",
  47115=>"111100101",
  47116=>"100000101",
  47117=>"101011100",
  47118=>"011011111",
  47119=>"101110010",
  47120=>"110111011",
  47121=>"101011010",
  47122=>"101000111",
  47123=>"111100011",
  47124=>"101100011",
  47125=>"100001101",
  47126=>"100111011",
  47127=>"001001000",
  47128=>"011111011",
  47129=>"110110110",
  47130=>"100010000",
  47131=>"001000100",
  47132=>"101101111",
  47133=>"111000011",
  47134=>"000000001",
  47135=>"010010001",
  47136=>"101100100",
  47137=>"110111110",
  47138=>"100100111",
  47139=>"000001101",
  47140=>"110001111",
  47141=>"100100101",
  47142=>"010101010",
  47143=>"010101000",
  47144=>"110011000",
  47145=>"100000101",
  47146=>"110111111",
  47147=>"110010101",
  47148=>"010011100",
  47149=>"001111110",
  47150=>"110000110",
  47151=>"100100011",
  47152=>"110010011",
  47153=>"111000000",
  47154=>"000000111",
  47155=>"010010011",
  47156=>"011011100",
  47157=>"010101101",
  47158=>"100010111",
  47159=>"111101101",
  47160=>"101101011",
  47161=>"000101000",
  47162=>"001010000",
  47163=>"001001001",
  47164=>"111110110",
  47165=>"111001001",
  47166=>"110110111",
  47167=>"001000110",
  47168=>"010000010",
  47169=>"000110101",
  47170=>"011101001",
  47171=>"101101110",
  47172=>"101001111",
  47173=>"111011100",
  47174=>"111110110",
  47175=>"001000001",
  47176=>"010110110",
  47177=>"111100100",
  47178=>"111000110",
  47179=>"110010111",
  47180=>"001001110",
  47181=>"101010111",
  47182=>"000001111",
  47183=>"000001000",
  47184=>"111110000",
  47185=>"100000000",
  47186=>"110010101",
  47187=>"100111101",
  47188=>"011011010",
  47189=>"101010000",
  47190=>"000010011",
  47191=>"001000001",
  47192=>"011010110",
  47193=>"000011000",
  47194=>"101110011",
  47195=>"000000101",
  47196=>"110111011",
  47197=>"100101111",
  47198=>"011101001",
  47199=>"011001000",
  47200=>"011111001",
  47201=>"000110000",
  47202=>"110011101",
  47203=>"000100011",
  47204=>"100101010",
  47205=>"010000010",
  47206=>"010100000",
  47207=>"001000010",
  47208=>"101001100",
  47209=>"110101001",
  47210=>"001010001",
  47211=>"000001001",
  47212=>"000110110",
  47213=>"010001001",
  47214=>"011110001",
  47215=>"110110100",
  47216=>"101011011",
  47217=>"010101101",
  47218=>"101001011",
  47219=>"011110111",
  47220=>"010101100",
  47221=>"010101110",
  47222=>"100011100",
  47223=>"101011000",
  47224=>"000011010",
  47225=>"001010011",
  47226=>"011011000",
  47227=>"010010101",
  47228=>"000101111",
  47229=>"101001011",
  47230=>"101100000",
  47231=>"010001111",
  47232=>"100111110",
  47233=>"101010001",
  47234=>"001111001",
  47235=>"000100010",
  47236=>"011011001",
  47237=>"010011110",
  47238=>"011001010",
  47239=>"000100000",
  47240=>"001010010",
  47241=>"111001101",
  47242=>"101100110",
  47243=>"011111000",
  47244=>"001001001",
  47245=>"100111111",
  47246=>"101001001",
  47247=>"111100100",
  47248=>"101101110",
  47249=>"000100111",
  47250=>"010001111",
  47251=>"000000100",
  47252=>"111110011",
  47253=>"000111111",
  47254=>"010011101",
  47255=>"110000100",
  47256=>"100001100",
  47257=>"010011001",
  47258=>"011001110",
  47259=>"110111110",
  47260=>"000110101",
  47261=>"101011010",
  47262=>"101010011",
  47263=>"101000000",
  47264=>"110001011",
  47265=>"110011011",
  47266=>"000111100",
  47267=>"100110001",
  47268=>"100011111",
  47269=>"010110010",
  47270=>"000101010",
  47271=>"010011011",
  47272=>"000100101",
  47273=>"011000110",
  47274=>"010100001",
  47275=>"111011000",
  47276=>"001110110",
  47277=>"100011000",
  47278=>"001010001",
  47279=>"010011111",
  47280=>"001001000",
  47281=>"111101001",
  47282=>"011010001",
  47283=>"110101010",
  47284=>"001111001",
  47285=>"111000000",
  47286=>"010010101",
  47287=>"000101111",
  47288=>"000000101",
  47289=>"000111011",
  47290=>"010101001",
  47291=>"011101001",
  47292=>"100011011",
  47293=>"001010011",
  47294=>"101101111",
  47295=>"110111001",
  47296=>"010101100",
  47297=>"001101000",
  47298=>"010010101",
  47299=>"011110111",
  47300=>"100100111",
  47301=>"011011010",
  47302=>"001100111",
  47303=>"001011011",
  47304=>"101010110",
  47305=>"001100111",
  47306=>"010101011",
  47307=>"001110010",
  47308=>"110110000",
  47309=>"100000101",
  47310=>"000010101",
  47311=>"001010000",
  47312=>"000111010",
  47313=>"000111110",
  47314=>"000101001",
  47315=>"111101101",
  47316=>"000011110",
  47317=>"011010111",
  47318=>"101001101",
  47319=>"100011110",
  47320=>"001110101",
  47321=>"000011101",
  47322=>"000110110",
  47323=>"000011001",
  47324=>"001000110",
  47325=>"100111100",
  47326=>"001010000",
  47327=>"101000111",
  47328=>"111110001",
  47329=>"100001111",
  47330=>"011010001",
  47331=>"011011000",
  47332=>"111111111",
  47333=>"110000111",
  47334=>"110000011",
  47335=>"101111000",
  47336=>"110001100",
  47337=>"000110001",
  47338=>"011001111",
  47339=>"001110111",
  47340=>"110110010",
  47341=>"010001101",
  47342=>"101001111",
  47343=>"000100111",
  47344=>"011000111",
  47345=>"110110111",
  47346=>"001010101",
  47347=>"000100111",
  47348=>"100000111",
  47349=>"101110000",
  47350=>"101000000",
  47351=>"000001111",
  47352=>"101101010",
  47353=>"000110110",
  47354=>"100011010",
  47355=>"000001111",
  47356=>"010001110",
  47357=>"011100001",
  47358=>"100111101",
  47359=>"010010000",
  47360=>"100000011",
  47361=>"011111011",
  47362=>"101001100",
  47363=>"011010011",
  47364=>"101101000",
  47365=>"000000100",
  47366=>"011101101",
  47367=>"111011101",
  47368=>"110111100",
  47369=>"110000000",
  47370=>"010110011",
  47371=>"001000100",
  47372=>"011011001",
  47373=>"011111101",
  47374=>"100110100",
  47375=>"000110010",
  47376=>"101110101",
  47377=>"000100010",
  47378=>"000111001",
  47379=>"111100001",
  47380=>"111000010",
  47381=>"110110010",
  47382=>"010101110",
  47383=>"100011001",
  47384=>"011011100",
  47385=>"010011111",
  47386=>"001100010",
  47387=>"100110101",
  47388=>"010101000",
  47389=>"001011111",
  47390=>"000001000",
  47391=>"100110101",
  47392=>"001111010",
  47393=>"000111010",
  47394=>"100111000",
  47395=>"001110101",
  47396=>"011100011",
  47397=>"111111001",
  47398=>"100010101",
  47399=>"101001111",
  47400=>"011111010",
  47401=>"111000010",
  47402=>"001011101",
  47403=>"111110111",
  47404=>"110101100",
  47405=>"101110010",
  47406=>"010101000",
  47407=>"101011111",
  47408=>"100101111",
  47409=>"100100001",
  47410=>"000000100",
  47411=>"011001001",
  47412=>"101000111",
  47413=>"101111111",
  47414=>"011001100",
  47415=>"111111101",
  47416=>"011010011",
  47417=>"111010001",
  47418=>"000110001",
  47419=>"010011111",
  47420=>"010101011",
  47421=>"101101101",
  47422=>"100010111",
  47423=>"010010110",
  47424=>"000110101",
  47425=>"011010001",
  47426=>"000101001",
  47427=>"110110100",
  47428=>"010101100",
  47429=>"110101001",
  47430=>"000101110",
  47431=>"011011111",
  47432=>"110111011",
  47433=>"101100100",
  47434=>"110011111",
  47435=>"101110111",
  47436=>"100101100",
  47437=>"011000101",
  47438=>"111100011",
  47439=>"111010001",
  47440=>"101011000",
  47441=>"001000000",
  47442=>"011101110",
  47443=>"001010100",
  47444=>"101101110",
  47445=>"010100110",
  47446=>"011101001",
  47447=>"100110001",
  47448=>"010110000",
  47449=>"000000000",
  47450=>"011011000",
  47451=>"111001111",
  47452=>"011011100",
  47453=>"111000101",
  47454=>"111001011",
  47455=>"000110000",
  47456=>"011110010",
  47457=>"111111001",
  47458=>"100010100",
  47459=>"010100001",
  47460=>"101001000",
  47461=>"100111010",
  47462=>"111110101",
  47463=>"111110000",
  47464=>"010001100",
  47465=>"000100010",
  47466=>"011111111",
  47467=>"110101010",
  47468=>"001101011",
  47469=>"011010001",
  47470=>"001011111",
  47471=>"100011101",
  47472=>"001000111",
  47473=>"110001010",
  47474=>"010111010",
  47475=>"110100000",
  47476=>"110111110",
  47477=>"001101000",
  47478=>"101100011",
  47479=>"001111000",
  47480=>"100100110",
  47481=>"011011001",
  47482=>"010110110",
  47483=>"011011111",
  47484=>"100011010",
  47485=>"111000101",
  47486=>"011000011",
  47487=>"100001111",
  47488=>"111101011",
  47489=>"010010100",
  47490=>"010011101",
  47491=>"000111010",
  47492=>"110111001",
  47493=>"101000000",
  47494=>"111001011",
  47495=>"000111100",
  47496=>"101111010",
  47497=>"110001111",
  47498=>"111011001",
  47499=>"000110100",
  47500=>"111100101",
  47501=>"100111011",
  47502=>"000100010",
  47503=>"111100111",
  47504=>"011001100",
  47505=>"011100111",
  47506=>"010101000",
  47507=>"011000100",
  47508=>"011010011",
  47509=>"110101011",
  47510=>"000000010",
  47511=>"111111111",
  47512=>"110100100",
  47513=>"111010111",
  47514=>"010100100",
  47515=>"010110001",
  47516=>"010011110",
  47517=>"010100000",
  47518=>"011001000",
  47519=>"000101000",
  47520=>"100101000",
  47521=>"010100001",
  47522=>"100001011",
  47523=>"101001001",
  47524=>"011010101",
  47525=>"001001000",
  47526=>"011110111",
  47527=>"111010101",
  47528=>"001100101",
  47529=>"100000000",
  47530=>"011011000",
  47531=>"101110000",
  47532=>"111001110",
  47533=>"000110001",
  47534=>"100101010",
  47535=>"000110000",
  47536=>"001011011",
  47537=>"100000110",
  47538=>"000111001",
  47539=>"001010111",
  47540=>"101111110",
  47541=>"000110101",
  47542=>"001111100",
  47543=>"110000110",
  47544=>"000101100",
  47545=>"001100100",
  47546=>"010000110",
  47547=>"010000000",
  47548=>"100001000",
  47549=>"001100001",
  47550=>"000110001",
  47551=>"011010011",
  47552=>"101000100",
  47553=>"100100000",
  47554=>"101010101",
  47555=>"000101101",
  47556=>"110010101",
  47557=>"010001110",
  47558=>"000000001",
  47559=>"111001110",
  47560=>"011001011",
  47561=>"110111001",
  47562=>"101011000",
  47563=>"110110110",
  47564=>"000111010",
  47565=>"101111001",
  47566=>"001111010",
  47567=>"100100100",
  47568=>"101101011",
  47569=>"001110111",
  47570=>"111101101",
  47571=>"011000010",
  47572=>"011100111",
  47573=>"011010010",
  47574=>"010110101",
  47575=>"110010110",
  47576=>"001001000",
  47577=>"110101010",
  47578=>"111001101",
  47579=>"101110010",
  47580=>"001001111",
  47581=>"001000111",
  47582=>"100011010",
  47583=>"011110000",
  47584=>"111110001",
  47585=>"101001011",
  47586=>"010010000",
  47587=>"111111011",
  47588=>"111000010",
  47589=>"101101011",
  47590=>"110100100",
  47591=>"011101011",
  47592=>"111111100",
  47593=>"001110011",
  47594=>"001000100",
  47595=>"000011100",
  47596=>"001100000",
  47597=>"101101111",
  47598=>"100010110",
  47599=>"110111011",
  47600=>"010110001",
  47601=>"101100000",
  47602=>"111100010",
  47603=>"101101111",
  47604=>"011100001",
  47605=>"001000000",
  47606=>"110001010",
  47607=>"010111010",
  47608=>"001011000",
  47609=>"110111100",
  47610=>"100101000",
  47611=>"010000111",
  47612=>"100100011",
  47613=>"011010001",
  47614=>"011110101",
  47615=>"110110111",
  47616=>"010011000",
  47617=>"010011100",
  47618=>"010010000",
  47619=>"101011111",
  47620=>"011000101",
  47621=>"101001101",
  47622=>"010011100",
  47623=>"011110100",
  47624=>"111001011",
  47625=>"010100001",
  47626=>"111100100",
  47627=>"000000001",
  47628=>"110100000",
  47629=>"000110100",
  47630=>"100000110",
  47631=>"101111110",
  47632=>"110000001",
  47633=>"110011111",
  47634=>"101011011",
  47635=>"101100000",
  47636=>"000010101",
  47637=>"010011011",
  47638=>"010110010",
  47639=>"010101011",
  47640=>"001111000",
  47641=>"100110000",
  47642=>"101011100",
  47643=>"101011011",
  47644=>"111011100",
  47645=>"000100101",
  47646=>"110101010",
  47647=>"011101111",
  47648=>"000101010",
  47649=>"110000101",
  47650=>"001011010",
  47651=>"101010000",
  47652=>"010001000",
  47653=>"111000000",
  47654=>"111101101",
  47655=>"010111101",
  47656=>"100000100",
  47657=>"101100101",
  47658=>"101001111",
  47659=>"001000000",
  47660=>"111111110",
  47661=>"000000001",
  47662=>"001110001",
  47663=>"011101010",
  47664=>"011001111",
  47665=>"000000111",
  47666=>"000110100",
  47667=>"000111101",
  47668=>"001101111",
  47669=>"011110010",
  47670=>"000110111",
  47671=>"110000100",
  47672=>"110101010",
  47673=>"100101010",
  47674=>"010010001",
  47675=>"000111101",
  47676=>"001101000",
  47677=>"110010000",
  47678=>"111111111",
  47679=>"101110111",
  47680=>"111111110",
  47681=>"100001011",
  47682=>"110110100",
  47683=>"011001110",
  47684=>"110000100",
  47685=>"100010010",
  47686=>"111111101",
  47687=>"011010000",
  47688=>"111010010",
  47689=>"101010000",
  47690=>"011010000",
  47691=>"000000101",
  47692=>"101011100",
  47693=>"001000010",
  47694=>"110100001",
  47695=>"100000010",
  47696=>"010110111",
  47697=>"100110111",
  47698=>"001100001",
  47699=>"000000111",
  47700=>"101111001",
  47701=>"011111110",
  47702=>"000100011",
  47703=>"111010101",
  47704=>"100011111",
  47705=>"011111010",
  47706=>"110101011",
  47707=>"111011011",
  47708=>"011000111",
  47709=>"000100101",
  47710=>"101011100",
  47711=>"111010010",
  47712=>"000010111",
  47713=>"001100000",
  47714=>"000011101",
  47715=>"100001101",
  47716=>"000100100",
  47717=>"000000110",
  47718=>"111010001",
  47719=>"010110010",
  47720=>"000111100",
  47721=>"000011010",
  47722=>"001100100",
  47723=>"001101110",
  47724=>"110110100",
  47725=>"110011101",
  47726=>"000000010",
  47727=>"110000110",
  47728=>"111100101",
  47729=>"000000001",
  47730=>"101110010",
  47731=>"000001100",
  47732=>"110000111",
  47733=>"000111110",
  47734=>"100001111",
  47735=>"101101010",
  47736=>"100010110",
  47737=>"000010101",
  47738=>"010001101",
  47739=>"000111100",
  47740=>"011111101",
  47741=>"111001101",
  47742=>"001111111",
  47743=>"101010100",
  47744=>"110010010",
  47745=>"000000000",
  47746=>"001100001",
  47747=>"100111001",
  47748=>"000111101",
  47749=>"000110001",
  47750=>"110010110",
  47751=>"010101111",
  47752=>"011000011",
  47753=>"001011011",
  47754=>"000110010",
  47755=>"000101000",
  47756=>"000110110",
  47757=>"101010000",
  47758=>"111001010",
  47759=>"000001100",
  47760=>"100100100",
  47761=>"001011001",
  47762=>"001011100",
  47763=>"011010110",
  47764=>"111010100",
  47765=>"000010000",
  47766=>"110010001",
  47767=>"000100101",
  47768=>"110101110",
  47769=>"011010100",
  47770=>"101001101",
  47771=>"111101110",
  47772=>"101011100",
  47773=>"111000111",
  47774=>"101000100",
  47775=>"000011010",
  47776=>"000101000",
  47777=>"001100011",
  47778=>"101111111",
  47779=>"010011101",
  47780=>"111100000",
  47781=>"111010011",
  47782=>"000001100",
  47783=>"000100110",
  47784=>"100011100",
  47785=>"000111000",
  47786=>"110001100",
  47787=>"111010010",
  47788=>"011110010",
  47789=>"111110011",
  47790=>"001001001",
  47791=>"011101011",
  47792=>"011111010",
  47793=>"110101000",
  47794=>"011000100",
  47795=>"000110011",
  47796=>"100100110",
  47797=>"001010111",
  47798=>"111100001",
  47799=>"000011011",
  47800=>"100111100",
  47801=>"100111010",
  47802=>"010001101",
  47803=>"010101001",
  47804=>"111010111",
  47805=>"011111101",
  47806=>"001011111",
  47807=>"100010001",
  47808=>"110001011",
  47809=>"011011111",
  47810=>"111100100",
  47811=>"111100011",
  47812=>"111101110",
  47813=>"010101011",
  47814=>"110000111",
  47815=>"011111000",
  47816=>"000000111",
  47817=>"010111110",
  47818=>"111111111",
  47819=>"001001011",
  47820=>"000100101",
  47821=>"111000111",
  47822=>"010011100",
  47823=>"000011001",
  47824=>"001010011",
  47825=>"110001011",
  47826=>"000110010",
  47827=>"000011000",
  47828=>"101010010",
  47829=>"000110100",
  47830=>"101101101",
  47831=>"101110010",
  47832=>"000100110",
  47833=>"111100000",
  47834=>"001111111",
  47835=>"111101110",
  47836=>"010001101",
  47837=>"110011100",
  47838=>"110110001",
  47839=>"010001100",
  47840=>"000000001",
  47841=>"010000101",
  47842=>"100001010",
  47843=>"000000001",
  47844=>"010010111",
  47845=>"101101100",
  47846=>"111100011",
  47847=>"111111101",
  47848=>"110101001",
  47849=>"011001001",
  47850=>"000100110",
  47851=>"010111010",
  47852=>"000001000",
  47853=>"110101010",
  47854=>"010011010",
  47855=>"000010010",
  47856=>"111011101",
  47857=>"111001011",
  47858=>"010101100",
  47859=>"001101001",
  47860=>"000010010",
  47861=>"101101111",
  47862=>"011010000",
  47863=>"001001011",
  47864=>"111111000",
  47865=>"000111111",
  47866=>"100010011",
  47867=>"100110000",
  47868=>"011111110",
  47869=>"110111110",
  47870=>"010110000",
  47871=>"111100000",
  47872=>"000011000",
  47873=>"100000001",
  47874=>"110100110",
  47875=>"111000101",
  47876=>"110011101",
  47877=>"100101110",
  47878=>"001001010",
  47879=>"001110010",
  47880=>"110101111",
  47881=>"111010001",
  47882=>"000100100",
  47883=>"000111001",
  47884=>"100110001",
  47885=>"001011000",
  47886=>"010100100",
  47887=>"001010100",
  47888=>"010001100",
  47889=>"100010011",
  47890=>"111101101",
  47891=>"100100001",
  47892=>"101001100",
  47893=>"100111011",
  47894=>"011110011",
  47895=>"011111110",
  47896=>"001101111",
  47897=>"001000000",
  47898=>"001110001",
  47899=>"000100110",
  47900=>"110000101",
  47901=>"001000101",
  47902=>"110010000",
  47903=>"111000100",
  47904=>"100101111",
  47905=>"100100011",
  47906=>"110000110",
  47907=>"001101100",
  47908=>"000001000",
  47909=>"000101100",
  47910=>"010101110",
  47911=>"010101110",
  47912=>"101100111",
  47913=>"111010001",
  47914=>"011001100",
  47915=>"100110111",
  47916=>"111000000",
  47917=>"000010001",
  47918=>"111001000",
  47919=>"111010101",
  47920=>"000001111",
  47921=>"111011001",
  47922=>"101011011",
  47923=>"111010110",
  47924=>"100000110",
  47925=>"010001000",
  47926=>"110101111",
  47927=>"100011100",
  47928=>"000001010",
  47929=>"101000000",
  47930=>"110111001",
  47931=>"011111100",
  47932=>"011100110",
  47933=>"101110101",
  47934=>"101001011",
  47935=>"001101110",
  47936=>"001100011",
  47937=>"011011011",
  47938=>"100101101",
  47939=>"011000000",
  47940=>"011011010",
  47941=>"100010111",
  47942=>"000110000",
  47943=>"111101000",
  47944=>"100110100",
  47945=>"010011001",
  47946=>"111101001",
  47947=>"101001111",
  47948=>"001001000",
  47949=>"010001110",
  47950=>"001000100",
  47951=>"101100011",
  47952=>"100010010",
  47953=>"010000000",
  47954=>"001000000",
  47955=>"110010010",
  47956=>"000111000",
  47957=>"000101101",
  47958=>"100000010",
  47959=>"100011000",
  47960=>"111110111",
  47961=>"111111011",
  47962=>"011011010",
  47963=>"101000011",
  47964=>"010011000",
  47965=>"101111111",
  47966=>"000101000",
  47967=>"000000000",
  47968=>"011011000",
  47969=>"101010100",
  47970=>"101110000",
  47971=>"001100011",
  47972=>"011110101",
  47973=>"110110010",
  47974=>"010101010",
  47975=>"001101110",
  47976=>"100010111",
  47977=>"011100110",
  47978=>"000110111",
  47979=>"001010110",
  47980=>"101100010",
  47981=>"101111000",
  47982=>"100100110",
  47983=>"001001000",
  47984=>"101111110",
  47985=>"001101010",
  47986=>"000011000",
  47987=>"010001000",
  47988=>"001110010",
  47989=>"010101010",
  47990=>"101101101",
  47991=>"110100110",
  47992=>"101101101",
  47993=>"001111111",
  47994=>"010001011",
  47995=>"001000011",
  47996=>"111101001",
  47997=>"010100100",
  47998=>"100011000",
  47999=>"100001111",
  48000=>"101111101",
  48001=>"011110101",
  48002=>"111111101",
  48003=>"111011010",
  48004=>"010110001",
  48005=>"101010000",
  48006=>"111000101",
  48007=>"111111001",
  48008=>"100010000",
  48009=>"111001111",
  48010=>"111100100",
  48011=>"001101100",
  48012=>"001111010",
  48013=>"101001111",
  48014=>"101101110",
  48015=>"111011001",
  48016=>"111100110",
  48017=>"011001000",
  48018=>"100101001",
  48019=>"000011111",
  48020=>"000010010",
  48021=>"011010011",
  48022=>"001101111",
  48023=>"110011100",
  48024=>"100001101",
  48025=>"100011001",
  48026=>"101000111",
  48027=>"100000011",
  48028=>"001101000",
  48029=>"111100000",
  48030=>"001010111",
  48031=>"100001000",
  48032=>"111100111",
  48033=>"100101111",
  48034=>"000110010",
  48035=>"001000101",
  48036=>"001101100",
  48037=>"010100101",
  48038=>"001111011",
  48039=>"110101111",
  48040=>"101011001",
  48041=>"100001011",
  48042=>"001100011",
  48043=>"101100001",
  48044=>"010001000",
  48045=>"010010011",
  48046=>"111111001",
  48047=>"010011111",
  48048=>"010000001",
  48049=>"111111100",
  48050=>"000101010",
  48051=>"100010100",
  48052=>"111110001",
  48053=>"110010011",
  48054=>"011100010",
  48055=>"010000001",
  48056=>"110101111",
  48057=>"110111110",
  48058=>"110111000",
  48059=>"000010001",
  48060=>"000101001",
  48061=>"111111111",
  48062=>"010010010",
  48063=>"100001101",
  48064=>"101101000",
  48065=>"110110001",
  48066=>"101100111",
  48067=>"001011000",
  48068=>"111100010",
  48069=>"001011010",
  48070=>"011011011",
  48071=>"111011111",
  48072=>"010101001",
  48073=>"000001111",
  48074=>"000010010",
  48075=>"111111101",
  48076=>"000101000",
  48077=>"010000100",
  48078=>"111100001",
  48079=>"110110011",
  48080=>"011111010",
  48081=>"001010001",
  48082=>"101000010",
  48083=>"110000010",
  48084=>"000101100",
  48085=>"011011100",
  48086=>"011111101",
  48087=>"110111010",
  48088=>"001011110",
  48089=>"100111110",
  48090=>"000001001",
  48091=>"000101010",
  48092=>"100101100",
  48093=>"110001100",
  48094=>"111001100",
  48095=>"111000000",
  48096=>"111011011",
  48097=>"100001101",
  48098=>"000100111",
  48099=>"111011010",
  48100=>"000011011",
  48101=>"000100011",
  48102=>"111001110",
  48103=>"101111000",
  48104=>"101100001",
  48105=>"010000111",
  48106=>"100110110",
  48107=>"010011011",
  48108=>"100011110",
  48109=>"110001000",
  48110=>"010011110",
  48111=>"000010010",
  48112=>"011011110",
  48113=>"100010011",
  48114=>"001001100",
  48115=>"000010011",
  48116=>"110001000",
  48117=>"010010000",
  48118=>"011100001",
  48119=>"000100001",
  48120=>"110001011",
  48121=>"101101111",
  48122=>"110011101",
  48123=>"010111100",
  48124=>"100000000",
  48125=>"001001000",
  48126=>"000101001",
  48127=>"011000011",
  48128=>"101111111",
  48129=>"001100101",
  48130=>"001001111",
  48131=>"001011011",
  48132=>"001100110",
  48133=>"100001010",
  48134=>"100110110",
  48135=>"111111110",
  48136=>"101101001",
  48137=>"000001110",
  48138=>"100011001",
  48139=>"110001000",
  48140=>"100000111",
  48141=>"000001100",
  48142=>"110010111",
  48143=>"111100011",
  48144=>"100001011",
  48145=>"010001100",
  48146=>"001011111",
  48147=>"010101011",
  48148=>"000010100",
  48149=>"100001111",
  48150=>"110110100",
  48151=>"001000110",
  48152=>"111000101",
  48153=>"000110101",
  48154=>"110011001",
  48155=>"101000000",
  48156=>"001000101",
  48157=>"110111101",
  48158=>"110100000",
  48159=>"111001111",
  48160=>"111111001",
  48161=>"000001011",
  48162=>"010000100",
  48163=>"100100101",
  48164=>"100111111",
  48165=>"010100000",
  48166=>"000100111",
  48167=>"101110101",
  48168=>"010110010",
  48169=>"011110100",
  48170=>"000100111",
  48171=>"000011111",
  48172=>"010100110",
  48173=>"000011101",
  48174=>"100111111",
  48175=>"110110110",
  48176=>"010011100",
  48177=>"010101000",
  48178=>"000110000",
  48179=>"101010011",
  48180=>"000101100",
  48181=>"011011011",
  48182=>"100111100",
  48183=>"111110101",
  48184=>"011001001",
  48185=>"001111001",
  48186=>"101111010",
  48187=>"100100100",
  48188=>"111010110",
  48189=>"111001011",
  48190=>"111011110",
  48191=>"001000100",
  48192=>"101100001",
  48193=>"010001010",
  48194=>"000001001",
  48195=>"110111111",
  48196=>"010000111",
  48197=>"111010001",
  48198=>"001111010",
  48199=>"111111101",
  48200=>"010110010",
  48201=>"001110101",
  48202=>"011110001",
  48203=>"101101000",
  48204=>"100011110",
  48205=>"111111111",
  48206=>"011010011",
  48207=>"001010100",
  48208=>"111010100",
  48209=>"011000000",
  48210=>"011111001",
  48211=>"111111111",
  48212=>"111111111",
  48213=>"010010011",
  48214=>"100100111",
  48215=>"101100110",
  48216=>"011011110",
  48217=>"010011000",
  48218=>"000011101",
  48219=>"000010011",
  48220=>"010000000",
  48221=>"101001101",
  48222=>"011101000",
  48223=>"100010000",
  48224=>"001101001",
  48225=>"001100001",
  48226=>"101110100",
  48227=>"000011101",
  48228=>"110001011",
  48229=>"111111010",
  48230=>"110110110",
  48231=>"001000010",
  48232=>"100101001",
  48233=>"101111001",
  48234=>"101010111",
  48235=>"000011111",
  48236=>"111111000",
  48237=>"001101000",
  48238=>"011100001",
  48239=>"001101110",
  48240=>"011011110",
  48241=>"110100100",
  48242=>"101000011",
  48243=>"100000000",
  48244=>"001000101",
  48245=>"110001011",
  48246=>"100000000",
  48247=>"111101000",
  48248=>"101000101",
  48249=>"111001001",
  48250=>"000111011",
  48251=>"110000100",
  48252=>"001010101",
  48253=>"100101101",
  48254=>"000000000",
  48255=>"000110010",
  48256=>"111111000",
  48257=>"001011011",
  48258=>"111110011",
  48259=>"011100000",
  48260=>"010111010",
  48261=>"101010110",
  48262=>"111101000",
  48263=>"100111001",
  48264=>"111000111",
  48265=>"001010011",
  48266=>"011000001",
  48267=>"000001100",
  48268=>"101101111",
  48269=>"000100100",
  48270=>"011100101",
  48271=>"000010111",
  48272=>"100100111",
  48273=>"101001111",
  48274=>"001001011",
  48275=>"110011100",
  48276=>"111001001",
  48277=>"111010011",
  48278=>"100000111",
  48279=>"101110001",
  48280=>"010000101",
  48281=>"111000111",
  48282=>"010000001",
  48283=>"101110011",
  48284=>"110110010",
  48285=>"010111000",
  48286=>"100000011",
  48287=>"101100011",
  48288=>"000000100",
  48289=>"110111011",
  48290=>"000000111",
  48291=>"111111110",
  48292=>"001010011",
  48293=>"111101100",
  48294=>"001011110",
  48295=>"001010111",
  48296=>"000100010",
  48297=>"111111011",
  48298=>"110001010",
  48299=>"010010001",
  48300=>"110101111",
  48301=>"011111111",
  48302=>"010100101",
  48303=>"110101100",
  48304=>"111110101",
  48305=>"001000001",
  48306=>"110011010",
  48307=>"000000111",
  48308=>"000010111",
  48309=>"000010001",
  48310=>"000001111",
  48311=>"100110111",
  48312=>"011001000",
  48313=>"010001111",
  48314=>"000100111",
  48315=>"001001100",
  48316=>"111011001",
  48317=>"100010011",
  48318=>"000001010",
  48319=>"111100000",
  48320=>"111000110",
  48321=>"001001111",
  48322=>"000111101",
  48323=>"000101000",
  48324=>"110100010",
  48325=>"010110011",
  48326=>"000000010",
  48327=>"110000010",
  48328=>"010001111",
  48329=>"000000111",
  48330=>"110010010",
  48331=>"111011101",
  48332=>"001001100",
  48333=>"111011101",
  48334=>"111110100",
  48335=>"011001100",
  48336=>"011001111",
  48337=>"011001011",
  48338=>"111000100",
  48339=>"101000110",
  48340=>"000110111",
  48341=>"101000010",
  48342=>"011110011",
  48343=>"000011001",
  48344=>"101100011",
  48345=>"111010010",
  48346=>"000000000",
  48347=>"010000000",
  48348=>"011100000",
  48349=>"001011011",
  48350=>"101010110",
  48351=>"110001111",
  48352=>"001000001",
  48353=>"000010010",
  48354=>"001101101",
  48355=>"101000011",
  48356=>"000010100",
  48357=>"000011000",
  48358=>"001111100",
  48359=>"100010110",
  48360=>"100100010",
  48361=>"110111011",
  48362=>"011000010",
  48363=>"100001100",
  48364=>"001011100",
  48365=>"100000111",
  48366=>"010011100",
  48367=>"010011100",
  48368=>"111001101",
  48369=>"110110001",
  48370=>"010011111",
  48371=>"111001100",
  48372=>"001110110",
  48373=>"111110100",
  48374=>"100111100",
  48375=>"010010110",
  48376=>"001001011",
  48377=>"110110110",
  48378=>"100100000",
  48379=>"110011000",
  48380=>"101111111",
  48381=>"010010101",
  48382=>"111010110",
  48383=>"000101111",
  48384=>"010011101",
  48385=>"111010010",
  48386=>"111100010",
  48387=>"000111101",
  48388=>"111111000",
  48389=>"101110110",
  48390=>"100001011",
  48391=>"111011100",
  48392=>"000010010",
  48393=>"010100110",
  48394=>"010111011",
  48395=>"111110100",
  48396=>"011011001",
  48397=>"010100111",
  48398=>"101001010",
  48399=>"010111101",
  48400=>"010010110",
  48401=>"101100110",
  48402=>"110111111",
  48403=>"100010110",
  48404=>"101100100",
  48405=>"111001000",
  48406=>"100111000",
  48407=>"101110110",
  48408=>"100000000",
  48409=>"111111101",
  48410=>"011101000",
  48411=>"100101101",
  48412=>"000111100",
  48413=>"101010101",
  48414=>"110010000",
  48415=>"101000111",
  48416=>"010000001",
  48417=>"000111101",
  48418=>"010001010",
  48419=>"101011000",
  48420=>"101001101",
  48421=>"101001111",
  48422=>"011010111",
  48423=>"101110001",
  48424=>"011100100",
  48425=>"011011111",
  48426=>"110110100",
  48427=>"110110101",
  48428=>"101101100",
  48429=>"111011000",
  48430=>"001100110",
  48431=>"010001000",
  48432=>"000111010",
  48433=>"000011001",
  48434=>"111111010",
  48435=>"110111110",
  48436=>"011011101",
  48437=>"000110101",
  48438=>"110110011",
  48439=>"100000010",
  48440=>"010111111",
  48441=>"010101101",
  48442=>"100101100",
  48443=>"000001101",
  48444=>"110010001",
  48445=>"001101010",
  48446=>"110011000",
  48447=>"010001001",
  48448=>"010011111",
  48449=>"011110010",
  48450=>"100110101",
  48451=>"100111011",
  48452=>"000100110",
  48453=>"110110011",
  48454=>"011100001",
  48455=>"101000000",
  48456=>"000111111",
  48457=>"011100001",
  48458=>"101100011",
  48459=>"110100110",
  48460=>"111111011",
  48461=>"000100110",
  48462=>"000010010",
  48463=>"110100101",
  48464=>"111111100",
  48465=>"010100100",
  48466=>"110011110",
  48467=>"000100110",
  48468=>"011110101",
  48469=>"010010101",
  48470=>"110011011",
  48471=>"111100010",
  48472=>"100001111",
  48473=>"101001101",
  48474=>"101000000",
  48475=>"011000000",
  48476=>"101011001",
  48477=>"100111001",
  48478=>"000001011",
  48479=>"100001011",
  48480=>"010110111",
  48481=>"110111111",
  48482=>"011101010",
  48483=>"000100101",
  48484=>"001010000",
  48485=>"111000010",
  48486=>"000001001",
  48487=>"011001101",
  48488=>"000000110",
  48489=>"110000111",
  48490=>"001001111",
  48491=>"111010110",
  48492=>"111110101",
  48493=>"011111110",
  48494=>"001010001",
  48495=>"111100001",
  48496=>"100100000",
  48497=>"001010000",
  48498=>"110101010",
  48499=>"111101110",
  48500=>"110010000",
  48501=>"010001001",
  48502=>"001100000",
  48503=>"101110000",
  48504=>"001101111",
  48505=>"101000011",
  48506=>"010010010",
  48507=>"110001010",
  48508=>"111001010",
  48509=>"100010011",
  48510=>"000110000",
  48511=>"101111000",
  48512=>"000100011",
  48513=>"001011101",
  48514=>"111101111",
  48515=>"011000011",
  48516=>"110101001",
  48517=>"000111110",
  48518=>"000000011",
  48519=>"000010100",
  48520=>"011011011",
  48521=>"000000011",
  48522=>"111001001",
  48523=>"100011011",
  48524=>"110010000",
  48525=>"100111011",
  48526=>"110100010",
  48527=>"111111100",
  48528=>"010110100",
  48529=>"100001000",
  48530=>"001011011",
  48531=>"011111001",
  48532=>"101010000",
  48533=>"001000000",
  48534=>"010101101",
  48535=>"101001101",
  48536=>"000101011",
  48537=>"100110100",
  48538=>"010101001",
  48539=>"100000111",
  48540=>"101110001",
  48541=>"001001000",
  48542=>"011011000",
  48543=>"100010001",
  48544=>"100011010",
  48545=>"100101000",
  48546=>"010000010",
  48547=>"001110101",
  48548=>"000101001",
  48549=>"110011110",
  48550=>"011000000",
  48551=>"000000101",
  48552=>"100001110",
  48553=>"000111111",
  48554=>"101100011",
  48555=>"100011011",
  48556=>"000011010",
  48557=>"101100111",
  48558=>"100010000",
  48559=>"111100111",
  48560=>"001110000",
  48561=>"000000000",
  48562=>"000000011",
  48563=>"111011100",
  48564=>"100000110",
  48565=>"011010111",
  48566=>"000100111",
  48567=>"000101111",
  48568=>"001100100",
  48569=>"000100011",
  48570=>"110111011",
  48571=>"110110000",
  48572=>"001001101",
  48573=>"101000001",
  48574=>"111110111",
  48575=>"000111010",
  48576=>"000011000",
  48577=>"110111000",
  48578=>"110110011",
  48579=>"111100000",
  48580=>"100011110",
  48581=>"000110000",
  48582=>"100000110",
  48583=>"111101000",
  48584=>"100010001",
  48585=>"010100000",
  48586=>"100000100",
  48587=>"101000010",
  48588=>"101010000",
  48589=>"101011010",
  48590=>"010111010",
  48591=>"101111001",
  48592=>"111100100",
  48593=>"000100011",
  48594=>"010010100",
  48595=>"110000001",
  48596=>"011111000",
  48597=>"000110111",
  48598=>"010001111",
  48599=>"111001010",
  48600=>"111001110",
  48601=>"110111100",
  48602=>"000011000",
  48603=>"001011001",
  48604=>"111111011",
  48605=>"101010101",
  48606=>"110010000",
  48607=>"010000100",
  48608=>"001100110",
  48609=>"100000101",
  48610=>"110110011",
  48611=>"110101101",
  48612=>"110111000",
  48613=>"111011111",
  48614=>"001011001",
  48615=>"110110011",
  48616=>"000110001",
  48617=>"011111111",
  48618=>"001001000",
  48619=>"100111100",
  48620=>"000110011",
  48621=>"111011010",
  48622=>"101010101",
  48623=>"010001101",
  48624=>"111100111",
  48625=>"111110111",
  48626=>"100001110",
  48627=>"110011010",
  48628=>"001011000",
  48629=>"011110000",
  48630=>"001011110",
  48631=>"110000001",
  48632=>"100101100",
  48633=>"011011001",
  48634=>"011011001",
  48635=>"100010010",
  48636=>"111010001",
  48637=>"001101010",
  48638=>"001001011",
  48639=>"101100000",
  48640=>"010011011",
  48641=>"111000010",
  48642=>"001001100",
  48643=>"011001111",
  48644=>"110000011",
  48645=>"010010111",
  48646=>"011111101",
  48647=>"101010111",
  48648=>"111010001",
  48649=>"101011110",
  48650=>"001001100",
  48651=>"000110010",
  48652=>"000000010",
  48653=>"101100110",
  48654=>"111010111",
  48655=>"110001110",
  48656=>"011100001",
  48657=>"111111001",
  48658=>"000110100",
  48659=>"011000011",
  48660=>"100100101",
  48661=>"010100100",
  48662=>"010000111",
  48663=>"100010011",
  48664=>"100000100",
  48665=>"001101001",
  48666=>"100110110",
  48667=>"000001000",
  48668=>"100101101",
  48669=>"111111101",
  48670=>"011001101",
  48671=>"011001100",
  48672=>"010010000",
  48673=>"100000100",
  48674=>"110100001",
  48675=>"100110100",
  48676=>"001111001",
  48677=>"000001111",
  48678=>"000011010",
  48679=>"101011101",
  48680=>"101010010",
  48681=>"010000101",
  48682=>"101000101",
  48683=>"100010000",
  48684=>"010111101",
  48685=>"110111011",
  48686=>"000011000",
  48687=>"001111101",
  48688=>"011100100",
  48689=>"001111011",
  48690=>"011000011",
  48691=>"100000100",
  48692=>"010000010",
  48693=>"101111111",
  48694=>"100111100",
  48695=>"001100101",
  48696=>"001001110",
  48697=>"000100001",
  48698=>"101010001",
  48699=>"111011111",
  48700=>"011011010",
  48701=>"000000000",
  48702=>"000101101",
  48703=>"011010011",
  48704=>"000111110",
  48705=>"001010110",
  48706=>"101000100",
  48707=>"000010001",
  48708=>"101110111",
  48709=>"110100111",
  48710=>"111111110",
  48711=>"000111100",
  48712=>"110001001",
  48713=>"110111000",
  48714=>"000101000",
  48715=>"011111100",
  48716=>"010000110",
  48717=>"000110111",
  48718=>"010100101",
  48719=>"011101100",
  48720=>"011010100",
  48721=>"001000001",
  48722=>"101011001",
  48723=>"110001100",
  48724=>"001011101",
  48725=>"010000011",
  48726=>"101111100",
  48727=>"100001111",
  48728=>"101000011",
  48729=>"111100000",
  48730=>"101110011",
  48731=>"111000101",
  48732=>"010000101",
  48733=>"011101111",
  48734=>"101110000",
  48735=>"100000000",
  48736=>"101001100",
  48737=>"110010101",
  48738=>"010010111",
  48739=>"100010111",
  48740=>"111101110",
  48741=>"110111001",
  48742=>"011101001",
  48743=>"000010001",
  48744=>"001111111",
  48745=>"101111111",
  48746=>"011000101",
  48747=>"000101110",
  48748=>"111000001",
  48749=>"110000001",
  48750=>"001000000",
  48751=>"010001110",
  48752=>"011100010",
  48753=>"011110110",
  48754=>"100010010",
  48755=>"010011011",
  48756=>"011110110",
  48757=>"110100011",
  48758=>"001100111",
  48759=>"010001101",
  48760=>"010011010",
  48761=>"111101110",
  48762=>"011101111",
  48763=>"101001110",
  48764=>"100011011",
  48765=>"101000000",
  48766=>"101100001",
  48767=>"100001001",
  48768=>"100001010",
  48769=>"001000000",
  48770=>"011000110",
  48771=>"011011110",
  48772=>"111001011",
  48773=>"011001000",
  48774=>"001111000",
  48775=>"011101011",
  48776=>"110111100",
  48777=>"000011000",
  48778=>"011010011",
  48779=>"100010100",
  48780=>"001110001",
  48781=>"100001011",
  48782=>"111011101",
  48783=>"010000101",
  48784=>"100110101",
  48785=>"011100111",
  48786=>"111010101",
  48787=>"111110100",
  48788=>"010011110",
  48789=>"101101100",
  48790=>"000100111",
  48791=>"110101001",
  48792=>"111110100",
  48793=>"001001101",
  48794=>"001011011",
  48795=>"010110110",
  48796=>"100001010",
  48797=>"100110010",
  48798=>"110000001",
  48799=>"110111111",
  48800=>"011110000",
  48801=>"101001111",
  48802=>"101111010",
  48803=>"101111101",
  48804=>"101100100",
  48805=>"011010001",
  48806=>"110000001",
  48807=>"111010011",
  48808=>"011101100",
  48809=>"110000011",
  48810=>"111111101",
  48811=>"000010000",
  48812=>"111111010",
  48813=>"001001100",
  48814=>"100000110",
  48815=>"010000101",
  48816=>"011110011",
  48817=>"101011100",
  48818=>"001000100",
  48819=>"000111011",
  48820=>"000010000",
  48821=>"011011001",
  48822=>"100101010",
  48823=>"110000010",
  48824=>"111101010",
  48825=>"010011111",
  48826=>"011110010",
  48827=>"101011111",
  48828=>"000001100",
  48829=>"011111110",
  48830=>"111101111",
  48831=>"110010100",
  48832=>"001110110",
  48833=>"101111011",
  48834=>"000100111",
  48835=>"000100010",
  48836=>"001100001",
  48837=>"111100011",
  48838=>"110011111",
  48839=>"111101110",
  48840=>"110110111",
  48841=>"100010100",
  48842=>"101011111",
  48843=>"000000111",
  48844=>"001101001",
  48845=>"110111100",
  48846=>"011101001",
  48847=>"010001110",
  48848=>"101110101",
  48849=>"010111011",
  48850=>"110111011",
  48851=>"111110001",
  48852=>"001000010",
  48853=>"111101100",
  48854=>"101100110",
  48855=>"100101101",
  48856=>"100000010",
  48857=>"101001110",
  48858=>"010000110",
  48859=>"001011100",
  48860=>"101111001",
  48861=>"001010011",
  48862=>"110110001",
  48863=>"010011000",
  48864=>"111111011",
  48865=>"101011100",
  48866=>"010100010",
  48867=>"111010001",
  48868=>"011011001",
  48869=>"100000110",
  48870=>"100110101",
  48871=>"100100010",
  48872=>"010101110",
  48873=>"110010010",
  48874=>"101111110",
  48875=>"111000111",
  48876=>"111011110",
  48877=>"101110011",
  48878=>"100000100",
  48879=>"010001100",
  48880=>"000111110",
  48881=>"111110010",
  48882=>"001110010",
  48883=>"000100011",
  48884=>"000001010",
  48885=>"100100100",
  48886=>"001001101",
  48887=>"101110000",
  48888=>"110100101",
  48889=>"010011011",
  48890=>"101100110",
  48891=>"111010100",
  48892=>"011011101",
  48893=>"000101101",
  48894=>"111001001",
  48895=>"110001011",
  48896=>"000001000",
  48897=>"000101101",
  48898=>"111010001",
  48899=>"000101000",
  48900=>"111001110",
  48901=>"110000100",
  48902=>"000101001",
  48903=>"010000010",
  48904=>"100001000",
  48905=>"010111110",
  48906=>"111111000",
  48907=>"000100001",
  48908=>"110001010",
  48909=>"110101101",
  48910=>"000100101",
  48911=>"000001001",
  48912=>"010100110",
  48913=>"001011000",
  48914=>"001111111",
  48915=>"101001111",
  48916=>"000101011",
  48917=>"100010101",
  48918=>"101011101",
  48919=>"001100000",
  48920=>"010110100",
  48921=>"010111010",
  48922=>"101101001",
  48923=>"000100100",
  48924=>"000100001",
  48925=>"111101001",
  48926=>"000010111",
  48927=>"111000010",
  48928=>"110110011",
  48929=>"111100001",
  48930=>"011110110",
  48931=>"101111111",
  48932=>"011011101",
  48933=>"100101000",
  48934=>"010011000",
  48935=>"010100110",
  48936=>"100011000",
  48937=>"000100111",
  48938=>"010100000",
  48939=>"100110011",
  48940=>"000000001",
  48941=>"101010101",
  48942=>"000001010",
  48943=>"000001000",
  48944=>"110101010",
  48945=>"010101101",
  48946=>"101111011",
  48947=>"101111101",
  48948=>"110101000",
  48949=>"111111010",
  48950=>"110111111",
  48951=>"111000101",
  48952=>"101011101",
  48953=>"001000111",
  48954=>"010000111",
  48955=>"001111101",
  48956=>"111000010",
  48957=>"101000100",
  48958=>"000100100",
  48959=>"000000000",
  48960=>"010100111",
  48961=>"101010010",
  48962=>"011100010",
  48963=>"011101111",
  48964=>"100111110",
  48965=>"010001111",
  48966=>"110101111",
  48967=>"001101000",
  48968=>"011010101",
  48969=>"010000000",
  48970=>"101100000",
  48971=>"000100100",
  48972=>"010000001",
  48973=>"110100011",
  48974=>"110000100",
  48975=>"000010010",
  48976=>"001000011",
  48977=>"111000001",
  48978=>"100000010",
  48979=>"110001100",
  48980=>"000111001",
  48981=>"110000110",
  48982=>"001100100",
  48983=>"101111101",
  48984=>"100001110",
  48985=>"000111001",
  48986=>"001001100",
  48987=>"111111010",
  48988=>"011010110",
  48989=>"011101010",
  48990=>"110000111",
  48991=>"000101010",
  48992=>"110000100",
  48993=>"000100101",
  48994=>"110000001",
  48995=>"011110011",
  48996=>"001110000",
  48997=>"000110000",
  48998=>"101110111",
  48999=>"110100010",
  49000=>"010000111",
  49001=>"101010100",
  49002=>"000111100",
  49003=>"101011101",
  49004=>"011101111",
  49005=>"010100100",
  49006=>"100100100",
  49007=>"010001101",
  49008=>"111100100",
  49009=>"000111111",
  49010=>"010000000",
  49011=>"001100111",
  49012=>"100011111",
  49013=>"001001111",
  49014=>"101010100",
  49015=>"011100111",
  49016=>"001001111",
  49017=>"001111000",
  49018=>"111100110",
  49019=>"001011110",
  49020=>"000010000",
  49021=>"110001001",
  49022=>"111110010",
  49023=>"010101111",
  49024=>"000010001",
  49025=>"011001111",
  49026=>"000010111",
  49027=>"011000000",
  49028=>"111010110",
  49029=>"110001001",
  49030=>"110001110",
  49031=>"111101010",
  49032=>"111000000",
  49033=>"001101100",
  49034=>"001111110",
  49035=>"101011111",
  49036=>"100000110",
  49037=>"111101001",
  49038=>"001111111",
  49039=>"000100001",
  49040=>"010110000",
  49041=>"010000110",
  49042=>"001000000",
  49043=>"100110011",
  49044=>"011001111",
  49045=>"110000100",
  49046=>"110110100",
  49047=>"001111110",
  49048=>"001110010",
  49049=>"000100011",
  49050=>"010111100",
  49051=>"000000101",
  49052=>"000110110",
  49053=>"000000110",
  49054=>"000100111",
  49055=>"010010000",
  49056=>"101000111",
  49057=>"100111000",
  49058=>"101111111",
  49059=>"100010000",
  49060=>"001100010",
  49061=>"101010110",
  49062=>"100000000",
  49063=>"000011000",
  49064=>"100000010",
  49065=>"101101101",
  49066=>"101010000",
  49067=>"001011001",
  49068=>"001111010",
  49069=>"010100100",
  49070=>"011010001",
  49071=>"000001111",
  49072=>"100101000",
  49073=>"111000010",
  49074=>"010011001",
  49075=>"101001010",
  49076=>"000010111",
  49077=>"000100000",
  49078=>"000101101",
  49079=>"011101000",
  49080=>"110010001",
  49081=>"111010100",
  49082=>"100010010",
  49083=>"111010001",
  49084=>"100001011",
  49085=>"000100100",
  49086=>"101001101",
  49087=>"010010111",
  49088=>"111111101",
  49089=>"011111010",
  49090=>"111001110",
  49091=>"010001110",
  49092=>"110010101",
  49093=>"101011100",
  49094=>"011111110",
  49095=>"110101011",
  49096=>"011000010",
  49097=>"111100110",
  49098=>"110001101",
  49099=>"011010011",
  49100=>"000001111",
  49101=>"011000110",
  49102=>"001010011",
  49103=>"111001000",
  49104=>"000001111",
  49105=>"100010111",
  49106=>"011000111",
  49107=>"100000000",
  49108=>"110011111",
  49109=>"010111100",
  49110=>"001001000",
  49111=>"101000001",
  49112=>"101000100",
  49113=>"111111111",
  49114=>"001111111",
  49115=>"111011001",
  49116=>"101011110",
  49117=>"111001011",
  49118=>"000010100",
  49119=>"100010000",
  49120=>"100111101",
  49121=>"010101001",
  49122=>"001111001",
  49123=>"000100110",
  49124=>"011000000",
  49125=>"000110001",
  49126=>"000010000",
  49127=>"100110100",
  49128=>"000100100",
  49129=>"110101100",
  49130=>"001100010",
  49131=>"000001100",
  49132=>"001101111",
  49133=>"011000010",
  49134=>"100010000",
  49135=>"000101011",
  49136=>"111010010",
  49137=>"000001100",
  49138=>"011011111",
  49139=>"010111010",
  49140=>"011100110",
  49141=>"000000001",
  49142=>"110000011",
  49143=>"100000011",
  49144=>"001010100",
  49145=>"100100100",
  49146=>"111110101",
  49147=>"000011011",
  49148=>"011000011",
  49149=>"010010101",
  49150=>"001100111",
  49151=>"010100101",
  49152=>"101101110",
  49153=>"001111100",
  49154=>"011110011",
  49155=>"001010111",
  49156=>"100001100",
  49157=>"000101001",
  49158=>"111111111",
  49159=>"111000111",
  49160=>"110101111",
  49161=>"110110000",
  49162=>"111011000",
  49163=>"111000110",
  49164=>"010011000",
  49165=>"100010111",
  49166=>"001000011",
  49167=>"111111010",
  49168=>"100011010",
  49169=>"100011101",
  49170=>"000011111",
  49171=>"010010100",
  49172=>"111011111",
  49173=>"001111011",
  49174=>"010000010",
  49175=>"011110011",
  49176=>"111100001",
  49177=>"001011110",
  49178=>"000010101",
  49179=>"000100011",
  49180=>"101000010",
  49181=>"010010101",
  49182=>"110000100",
  49183=>"110001011",
  49184=>"100100111",
  49185=>"010000110",
  49186=>"110001110",
  49187=>"101111010",
  49188=>"010001011",
  49189=>"000100110",
  49190=>"101100010",
  49191=>"010101010",
  49192=>"001010110",
  49193=>"001001011",
  49194=>"100100111",
  49195=>"000111111",
  49196=>"110101111",
  49197=>"011101010",
  49198=>"100111011",
  49199=>"100110110",
  49200=>"101001011",
  49201=>"011110100",
  49202=>"101000110",
  49203=>"001000001",
  49204=>"100101100",
  49205=>"101001011",
  49206=>"011010001",
  49207=>"000000000",
  49208=>"001110000",
  49209=>"101100100",
  49210=>"100100010",
  49211=>"011100000",
  49212=>"101100101",
  49213=>"011110010",
  49214=>"110110000",
  49215=>"001011011",
  49216=>"010101010",
  49217=>"001010000",
  49218=>"010110000",
  49219=>"101100101",
  49220=>"100110110",
  49221=>"001010101",
  49222=>"111101100",
  49223=>"011101101",
  49224=>"011101111",
  49225=>"111010110",
  49226=>"100000101",
  49227=>"001001111",
  49228=>"100000110",
  49229=>"101000100",
  49230=>"111011010",
  49231=>"110001100",
  49232=>"001000100",
  49233=>"000001010",
  49234=>"011000011",
  49235=>"001000100",
  49236=>"111011100",
  49237=>"000000011",
  49238=>"100001001",
  49239=>"011010011",
  49240=>"011010111",
  49241=>"011001101",
  49242=>"010011101",
  49243=>"111000010",
  49244=>"100110101",
  49245=>"011011010",
  49246=>"001001110",
  49247=>"001000011",
  49248=>"011110000",
  49249=>"011100100",
  49250=>"001100010",
  49251=>"010001011",
  49252=>"011000011",
  49253=>"011100101",
  49254=>"110100111",
  49255=>"111100111",
  49256=>"010111101",
  49257=>"111000101",
  49258=>"001110111",
  49259=>"110011000",
  49260=>"010110001",
  49261=>"100000101",
  49262=>"010000011",
  49263=>"000100000",
  49264=>"010101111",
  49265=>"110111100",
  49266=>"110001110",
  49267=>"010100001",
  49268=>"101111110",
  49269=>"101010101",
  49270=>"010010011",
  49271=>"011111010",
  49272=>"111001011",
  49273=>"101000001",
  49274=>"101010101",
  49275=>"000111000",
  49276=>"101011100",
  49277=>"010000000",
  49278=>"111001111",
  49279=>"001010000",
  49280=>"100000100",
  49281=>"001100000",
  49282=>"100011101",
  49283=>"011000010",
  49284=>"101000000",
  49285=>"110100110",
  49286=>"101000000",
  49287=>"011110101",
  49288=>"100111111",
  49289=>"110001111",
  49290=>"110000011",
  49291=>"001111011",
  49292=>"100100011",
  49293=>"000000101",
  49294=>"001110111",
  49295=>"011000101",
  49296=>"000111000",
  49297=>"100101000",
  49298=>"011000100",
  49299=>"100000000",
  49300=>"111010100",
  49301=>"001111111",
  49302=>"010000000",
  49303=>"010101111",
  49304=>"100011011",
  49305=>"111010000",
  49306=>"110010101",
  49307=>"111110000",
  49308=>"001110011",
  49309=>"000111011",
  49310=>"001111110",
  49311=>"000001101",
  49312=>"011011001",
  49313=>"110011111",
  49314=>"111111001",
  49315=>"100000000",
  49316=>"001000111",
  49317=>"001011111",
  49318=>"001101111",
  49319=>"010100001",
  49320=>"011000101",
  49321=>"111011000",
  49322=>"011011001",
  49323=>"110010000",
  49324=>"001011100",
  49325=>"101000100",
  49326=>"011001101",
  49327=>"001011011",
  49328=>"111111110",
  49329=>"010001010",
  49330=>"000101011",
  49331=>"001111111",
  49332=>"010110001",
  49333=>"010010010",
  49334=>"100110010",
  49335=>"100011100",
  49336=>"011110000",
  49337=>"110100000",
  49338=>"010000111",
  49339=>"011100100",
  49340=>"000100100",
  49341=>"100001100",
  49342=>"011101011",
  49343=>"000111001",
  49344=>"011101110",
  49345=>"100110100",
  49346=>"100011000",
  49347=>"101010001",
  49348=>"000110100",
  49349=>"010011100",
  49350=>"101000111",
  49351=>"000100010",
  49352=>"111100010",
  49353=>"000101001",
  49354=>"110010111",
  49355=>"111011001",
  49356=>"110111001",
  49357=>"011001111",
  49358=>"010000101",
  49359=>"000101001",
  49360=>"100011000",
  49361=>"111010100",
  49362=>"100010010",
  49363=>"111011110",
  49364=>"000010010",
  49365=>"000001111",
  49366=>"101011100",
  49367=>"010100001",
  49368=>"011110100",
  49369=>"111110010",
  49370=>"100000111",
  49371=>"100111101",
  49372=>"101011001",
  49373=>"011000010",
  49374=>"000000111",
  49375=>"000000011",
  49376=>"110001000",
  49377=>"000101111",
  49378=>"010101000",
  49379=>"001011101",
  49380=>"000110100",
  49381=>"000100001",
  49382=>"100100111",
  49383=>"001000011",
  49384=>"110100010",
  49385=>"001100111",
  49386=>"000010001",
  49387=>"001011011",
  49388=>"111011001",
  49389=>"001010000",
  49390=>"111100100",
  49391=>"011100111",
  49392=>"110101011",
  49393=>"101000001",
  49394=>"011010110",
  49395=>"000001001",
  49396=>"010110100",
  49397=>"101000001",
  49398=>"101010010",
  49399=>"000111010",
  49400=>"000100000",
  49401=>"011000001",
  49402=>"100101001",
  49403=>"100101001",
  49404=>"110001000",
  49405=>"011011010",
  49406=>"110000100",
  49407=>"011011101",
  49408=>"110100111",
  49409=>"010010101",
  49410=>"000110000",
  49411=>"010000000",
  49412=>"010010100",
  49413=>"100101010",
  49414=>"001110011",
  49415=>"011100011",
  49416=>"111111110",
  49417=>"111101010",
  49418=>"101001000",
  49419=>"001101001",
  49420=>"101110011",
  49421=>"001111101",
  49422=>"101110110",
  49423=>"000101010",
  49424=>"110110001",
  49425=>"000010000",
  49426=>"000111100",
  49427=>"001010110",
  49428=>"110101100",
  49429=>"101000001",
  49430=>"000001010",
  49431=>"001011101",
  49432=>"110010100",
  49433=>"011101011",
  49434=>"111001010",
  49435=>"011001001",
  49436=>"001110001",
  49437=>"010000110",
  49438=>"010111010",
  49439=>"101101000",
  49440=>"111000011",
  49441=>"100110100",
  49442=>"110100010",
  49443=>"010101000",
  49444=>"010100000",
  49445=>"101110110",
  49446=>"000111111",
  49447=>"000111110",
  49448=>"000110100",
  49449=>"100111000",
  49450=>"111010010",
  49451=>"111100011",
  49452=>"100001101",
  49453=>"001111001",
  49454=>"111001010",
  49455=>"010010010",
  49456=>"100111000",
  49457=>"101010100",
  49458=>"101111110",
  49459=>"110111010",
  49460=>"100101011",
  49461=>"000100000",
  49462=>"011101000",
  49463=>"000111111",
  49464=>"101111010",
  49465=>"001010011",
  49466=>"111011001",
  49467=>"001011111",
  49468=>"001000111",
  49469=>"010110000",
  49470=>"010010010",
  49471=>"010101010",
  49472=>"111011100",
  49473=>"111011000",
  49474=>"010110001",
  49475=>"100111100",
  49476=>"010111110",
  49477=>"000010111",
  49478=>"010100100",
  49479=>"010110110",
  49480=>"011100001",
  49481=>"010010101",
  49482=>"010001011",
  49483=>"000110110",
  49484=>"111100000",
  49485=>"101000000",
  49486=>"010111100",
  49487=>"111011111",
  49488=>"010010001",
  49489=>"011100100",
  49490=>"010100000",
  49491=>"101100100",
  49492=>"010101001",
  49493=>"100101000",
  49494=>"000111001",
  49495=>"010100011",
  49496=>"111001111",
  49497=>"011100011",
  49498=>"110110010",
  49499=>"011110101",
  49500=>"010100110",
  49501=>"000100111",
  49502=>"000010101",
  49503=>"011111011",
  49504=>"011011110",
  49505=>"111110110",
  49506=>"000011011",
  49507=>"111110010",
  49508=>"000000010",
  49509=>"101100000",
  49510=>"100110000",
  49511=>"111100000",
  49512=>"111100100",
  49513=>"001001110",
  49514=>"000010000",
  49515=>"111101101",
  49516=>"111001110",
  49517=>"111110101",
  49518=>"100111000",
  49519=>"100010001",
  49520=>"000011010",
  49521=>"010001000",
  49522=>"001001110",
  49523=>"001111010",
  49524=>"100001001",
  49525=>"010001010",
  49526=>"110100011",
  49527=>"001001000",
  49528=>"110110100",
  49529=>"100110100",
  49530=>"000000110",
  49531=>"010000101",
  49532=>"000101010",
  49533=>"010010011",
  49534=>"110110001",
  49535=>"000000101",
  49536=>"000010010",
  49537=>"000011001",
  49538=>"111011010",
  49539=>"100011000",
  49540=>"110100101",
  49541=>"110001000",
  49542=>"000111110",
  49543=>"101000010",
  49544=>"110001101",
  49545=>"000110100",
  49546=>"000011111",
  49547=>"001011100",
  49548=>"100111100",
  49549=>"000001000",
  49550=>"100100111",
  49551=>"010100111",
  49552=>"001111100",
  49553=>"011000001",
  49554=>"111010110",
  49555=>"101000011",
  49556=>"011100110",
  49557=>"000001001",
  49558=>"000001111",
  49559=>"111111001",
  49560=>"101111111",
  49561=>"111010010",
  49562=>"111111111",
  49563=>"101010110",
  49564=>"101100111",
  49565=>"001011000",
  49566=>"111010000",
  49567=>"111111100",
  49568=>"100100101",
  49569=>"111110001",
  49570=>"000000000",
  49571=>"011001001",
  49572=>"000011001",
  49573=>"101011100",
  49574=>"100001000",
  49575=>"110110101",
  49576=>"001000100",
  49577=>"110110100",
  49578=>"111101111",
  49579=>"111100101",
  49580=>"000000001",
  49581=>"001000010",
  49582=>"001100101",
  49583=>"010110111",
  49584=>"101101110",
  49585=>"100100101",
  49586=>"010101011",
  49587=>"001001100",
  49588=>"110100111",
  49589=>"011010011",
  49590=>"000000111",
  49591=>"101000011",
  49592=>"111001101",
  49593=>"010000001",
  49594=>"101101101",
  49595=>"100111000",
  49596=>"101011111",
  49597=>"010010100",
  49598=>"101001011",
  49599=>"001001100",
  49600=>"001101000",
  49601=>"001101000",
  49602=>"110110100",
  49603=>"010101101",
  49604=>"000010000",
  49605=>"101100110",
  49606=>"100000100",
  49607=>"101001101",
  49608=>"101110100",
  49609=>"111110110",
  49610=>"011101010",
  49611=>"011110011",
  49612=>"101111100",
  49613=>"100011100",
  49614=>"100111111",
  49615=>"100010001",
  49616=>"100111100",
  49617=>"110001000",
  49618=>"100010100",
  49619=>"101111011",
  49620=>"111010110",
  49621=>"010101110",
  49622=>"001011101",
  49623=>"000010110",
  49624=>"010111110",
  49625=>"000100010",
  49626=>"000010111",
  49627=>"110101111",
  49628=>"111101101",
  49629=>"000110100",
  49630=>"110110100",
  49631=>"110101000",
  49632=>"000011101",
  49633=>"001000111",
  49634=>"110011110",
  49635=>"001101111",
  49636=>"100100011",
  49637=>"100100111",
  49638=>"100000101",
  49639=>"110110100",
  49640=>"100011110",
  49641=>"001001101",
  49642=>"001011000",
  49643=>"110111000",
  49644=>"110111101",
  49645=>"111101001",
  49646=>"100000000",
  49647=>"100010111",
  49648=>"001111110",
  49649=>"100101101",
  49650=>"110110010",
  49651=>"001000000",
  49652=>"000010001",
  49653=>"000011010",
  49654=>"011000001",
  49655=>"110010010",
  49656=>"101001001",
  49657=>"110010000",
  49658=>"001000000",
  49659=>"110001111",
  49660=>"111011111",
  49661=>"101011010",
  49662=>"111001111",
  49663=>"111110000",
  49664=>"011110111",
  49665=>"011111010",
  49666=>"101101101",
  49667=>"000001000",
  49668=>"000111001",
  49669=>"000001111",
  49670=>"100111110",
  49671=>"011111111",
  49672=>"110011101",
  49673=>"100111110",
  49674=>"000010010",
  49675=>"111010100",
  49676=>"000011000",
  49677=>"000001110",
  49678=>"010001110",
  49679=>"100110010",
  49680=>"100000001",
  49681=>"011100101",
  49682=>"010101000",
  49683=>"110100000",
  49684=>"001011111",
  49685=>"011010010",
  49686=>"010100001",
  49687=>"001100000",
  49688=>"000110111",
  49689=>"000010101",
  49690=>"101010110",
  49691=>"101000001",
  49692=>"100001110",
  49693=>"111011011",
  49694=>"000101000",
  49695=>"111000111",
  49696=>"100111100",
  49697=>"101100010",
  49698=>"001011110",
  49699=>"111011101",
  49700=>"100101111",
  49701=>"101101011",
  49702=>"010001011",
  49703=>"010100000",
  49704=>"000010111",
  49705=>"111000101",
  49706=>"101101110",
  49707=>"100011100",
  49708=>"000011000",
  49709=>"101101110",
  49710=>"101100011",
  49711=>"100010010",
  49712=>"011011100",
  49713=>"011010010",
  49714=>"010010011",
  49715=>"011110010",
  49716=>"000001010",
  49717=>"001101100",
  49718=>"000011101",
  49719=>"111110011",
  49720=>"111001001",
  49721=>"100011011",
  49722=>"011000111",
  49723=>"111011101",
  49724=>"000011010",
  49725=>"000101101",
  49726=>"101101000",
  49727=>"101100000",
  49728=>"110101101",
  49729=>"010011001",
  49730=>"101000111",
  49731=>"101010000",
  49732=>"110100001",
  49733=>"110101101",
  49734=>"010001110",
  49735=>"001001101",
  49736=>"100101111",
  49737=>"011100001",
  49738=>"101001110",
  49739=>"010110101",
  49740=>"010010111",
  49741=>"001000100",
  49742=>"101110011",
  49743=>"010001101",
  49744=>"110000000",
  49745=>"000001101",
  49746=>"000111111",
  49747=>"101001111",
  49748=>"010101110",
  49749=>"100001001",
  49750=>"111100000",
  49751=>"010001010",
  49752=>"011001110",
  49753=>"010010001",
  49754=>"110110110",
  49755=>"101001111",
  49756=>"100000001",
  49757=>"110101101",
  49758=>"111110111",
  49759=>"010010011",
  49760=>"000011011",
  49761=>"011101101",
  49762=>"101000001",
  49763=>"111101100",
  49764=>"111111111",
  49765=>"000010110",
  49766=>"001100010",
  49767=>"101001011",
  49768=>"000000001",
  49769=>"001100000",
  49770=>"001100011",
  49771=>"100000000",
  49772=>"111111110",
  49773=>"110001011",
  49774=>"010111001",
  49775=>"110111100",
  49776=>"111111111",
  49777=>"101110101",
  49778=>"110101100",
  49779=>"001010100",
  49780=>"100110001",
  49781=>"000001010",
  49782=>"011101100",
  49783=>"101111101",
  49784=>"010110000",
  49785=>"110111011",
  49786=>"100010110",
  49787=>"111010111",
  49788=>"111010010",
  49789=>"110110010",
  49790=>"111111011",
  49791=>"100101100",
  49792=>"000000101",
  49793=>"101110111",
  49794=>"011100111",
  49795=>"001000101",
  49796=>"011000101",
  49797=>"010011010",
  49798=>"001000100",
  49799=>"000100001",
  49800=>"101010010",
  49801=>"001000011",
  49802=>"111110011",
  49803=>"001110001",
  49804=>"111111100",
  49805=>"101001011",
  49806=>"010100010",
  49807=>"111101111",
  49808=>"010111101",
  49809=>"101001111",
  49810=>"101110110",
  49811=>"010001100",
  49812=>"111101101",
  49813=>"011000001",
  49814=>"001000011",
  49815=>"011001000",
  49816=>"101101111",
  49817=>"010010101",
  49818=>"000100000",
  49819=>"000110001",
  49820=>"000010010",
  49821=>"110101110",
  49822=>"100101111",
  49823=>"100000100",
  49824=>"110110000",
  49825=>"001100000",
  49826=>"000100001",
  49827=>"100101000",
  49828=>"010010000",
  49829=>"000011001",
  49830=>"101010110",
  49831=>"010111000",
  49832=>"100111110",
  49833=>"001000011",
  49834=>"001111111",
  49835=>"001000111",
  49836=>"111010100",
  49837=>"101110101",
  49838=>"001100010",
  49839=>"110101110",
  49840=>"100100100",
  49841=>"111101010",
  49842=>"100111101",
  49843=>"011011010",
  49844=>"000000000",
  49845=>"111000000",
  49846=>"110100010",
  49847=>"001000011",
  49848=>"011011011",
  49849=>"110110001",
  49850=>"110011011",
  49851=>"101000000",
  49852=>"001001000",
  49853=>"011111010",
  49854=>"100110111",
  49855=>"111110111",
  49856=>"000110110",
  49857=>"100110110",
  49858=>"100100010",
  49859=>"110001101",
  49860=>"101011101",
  49861=>"000000010",
  49862=>"100110010",
  49863=>"011001110",
  49864=>"101001110",
  49865=>"011010111",
  49866=>"111000001",
  49867=>"110011111",
  49868=>"010100001",
  49869=>"010010100",
  49870=>"001101000",
  49871=>"010001010",
  49872=>"000010110",
  49873=>"011111101",
  49874=>"011101101",
  49875=>"111111001",
  49876=>"010100011",
  49877=>"011100110",
  49878=>"010011101",
  49879=>"010000100",
  49880=>"100111111",
  49881=>"101110110",
  49882=>"111100110",
  49883=>"010001101",
  49884=>"110110001",
  49885=>"101100011",
  49886=>"111100111",
  49887=>"001100110",
  49888=>"001111111",
  49889=>"111011011",
  49890=>"111001000",
  49891=>"011111111",
  49892=>"000001000",
  49893=>"001110001",
  49894=>"001011011",
  49895=>"000111011",
  49896=>"100101101",
  49897=>"001011001",
  49898=>"001101000",
  49899=>"100101111",
  49900=>"000100000",
  49901=>"010110111",
  49902=>"101101011",
  49903=>"101110100",
  49904=>"111111011",
  49905=>"101011011",
  49906=>"011111110",
  49907=>"010101001",
  49908=>"110000101",
  49909=>"111110110",
  49910=>"101000110",
  49911=>"100001111",
  49912=>"111101010",
  49913=>"000011000",
  49914=>"000010001",
  49915=>"010000100",
  49916=>"000110001",
  49917=>"001110111",
  49918=>"010001110",
  49919=>"101111001",
  49920=>"011010000",
  49921=>"000011011",
  49922=>"100010111",
  49923=>"010100110",
  49924=>"111000001",
  49925=>"111000111",
  49926=>"001010011",
  49927=>"111010000",
  49928=>"011001000",
  49929=>"011100101",
  49930=>"010001110",
  49931=>"111000001",
  49932=>"101100110",
  49933=>"101000000",
  49934=>"001000001",
  49935=>"011110010",
  49936=>"001011000",
  49937=>"011101010",
  49938=>"110111011",
  49939=>"100100100",
  49940=>"000110000",
  49941=>"011000001",
  49942=>"100001000",
  49943=>"110101011",
  49944=>"111111100",
  49945=>"010111010",
  49946=>"000111010",
  49947=>"101011111",
  49948=>"010101001",
  49949=>"100111000",
  49950=>"000001010",
  49951=>"001110001",
  49952=>"101000101",
  49953=>"000101100",
  49954=>"100100001",
  49955=>"000001111",
  49956=>"000110001",
  49957=>"101011011",
  49958=>"110110101",
  49959=>"011011111",
  49960=>"001000100",
  49961=>"000011011",
  49962=>"011111011",
  49963=>"000100100",
  49964=>"011001111",
  49965=>"101111111",
  49966=>"000000000",
  49967=>"101101101",
  49968=>"111101000",
  49969=>"000010010",
  49970=>"101001011",
  49971=>"001100011",
  49972=>"111101000",
  49973=>"000101000",
  49974=>"101010011",
  49975=>"110011101",
  49976=>"110000110",
  49977=>"101111001",
  49978=>"001111111",
  49979=>"110100100",
  49980=>"111001011",
  49981=>"011000011",
  49982=>"110101010",
  49983=>"001001011",
  49984=>"110010011",
  49985=>"101100001",
  49986=>"100000010",
  49987=>"011111001",
  49988=>"001000010",
  49989=>"110011000",
  49990=>"011111000",
  49991=>"110101010",
  49992=>"001111001",
  49993=>"111101110",
  49994=>"101110011",
  49995=>"110100100",
  49996=>"101100010",
  49997=>"111001101",
  49998=>"000011111",
  49999=>"100000110",
  50000=>"101001101",
  50001=>"101001111",
  50002=>"110001010",
  50003=>"101000110",
  50004=>"010111001",
  50005=>"011110111",
  50006=>"100101110",
  50007=>"101010111",
  50008=>"010111001",
  50009=>"100101001",
  50010=>"100111000",
  50011=>"001011011",
  50012=>"000011101",
  50013=>"010000100",
  50014=>"000101110",
  50015=>"000010110",
  50016=>"011000001",
  50017=>"010010110",
  50018=>"001110000",
  50019=>"111010000",
  50020=>"011110100",
  50021=>"111100101",
  50022=>"101111111",
  50023=>"111100001",
  50024=>"110110000",
  50025=>"101101010",
  50026=>"110011000",
  50027=>"110110000",
  50028=>"011100011",
  50029=>"100111101",
  50030=>"110010001",
  50031=>"010111110",
  50032=>"110001101",
  50033=>"000000001",
  50034=>"010011011",
  50035=>"000101010",
  50036=>"011110110",
  50037=>"100100010",
  50038=>"001110011",
  50039=>"010101010",
  50040=>"000010011",
  50041=>"010001000",
  50042=>"101011101",
  50043=>"111111101",
  50044=>"011111001",
  50045=>"111010011",
  50046=>"000100100",
  50047=>"101101000",
  50048=>"101101011",
  50049=>"010010011",
  50050=>"110000001",
  50051=>"111000111",
  50052=>"010000000",
  50053=>"111000001",
  50054=>"000001000",
  50055=>"101011111",
  50056=>"101111101",
  50057=>"000101100",
  50058=>"110110110",
  50059=>"100110110",
  50060=>"000101100",
  50061=>"100011000",
  50062=>"111111100",
  50063=>"100101001",
  50064=>"110010111",
  50065=>"010101010",
  50066=>"001101101",
  50067=>"000001111",
  50068=>"101011001",
  50069=>"101010001",
  50070=>"110111110",
  50071=>"100000010",
  50072=>"110111100",
  50073=>"001110011",
  50074=>"111101011",
  50075=>"011011110",
  50076=>"000100100",
  50077=>"100001011",
  50078=>"101111010",
  50079=>"001101100",
  50080=>"010101001",
  50081=>"110110000",
  50082=>"010000000",
  50083=>"111111111",
  50084=>"001011011",
  50085=>"010110010",
  50086=>"011101011",
  50087=>"111111101",
  50088=>"110111111",
  50089=>"010000100",
  50090=>"011010000",
  50091=>"010101000",
  50092=>"101101101",
  50093=>"110001111",
  50094=>"000011010",
  50095=>"100000001",
  50096=>"101111100",
  50097=>"110110100",
  50098=>"100100000",
  50099=>"110011001",
  50100=>"101101110",
  50101=>"011001100",
  50102=>"001001000",
  50103=>"111110000",
  50104=>"100011000",
  50105=>"110010010",
  50106=>"110011100",
  50107=>"110011100",
  50108=>"111101111",
  50109=>"001000000",
  50110=>"101101110",
  50111=>"001111011",
  50112=>"000011110",
  50113=>"111000000",
  50114=>"111110011",
  50115=>"011101101",
  50116=>"000111100",
  50117=>"001110111",
  50118=>"100101010",
  50119=>"010111111",
  50120=>"101001011",
  50121=>"111011001",
  50122=>"011111011",
  50123=>"110101011",
  50124=>"011000111",
  50125=>"010001010",
  50126=>"011100110",
  50127=>"000111010",
  50128=>"000010001",
  50129=>"000110100",
  50130=>"010001000",
  50131=>"000001100",
  50132=>"010011110",
  50133=>"110011111",
  50134=>"010111101",
  50135=>"000011111",
  50136=>"010000101",
  50137=>"000110000",
  50138=>"110001000",
  50139=>"010101001",
  50140=>"101001101",
  50141=>"000111101",
  50142=>"010101000",
  50143=>"101111111",
  50144=>"110000110",
  50145=>"000010000",
  50146=>"000000110",
  50147=>"101111101",
  50148=>"110011010",
  50149=>"000001101",
  50150=>"000011010",
  50151=>"101101001",
  50152=>"101010101",
  50153=>"011000011",
  50154=>"111011011",
  50155=>"111010100",
  50156=>"010100010",
  50157=>"000010101",
  50158=>"111000010",
  50159=>"010010110",
  50160=>"100010100",
  50161=>"000011110",
  50162=>"100001010",
  50163=>"010101010",
  50164=>"100010010",
  50165=>"000000101",
  50166=>"010111010",
  50167=>"011011111",
  50168=>"000011010",
  50169=>"000110000",
  50170=>"001011001",
  50171=>"100101001",
  50172=>"111110011",
  50173=>"000101010",
  50174=>"001111011",
  50175=>"010011011",
  50176=>"010000111",
  50177=>"001101011",
  50178=>"010101010",
  50179=>"111101011",
  50180=>"101011101",
  50181=>"111011011",
  50182=>"011111101",
  50183=>"001011111",
  50184=>"011000101",
  50185=>"110111010",
  50186=>"100101010",
  50187=>"011100001",
  50188=>"000111101",
  50189=>"100101011",
  50190=>"101100110",
  50191=>"001000000",
  50192=>"001110011",
  50193=>"110100000",
  50194=>"110000001",
  50195=>"101110110",
  50196=>"000010000",
  50197=>"001100100",
  50198=>"001110110",
  50199=>"101111010",
  50200=>"101100000",
  50201=>"100000101",
  50202=>"011011011",
  50203=>"111011000",
  50204=>"001101000",
  50205=>"000000111",
  50206=>"110110000",
  50207=>"011011100",
  50208=>"000011111",
  50209=>"101101000",
  50210=>"100001111",
  50211=>"101010101",
  50212=>"010010111",
  50213=>"111110011",
  50214=>"001110001",
  50215=>"101111010",
  50216=>"011001001",
  50217=>"000011110",
  50218=>"100100011",
  50219=>"011000001",
  50220=>"101000100",
  50221=>"101100110",
  50222=>"011011111",
  50223=>"000011111",
  50224=>"011011001",
  50225=>"011100001",
  50226=>"101101001",
  50227=>"000001000",
  50228=>"010000110",
  50229=>"010010011",
  50230=>"110110101",
  50231=>"111010110",
  50232=>"111101010",
  50233=>"001001011",
  50234=>"011010110",
  50235=>"101111011",
  50236=>"101010100",
  50237=>"100111000",
  50238=>"110101101",
  50239=>"101000000",
  50240=>"000011101",
  50241=>"000101110",
  50242=>"001101110",
  50243=>"010110010",
  50244=>"001110000",
  50245=>"011000110",
  50246=>"110111100",
  50247=>"000000000",
  50248=>"000010011",
  50249=>"111000001",
  50250=>"010101111",
  50251=>"000101000",
  50252=>"111001101",
  50253=>"110110111",
  50254=>"000000000",
  50255=>"101111110",
  50256=>"111001111",
  50257=>"001111110",
  50258=>"001101010",
  50259=>"010001111",
  50260=>"011000111",
  50261=>"111011101",
  50262=>"011110010",
  50263=>"001111111",
  50264=>"110111001",
  50265=>"111111000",
  50266=>"111010010",
  50267=>"100001111",
  50268=>"111011010",
  50269=>"010010011",
  50270=>"110111001",
  50271=>"010100110",
  50272=>"000000111",
  50273=>"101101100",
  50274=>"100001100",
  50275=>"011100011",
  50276=>"111111000",
  50277=>"100110111",
  50278=>"101011011",
  50279=>"100000011",
  50280=>"000000000",
  50281=>"100010000",
  50282=>"100010100",
  50283=>"110111101",
  50284=>"001011101",
  50285=>"101010000",
  50286=>"011110100",
  50287=>"101001011",
  50288=>"001000000",
  50289=>"000001101",
  50290=>"000110001",
  50291=>"000111111",
  50292=>"011001000",
  50293=>"001111010",
  50294=>"101001010",
  50295=>"011110110",
  50296=>"101100000",
  50297=>"001011110",
  50298=>"100001100",
  50299=>"000111111",
  50300=>"100101110",
  50301=>"110101110",
  50302=>"111010111",
  50303=>"001010110",
  50304=>"010101101",
  50305=>"011100110",
  50306=>"011001001",
  50307=>"010110101",
  50308=>"000010101",
  50309=>"011001000",
  50310=>"010110011",
  50311=>"000111010",
  50312=>"011010110",
  50313=>"101100000",
  50314=>"000000101",
  50315=>"101110010",
  50316=>"011100001",
  50317=>"110001010",
  50318=>"110110111",
  50319=>"010001010",
  50320=>"011011111",
  50321=>"001010111",
  50322=>"111100111",
  50323=>"101011000",
  50324=>"000101110",
  50325=>"100000010",
  50326=>"010101111",
  50327=>"100000001",
  50328=>"011001011",
  50329=>"010001100",
  50330=>"110001000",
  50331=>"110001100",
  50332=>"110011100",
  50333=>"110001110",
  50334=>"001010100",
  50335=>"011100101",
  50336=>"001111111",
  50337=>"100111010",
  50338=>"000110000",
  50339=>"111101000",
  50340=>"010111000",
  50341=>"101010001",
  50342=>"100101011",
  50343=>"000110101",
  50344=>"110101100",
  50345=>"110001011",
  50346=>"000101010",
  50347=>"111100110",
  50348=>"000010100",
  50349=>"100110011",
  50350=>"100010100",
  50351=>"101100001",
  50352=>"101000011",
  50353=>"110011011",
  50354=>"000100110",
  50355=>"011000100",
  50356=>"000000001",
  50357=>"011110100",
  50358=>"010000001",
  50359=>"001110100",
  50360=>"111111010",
  50361=>"001011001",
  50362=>"100011010",
  50363=>"001001010",
  50364=>"000101110",
  50365=>"000001110",
  50366=>"011010010",
  50367=>"010111101",
  50368=>"001100110",
  50369=>"101100010",
  50370=>"110100000",
  50371=>"001011000",
  50372=>"000010011",
  50373=>"101111111",
  50374=>"100000011",
  50375=>"110010110",
  50376=>"111111010",
  50377=>"101100100",
  50378=>"000100010",
  50379=>"111110000",
  50380=>"011001111",
  50381=>"010010111",
  50382=>"010000010",
  50383=>"001100000",
  50384=>"000000010",
  50385=>"101011100",
  50386=>"111000010",
  50387=>"010101100",
  50388=>"111100110",
  50389=>"100110100",
  50390=>"101101011",
  50391=>"010111101",
  50392=>"100111001",
  50393=>"001111110",
  50394=>"000001110",
  50395=>"000011000",
  50396=>"010110000",
  50397=>"101111100",
  50398=>"001011111",
  50399=>"101000000",
  50400=>"111000100",
  50401=>"100101010",
  50402=>"111001110",
  50403=>"011000110",
  50404=>"011110101",
  50405=>"101010011",
  50406=>"110110011",
  50407=>"111100111",
  50408=>"100000111",
  50409=>"001110010",
  50410=>"000001000",
  50411=>"111100111",
  50412=>"110110100",
  50413=>"010010011",
  50414=>"011001000",
  50415=>"011000010",
  50416=>"111110110",
  50417=>"101101101",
  50418=>"000101001",
  50419=>"001010011",
  50420=>"101101110",
  50421=>"011001111",
  50422=>"100010111",
  50423=>"100101001",
  50424=>"001001011",
  50425=>"101101110",
  50426=>"000000001",
  50427=>"000010001",
  50428=>"111011110",
  50429=>"101101000",
  50430=>"010001101",
  50431=>"100111001",
  50432=>"010010101",
  50433=>"110110000",
  50434=>"010111111",
  50435=>"110010010",
  50436=>"111010000",
  50437=>"100111111",
  50438=>"101111111",
  50439=>"011000111",
  50440=>"001010101",
  50441=>"000110111",
  50442=>"000111110",
  50443=>"111010000",
  50444=>"110101001",
  50445=>"011000111",
  50446=>"001101111",
  50447=>"010010011",
  50448=>"011010101",
  50449=>"011001010",
  50450=>"101011110",
  50451=>"011010110",
  50452=>"010000101",
  50453=>"100101001",
  50454=>"100000111",
  50455=>"111101101",
  50456=>"010101010",
  50457=>"101011110",
  50458=>"110111000",
  50459=>"000110111",
  50460=>"111111110",
  50461=>"110001011",
  50462=>"010011010",
  50463=>"000011110",
  50464=>"000101101",
  50465=>"000000111",
  50466=>"101011011",
  50467=>"111010110",
  50468=>"010110001",
  50469=>"010000100",
  50470=>"110111010",
  50471=>"000011111",
  50472=>"111101000",
  50473=>"010101110",
  50474=>"110001100",
  50475=>"010111110",
  50476=>"010000110",
  50477=>"110010000",
  50478=>"101101011",
  50479=>"000010000",
  50480=>"100011101",
  50481=>"000100010",
  50482=>"010001101",
  50483=>"111100011",
  50484=>"000110001",
  50485=>"110001101",
  50486=>"010000001",
  50487=>"010001010",
  50488=>"011000011",
  50489=>"000011010",
  50490=>"000100011",
  50491=>"110000100",
  50492=>"010110111",
  50493=>"110001110",
  50494=>"110110011",
  50495=>"011111111",
  50496=>"010101010",
  50497=>"100000111",
  50498=>"110010011",
  50499=>"101010011",
  50500=>"011000010",
  50501=>"100000111",
  50502=>"011000111",
  50503=>"110111100",
  50504=>"111100000",
  50505=>"001001100",
  50506=>"101111100",
  50507=>"011000001",
  50508=>"001100101",
  50509=>"011011101",
  50510=>"010111110",
  50511=>"110000001",
  50512=>"111011101",
  50513=>"101000100",
  50514=>"000000110",
  50515=>"010110111",
  50516=>"101000000",
  50517=>"000100010",
  50518=>"001101000",
  50519=>"011000010",
  50520=>"011101100",
  50521=>"100001100",
  50522=>"100110010",
  50523=>"101101101",
  50524=>"011111110",
  50525=>"111101101",
  50526=>"011011001",
  50527=>"111101110",
  50528=>"110101010",
  50529=>"011110001",
  50530=>"110111101",
  50531=>"011100010",
  50532=>"100000110",
  50533=>"000000101",
  50534=>"011001101",
  50535=>"101001101",
  50536=>"101100010",
  50537=>"000110000",
  50538=>"011011101",
  50539=>"001000011",
  50540=>"011111111",
  50541=>"101010110",
  50542=>"101101110",
  50543=>"101101111",
  50544=>"000001110",
  50545=>"000011010",
  50546=>"000000001",
  50547=>"010111011",
  50548=>"000101110",
  50549=>"110101100",
  50550=>"010110011",
  50551=>"010111110",
  50552=>"001111100",
  50553=>"101110011",
  50554=>"010101011",
  50555=>"010101001",
  50556=>"000011110",
  50557=>"111111111",
  50558=>"011010101",
  50559=>"011111111",
  50560=>"111101010",
  50561=>"111111101",
  50562=>"011101101",
  50563=>"010101110",
  50564=>"010000011",
  50565=>"111101001",
  50566=>"111001111",
  50567=>"111110011",
  50568=>"101011001",
  50569=>"111111011",
  50570=>"010011110",
  50571=>"110110010",
  50572=>"000110101",
  50573=>"111010111",
  50574=>"001101000",
  50575=>"011111010",
  50576=>"101010000",
  50577=>"010011100",
  50578=>"110010111",
  50579=>"000111001",
  50580=>"001100100",
  50581=>"101110101",
  50582=>"001010101",
  50583=>"110001011",
  50584=>"110110000",
  50585=>"110100110",
  50586=>"101100100",
  50587=>"001001010",
  50588=>"010000101",
  50589=>"100101011",
  50590=>"110101001",
  50591=>"000000111",
  50592=>"000100000",
  50593=>"100011000",
  50594=>"010000101",
  50595=>"110001110",
  50596=>"110001011",
  50597=>"010010110",
  50598=>"100000100",
  50599=>"100111100",
  50600=>"000111101",
  50601=>"011000010",
  50602=>"011001011",
  50603=>"110011010",
  50604=>"110011010",
  50605=>"110111101",
  50606=>"011100100",
  50607=>"000111001",
  50608=>"001010010",
  50609=>"000000111",
  50610=>"010111100",
  50611=>"110111010",
  50612=>"100101110",
  50613=>"101110100",
  50614=>"001100110",
  50615=>"101100011",
  50616=>"110010100",
  50617=>"001001010",
  50618=>"000010110",
  50619=>"011110110",
  50620=>"111110111",
  50621=>"000000011",
  50622=>"001110000",
  50623=>"101011010",
  50624=>"001000110",
  50625=>"101100001",
  50626=>"100100111",
  50627=>"011111000",
  50628=>"001100101",
  50629=>"100101100",
  50630=>"011000110",
  50631=>"100101111",
  50632=>"101000010",
  50633=>"010100000",
  50634=>"110101000",
  50635=>"100110011",
  50636=>"001110100",
  50637=>"011111101",
  50638=>"000100110",
  50639=>"001000100",
  50640=>"101001010",
  50641=>"111110101",
  50642=>"011001000",
  50643=>"010111100",
  50644=>"101011100",
  50645=>"011010011",
  50646=>"101111011",
  50647=>"111111111",
  50648=>"111110000",
  50649=>"010100100",
  50650=>"000100000",
  50651=>"110011110",
  50652=>"011101000",
  50653=>"110101001",
  50654=>"111101101",
  50655=>"100011011",
  50656=>"011001101",
  50657=>"001011011",
  50658=>"001100101",
  50659=>"011011001",
  50660=>"111100001",
  50661=>"100101011",
  50662=>"110111100",
  50663=>"000010100",
  50664=>"110111011",
  50665=>"101110100",
  50666=>"000111010",
  50667=>"011110101",
  50668=>"111000001",
  50669=>"010100100",
  50670=>"111001011",
  50671=>"100101100",
  50672=>"100010110",
  50673=>"011010100",
  50674=>"011111101",
  50675=>"100001111",
  50676=>"110110101",
  50677=>"100000000",
  50678=>"101010011",
  50679=>"000111011",
  50680=>"001000011",
  50681=>"010010000",
  50682=>"111010001",
  50683=>"001010110",
  50684=>"000000011",
  50685=>"111111110",
  50686=>"101110011",
  50687=>"011011111",
  50688=>"111000011",
  50689=>"101011101",
  50690=>"101000011",
  50691=>"101111001",
  50692=>"111111011",
  50693=>"000000100",
  50694=>"010100100",
  50695=>"001010110",
  50696=>"001100011",
  50697=>"111010101",
  50698=>"000111011",
  50699=>"001010001",
  50700=>"100001000",
  50701=>"110110111",
  50702=>"000011000",
  50703=>"011110001",
  50704=>"000111100",
  50705=>"011110001",
  50706=>"111011111",
  50707=>"010100101",
  50708=>"010011010",
  50709=>"101000101",
  50710=>"110111111",
  50711=>"101111101",
  50712=>"011101001",
  50713=>"100111001",
  50714=>"100001000",
  50715=>"011001101",
  50716=>"101100111",
  50717=>"011010101",
  50718=>"101101111",
  50719=>"000101110",
  50720=>"001001000",
  50721=>"101110111",
  50722=>"000001010",
  50723=>"001010100",
  50724=>"001111100",
  50725=>"111100000",
  50726=>"010011010",
  50727=>"101011100",
  50728=>"101000101",
  50729=>"101100011",
  50730=>"110101011",
  50731=>"111110111",
  50732=>"101011000",
  50733=>"001101000",
  50734=>"101000001",
  50735=>"011111010",
  50736=>"001100100",
  50737=>"001001000",
  50738=>"100001000",
  50739=>"110000100",
  50740=>"010001011",
  50741=>"111100000",
  50742=>"111101010",
  50743=>"000110000",
  50744=>"001101101",
  50745=>"101111110",
  50746=>"001000100",
  50747=>"011011010",
  50748=>"100100110",
  50749=>"011001111",
  50750=>"100011011",
  50751=>"000010110",
  50752=>"000001100",
  50753=>"001011000",
  50754=>"110010010",
  50755=>"101000001",
  50756=>"010000100",
  50757=>"100001010",
  50758=>"010100110",
  50759=>"110101100",
  50760=>"001011100",
  50761=>"101111101",
  50762=>"101010110",
  50763=>"101101111",
  50764=>"001010001",
  50765=>"100110000",
  50766=>"110111001",
  50767=>"011101110",
  50768=>"011110011",
  50769=>"100000000",
  50770=>"111010100",
  50771=>"000100000",
  50772=>"111000000",
  50773=>"111000100",
  50774=>"001100001",
  50775=>"000000011",
  50776=>"110101100",
  50777=>"001111010",
  50778=>"110100110",
  50779=>"110001100",
  50780=>"010101111",
  50781=>"000110000",
  50782=>"000101000",
  50783=>"010000101",
  50784=>"010101001",
  50785=>"001110000",
  50786=>"100000011",
  50787=>"100001100",
  50788=>"000110100",
  50789=>"111110011",
  50790=>"100000101",
  50791=>"111110101",
  50792=>"000111010",
  50793=>"110000010",
  50794=>"000110100",
  50795=>"101011101",
  50796=>"011111100",
  50797=>"011010010",
  50798=>"101111100",
  50799=>"111101110",
  50800=>"110101101",
  50801=>"000010000",
  50802=>"001111011",
  50803=>"010001101",
  50804=>"011110001",
  50805=>"101000111",
  50806=>"010100110",
  50807=>"100110101",
  50808=>"110000001",
  50809=>"000000010",
  50810=>"110111000",
  50811=>"011000000",
  50812=>"011001101",
  50813=>"111001010",
  50814=>"100001101",
  50815=>"110011111",
  50816=>"100011011",
  50817=>"101111110",
  50818=>"111101111",
  50819=>"010111101",
  50820=>"000110110",
  50821=>"000111000",
  50822=>"010101001",
  50823=>"011101001",
  50824=>"001111101",
  50825=>"000001001",
  50826=>"100011111",
  50827=>"110110011",
  50828=>"001110101",
  50829=>"101110101",
  50830=>"100011001",
  50831=>"010010110",
  50832=>"110000010",
  50833=>"010100000",
  50834=>"011110100",
  50835=>"001000111",
  50836=>"010011110",
  50837=>"000101001",
  50838=>"111101100",
  50839=>"101000110",
  50840=>"000000110",
  50841=>"100100100",
  50842=>"110110111",
  50843=>"000001110",
  50844=>"000100010",
  50845=>"100010011",
  50846=>"110011000",
  50847=>"010111111",
  50848=>"110001111",
  50849=>"011100010",
  50850=>"101000011",
  50851=>"100100001",
  50852=>"010010101",
  50853=>"000000001",
  50854=>"110110101",
  50855=>"111010010",
  50856=>"001010010",
  50857=>"110110001",
  50858=>"110010000",
  50859=>"011101000",
  50860=>"110011000",
  50861=>"000010010",
  50862=>"010000101",
  50863=>"010100101",
  50864=>"110000100",
  50865=>"011001110",
  50866=>"000011000",
  50867=>"101100100",
  50868=>"001000001",
  50869=>"100111010",
  50870=>"111100100",
  50871=>"110011011",
  50872=>"010111010",
  50873=>"110011010",
  50874=>"000000001",
  50875=>"111011111",
  50876=>"011100110",
  50877=>"111111001",
  50878=>"000001011",
  50879=>"000100011",
  50880=>"000000000",
  50881=>"001110000",
  50882=>"101111101",
  50883=>"010001111",
  50884=>"001000111",
  50885=>"100001110",
  50886=>"001000110",
  50887=>"001000110",
  50888=>"011011011",
  50889=>"100011110",
  50890=>"111110101",
  50891=>"101100101",
  50892=>"110101010",
  50893=>"110011001",
  50894=>"000110110",
  50895=>"111101010",
  50896=>"101000001",
  50897=>"000000010",
  50898=>"000101000",
  50899=>"101010010",
  50900=>"100111011",
  50901=>"001010101",
  50902=>"100100100",
  50903=>"110110000",
  50904=>"110111100",
  50905=>"000110110",
  50906=>"001000111",
  50907=>"000011000",
  50908=>"001000000",
  50909=>"101001111",
  50910=>"001101011",
  50911=>"110001101",
  50912=>"110010111",
  50913=>"110100101",
  50914=>"101111110",
  50915=>"011100011",
  50916=>"001101101",
  50917=>"101100101",
  50918=>"001100000",
  50919=>"001110000",
  50920=>"010000000",
  50921=>"111001011",
  50922=>"011000011",
  50923=>"000101010",
  50924=>"001100010",
  50925=>"110101110",
  50926=>"111110111",
  50927=>"010100111",
  50928=>"100010010",
  50929=>"001000010",
  50930=>"000000110",
  50931=>"000100010",
  50932=>"101100011",
  50933=>"100000100",
  50934=>"010100111",
  50935=>"001011000",
  50936=>"000001001",
  50937=>"111101001",
  50938=>"101100010",
  50939=>"100111011",
  50940=>"110000001",
  50941=>"100110101",
  50942=>"111100001",
  50943=>"001010000",
  50944=>"101000001",
  50945=>"000101000",
  50946=>"010001101",
  50947=>"111001100",
  50948=>"110111001",
  50949=>"001011111",
  50950=>"111010110",
  50951=>"111100101",
  50952=>"100100011",
  50953=>"100011011",
  50954=>"110101110",
  50955=>"110111101",
  50956=>"100101110",
  50957=>"100010011",
  50958=>"001010110",
  50959=>"101001111",
  50960=>"010111101",
  50961=>"111111101",
  50962=>"010000101",
  50963=>"101000011",
  50964=>"100111010",
  50965=>"101001111",
  50966=>"010100011",
  50967=>"010011010",
  50968=>"101001100",
  50969=>"001001110",
  50970=>"010101000",
  50971=>"101000101",
  50972=>"000100010",
  50973=>"010010111",
  50974=>"100110110",
  50975=>"010100011",
  50976=>"101110010",
  50977=>"011100101",
  50978=>"101100101",
  50979=>"000011110",
  50980=>"000101100",
  50981=>"000010000",
  50982=>"101010111",
  50983=>"111101010",
  50984=>"101101001",
  50985=>"011100011",
  50986=>"001011110",
  50987=>"111011010",
  50988=>"011111010",
  50989=>"111100110",
  50990=>"001001001",
  50991=>"110010100",
  50992=>"010011000",
  50993=>"001010000",
  50994=>"001101100",
  50995=>"011101110",
  50996=>"101110011",
  50997=>"011111111",
  50998=>"000000010",
  50999=>"010111110",
  51000=>"111010100",
  51001=>"100100111",
  51002=>"101000110",
  51003=>"001010100",
  51004=>"001110000",
  51005=>"100010000",
  51006=>"110110010",
  51007=>"110110100",
  51008=>"010011001",
  51009=>"000110101",
  51010=>"001011111",
  51011=>"111111000",
  51012=>"011100001",
  51013=>"111000000",
  51014=>"011001001",
  51015=>"101001101",
  51016=>"101111101",
  51017=>"000011010",
  51018=>"110001010",
  51019=>"011010011",
  51020=>"001000011",
  51021=>"011011101",
  51022=>"100000110",
  51023=>"111100101",
  51024=>"100111101",
  51025=>"011100000",
  51026=>"100101111",
  51027=>"000100110",
  51028=>"100001010",
  51029=>"001111110",
  51030=>"101110110",
  51031=>"011001010",
  51032=>"010000010",
  51033=>"111000111",
  51034=>"100001000",
  51035=>"001001010",
  51036=>"111111111",
  51037=>"110001111",
  51038=>"010111100",
  51039=>"000100001",
  51040=>"101111010",
  51041=>"111111011",
  51042=>"111001110",
  51043=>"100100110",
  51044=>"011001001",
  51045=>"101000111",
  51046=>"100100000",
  51047=>"010011100",
  51048=>"101101000",
  51049=>"101010011",
  51050=>"111000000",
  51051=>"001100010",
  51052=>"000000000",
  51053=>"010001010",
  51054=>"100011000",
  51055=>"010001011",
  51056=>"000011010",
  51057=>"000010110",
  51058=>"111111000",
  51059=>"111011001",
  51060=>"000001000",
  51061=>"110001101",
  51062=>"110101000",
  51063=>"011110000",
  51064=>"111010011",
  51065=>"000011001",
  51066=>"110010111",
  51067=>"110010011",
  51068=>"101111111",
  51069=>"110101100",
  51070=>"101101010",
  51071=>"011101001",
  51072=>"100101100",
  51073=>"000101100",
  51074=>"101000010",
  51075=>"001100011",
  51076=>"010010010",
  51077=>"110000101",
  51078=>"011111011",
  51079=>"010011000",
  51080=>"110111010",
  51081=>"100110000",
  51082=>"001111001",
  51083=>"111101010",
  51084=>"101100011",
  51085=>"011010010",
  51086=>"000100000",
  51087=>"000100101",
  51088=>"100111111",
  51089=>"011011111",
  51090=>"001110000",
  51091=>"110001101",
  51092=>"010010000",
  51093=>"101101110",
  51094=>"100001010",
  51095=>"001100100",
  51096=>"111100101",
  51097=>"010111011",
  51098=>"010010001",
  51099=>"100101100",
  51100=>"100010111",
  51101=>"010110000",
  51102=>"101111110",
  51103=>"100001101",
  51104=>"100100111",
  51105=>"000011101",
  51106=>"100110001",
  51107=>"010110000",
  51108=>"000100000",
  51109=>"101111101",
  51110=>"011011000",
  51111=>"011010111",
  51112=>"011001001",
  51113=>"001111101",
  51114=>"101000001",
  51115=>"011111010",
  51116=>"000001111",
  51117=>"011100010",
  51118=>"010011110",
  51119=>"100110010",
  51120=>"010100110",
  51121=>"110011101",
  51122=>"010111000",
  51123=>"000000001",
  51124=>"100000000",
  51125=>"110100111",
  51126=>"101110110",
  51127=>"001001111",
  51128=>"110100000",
  51129=>"000010011",
  51130=>"100111011",
  51131=>"001000001",
  51132=>"000110100",
  51133=>"001111011",
  51134=>"111110010",
  51135=>"100000000",
  51136=>"101100111",
  51137=>"001000110",
  51138=>"100011110",
  51139=>"101001001",
  51140=>"011000100",
  51141=>"001100011",
  51142=>"101110100",
  51143=>"111011111",
  51144=>"000010000",
  51145=>"001111111",
  51146=>"101111010",
  51147=>"101110111",
  51148=>"111000010",
  51149=>"001110110",
  51150=>"010111100",
  51151=>"111111101",
  51152=>"111111110",
  51153=>"101011000",
  51154=>"110110111",
  51155=>"000000111",
  51156=>"000000000",
  51157=>"000010101",
  51158=>"110001101",
  51159=>"100000110",
  51160=>"000100110",
  51161=>"111101011",
  51162=>"111101011",
  51163=>"011010110",
  51164=>"010011100",
  51165=>"111010101",
  51166=>"000010100",
  51167=>"011111101",
  51168=>"000111010",
  51169=>"000111010",
  51170=>"011111011",
  51171=>"101110101",
  51172=>"001111001",
  51173=>"111011011",
  51174=>"101000011",
  51175=>"010101101",
  51176=>"000100010",
  51177=>"100001010",
  51178=>"010011010",
  51179=>"001110000",
  51180=>"011111101",
  51181=>"101000010",
  51182=>"001100001",
  51183=>"000110100",
  51184=>"000001000",
  51185=>"111001011",
  51186=>"000011001",
  51187=>"110101001",
  51188=>"110111011",
  51189=>"001001000",
  51190=>"110001101",
  51191=>"011101110",
  51192=>"100100111",
  51193=>"010110010",
  51194=>"100000000",
  51195=>"110101010",
  51196=>"001000100",
  51197=>"000001100",
  51198=>"100010011",
  51199=>"111001110",
  51200=>"111011011",
  51201=>"110010010",
  51202=>"100110101",
  51203=>"100101010",
  51204=>"100001001",
  51205=>"100000010",
  51206=>"110010001",
  51207=>"111001010",
  51208=>"000111100",
  51209=>"011000111",
  51210=>"000101000",
  51211=>"010010100",
  51212=>"111100001",
  51213=>"011000110",
  51214=>"101010010",
  51215=>"110110000",
  51216=>"111101111",
  51217=>"111011000",
  51218=>"111000111",
  51219=>"101010001",
  51220=>"101001010",
  51221=>"010111011",
  51222=>"001101111",
  51223=>"010010110",
  51224=>"110101011",
  51225=>"100100001",
  51226=>"001111010",
  51227=>"101011011",
  51228=>"011111010",
  51229=>"110101011",
  51230=>"101011001",
  51231=>"101110000",
  51232=>"111101000",
  51233=>"100100001",
  51234=>"010000111",
  51235=>"001101100",
  51236=>"000101101",
  51237=>"100111100",
  51238=>"010000010",
  51239=>"001111110",
  51240=>"111101101",
  51241=>"101101011",
  51242=>"001110100",
  51243=>"001110011",
  51244=>"011101100",
  51245=>"111111010",
  51246=>"101111111",
  51247=>"110001010",
  51248=>"111110100",
  51249=>"011100010",
  51250=>"010001111",
  51251=>"111111010",
  51252=>"101110000",
  51253=>"110000000",
  51254=>"000010011",
  51255=>"101011100",
  51256=>"010010000",
  51257=>"001110111",
  51258=>"010011101",
  51259=>"001011001",
  51260=>"001100110",
  51261=>"111101001",
  51262=>"011000011",
  51263=>"001000100",
  51264=>"000000010",
  51265=>"101000011",
  51266=>"101101000",
  51267=>"101011001",
  51268=>"101001110",
  51269=>"001000110",
  51270=>"111100100",
  51271=>"010100001",
  51272=>"001000000",
  51273=>"001100110",
  51274=>"000000001",
  51275=>"110100011",
  51276=>"101000100",
  51277=>"110111100",
  51278=>"111101101",
  51279=>"011101100",
  51280=>"011010100",
  51281=>"110111110",
  51282=>"000011100",
  51283=>"101111010",
  51284=>"111001010",
  51285=>"001000011",
  51286=>"110101000",
  51287=>"110001001",
  51288=>"100011110",
  51289=>"001100011",
  51290=>"001001000",
  51291=>"010111010",
  51292=>"010010110",
  51293=>"000101001",
  51294=>"010010011",
  51295=>"101001011",
  51296=>"101001111",
  51297=>"100101111",
  51298=>"110110111",
  51299=>"100001000",
  51300=>"101010000",
  51301=>"001000110",
  51302=>"110000110",
  51303=>"011000011",
  51304=>"000110010",
  51305=>"110001000",
  51306=>"000000111",
  51307=>"001110100",
  51308=>"110010010",
  51309=>"001011100",
  51310=>"100000011",
  51311=>"010011010",
  51312=>"100101010",
  51313=>"001011001",
  51314=>"000010001",
  51315=>"001101101",
  51316=>"000000010",
  51317=>"100011100",
  51318=>"101110010",
  51319=>"111101111",
  51320=>"010101001",
  51321=>"110111000",
  51322=>"000000100",
  51323=>"100000110",
  51324=>"011111110",
  51325=>"111011000",
  51326=>"110010001",
  51327=>"011111111",
  51328=>"010001100",
  51329=>"110100010",
  51330=>"110001001",
  51331=>"010111100",
  51332=>"101110011",
  51333=>"110111100",
  51334=>"110111111",
  51335=>"111101011",
  51336=>"100110110",
  51337=>"110100010",
  51338=>"101001011",
  51339=>"000110001",
  51340=>"001000100",
  51341=>"100001010",
  51342=>"110010011",
  51343=>"010001110",
  51344=>"000101101",
  51345=>"100000010",
  51346=>"011101000",
  51347=>"101001011",
  51348=>"010111011",
  51349=>"010100100",
  51350=>"101101000",
  51351=>"110110010",
  51352=>"001011101",
  51353=>"000010001",
  51354=>"000001101",
  51355=>"101111101",
  51356=>"100000110",
  51357=>"100001110",
  51358=>"000001000",
  51359=>"111101010",
  51360=>"000100010",
  51361=>"101010110",
  51362=>"000000011",
  51363=>"001111100",
  51364=>"101000011",
  51365=>"000101111",
  51366=>"001111000",
  51367=>"101100101",
  51368=>"100100001",
  51369=>"111101001",
  51370=>"111001101",
  51371=>"110001101",
  51372=>"100101010",
  51373=>"000110000",
  51374=>"010010100",
  51375=>"011011001",
  51376=>"011011111",
  51377=>"001101000",
  51378=>"010110011",
  51379=>"111110000",
  51380=>"111001010",
  51381=>"101000101",
  51382=>"101100100",
  51383=>"010001001",
  51384=>"001101000",
  51385=>"000010101",
  51386=>"011011101",
  51387=>"100111101",
  51388=>"001001001",
  51389=>"100001010",
  51390=>"111001010",
  51391=>"110011011",
  51392=>"101011000",
  51393=>"101011101",
  51394=>"100000111",
  51395=>"011001101",
  51396=>"001100111",
  51397=>"001100010",
  51398=>"000101110",
  51399=>"100001000",
  51400=>"111010011",
  51401=>"000110101",
  51402=>"100110101",
  51403=>"010101001",
  51404=>"110010101",
  51405=>"000110110",
  51406=>"000011001",
  51407=>"010101010",
  51408=>"011111001",
  51409=>"100100011",
  51410=>"010001111",
  51411=>"011101000",
  51412=>"111001100",
  51413=>"111111101",
  51414=>"111001011",
  51415=>"001011101",
  51416=>"000011011",
  51417=>"111001110",
  51418=>"011001011",
  51419=>"100010010",
  51420=>"000111100",
  51421=>"101111111",
  51422=>"110010110",
  51423=>"000100100",
  51424=>"111101110",
  51425=>"100110001",
  51426=>"101101000",
  51427=>"000011110",
  51428=>"010111100",
  51429=>"101000111",
  51430=>"100110000",
  51431=>"010000011",
  51432=>"000000101",
  51433=>"100011010",
  51434=>"100010010",
  51435=>"010100111",
  51436=>"000100010",
  51437=>"000001100",
  51438=>"110010011",
  51439=>"011110010",
  51440=>"110111011",
  51441=>"000001000",
  51442=>"101000000",
  51443=>"000011110",
  51444=>"000101011",
  51445=>"111110111",
  51446=>"001100011",
  51447=>"001000100",
  51448=>"000000101",
  51449=>"011101100",
  51450=>"101100001",
  51451=>"111000000",
  51452=>"001011001",
  51453=>"010001111",
  51454=>"111011000",
  51455=>"100010001",
  51456=>"010111110",
  51457=>"110111101",
  51458=>"011100011",
  51459=>"010011011",
  51460=>"000101101",
  51461=>"111000011",
  51462=>"010101000",
  51463=>"010111101",
  51464=>"000010101",
  51465=>"000100100",
  51466=>"001100011",
  51467=>"101101101",
  51468=>"101000000",
  51469=>"110001100",
  51470=>"101011010",
  51471=>"001100111",
  51472=>"101011111",
  51473=>"110100100",
  51474=>"001100101",
  51475=>"000101111",
  51476=>"000000110",
  51477=>"111000001",
  51478=>"110000100",
  51479=>"010100011",
  51480=>"101100000",
  51481=>"111001111",
  51482=>"011101101",
  51483=>"011100111",
  51484=>"101010100",
  51485=>"001101111",
  51486=>"000001101",
  51487=>"100010001",
  51488=>"100100101",
  51489=>"011000000",
  51490=>"000010100",
  51491=>"100100111",
  51492=>"110110010",
  51493=>"000010010",
  51494=>"000000100",
  51495=>"011110101",
  51496=>"011000011",
  51497=>"110001110",
  51498=>"001110111",
  51499=>"100000011",
  51500=>"001100000",
  51501=>"110010111",
  51502=>"101111000",
  51503=>"101111010",
  51504=>"110011011",
  51505=>"111111001",
  51506=>"110000100",
  51507=>"100110110",
  51508=>"100011100",
  51509=>"100000000",
  51510=>"101011011",
  51511=>"111111111",
  51512=>"001000100",
  51513=>"110110010",
  51514=>"101111010",
  51515=>"101000011",
  51516=>"011000110",
  51517=>"010010010",
  51518=>"111111100",
  51519=>"000100011",
  51520=>"000100101",
  51521=>"111000001",
  51522=>"010010010",
  51523=>"111110110",
  51524=>"001000111",
  51525=>"111111101",
  51526=>"111000011",
  51527=>"011110101",
  51528=>"011000001",
  51529=>"100000001",
  51530=>"111101000",
  51531=>"100000011",
  51532=>"011010000",
  51533=>"101110001",
  51534=>"111011100",
  51535=>"101100001",
  51536=>"100100010",
  51537=>"101000011",
  51538=>"000000010",
  51539=>"001010100",
  51540=>"010101001",
  51541=>"110111111",
  51542=>"101010001",
  51543=>"001100010",
  51544=>"111000101",
  51545=>"011011111",
  51546=>"110100011",
  51547=>"100100101",
  51548=>"000111110",
  51549=>"100100100",
  51550=>"100010110",
  51551=>"011010011",
  51552=>"000101110",
  51553=>"100100010",
  51554=>"000101000",
  51555=>"111000000",
  51556=>"010010010",
  51557=>"110001111",
  51558=>"000101110",
  51559=>"111000000",
  51560=>"111111101",
  51561=>"011000010",
  51562=>"010111010",
  51563=>"001110100",
  51564=>"010001001",
  51565=>"111000011",
  51566=>"111000111",
  51567=>"001011001",
  51568=>"000010100",
  51569=>"010101111",
  51570=>"111010001",
  51571=>"110110010",
  51572=>"011110111",
  51573=>"100001011",
  51574=>"011010011",
  51575=>"111100000",
  51576=>"000110001",
  51577=>"011110110",
  51578=>"011001100",
  51579=>"011111111",
  51580=>"010101011",
  51581=>"111011010",
  51582=>"110111001",
  51583=>"011101111",
  51584=>"101001000",
  51585=>"100101001",
  51586=>"010010100",
  51587=>"000000010",
  51588=>"111110000",
  51589=>"000011000",
  51590=>"111100010",
  51591=>"011110001",
  51592=>"010111001",
  51593=>"001101100",
  51594=>"100010011",
  51595=>"000010110",
  51596=>"100000000",
  51597=>"011111001",
  51598=>"100010100",
  51599=>"011001110",
  51600=>"000110001",
  51601=>"011010101",
  51602=>"001000101",
  51603=>"111110001",
  51604=>"010101101",
  51605=>"111000000",
  51606=>"101110010",
  51607=>"111011011",
  51608=>"010101111",
  51609=>"100000000",
  51610=>"110001101",
  51611=>"010001110",
  51612=>"110111111",
  51613=>"001000001",
  51614=>"010100000",
  51615=>"000101100",
  51616=>"101100010",
  51617=>"100000101",
  51618=>"111010011",
  51619=>"100001010",
  51620=>"000100111",
  51621=>"011010010",
  51622=>"111010100",
  51623=>"001011000",
  51624=>"001000011",
  51625=>"110100100",
  51626=>"111001000",
  51627=>"011001100",
  51628=>"010001110",
  51629=>"011000010",
  51630=>"011111010",
  51631=>"010111110",
  51632=>"100111000",
  51633=>"101001000",
  51634=>"000011101",
  51635=>"001010111",
  51636=>"110111101",
  51637=>"011110110",
  51638=>"100111011",
  51639=>"100010111",
  51640=>"111100111",
  51641=>"100001111",
  51642=>"000111001",
  51643=>"001101110",
  51644=>"011010111",
  51645=>"001001101",
  51646=>"000100100",
  51647=>"100101101",
  51648=>"010100011",
  51649=>"001011100",
  51650=>"001101110",
  51651=>"110010001",
  51652=>"010111000",
  51653=>"111110010",
  51654=>"010001111",
  51655=>"011100000",
  51656=>"110000000",
  51657=>"001110100",
  51658=>"111001110",
  51659=>"000100100",
  51660=>"000001100",
  51661=>"011010010",
  51662=>"010001111",
  51663=>"111111000",
  51664=>"000000010",
  51665=>"101001000",
  51666=>"011100000",
  51667=>"000011001",
  51668=>"110100100",
  51669=>"001011001",
  51670=>"100011010",
  51671=>"000100010",
  51672=>"011000110",
  51673=>"111101101",
  51674=>"111010010",
  51675=>"110001100",
  51676=>"000000111",
  51677=>"110101100",
  51678=>"110111111",
  51679=>"111011100",
  51680=>"000101110",
  51681=>"000010011",
  51682=>"110101011",
  51683=>"101101001",
  51684=>"001010111",
  51685=>"110110101",
  51686=>"110101000",
  51687=>"001001010",
  51688=>"001101100",
  51689=>"001010110",
  51690=>"100001110",
  51691=>"010000001",
  51692=>"111000110",
  51693=>"111111110",
  51694=>"100111111",
  51695=>"010010010",
  51696=>"010011000",
  51697=>"111110111",
  51698=>"000101011",
  51699=>"101100110",
  51700=>"110110100",
  51701=>"111001000",
  51702=>"100010110",
  51703=>"000101101",
  51704=>"111010101",
  51705=>"101111101",
  51706=>"010001111",
  51707=>"000101001",
  51708=>"001010111",
  51709=>"110111100",
  51710=>"111101111",
  51711=>"110000100",
  51712=>"011011000",
  51713=>"011000001",
  51714=>"110000110",
  51715=>"100110010",
  51716=>"110010111",
  51717=>"001110000",
  51718=>"010101010",
  51719=>"101100010",
  51720=>"010110010",
  51721=>"000001010",
  51722=>"100110011",
  51723=>"000001101",
  51724=>"000001101",
  51725=>"001110101",
  51726=>"010100000",
  51727=>"010111001",
  51728=>"001010011",
  51729=>"000101000",
  51730=>"011110110",
  51731=>"100001011",
  51732=>"100000101",
  51733=>"100011001",
  51734=>"101010001",
  51735=>"011101011",
  51736=>"111100101",
  51737=>"110010011",
  51738=>"010001110",
  51739=>"001010001",
  51740=>"001010000",
  51741=>"011011011",
  51742=>"011010001",
  51743=>"100000100",
  51744=>"011110001",
  51745=>"011010000",
  51746=>"000100001",
  51747=>"101110001",
  51748=>"111100000",
  51749=>"100100001",
  51750=>"101010101",
  51751=>"110110101",
  51752=>"001000001",
  51753=>"101000011",
  51754=>"000000100",
  51755=>"011110100",
  51756=>"100001011",
  51757=>"010101011",
  51758=>"001111111",
  51759=>"101100000",
  51760=>"100001000",
  51761=>"011100111",
  51762=>"000101011",
  51763=>"111000010",
  51764=>"001011001",
  51765=>"100110000",
  51766=>"101001000",
  51767=>"111101111",
  51768=>"010100111",
  51769=>"110111111",
  51770=>"001011111",
  51771=>"111110010",
  51772=>"000000011",
  51773=>"001000000",
  51774=>"010001001",
  51775=>"111110010",
  51776=>"101000110",
  51777=>"101000011",
  51778=>"011001110",
  51779=>"111001011",
  51780=>"000001100",
  51781=>"011101001",
  51782=>"011111010",
  51783=>"010001101",
  51784=>"100001101",
  51785=>"110111001",
  51786=>"111110000",
  51787=>"001010010",
  51788=>"010111111",
  51789=>"011110110",
  51790=>"101000010",
  51791=>"100110000",
  51792=>"111110110",
  51793=>"001001110",
  51794=>"100100001",
  51795=>"011100110",
  51796=>"001011011",
  51797=>"110000000",
  51798=>"101010001",
  51799=>"100111110",
  51800=>"011010001",
  51801=>"010001110",
  51802=>"011111011",
  51803=>"100000000",
  51804=>"100101111",
  51805=>"010010101",
  51806=>"100001111",
  51807=>"101111011",
  51808=>"100000111",
  51809=>"110111000",
  51810=>"110110011",
  51811=>"111111000",
  51812=>"011011000",
  51813=>"111110110",
  51814=>"111111011",
  51815=>"111001000",
  51816=>"110000111",
  51817=>"000000011",
  51818=>"011110110",
  51819=>"111011100",
  51820=>"011000111",
  51821=>"110100011",
  51822=>"111001000",
  51823=>"110000111",
  51824=>"010101001",
  51825=>"001100000",
  51826=>"111011111",
  51827=>"000111110",
  51828=>"110011011",
  51829=>"100011010",
  51830=>"110110000",
  51831=>"011011111",
  51832=>"101111100",
  51833=>"100111110",
  51834=>"110000010",
  51835=>"100101010",
  51836=>"111111000",
  51837=>"101100111",
  51838=>"111110110",
  51839=>"111101000",
  51840=>"100011110",
  51841=>"011111001",
  51842=>"010001000",
  51843=>"100000001",
  51844=>"110011100",
  51845=>"110000111",
  51846=>"010011110",
  51847=>"001100101",
  51848=>"001100010",
  51849=>"101101110",
  51850=>"100111101",
  51851=>"010100001",
  51852=>"001101010",
  51853=>"011000101",
  51854=>"101001000",
  51855=>"110000110",
  51856=>"100000111",
  51857=>"010000011",
  51858=>"100011111",
  51859=>"111011111",
  51860=>"101011011",
  51861=>"111011000",
  51862=>"010110000",
  51863=>"110001010",
  51864=>"110100010",
  51865=>"100100100",
  51866=>"110001110",
  51867=>"001101010",
  51868=>"101100010",
  51869=>"101101011",
  51870=>"000001000",
  51871=>"111100100",
  51872=>"111000110",
  51873=>"001101000",
  51874=>"101100101",
  51875=>"101010100",
  51876=>"010000000",
  51877=>"001010110",
  51878=>"111001111",
  51879=>"011011000",
  51880=>"110110010",
  51881=>"110011110",
  51882=>"111011001",
  51883=>"111000000",
  51884=>"101010000",
  51885=>"111011001",
  51886=>"110000011",
  51887=>"100100100",
  51888=>"000010001",
  51889=>"101111001",
  51890=>"000100101",
  51891=>"111111111",
  51892=>"101101111",
  51893=>"011110000",
  51894=>"101010010",
  51895=>"010110100",
  51896=>"100100001",
  51897=>"100000110",
  51898=>"010110111",
  51899=>"010000001",
  51900=>"110001100",
  51901=>"001101010",
  51902=>"010001000",
  51903=>"010101110",
  51904=>"111101100",
  51905=>"000111101",
  51906=>"111010111",
  51907=>"100010000",
  51908=>"010001011",
  51909=>"011111001",
  51910=>"101101101",
  51911=>"110010010",
  51912=>"000111000",
  51913=>"100011101",
  51914=>"101000001",
  51915=>"101000001",
  51916=>"110000110",
  51917=>"111000001",
  51918=>"010010000",
  51919=>"001000111",
  51920=>"101000100",
  51921=>"001111111",
  51922=>"101000110",
  51923=>"001010110",
  51924=>"010111000",
  51925=>"000100001",
  51926=>"101101100",
  51927=>"000100000",
  51928=>"001110000",
  51929=>"111101000",
  51930=>"110001011",
  51931=>"111100011",
  51932=>"110000110",
  51933=>"111111011",
  51934=>"110101000",
  51935=>"111101101",
  51936=>"100010100",
  51937=>"011101111",
  51938=>"101111011",
  51939=>"110101100",
  51940=>"101000011",
  51941=>"110100110",
  51942=>"001000000",
  51943=>"101000000",
  51944=>"000011001",
  51945=>"101011011",
  51946=>"000101111",
  51947=>"100010001",
  51948=>"110000010",
  51949=>"011000101",
  51950=>"000111001",
  51951=>"001000111",
  51952=>"101111111",
  51953=>"010000000",
  51954=>"101011011",
  51955=>"001101100",
  51956=>"101111111",
  51957=>"011000110",
  51958=>"110100101",
  51959=>"011011101",
  51960=>"000001010",
  51961=>"011111001",
  51962=>"111010001",
  51963=>"001101110",
  51964=>"100100111",
  51965=>"100001011",
  51966=>"011111110",
  51967=>"010101001",
  51968=>"001010010",
  51969=>"110101001",
  51970=>"010101000",
  51971=>"000010011",
  51972=>"101011011",
  51973=>"010111000",
  51974=>"010001111",
  51975=>"101101111",
  51976=>"011011010",
  51977=>"010001101",
  51978=>"111010111",
  51979=>"001111010",
  51980=>"010001101",
  51981=>"010010010",
  51982=>"001101100",
  51983=>"010110100",
  51984=>"110000101",
  51985=>"110000111",
  51986=>"111101010",
  51987=>"001011111",
  51988=>"101000100",
  51989=>"010111101",
  51990=>"111110010",
  51991=>"111001001",
  51992=>"110110010",
  51993=>"011000111",
  51994=>"000011111",
  51995=>"000010110",
  51996=>"100001001",
  51997=>"001001100",
  51998=>"111100011",
  51999=>"001101101",
  52000=>"100111111",
  52001=>"111001100",
  52002=>"101110100",
  52003=>"110001110",
  52004=>"000001100",
  52005=>"111111110",
  52006=>"010001110",
  52007=>"111011011",
  52008=>"011001101",
  52009=>"001001111",
  52010=>"110101111",
  52011=>"011111110",
  52012=>"111110110",
  52013=>"100011100",
  52014=>"100100101",
  52015=>"110000111",
  52016=>"101000001",
  52017=>"000001110",
  52018=>"000100001",
  52019=>"001000000",
  52020=>"011000110",
  52021=>"000101101",
  52022=>"010000111",
  52023=>"111001001",
  52024=>"110101010",
  52025=>"100110010",
  52026=>"000101101",
  52027=>"100011101",
  52028=>"001000100",
  52029=>"100011000",
  52030=>"011001010",
  52031=>"000111110",
  52032=>"100101000",
  52033=>"101110011",
  52034=>"110010110",
  52035=>"001000000",
  52036=>"101000111",
  52037=>"010110001",
  52038=>"111110000",
  52039=>"101000100",
  52040=>"101010110",
  52041=>"000001100",
  52042=>"101010011",
  52043=>"001000001",
  52044=>"010100111",
  52045=>"110010110",
  52046=>"111010100",
  52047=>"101011101",
  52048=>"010101110",
  52049=>"000011011",
  52050=>"111010001",
  52051=>"110000011",
  52052=>"010000010",
  52053=>"001001001",
  52054=>"001011001",
  52055=>"111011001",
  52056=>"010001001",
  52057=>"011110110",
  52058=>"010000001",
  52059=>"010011010",
  52060=>"100001010",
  52061=>"001101010",
  52062=>"011000001",
  52063=>"000001111",
  52064=>"000000000",
  52065=>"010111010",
  52066=>"001011100",
  52067=>"000010101",
  52068=>"111010000",
  52069=>"011010010",
  52070=>"010001100",
  52071=>"110111011",
  52072=>"110111100",
  52073=>"000001011",
  52074=>"010001011",
  52075=>"000011010",
  52076=>"111111111",
  52077=>"000001000",
  52078=>"110100110",
  52079=>"010111010",
  52080=>"001100011",
  52081=>"011010011",
  52082=>"100101100",
  52083=>"010111110",
  52084=>"111010100",
  52085=>"010000010",
  52086=>"011100110",
  52087=>"101011101",
  52088=>"011100100",
  52089=>"000011101",
  52090=>"001001101",
  52091=>"111001001",
  52092=>"000010010",
  52093=>"011010100",
  52094=>"101011011",
  52095=>"110000111",
  52096=>"011101101",
  52097=>"111011111",
  52098=>"011001011",
  52099=>"101110110",
  52100=>"001111110",
  52101=>"111001111",
  52102=>"011010001",
  52103=>"010100000",
  52104=>"010001001",
  52105=>"110100100",
  52106=>"000010111",
  52107=>"011010000",
  52108=>"000000001",
  52109=>"110101011",
  52110=>"001001111",
  52111=>"011111000",
  52112=>"100101001",
  52113=>"010001111",
  52114=>"110000100",
  52115=>"100001011",
  52116=>"010011001",
  52117=>"111111111",
  52118=>"010011011",
  52119=>"101101001",
  52120=>"100100001",
  52121=>"010100000",
  52122=>"000010000",
  52123=>"000000111",
  52124=>"001101011",
  52125=>"001100101",
  52126=>"010011000",
  52127=>"000000110",
  52128=>"110000010",
  52129=>"110100011",
  52130=>"110000000",
  52131=>"010100100",
  52132=>"010000100",
  52133=>"101100000",
  52134=>"000000111",
  52135=>"111010001",
  52136=>"000000000",
  52137=>"001000110",
  52138=>"011011111",
  52139=>"001010000",
  52140=>"000010101",
  52141=>"010000101",
  52142=>"110101001",
  52143=>"101100010",
  52144=>"010110010",
  52145=>"110010110",
  52146=>"100111111",
  52147=>"100110011",
  52148=>"011000110",
  52149=>"011110101",
  52150=>"011101001",
  52151=>"010010001",
  52152=>"100101111",
  52153=>"111110010",
  52154=>"001110010",
  52155=>"101010000",
  52156=>"100100111",
  52157=>"101011001",
  52158=>"010100001",
  52159=>"010100001",
  52160=>"010011010",
  52161=>"111000110",
  52162=>"101111101",
  52163=>"110010111",
  52164=>"011011100",
  52165=>"010010011",
  52166=>"100111100",
  52167=>"110100100",
  52168=>"100000011",
  52169=>"111111111",
  52170=>"111111011",
  52171=>"110111111",
  52172=>"011101100",
  52173=>"010110111",
  52174=>"010100110",
  52175=>"011001010",
  52176=>"010010111",
  52177=>"100111000",
  52178=>"000110010",
  52179=>"110011000",
  52180=>"100010001",
  52181=>"000000000",
  52182=>"100101101",
  52183=>"000010011",
  52184=>"000001010",
  52185=>"100111010",
  52186=>"110100100",
  52187=>"000000000",
  52188=>"010000000",
  52189=>"000000100",
  52190=>"111100100",
  52191=>"011110011",
  52192=>"000010010",
  52193=>"110010110",
  52194=>"011010011",
  52195=>"111100000",
  52196=>"110001000",
  52197=>"100101010",
  52198=>"010001011",
  52199=>"100100100",
  52200=>"111001010",
  52201=>"000001110",
  52202=>"000011011",
  52203=>"011100011",
  52204=>"011101110",
  52205=>"101100001",
  52206=>"111010000",
  52207=>"010001100",
  52208=>"011101100",
  52209=>"101100000",
  52210=>"001111100",
  52211=>"110101100",
  52212=>"010111011",
  52213=>"010101000",
  52214=>"001001000",
  52215=>"110010001",
  52216=>"010100011",
  52217=>"101110010",
  52218=>"110011011",
  52219=>"100111011",
  52220=>"010011000",
  52221=>"101101001",
  52222=>"101101111",
  52223=>"000011110",
  52224=>"101101100",
  52225=>"100001111",
  52226=>"111010001",
  52227=>"001110011",
  52228=>"010000100",
  52229=>"010011011",
  52230=>"001101000",
  52231=>"100101111",
  52232=>"001001100",
  52233=>"000010101",
  52234=>"111000101",
  52235=>"001101110",
  52236=>"111000111",
  52237=>"000111100",
  52238=>"110110011",
  52239=>"000000000",
  52240=>"101101000",
  52241=>"110010001",
  52242=>"110011100",
  52243=>"010010111",
  52244=>"000001000",
  52245=>"010101011",
  52246=>"010010000",
  52247=>"000000001",
  52248=>"000101110",
  52249=>"000001001",
  52250=>"111101100",
  52251=>"111011111",
  52252=>"001101100",
  52253=>"100010010",
  52254=>"100010101",
  52255=>"010110000",
  52256=>"010100101",
  52257=>"000101110",
  52258=>"111110100",
  52259=>"000000010",
  52260=>"010001100",
  52261=>"011110000",
  52262=>"011000011",
  52263=>"001010011",
  52264=>"101010000",
  52265=>"110010100",
  52266=>"101100001",
  52267=>"110000011",
  52268=>"100111000",
  52269=>"001100010",
  52270=>"111011001",
  52271=>"001011011",
  52272=>"111011101",
  52273=>"010101011",
  52274=>"000001100",
  52275=>"111001101",
  52276=>"101101011",
  52277=>"100100100",
  52278=>"011110111",
  52279=>"011100110",
  52280=>"010010010",
  52281=>"000010101",
  52282=>"000001010",
  52283=>"010000110",
  52284=>"101010110",
  52285=>"011111001",
  52286=>"010011101",
  52287=>"000100010",
  52288=>"100001101",
  52289=>"000000000",
  52290=>"100000110",
  52291=>"000001000",
  52292=>"010001000",
  52293=>"100100011",
  52294=>"011111011",
  52295=>"101111010",
  52296=>"000111101",
  52297=>"011110100",
  52298=>"000000010",
  52299=>"001011011",
  52300=>"110111110",
  52301=>"001001011",
  52302=>"011110110",
  52303=>"100010011",
  52304=>"011111011",
  52305=>"100110101",
  52306=>"101011101",
  52307=>"111101011",
  52308=>"111011000",
  52309=>"000001100",
  52310=>"111011101",
  52311=>"100000110",
  52312=>"111100110",
  52313=>"111001101",
  52314=>"010100101",
  52315=>"001000101",
  52316=>"001011010",
  52317=>"000010111",
  52318=>"001000001",
  52319=>"100101110",
  52320=>"111000110",
  52321=>"000000000",
  52322=>"000011001",
  52323=>"110100101",
  52324=>"110101111",
  52325=>"111111101",
  52326=>"001000000",
  52327=>"001000111",
  52328=>"110101001",
  52329=>"111010101",
  52330=>"001010010",
  52331=>"000101010",
  52332=>"110000101",
  52333=>"101011110",
  52334=>"011100101",
  52335=>"111100101",
  52336=>"100101010",
  52337=>"110001000",
  52338=>"110011101",
  52339=>"100000110",
  52340=>"011111011",
  52341=>"001111000",
  52342=>"111101101",
  52343=>"100001110",
  52344=>"001010000",
  52345=>"110101111",
  52346=>"010110011",
  52347=>"000001100",
  52348=>"011110110",
  52349=>"110101100",
  52350=>"000001100",
  52351=>"011000001",
  52352=>"001101111",
  52353=>"010010011",
  52354=>"111111001",
  52355=>"111101110",
  52356=>"101100010",
  52357=>"110000100",
  52358=>"011010101",
  52359=>"110010111",
  52360=>"011100001",
  52361=>"110110110",
  52362=>"010010010",
  52363=>"111010001",
  52364=>"000001100",
  52365=>"010010111",
  52366=>"011011111",
  52367=>"011111011",
  52368=>"100110011",
  52369=>"011011011",
  52370=>"111101010",
  52371=>"000111010",
  52372=>"011000000",
  52373=>"000100110",
  52374=>"111010011",
  52375=>"111111111",
  52376=>"000111101",
  52377=>"001000000",
  52378=>"011000011",
  52379=>"011110001",
  52380=>"000100110",
  52381=>"001010011",
  52382=>"110111010",
  52383=>"101000010",
  52384=>"110010011",
  52385=>"111011100",
  52386=>"110011011",
  52387=>"001010101",
  52388=>"111110000",
  52389=>"101011101",
  52390=>"001101011",
  52391=>"000000100",
  52392=>"100111010",
  52393=>"100101100",
  52394=>"010011000",
  52395=>"000111001",
  52396=>"100001110",
  52397=>"111100000",
  52398=>"000001110",
  52399=>"010001111",
  52400=>"000110010",
  52401=>"100100010",
  52402=>"001010111",
  52403=>"000010000",
  52404=>"110000000",
  52405=>"000001001",
  52406=>"111000001",
  52407=>"110010101",
  52408=>"100101110",
  52409=>"010010110",
  52410=>"001101011",
  52411=>"111010100",
  52412=>"000110011",
  52413=>"110101101",
  52414=>"010010111",
  52415=>"110001010",
  52416=>"000010010",
  52417=>"100011011",
  52418=>"111000000",
  52419=>"101110111",
  52420=>"001111111",
  52421=>"000010011",
  52422=>"011011011",
  52423=>"000010100",
  52424=>"100111000",
  52425=>"000101011",
  52426=>"100010110",
  52427=>"010100110",
  52428=>"011110111",
  52429=>"000001110",
  52430=>"001000110",
  52431=>"000011001",
  52432=>"011101010",
  52433=>"001001110",
  52434=>"000101001",
  52435=>"001001100",
  52436=>"101101000",
  52437=>"000101100",
  52438=>"100110100",
  52439=>"011111111",
  52440=>"001101100",
  52441=>"001101110",
  52442=>"000110000",
  52443=>"111100110",
  52444=>"011101111",
  52445=>"011000110",
  52446=>"111111110",
  52447=>"110011010",
  52448=>"101100001",
  52449=>"001010010",
  52450=>"000100000",
  52451=>"001000001",
  52452=>"110010000",
  52453=>"011100000",
  52454=>"001000010",
  52455=>"111001010",
  52456=>"100100110",
  52457=>"100110000",
  52458=>"001001110",
  52459=>"000110011",
  52460=>"010011011",
  52461=>"101110110",
  52462=>"000010001",
  52463=>"110110111",
  52464=>"110010001",
  52465=>"000010000",
  52466=>"000000011",
  52467=>"000100111",
  52468=>"110100011",
  52469=>"011000100",
  52470=>"101110101",
  52471=>"110100010",
  52472=>"110000010",
  52473=>"000001010",
  52474=>"000101001",
  52475=>"000010001",
  52476=>"000001110",
  52477=>"011000010",
  52478=>"000101111",
  52479=>"000011101",
  52480=>"010110000",
  52481=>"010110010",
  52482=>"110010101",
  52483=>"010001100",
  52484=>"001010100",
  52485=>"010101111",
  52486=>"010110001",
  52487=>"111110101",
  52488=>"011011000",
  52489=>"101010110",
  52490=>"000010110",
  52491=>"101001111",
  52492=>"000111001",
  52493=>"111110011",
  52494=>"010001100",
  52495=>"011001110",
  52496=>"001101001",
  52497=>"001000110",
  52498=>"111101010",
  52499=>"000110101",
  52500=>"000111011",
  52501=>"010010110",
  52502=>"010010010",
  52503=>"010101011",
  52504=>"011110100",
  52505=>"001010000",
  52506=>"111111011",
  52507=>"010101011",
  52508=>"111111111",
  52509=>"101000100",
  52510=>"001011001",
  52511=>"010000100",
  52512=>"000010110",
  52513=>"101110001",
  52514=>"110111100",
  52515=>"001011110",
  52516=>"111000100",
  52517=>"110111101",
  52518=>"011111101",
  52519=>"011000001",
  52520=>"001001000",
  52521=>"001010111",
  52522=>"001010111",
  52523=>"101100100",
  52524=>"001110011",
  52525=>"001111111",
  52526=>"000100111",
  52527=>"100000111",
  52528=>"101100100",
  52529=>"100010011",
  52530=>"110000101",
  52531=>"101101010",
  52532=>"111000001",
  52533=>"111010011",
  52534=>"001000100",
  52535=>"111100011",
  52536=>"110000000",
  52537=>"000100101",
  52538=>"101010110",
  52539=>"011000100",
  52540=>"011010010",
  52541=>"101001111",
  52542=>"000010000",
  52543=>"001100010",
  52544=>"001000001",
  52545=>"000111010",
  52546=>"011101111",
  52547=>"010001010",
  52548=>"101001000",
  52549=>"010100000",
  52550=>"111001110",
  52551=>"100000111",
  52552=>"111010100",
  52553=>"000100010",
  52554=>"111111100",
  52555=>"110010001",
  52556=>"011101111",
  52557=>"011101000",
  52558=>"010010101",
  52559=>"001110101",
  52560=>"101010001",
  52561=>"001111001",
  52562=>"001000000",
  52563=>"011001010",
  52564=>"110111000",
  52565=>"111110010",
  52566=>"101100101",
  52567=>"011011100",
  52568=>"101101111",
  52569=>"110001010",
  52570=>"100001000",
  52571=>"000000010",
  52572=>"100110011",
  52573=>"011001110",
  52574=>"011111001",
  52575=>"010100100",
  52576=>"110000010",
  52577=>"001011100",
  52578=>"101101001",
  52579=>"000000101",
  52580=>"001111110",
  52581=>"010110001",
  52582=>"010010000",
  52583=>"010111000",
  52584=>"010001010",
  52585=>"001001011",
  52586=>"111111010",
  52587=>"000001000",
  52588=>"010100001",
  52589=>"110101111",
  52590=>"000001000",
  52591=>"100000010",
  52592=>"100000010",
  52593=>"001111010",
  52594=>"110001000",
  52595=>"110100000",
  52596=>"010100001",
  52597=>"000000101",
  52598=>"010101001",
  52599=>"110011000",
  52600=>"100001011",
  52601=>"110100011",
  52602=>"000000001",
  52603=>"011000111",
  52604=>"001110011",
  52605=>"010001000",
  52606=>"111010011",
  52607=>"000000000",
  52608=>"101001001",
  52609=>"010001011",
  52610=>"101011101",
  52611=>"001110010",
  52612=>"001000111",
  52613=>"010100010",
  52614=>"110111010",
  52615=>"000100011",
  52616=>"101110101",
  52617=>"010011101",
  52618=>"000000101",
  52619=>"110000111",
  52620=>"100000111",
  52621=>"100000111",
  52622=>"110100111",
  52623=>"000100001",
  52624=>"110101110",
  52625=>"010101111",
  52626=>"001110001",
  52627=>"111000111",
  52628=>"001110100",
  52629=>"000000100",
  52630=>"110000000",
  52631=>"101110011",
  52632=>"000110110",
  52633=>"000001000",
  52634=>"101001110",
  52635=>"111000111",
  52636=>"001000101",
  52637=>"111100000",
  52638=>"010110111",
  52639=>"101101001",
  52640=>"110110110",
  52641=>"111001101",
  52642=>"111011100",
  52643=>"001010111",
  52644=>"100000010",
  52645=>"000100010",
  52646=>"111001101",
  52647=>"011111000",
  52648=>"001010111",
  52649=>"001001101",
  52650=>"010011010",
  52651=>"111110100",
  52652=>"001101101",
  52653=>"000111001",
  52654=>"101000010",
  52655=>"111111110",
  52656=>"000010010",
  52657=>"010010000",
  52658=>"001110101",
  52659=>"110101011",
  52660=>"110100001",
  52661=>"111000101",
  52662=>"110111000",
  52663=>"000110010",
  52664=>"000100100",
  52665=>"100000111",
  52666=>"101000101",
  52667=>"001110011",
  52668=>"000110000",
  52669=>"010100111",
  52670=>"011000111",
  52671=>"010000000",
  52672=>"100000101",
  52673=>"011001011",
  52674=>"011011001",
  52675=>"111100111",
  52676=>"011011111",
  52677=>"101100000",
  52678=>"111100101",
  52679=>"111110000",
  52680=>"010010101",
  52681=>"111000001",
  52682=>"010001111",
  52683=>"001111110",
  52684=>"111000001",
  52685=>"110110010",
  52686=>"000011000",
  52687=>"100011101",
  52688=>"001101010",
  52689=>"001111001",
  52690=>"000101100",
  52691=>"000101100",
  52692=>"101110010",
  52693=>"011011001",
  52694=>"011001100",
  52695=>"100110011",
  52696=>"111100010",
  52697=>"010100100",
  52698=>"111111101",
  52699=>"110000000",
  52700=>"110110001",
  52701=>"011101100",
  52702=>"101000001",
  52703=>"100011011",
  52704=>"110100000",
  52705=>"011001010",
  52706=>"001001010",
  52707=>"000110101",
  52708=>"101010001",
  52709=>"100110010",
  52710=>"001100000",
  52711=>"101000111",
  52712=>"111110111",
  52713=>"100111110",
  52714=>"011001011",
  52715=>"001011010",
  52716=>"001100001",
  52717=>"000000111",
  52718=>"010000100",
  52719=>"011011011",
  52720=>"111010000",
  52721=>"110000011",
  52722=>"000001010",
  52723=>"101110110",
  52724=>"000111001",
  52725=>"000100111",
  52726=>"010011000",
  52727=>"010100000",
  52728=>"000000000",
  52729=>"111001111",
  52730=>"010100001",
  52731=>"100001100",
  52732=>"010110010",
  52733=>"010101100",
  52734=>"101101001",
  52735=>"101100011",
  52736=>"001010001",
  52737=>"111010010",
  52738=>"011011010",
  52739=>"100110010",
  52740=>"110110110",
  52741=>"101011101",
  52742=>"110110111",
  52743=>"000010101",
  52744=>"001011010",
  52745=>"001111110",
  52746=>"001111001",
  52747=>"000000010",
  52748=>"010011111",
  52749=>"100100101",
  52750=>"010001010",
  52751=>"011111101",
  52752=>"110001011",
  52753=>"100111110",
  52754=>"111111101",
  52755=>"101011101",
  52756=>"001001110",
  52757=>"100111011",
  52758=>"001100011",
  52759=>"101010100",
  52760=>"010000110",
  52761=>"011110100",
  52762=>"100010000",
  52763=>"101010011",
  52764=>"000001000",
  52765=>"110001011",
  52766=>"111100001",
  52767=>"101010111",
  52768=>"001011001",
  52769=>"101010010",
  52770=>"011101101",
  52771=>"101000000",
  52772=>"110101100",
  52773=>"101001110",
  52774=>"101100111",
  52775=>"111111100",
  52776=>"011110010",
  52777=>"000100110",
  52778=>"001111110",
  52779=>"101110000",
  52780=>"100000000",
  52781=>"000101101",
  52782=>"010111000",
  52783=>"011000011",
  52784=>"111001010",
  52785=>"011100000",
  52786=>"111111000",
  52787=>"000000100",
  52788=>"111000100",
  52789=>"001000111",
  52790=>"001010111",
  52791=>"010100111",
  52792=>"100001011",
  52793=>"000001100",
  52794=>"001100101",
  52795=>"101001110",
  52796=>"010011111",
  52797=>"010101110",
  52798=>"011011110",
  52799=>"001010110",
  52800=>"010000110",
  52801=>"011001000",
  52802=>"000001011",
  52803=>"100011011",
  52804=>"111010001",
  52805=>"000010101",
  52806=>"010101000",
  52807=>"110101000",
  52808=>"111101011",
  52809=>"101100100",
  52810=>"001000000",
  52811=>"010011000",
  52812=>"000101010",
  52813=>"100001010",
  52814=>"000100010",
  52815=>"001000111",
  52816=>"000000000",
  52817=>"110110010",
  52818=>"011111011",
  52819=>"000101011",
  52820=>"000111101",
  52821=>"000100011",
  52822=>"101010111",
  52823=>"010001111",
  52824=>"111011001",
  52825=>"111000001",
  52826=>"001100010",
  52827=>"010011101",
  52828=>"100001011",
  52829=>"010010010",
  52830=>"001000010",
  52831=>"001111101",
  52832=>"100110111",
  52833=>"001011010",
  52834=>"100101000",
  52835=>"100101011",
  52836=>"010110100",
  52837=>"110100011",
  52838=>"101010010",
  52839=>"101110011",
  52840=>"100111001",
  52841=>"011001011",
  52842=>"000101001",
  52843=>"000010110",
  52844=>"011001100",
  52845=>"010010000",
  52846=>"111011101",
  52847=>"011011011",
  52848=>"110001000",
  52849=>"001100010",
  52850=>"001100010",
  52851=>"110101110",
  52852=>"001001000",
  52853=>"010111111",
  52854=>"000000001",
  52855=>"001011110",
  52856=>"111110000",
  52857=>"010010001",
  52858=>"111011011",
  52859=>"100101100",
  52860=>"101111000",
  52861=>"001011010",
  52862=>"011110011",
  52863=>"001100010",
  52864=>"000011110",
  52865=>"100100101",
  52866=>"000001011",
  52867=>"001011111",
  52868=>"011101101",
  52869=>"110100011",
  52870=>"110101000",
  52871=>"111111111",
  52872=>"100100101",
  52873=>"100100010",
  52874=>"111111010",
  52875=>"011011101",
  52876=>"010110000",
  52877=>"001100011",
  52878=>"101111111",
  52879=>"001000000",
  52880=>"111100100",
  52881=>"011001001",
  52882=>"101011100",
  52883=>"101101101",
  52884=>"110010010",
  52885=>"010111111",
  52886=>"011100101",
  52887=>"110010110",
  52888=>"000010011",
  52889=>"111000000",
  52890=>"010100011",
  52891=>"101010011",
  52892=>"110110000",
  52893=>"000001001",
  52894=>"101011000",
  52895=>"011000010",
  52896=>"000000000",
  52897=>"001111001",
  52898=>"111110011",
  52899=>"101101110",
  52900=>"111001001",
  52901=>"010011011",
  52902=>"110000011",
  52903=>"000111000",
  52904=>"100001001",
  52905=>"111101110",
  52906=>"010001000",
  52907=>"101000111",
  52908=>"000001000",
  52909=>"000001000",
  52910=>"000100011",
  52911=>"110001000",
  52912=>"000000100",
  52913=>"010101001",
  52914=>"000111110",
  52915=>"101101010",
  52916=>"000010101",
  52917=>"001010010",
  52918=>"000100001",
  52919=>"000001111",
  52920=>"000111111",
  52921=>"000011111",
  52922=>"111010101",
  52923=>"101110011",
  52924=>"111011111",
  52925=>"000010100",
  52926=>"011001000",
  52927=>"000000101",
  52928=>"100010010",
  52929=>"011000110",
  52930=>"100011001",
  52931=>"110010100",
  52932=>"001111101",
  52933=>"010111011",
  52934=>"101011100",
  52935=>"100101100",
  52936=>"110000000",
  52937=>"010100111",
  52938=>"000100101",
  52939=>"010001110",
  52940=>"001010001",
  52941=>"010001111",
  52942=>"100100111",
  52943=>"110011111",
  52944=>"001110010",
  52945=>"101000101",
  52946=>"001110010",
  52947=>"100110111",
  52948=>"010001001",
  52949=>"100000111",
  52950=>"000011000",
  52951=>"001000001",
  52952=>"010000000",
  52953=>"100100111",
  52954=>"111000010",
  52955=>"101011011",
  52956=>"101100100",
  52957=>"111111110",
  52958=>"010101010",
  52959=>"100110101",
  52960=>"111111111",
  52961=>"010000111",
  52962=>"100001010",
  52963=>"001011001",
  52964=>"111001010",
  52965=>"110000111",
  52966=>"011001110",
  52967=>"110010111",
  52968=>"000001000",
  52969=>"101011110",
  52970=>"011001110",
  52971=>"011110000",
  52972=>"100000011",
  52973=>"100010101",
  52974=>"110100101",
  52975=>"101000000",
  52976=>"000001000",
  52977=>"100010001",
  52978=>"000001001",
  52979=>"010110011",
  52980=>"101011110",
  52981=>"000001011",
  52982=>"110100111",
  52983=>"100111100",
  52984=>"010010000",
  52985=>"100100110",
  52986=>"000000111",
  52987=>"010001001",
  52988=>"111000110",
  52989=>"001101111",
  52990=>"101100111",
  52991=>"011000000",
  52992=>"001110111",
  52993=>"000111010",
  52994=>"101111111",
  52995=>"100011001",
  52996=>"010100000",
  52997=>"101110110",
  52998=>"000100001",
  52999=>"011011000",
  53000=>"110001100",
  53001=>"011000001",
  53002=>"001010110",
  53003=>"100000100",
  53004=>"001100010",
  53005=>"110001001",
  53006=>"001110010",
  53007=>"000010100",
  53008=>"110011011",
  53009=>"011101011",
  53010=>"011100101",
  53011=>"100101100",
  53012=>"010001110",
  53013=>"101111001",
  53014=>"010010000",
  53015=>"111000101",
  53016=>"001001010",
  53017=>"000000000",
  53018=>"100001001",
  53019=>"100100010",
  53020=>"101011011",
  53021=>"001000110",
  53022=>"001011000",
  53023=>"101000011",
  53024=>"110011011",
  53025=>"011101010",
  53026=>"011011011",
  53027=>"110010110",
  53028=>"010000100",
  53029=>"010111010",
  53030=>"100110110",
  53031=>"000110110",
  53032=>"101010110",
  53033=>"000001111",
  53034=>"000111010",
  53035=>"010111010",
  53036=>"111000011",
  53037=>"000001010",
  53038=>"010100111",
  53039=>"011000100",
  53040=>"100000111",
  53041=>"000100011",
  53042=>"000011110",
  53043=>"111010011",
  53044=>"010100000",
  53045=>"000111000",
  53046=>"010011100",
  53047=>"100001100",
  53048=>"110111111",
  53049=>"100010110",
  53050=>"011101010",
  53051=>"011010000",
  53052=>"010010011",
  53053=>"100110011",
  53054=>"110010111",
  53055=>"011111101",
  53056=>"111011111",
  53057=>"110110000",
  53058=>"010000111",
  53059=>"110000110",
  53060=>"000000111",
  53061=>"001001000",
  53062=>"100110101",
  53063=>"010100010",
  53064=>"010110111",
  53065=>"100101111",
  53066=>"111001001",
  53067=>"001100101",
  53068=>"001110110",
  53069=>"110001100",
  53070=>"010010101",
  53071=>"110110111",
  53072=>"110000110",
  53073=>"111110110",
  53074=>"010010000",
  53075=>"001000111",
  53076=>"100010000",
  53077=>"100101000",
  53078=>"010010001",
  53079=>"111011010",
  53080=>"100010001",
  53081=>"010111001",
  53082=>"011001101",
  53083=>"011010010",
  53084=>"110101101",
  53085=>"101010111",
  53086=>"000000001",
  53087=>"000001010",
  53088=>"110100001",
  53089=>"010011000",
  53090=>"100010011",
  53091=>"011010001",
  53092=>"111000110",
  53093=>"000010010",
  53094=>"000000010",
  53095=>"011000001",
  53096=>"101001100",
  53097=>"100000111",
  53098=>"010000110",
  53099=>"011011110",
  53100=>"010100111",
  53101=>"010110010",
  53102=>"011000110",
  53103=>"001010101",
  53104=>"101101101",
  53105=>"000100001",
  53106=>"100010011",
  53107=>"100000111",
  53108=>"000000000",
  53109=>"000111011",
  53110=>"110010110",
  53111=>"110011100",
  53112=>"111010000",
  53113=>"011101010",
  53114=>"000101000",
  53115=>"100010101",
  53116=>"000000000",
  53117=>"100010111",
  53118=>"110010110",
  53119=>"101100010",
  53120=>"010111110",
  53121=>"001101100",
  53122=>"001011110",
  53123=>"011000111",
  53124=>"011010000",
  53125=>"111101111",
  53126=>"110100110",
  53127=>"000001100",
  53128=>"111001001",
  53129=>"110100111",
  53130=>"100000111",
  53131=>"100001100",
  53132=>"110010000",
  53133=>"011110110",
  53134=>"011111110",
  53135=>"010110100",
  53136=>"101111010",
  53137=>"100110111",
  53138=>"010110011",
  53139=>"010101110",
  53140=>"000101000",
  53141=>"010001100",
  53142=>"001000000",
  53143=>"110101110",
  53144=>"000000111",
  53145=>"001110010",
  53146=>"100110011",
  53147=>"110110001",
  53148=>"011110111",
  53149=>"100000110",
  53150=>"101011111",
  53151=>"111001001",
  53152=>"010010101",
  53153=>"000101101",
  53154=>"010110110",
  53155=>"101010010",
  53156=>"100010011",
  53157=>"111001100",
  53158=>"101011110",
  53159=>"011010111",
  53160=>"111101110",
  53161=>"010001010",
  53162=>"001101101",
  53163=>"100011010",
  53164=>"000011000",
  53165=>"001110110",
  53166=>"101100011",
  53167=>"101000000",
  53168=>"000111011",
  53169=>"000110111",
  53170=>"110110011",
  53171=>"100110000",
  53172=>"001100110",
  53173=>"100000011",
  53174=>"101111110",
  53175=>"110111111",
  53176=>"011000100",
  53177=>"100010110",
  53178=>"000101011",
  53179=>"110111100",
  53180=>"110100110",
  53181=>"001010110",
  53182=>"110001101",
  53183=>"101100110",
  53184=>"000100110",
  53185=>"101001011",
  53186=>"101100000",
  53187=>"100010000",
  53188=>"110010010",
  53189=>"101000011",
  53190=>"011111010",
  53191=>"001101100",
  53192=>"010100110",
  53193=>"010110001",
  53194=>"001110000",
  53195=>"110000010",
  53196=>"010110001",
  53197=>"010001000",
  53198=>"000000111",
  53199=>"100000101",
  53200=>"100110101",
  53201=>"001100010",
  53202=>"001000110",
  53203=>"101101011",
  53204=>"111001011",
  53205=>"001010010",
  53206=>"010001000",
  53207=>"000111000",
  53208=>"000000100",
  53209=>"110001100",
  53210=>"010001000",
  53211=>"010010111",
  53212=>"111100000",
  53213=>"111101000",
  53214=>"011100101",
  53215=>"011010011",
  53216=>"010100000",
  53217=>"111001101",
  53218=>"100100111",
  53219=>"100100100",
  53220=>"100000010",
  53221=>"100000100",
  53222=>"100001111",
  53223=>"001000011",
  53224=>"110111100",
  53225=>"010101010",
  53226=>"011100101",
  53227=>"010000101",
  53228=>"110001010",
  53229=>"000001001",
  53230=>"000110010",
  53231=>"010010011",
  53232=>"111111101",
  53233=>"001011101",
  53234=>"110000110",
  53235=>"100011101",
  53236=>"010001000",
  53237=>"001010010",
  53238=>"001101111",
  53239=>"111101001",
  53240=>"001011001",
  53241=>"100111001",
  53242=>"000110110",
  53243=>"101101100",
  53244=>"000100010",
  53245=>"100101000",
  53246=>"010001111",
  53247=>"110100001",
  53248=>"111111000",
  53249=>"110010111",
  53250=>"111101000",
  53251=>"001000001",
  53252=>"000001110",
  53253=>"000100110",
  53254=>"010001101",
  53255=>"011000001",
  53256=>"000101001",
  53257=>"011110101",
  53258=>"000001100",
  53259=>"001101100",
  53260=>"100011101",
  53261=>"000011010",
  53262=>"111011100",
  53263=>"001000101",
  53264=>"110011110",
  53265=>"001011111",
  53266=>"110001111",
  53267=>"100101110",
  53268=>"101111011",
  53269=>"000100000",
  53270=>"100011011",
  53271=>"000111010",
  53272=>"101000101",
  53273=>"101011001",
  53274=>"110010100",
  53275=>"100010101",
  53276=>"011110110",
  53277=>"000011000",
  53278=>"000111111",
  53279=>"011101111",
  53280=>"010001100",
  53281=>"000100000",
  53282=>"011111111",
  53283=>"110001110",
  53284=>"010001000",
  53285=>"110110100",
  53286=>"001111010",
  53287=>"000011110",
  53288=>"100011011",
  53289=>"001100001",
  53290=>"101100011",
  53291=>"111101011",
  53292=>"010101110",
  53293=>"101101000",
  53294=>"100100001",
  53295=>"000110001",
  53296=>"111111011",
  53297=>"000110111",
  53298=>"110011110",
  53299=>"011111100",
  53300=>"001010000",
  53301=>"101000110",
  53302=>"111011101",
  53303=>"100111100",
  53304=>"001100110",
  53305=>"110001000",
  53306=>"000111000",
  53307=>"111010111",
  53308=>"101001001",
  53309=>"100001100",
  53310=>"001111011",
  53311=>"010010011",
  53312=>"111110110",
  53313=>"011101111",
  53314=>"011101000",
  53315=>"011101110",
  53316=>"010101111",
  53317=>"111110111",
  53318=>"010000001",
  53319=>"000000101",
  53320=>"110001111",
  53321=>"111101011",
  53322=>"001100010",
  53323=>"011100001",
  53324=>"001001101",
  53325=>"000001110",
  53326=>"000101001",
  53327=>"111010110",
  53328=>"110000001",
  53329=>"001101110",
  53330=>"010101101",
  53331=>"110000110",
  53332=>"000100010",
  53333=>"100100000",
  53334=>"100110101",
  53335=>"011010101",
  53336=>"010111011",
  53337=>"010110100",
  53338=>"000101010",
  53339=>"001011000",
  53340=>"011100000",
  53341=>"000001001",
  53342=>"000011011",
  53343=>"000000000",
  53344=>"001100011",
  53345=>"111010111",
  53346=>"101101000",
  53347=>"000001010",
  53348=>"111001001",
  53349=>"000010110",
  53350=>"111100011",
  53351=>"100011000",
  53352=>"100011110",
  53353=>"110001010",
  53354=>"100001000",
  53355=>"001000101",
  53356=>"101000001",
  53357=>"010011111",
  53358=>"101000110",
  53359=>"101001001",
  53360=>"110000000",
  53361=>"000110111",
  53362=>"110000000",
  53363=>"101100101",
  53364=>"111010100",
  53365=>"000001100",
  53366=>"110001111",
  53367=>"010110100",
  53368=>"101111101",
  53369=>"110011010",
  53370=>"010010011",
  53371=>"000000000",
  53372=>"001110110",
  53373=>"101001010",
  53374=>"000010000",
  53375=>"001111000",
  53376=>"010000001",
  53377=>"110010011",
  53378=>"010111000",
  53379=>"100010001",
  53380=>"100000101",
  53381=>"100111111",
  53382=>"100101000",
  53383=>"111110111",
  53384=>"100000010",
  53385=>"010101111",
  53386=>"000110001",
  53387=>"110111111",
  53388=>"001000101",
  53389=>"001001001",
  53390=>"111011101",
  53391=>"000011000",
  53392=>"111000000",
  53393=>"110010011",
  53394=>"001101010",
  53395=>"110000101",
  53396=>"000000100",
  53397=>"110100101",
  53398=>"100111011",
  53399=>"000110110",
  53400=>"011011000",
  53401=>"110011010",
  53402=>"011100111",
  53403=>"010110000",
  53404=>"101111100",
  53405=>"101000000",
  53406=>"000010100",
  53407=>"111101011",
  53408=>"011010011",
  53409=>"100011110",
  53410=>"011110001",
  53411=>"101110010",
  53412=>"000111100",
  53413=>"001001110",
  53414=>"000011100",
  53415=>"000010111",
  53416=>"101101100",
  53417=>"000000000",
  53418=>"001000110",
  53419=>"011111010",
  53420=>"000110101",
  53421=>"010100011",
  53422=>"100111011",
  53423=>"000011101",
  53424=>"000111000",
  53425=>"001011010",
  53426=>"010100000",
  53427=>"100101101",
  53428=>"101000000",
  53429=>"001001111",
  53430=>"010010101",
  53431=>"110111101",
  53432=>"001000010",
  53433=>"001100010",
  53434=>"101100101",
  53435=>"010101111",
  53436=>"011010011",
  53437=>"001000110",
  53438=>"001001001",
  53439=>"101000000",
  53440=>"110011011",
  53441=>"010111000",
  53442=>"011011111",
  53443=>"101010010",
  53444=>"110101010",
  53445=>"100111010",
  53446=>"000100101",
  53447=>"001111101",
  53448=>"100011010",
  53449=>"000111111",
  53450=>"001110001",
  53451=>"000111100",
  53452=>"010101010",
  53453=>"111110111",
  53454=>"101111101",
  53455=>"000011110",
  53456=>"101100000",
  53457=>"101010110",
  53458=>"101110000",
  53459=>"001001001",
  53460=>"110001000",
  53461=>"000101000",
  53462=>"101101010",
  53463=>"100110000",
  53464=>"101010000",
  53465=>"110111000",
  53466=>"010000110",
  53467=>"110011100",
  53468=>"011001100",
  53469=>"100110001",
  53470=>"011001110",
  53471=>"011110000",
  53472=>"011110000",
  53473=>"111001011",
  53474=>"110100011",
  53475=>"111011100",
  53476=>"001100100",
  53477=>"110001111",
  53478=>"111000000",
  53479=>"001010000",
  53480=>"011110010",
  53481=>"100110101",
  53482=>"011011101",
  53483=>"001001100",
  53484=>"101100110",
  53485=>"010010101",
  53486=>"111001100",
  53487=>"101100101",
  53488=>"010001100",
  53489=>"101110011",
  53490=>"011000010",
  53491=>"000110110",
  53492=>"111011111",
  53493=>"011101110",
  53494=>"111110001",
  53495=>"001010011",
  53496=>"111011100",
  53497=>"011110010",
  53498=>"011111110",
  53499=>"100001000",
  53500=>"001011100",
  53501=>"001000100",
  53502=>"001010100",
  53503=>"110010010",
  53504=>"110101110",
  53505=>"001111001",
  53506=>"100001100",
  53507=>"000000100",
  53508=>"111111101",
  53509=>"001100100",
  53510=>"101000010",
  53511=>"111110001",
  53512=>"010110011",
  53513=>"011101010",
  53514=>"010110101",
  53515=>"101100110",
  53516=>"000111100",
  53517=>"001111000",
  53518=>"011111010",
  53519=>"010111100",
  53520=>"101010111",
  53521=>"101011101",
  53522=>"111010100",
  53523=>"000101100",
  53524=>"101001000",
  53525=>"001101010",
  53526=>"101110010",
  53527=>"000100000",
  53528=>"111111010",
  53529=>"011110001",
  53530=>"011110100",
  53531=>"011110001",
  53532=>"011011110",
  53533=>"110100100",
  53534=>"010000001",
  53535=>"110111001",
  53536=>"100011110",
  53537=>"010010110",
  53538=>"111110000",
  53539=>"100010110",
  53540=>"110110010",
  53541=>"011110011",
  53542=>"110011001",
  53543=>"110001110",
  53544=>"000101010",
  53545=>"000001100",
  53546=>"000000010",
  53547=>"000010011",
  53548=>"011000010",
  53549=>"010101000",
  53550=>"000100000",
  53551=>"111111101",
  53552=>"111101011",
  53553=>"000110110",
  53554=>"111011000",
  53555=>"110101000",
  53556=>"011000011",
  53557=>"011101111",
  53558=>"111101110",
  53559=>"101111111",
  53560=>"101100011",
  53561=>"100011100",
  53562=>"110101000",
  53563=>"110010111",
  53564=>"100001100",
  53565=>"100110101",
  53566=>"101101111",
  53567=>"001111011",
  53568=>"111100100",
  53569=>"111100001",
  53570=>"010111101",
  53571=>"011101111",
  53572=>"101001110",
  53573=>"100011101",
  53574=>"000111100",
  53575=>"100011011",
  53576=>"011010001",
  53577=>"001010111",
  53578=>"000110000",
  53579=>"001111110",
  53580=>"000011011",
  53581=>"000111011",
  53582=>"011000001",
  53583=>"100010010",
  53584=>"101001000",
  53585=>"100010110",
  53586=>"001110001",
  53587=>"111101110",
  53588=>"010010001",
  53589=>"011111111",
  53590=>"111011000",
  53591=>"001111111",
  53592=>"001011111",
  53593=>"100000011",
  53594=>"000011000",
  53595=>"100001000",
  53596=>"011101111",
  53597=>"011101001",
  53598=>"101011100",
  53599=>"001001101",
  53600=>"111100001",
  53601=>"101000001",
  53602=>"001110111",
  53603=>"001111001",
  53604=>"101000110",
  53605=>"001100001",
  53606=>"111011111",
  53607=>"100011101",
  53608=>"101001000",
  53609=>"000001000",
  53610=>"010101001",
  53611=>"101111001",
  53612=>"100001001",
  53613=>"101000000",
  53614=>"000100000",
  53615=>"010010011",
  53616=>"110110011",
  53617=>"011011101",
  53618=>"010011111",
  53619=>"010111000",
  53620=>"111100111",
  53621=>"010010101",
  53622=>"001000000",
  53623=>"001110000",
  53624=>"000111011",
  53625=>"000010101",
  53626=>"001100011",
  53627=>"000101000",
  53628=>"100111111",
  53629=>"111111110",
  53630=>"110010110",
  53631=>"010011011",
  53632=>"111101111",
  53633=>"000010100",
  53634=>"110011011",
  53635=>"001110111",
  53636=>"001001011",
  53637=>"100001101",
  53638=>"101011101",
  53639=>"110111011",
  53640=>"100101011",
  53641=>"100011100",
  53642=>"010010101",
  53643=>"001001000",
  53644=>"111101100",
  53645=>"000101100",
  53646=>"011011001",
  53647=>"000001010",
  53648=>"111111011",
  53649=>"100010001",
  53650=>"101001011",
  53651=>"111110000",
  53652=>"010010010",
  53653=>"101011100",
  53654=>"001010000",
  53655=>"011010011",
  53656=>"001001100",
  53657=>"001010001",
  53658=>"100011101",
  53659=>"101101111",
  53660=>"000011001",
  53661=>"010000000",
  53662=>"000100011",
  53663=>"110011001",
  53664=>"101100101",
  53665=>"000010001",
  53666=>"111010000",
  53667=>"000100010",
  53668=>"110111101",
  53669=>"011100000",
  53670=>"111000001",
  53671=>"111000111",
  53672=>"010111111",
  53673=>"010000001",
  53674=>"011110001",
  53675=>"010001001",
  53676=>"000100010",
  53677=>"101000100",
  53678=>"110010101",
  53679=>"000000001",
  53680=>"111111011",
  53681=>"000101001",
  53682=>"011000001",
  53683=>"110010001",
  53684=>"000001011",
  53685=>"011101001",
  53686=>"011001000",
  53687=>"111011101",
  53688=>"001001011",
  53689=>"100111101",
  53690=>"010101000",
  53691=>"101010110",
  53692=>"010100000",
  53693=>"110111100",
  53694=>"001011010",
  53695=>"010000110",
  53696=>"101110111",
  53697=>"000010010",
  53698=>"010111011",
  53699=>"001101000",
  53700=>"000000111",
  53701=>"001010000",
  53702=>"011011101",
  53703=>"100000000",
  53704=>"100000101",
  53705=>"010011010",
  53706=>"011010100",
  53707=>"000101101",
  53708=>"010011000",
  53709=>"110010011",
  53710=>"111100010",
  53711=>"101100110",
  53712=>"011110010",
  53713=>"000011001",
  53714=>"111001111",
  53715=>"001111110",
  53716=>"011110101",
  53717=>"111101001",
  53718=>"011110011",
  53719=>"000111011",
  53720=>"010000001",
  53721=>"101100010",
  53722=>"011010101",
  53723=>"011001001",
  53724=>"101010000",
  53725=>"111101100",
  53726=>"001100011",
  53727=>"111111111",
  53728=>"101101101",
  53729=>"000100011",
  53730=>"001001010",
  53731=>"000100101",
  53732=>"010010110",
  53733=>"101101100",
  53734=>"011110111",
  53735=>"001011000",
  53736=>"010000100",
  53737=>"100101110",
  53738=>"011100000",
  53739=>"100001000",
  53740=>"001001000",
  53741=>"110010110",
  53742=>"010010011",
  53743=>"000100010",
  53744=>"001010000",
  53745=>"101101000",
  53746=>"110011110",
  53747=>"011101011",
  53748=>"101111110",
  53749=>"010000010",
  53750=>"101011101",
  53751=>"100100100",
  53752=>"011111101",
  53753=>"111000111",
  53754=>"010111001",
  53755=>"011100010",
  53756=>"110111110",
  53757=>"001110001",
  53758=>"111101010",
  53759=>"100101011",
  53760=>"111010111",
  53761=>"010111100",
  53762=>"111100001",
  53763=>"100101000",
  53764=>"101001000",
  53765=>"110111110",
  53766=>"110011101",
  53767=>"010100100",
  53768=>"000000000",
  53769=>"011010101",
  53770=>"010111110",
  53771=>"101001100",
  53772=>"011001100",
  53773=>"010111011",
  53774=>"011001111",
  53775=>"100000100",
  53776=>"000010101",
  53777=>"001011110",
  53778=>"001000000",
  53779=>"101100111",
  53780=>"010011100",
  53781=>"110011110",
  53782=>"001111101",
  53783=>"100101110",
  53784=>"111100000",
  53785=>"100101100",
  53786=>"111111101",
  53787=>"000011111",
  53788=>"110001000",
  53789=>"110101100",
  53790=>"010100001",
  53791=>"101110001",
  53792=>"100110110",
  53793=>"000000101",
  53794=>"000110010",
  53795=>"110100110",
  53796=>"110001011",
  53797=>"101000000",
  53798=>"111111101",
  53799=>"011000100",
  53800=>"110000011",
  53801=>"001111000",
  53802=>"100100110",
  53803=>"001111100",
  53804=>"111100110",
  53805=>"010011000",
  53806=>"101101111",
  53807=>"001000010",
  53808=>"010010111",
  53809=>"111111111",
  53810=>"011111100",
  53811=>"100011010",
  53812=>"011000110",
  53813=>"100001101",
  53814=>"010110111",
  53815=>"111010000",
  53816=>"110100000",
  53817=>"101110101",
  53818=>"001100011",
  53819=>"100011110",
  53820=>"101101001",
  53821=>"011011110",
  53822=>"000000001",
  53823=>"000011100",
  53824=>"110010001",
  53825=>"011001001",
  53826=>"000100110",
  53827=>"101000010",
  53828=>"110110000",
  53829=>"100110000",
  53830=>"001100101",
  53831=>"000010101",
  53832=>"011110100",
  53833=>"011100110",
  53834=>"010111101",
  53835=>"110111101",
  53836=>"000101011",
  53837=>"111101100",
  53838=>"101010111",
  53839=>"101111000",
  53840=>"101100110",
  53841=>"011101101",
  53842=>"010101011",
  53843=>"011010000",
  53844=>"100101011",
  53845=>"100000101",
  53846=>"101010010",
  53847=>"011111010",
  53848=>"011010000",
  53849=>"100111001",
  53850=>"100010101",
  53851=>"110111111",
  53852=>"010010000",
  53853=>"000100001",
  53854=>"001001001",
  53855=>"010110111",
  53856=>"010011010",
  53857=>"100100001",
  53858=>"011111000",
  53859=>"001001111",
  53860=>"101111011",
  53861=>"110001010",
  53862=>"111001110",
  53863=>"001010111",
  53864=>"000000001",
  53865=>"000110001",
  53866=>"000010001",
  53867=>"010011101",
  53868=>"000010101",
  53869=>"011110101",
  53870=>"100001101",
  53871=>"011100100",
  53872=>"011111010",
  53873=>"000001000",
  53874=>"001100110",
  53875=>"001111111",
  53876=>"000000110",
  53877=>"101101111",
  53878=>"101010011",
  53879=>"100000110",
  53880=>"011100111",
  53881=>"110010011",
  53882=>"110010001",
  53883=>"110110100",
  53884=>"011101110",
  53885=>"010010001",
  53886=>"101111011",
  53887=>"011011100",
  53888=>"001101010",
  53889=>"000000010",
  53890=>"011011010",
  53891=>"011000011",
  53892=>"101011010",
  53893=>"101101111",
  53894=>"000110100",
  53895=>"100100000",
  53896=>"110110111",
  53897=>"111001000",
  53898=>"111111000",
  53899=>"101001100",
  53900=>"110101000",
  53901=>"010110011",
  53902=>"111001110",
  53903=>"000101010",
  53904=>"101001010",
  53905=>"011010111",
  53906=>"110101101",
  53907=>"101100000",
  53908=>"100101001",
  53909=>"100011010",
  53910=>"110101111",
  53911=>"101001001",
  53912=>"010100001",
  53913=>"000001110",
  53914=>"101000000",
  53915=>"010101001",
  53916=>"011010000",
  53917=>"010010101",
  53918=>"000111010",
  53919=>"110111111",
  53920=>"101010000",
  53921=>"100111100",
  53922=>"110110001",
  53923=>"101000000",
  53924=>"011001100",
  53925=>"111101101",
  53926=>"110100011",
  53927=>"101111000",
  53928=>"010101010",
  53929=>"011100111",
  53930=>"001111111",
  53931=>"000000111",
  53932=>"000010100",
  53933=>"000011100",
  53934=>"100010101",
  53935=>"001111110",
  53936=>"010101000",
  53937=>"000011001",
  53938=>"010110011",
  53939=>"101010100",
  53940=>"011001100",
  53941=>"101110110",
  53942=>"111011000",
  53943=>"111110001",
  53944=>"111111001",
  53945=>"010100011",
  53946=>"000011100",
  53947=>"110110100",
  53948=>"101111010",
  53949=>"000010011",
  53950=>"110001000",
  53951=>"010001101",
  53952=>"100101111",
  53953=>"010110111",
  53954=>"001111011",
  53955=>"111001110",
  53956=>"011111110",
  53957=>"000111010",
  53958=>"110111000",
  53959=>"111001111",
  53960=>"110111010",
  53961=>"100000011",
  53962=>"010010010",
  53963=>"011100000",
  53964=>"000000001",
  53965=>"010000011",
  53966=>"001111111",
  53967=>"010001001",
  53968=>"100011111",
  53969=>"001011110",
  53970=>"001000011",
  53971=>"111101000",
  53972=>"110100000",
  53973=>"001001000",
  53974=>"111100011",
  53975=>"100000101",
  53976=>"010110010",
  53977=>"011000101",
  53978=>"101100001",
  53979=>"001000001",
  53980=>"101110111",
  53981=>"111110101",
  53982=>"000100000",
  53983=>"111011111",
  53984=>"001100101",
  53985=>"011100111",
  53986=>"001101101",
  53987=>"000101001",
  53988=>"011101111",
  53989=>"011110100",
  53990=>"001101011",
  53991=>"001001011",
  53992=>"111110010",
  53993=>"000010101",
  53994=>"111001000",
  53995=>"010001101",
  53996=>"000011000",
  53997=>"011100110",
  53998=>"011000000",
  53999=>"000101100",
  54000=>"010000011",
  54001=>"011111001",
  54002=>"010110110",
  54003=>"100010101",
  54004=>"000010100",
  54005=>"100010000",
  54006=>"101110010",
  54007=>"011110100",
  54008=>"100010111",
  54009=>"111111111",
  54010=>"000001000",
  54011=>"011011000",
  54012=>"000101100",
  54013=>"100000011",
  54014=>"000010001",
  54015=>"000110101",
  54016=>"010100001",
  54017=>"111010000",
  54018=>"110111101",
  54019=>"101100101",
  54020=>"100010100",
  54021=>"110101011",
  54022=>"110110001",
  54023=>"000111000",
  54024=>"000010011",
  54025=>"010110001",
  54026=>"000010110",
  54027=>"010110110",
  54028=>"111000110",
  54029=>"010111011",
  54030=>"010011100",
  54031=>"010010000",
  54032=>"100100011",
  54033=>"000101111",
  54034=>"111010000",
  54035=>"011011111",
  54036=>"111001110",
  54037=>"010011111",
  54038=>"010100111",
  54039=>"100110011",
  54040=>"010100101",
  54041=>"000010111",
  54042=>"000010101",
  54043=>"101000010",
  54044=>"101010110",
  54045=>"001110100",
  54046=>"100100101",
  54047=>"010101010",
  54048=>"101110100",
  54049=>"111111011",
  54050=>"100001111",
  54051=>"001011011",
  54052=>"001101000",
  54053=>"001010011",
  54054=>"111101011",
  54055=>"000101000",
  54056=>"011101101",
  54057=>"100001110",
  54058=>"010000101",
  54059=>"010110110",
  54060=>"110010001",
  54061=>"010100101",
  54062=>"001011001",
  54063=>"000010111",
  54064=>"101111100",
  54065=>"100111000",
  54066=>"010110000",
  54067=>"000001010",
  54068=>"111101101",
  54069=>"101011011",
  54070=>"111010000",
  54071=>"101001101",
  54072=>"111100100",
  54073=>"011010010",
  54074=>"000111001",
  54075=>"111110101",
  54076=>"100011110",
  54077=>"110111001",
  54078=>"001101110",
  54079=>"101100101",
  54080=>"011110000",
  54081=>"100011011",
  54082=>"001101011",
  54083=>"111011111",
  54084=>"011001101",
  54085=>"111110010",
  54086=>"100011010",
  54087=>"111111101",
  54088=>"110110001",
  54089=>"111101110",
  54090=>"011100101",
  54091=>"001011000",
  54092=>"000010100",
  54093=>"101111000",
  54094=>"100100111",
  54095=>"011010000",
  54096=>"101100111",
  54097=>"100111000",
  54098=>"000100110",
  54099=>"111000101",
  54100=>"101100001",
  54101=>"000100001",
  54102=>"010000001",
  54103=>"100110000",
  54104=>"111001100",
  54105=>"000010011",
  54106=>"111111001",
  54107=>"000000100",
  54108=>"111101001",
  54109=>"111110011",
  54110=>"111100100",
  54111=>"011000000",
  54112=>"101110010",
  54113=>"101110111",
  54114=>"100000011",
  54115=>"101100011",
  54116=>"011001011",
  54117=>"110011010",
  54118=>"101111000",
  54119=>"111011101",
  54120=>"001100101",
  54121=>"011010001",
  54122=>"011011101",
  54123=>"111010000",
  54124=>"101100001",
  54125=>"110010001",
  54126=>"110010100",
  54127=>"001001010",
  54128=>"101010010",
  54129=>"110010111",
  54130=>"000101111",
  54131=>"110100110",
  54132=>"111011000",
  54133=>"100100100",
  54134=>"011101100",
  54135=>"011000010",
  54136=>"111111101",
  54137=>"110000011",
  54138=>"011000101",
  54139=>"000000101",
  54140=>"011011001",
  54141=>"001101111",
  54142=>"100001110",
  54143=>"010011001",
  54144=>"100111111",
  54145=>"101101110",
  54146=>"011000010",
  54147=>"010101000",
  54148=>"011011001",
  54149=>"110000101",
  54150=>"010011101",
  54151=>"101011001",
  54152=>"000010100",
  54153=>"011110001",
  54154=>"110010010",
  54155=>"000010001",
  54156=>"010110010",
  54157=>"010010001",
  54158=>"111101100",
  54159=>"111101110",
  54160=>"100011100",
  54161=>"100001101",
  54162=>"100001111",
  54163=>"101001001",
  54164=>"110001010",
  54165=>"011000010",
  54166=>"101001000",
  54167=>"110011110",
  54168=>"111100101",
  54169=>"001111001",
  54170=>"000001111",
  54171=>"100110110",
  54172=>"110111000",
  54173=>"000001010",
  54174=>"000111001",
  54175=>"010000000",
  54176=>"101101000",
  54177=>"001001111",
  54178=>"101001110",
  54179=>"000111011",
  54180=>"111010000",
  54181=>"110000000",
  54182=>"001000110",
  54183=>"011010011",
  54184=>"100101110",
  54185=>"100101111",
  54186=>"111111110",
  54187=>"000010010",
  54188=>"001010110",
  54189=>"110111010",
  54190=>"101011111",
  54191=>"101000011",
  54192=>"000100101",
  54193=>"111111111",
  54194=>"001001001",
  54195=>"000101011",
  54196=>"110000110",
  54197=>"101110010",
  54198=>"010011111",
  54199=>"101111011",
  54200=>"001100000",
  54201=>"001001111",
  54202=>"001111111",
  54203=>"000111100",
  54204=>"100111100",
  54205=>"101001101",
  54206=>"111000101",
  54207=>"011000000",
  54208=>"001010101",
  54209=>"101011001",
  54210=>"111001000",
  54211=>"101000111",
  54212=>"110100010",
  54213=>"100111101",
  54214=>"011001111",
  54215=>"100111010",
  54216=>"010010100",
  54217=>"000101001",
  54218=>"100001011",
  54219=>"001011000",
  54220=>"100100100",
  54221=>"100111100",
  54222=>"111011001",
  54223=>"100010000",
  54224=>"011001111",
  54225=>"010100110",
  54226=>"010000010",
  54227=>"010011000",
  54228=>"011000101",
  54229=>"100011010",
  54230=>"001011111",
  54231=>"111101111",
  54232=>"010111110",
  54233=>"111111100",
  54234=>"000001011",
  54235=>"011110011",
  54236=>"000001011",
  54237=>"000100101",
  54238=>"000000101",
  54239=>"111111100",
  54240=>"101100000",
  54241=>"100111111",
  54242=>"010001111",
  54243=>"110110101",
  54244=>"011010011",
  54245=>"100011100",
  54246=>"011011010",
  54247=>"001010010",
  54248=>"000100010",
  54249=>"110100101",
  54250=>"101111111",
  54251=>"111100010",
  54252=>"001010110",
  54253=>"011011100",
  54254=>"100010110",
  54255=>"110000110",
  54256=>"000000111",
  54257=>"100110000",
  54258=>"001011001",
  54259=>"101010010",
  54260=>"101010011",
  54261=>"010000000",
  54262=>"010010111",
  54263=>"110111100",
  54264=>"011001010",
  54265=>"001001110",
  54266=>"001111010",
  54267=>"111110101",
  54268=>"001011000",
  54269=>"101100100",
  54270=>"000100010",
  54271=>"100010001",
  54272=>"100010010",
  54273=>"100111001",
  54274=>"011010001",
  54275=>"101101101",
  54276=>"111001101",
  54277=>"000000111",
  54278=>"110110001",
  54279=>"000110101",
  54280=>"011010111",
  54281=>"110010101",
  54282=>"010010000",
  54283=>"110100001",
  54284=>"110001000",
  54285=>"111000001",
  54286=>"000001111",
  54287=>"100011101",
  54288=>"100010100",
  54289=>"101110100",
  54290=>"111010000",
  54291=>"100101101",
  54292=>"111100001",
  54293=>"001111110",
  54294=>"101100010",
  54295=>"111111111",
  54296=>"110001010",
  54297=>"101011011",
  54298=>"011010100",
  54299=>"001001101",
  54300=>"000001000",
  54301=>"010010111",
  54302=>"111001010",
  54303=>"100011111",
  54304=>"010011000",
  54305=>"100111010",
  54306=>"110101010",
  54307=>"110111001",
  54308=>"111000001",
  54309=>"000110111",
  54310=>"001000011",
  54311=>"010011000",
  54312=>"000111011",
  54313=>"111001001",
  54314=>"011001000",
  54315=>"100101101",
  54316=>"001110101",
  54317=>"011011101",
  54318=>"010000100",
  54319=>"111011011",
  54320=>"110011101",
  54321=>"101111111",
  54322=>"100011101",
  54323=>"100011000",
  54324=>"011111000",
  54325=>"101100101",
  54326=>"000011100",
  54327=>"110001110",
  54328=>"111101111",
  54329=>"110110010",
  54330=>"011000110",
  54331=>"110000111",
  54332=>"010000011",
  54333=>"011011110",
  54334=>"000101001",
  54335=>"111001111",
  54336=>"011011000",
  54337=>"110000001",
  54338=>"100110100",
  54339=>"010000001",
  54340=>"101001001",
  54341=>"000000100",
  54342=>"111000110",
  54343=>"111001011",
  54344=>"100100100",
  54345=>"000000111",
  54346=>"010100011",
  54347=>"001001000",
  54348=>"011100111",
  54349=>"110111111",
  54350=>"001100011",
  54351=>"110100100",
  54352=>"100001111",
  54353=>"010010001",
  54354=>"010110100",
  54355=>"010011100",
  54356=>"010000110",
  54357=>"101101111",
  54358=>"100000001",
  54359=>"000100000",
  54360=>"010111100",
  54361=>"111110111",
  54362=>"101110011",
  54363=>"011001110",
  54364=>"000000011",
  54365=>"111000011",
  54366=>"010010000",
  54367=>"101000111",
  54368=>"010100001",
  54369=>"011000110",
  54370=>"010110111",
  54371=>"000001011",
  54372=>"110000100",
  54373=>"110100011",
  54374=>"101000111",
  54375=>"111001111",
  54376=>"001100111",
  54377=>"110101111",
  54378=>"010100111",
  54379=>"010010100",
  54380=>"000100011",
  54381=>"110100011",
  54382=>"000111110",
  54383=>"011000010",
  54384=>"111110001",
  54385=>"001101001",
  54386=>"111010100",
  54387=>"000000111",
  54388=>"010101000",
  54389=>"010110110",
  54390=>"010101101",
  54391=>"001001000",
  54392=>"101000000",
  54393=>"010000010",
  54394=>"111111010",
  54395=>"000000101",
  54396=>"100010100",
  54397=>"101000110",
  54398=>"111010000",
  54399=>"110011101",
  54400=>"100100000",
  54401=>"110101010",
  54402=>"111101010",
  54403=>"001101101",
  54404=>"010111000",
  54405=>"011010011",
  54406=>"100100110",
  54407=>"001010000",
  54408=>"000000000",
  54409=>"000110010",
  54410=>"000111110",
  54411=>"001100011",
  54412=>"110000011",
  54413=>"001001100",
  54414=>"000100001",
  54415=>"100101101",
  54416=>"001011111",
  54417=>"001101010",
  54418=>"000000011",
  54419=>"101101000",
  54420=>"001101000",
  54421=>"010010000",
  54422=>"100001010",
  54423=>"111110111",
  54424=>"100001111",
  54425=>"101010000",
  54426=>"010011000",
  54427=>"010010001",
  54428=>"000100100",
  54429=>"111111101",
  54430=>"001111111",
  54431=>"001100100",
  54432=>"011010000",
  54433=>"101010010",
  54434=>"100010001",
  54435=>"001000011",
  54436=>"110111110",
  54437=>"001010010",
  54438=>"101001110",
  54439=>"001010100",
  54440=>"011101101",
  54441=>"011011010",
  54442=>"000010011",
  54443=>"110110110",
  54444=>"100100001",
  54445=>"001110011",
  54446=>"111011100",
  54447=>"100011101",
  54448=>"100110001",
  54449=>"011001111",
  54450=>"000100001",
  54451=>"100111010",
  54452=>"111100000",
  54453=>"101000101",
  54454=>"101101111",
  54455=>"101111101",
  54456=>"101011000",
  54457=>"011101101",
  54458=>"101101000",
  54459=>"001110000",
  54460=>"001001100",
  54461=>"010000100",
  54462=>"111101011",
  54463=>"101101110",
  54464=>"111001111",
  54465=>"000101010",
  54466=>"010100100",
  54467=>"100000100",
  54468=>"101110100",
  54469=>"111101001",
  54470=>"011010010",
  54471=>"101100110",
  54472=>"100000000",
  54473=>"001010010",
  54474=>"100010010",
  54475=>"001001011",
  54476=>"110111110",
  54477=>"000111001",
  54478=>"101111100",
  54479=>"101111100",
  54480=>"010110010",
  54481=>"100101010",
  54482=>"110001110",
  54483=>"001110101",
  54484=>"000001011",
  54485=>"011011110",
  54486=>"010111010",
  54487=>"001010010",
  54488=>"000000101",
  54489=>"101110110",
  54490=>"111111010",
  54491=>"100110011",
  54492=>"000010011",
  54493=>"100010011",
  54494=>"001110101",
  54495=>"010100010",
  54496=>"011110001",
  54497=>"011111110",
  54498=>"111011111",
  54499=>"011000110",
  54500=>"110111010",
  54501=>"100111101",
  54502=>"000100001",
  54503=>"100111010",
  54504=>"110000100",
  54505=>"101001100",
  54506=>"101001101",
  54507=>"011100111",
  54508=>"010100100",
  54509=>"111010100",
  54510=>"111000100",
  54511=>"000101010",
  54512=>"010000010",
  54513=>"000101000",
  54514=>"110110000",
  54515=>"001000001",
  54516=>"000011001",
  54517=>"000010001",
  54518=>"101100111",
  54519=>"001100000",
  54520=>"111010011",
  54521=>"001010011",
  54522=>"110010011",
  54523=>"001111000",
  54524=>"000000010",
  54525=>"110001001",
  54526=>"111011000",
  54527=>"111101101",
  54528=>"001111110",
  54529=>"111010101",
  54530=>"000111110",
  54531=>"010111011",
  54532=>"000010101",
  54533=>"111110100",
  54534=>"111011111",
  54535=>"110101011",
  54536=>"111001001",
  54537=>"000010010",
  54538=>"111011011",
  54539=>"101000101",
  54540=>"111011101",
  54541=>"101110101",
  54542=>"001001110",
  54543=>"101110110",
  54544=>"000001110",
  54545=>"100111110",
  54546=>"111101111",
  54547=>"000010010",
  54548=>"100001101",
  54549=>"110101000",
  54550=>"000001010",
  54551=>"110111110",
  54552=>"110000101",
  54553=>"111111010",
  54554=>"000100011",
  54555=>"001100100",
  54556=>"010000101",
  54557=>"101111011",
  54558=>"011011100",
  54559=>"000000110",
  54560=>"011000000",
  54561=>"101111011",
  54562=>"111011100",
  54563=>"000111101",
  54564=>"000000000",
  54565=>"011010000",
  54566=>"100001001",
  54567=>"101100101",
  54568=>"010011001",
  54569=>"000100001",
  54570=>"101001001",
  54571=>"110010111",
  54572=>"100011001",
  54573=>"000010100",
  54574=>"101000110",
  54575=>"001110001",
  54576=>"111100101",
  54577=>"101100011",
  54578=>"100111111",
  54579=>"111000010",
  54580=>"001000010",
  54581=>"000111010",
  54582=>"011110101",
  54583=>"000111111",
  54584=>"101001000",
  54585=>"100010011",
  54586=>"101000101",
  54587=>"111111000",
  54588=>"100001110",
  54589=>"111101000",
  54590=>"110100011",
  54591=>"101000000",
  54592=>"100011101",
  54593=>"110001010",
  54594=>"010010111",
  54595=>"100000111",
  54596=>"000110000",
  54597=>"000010010",
  54598=>"110000011",
  54599=>"100000100",
  54600=>"100001000",
  54601=>"110101100",
  54602=>"000110111",
  54603=>"000000111",
  54604=>"100011110",
  54605=>"000001100",
  54606=>"100101110",
  54607=>"011110011",
  54608=>"100001010",
  54609=>"100000111",
  54610=>"001001000",
  54611=>"001001000",
  54612=>"111110011",
  54613=>"100100110",
  54614=>"001000101",
  54615=>"100111010",
  54616=>"110011100",
  54617=>"010010011",
  54618=>"010001010",
  54619=>"000101101",
  54620=>"001100110",
  54621=>"100011100",
  54622=>"111110100",
  54623=>"111010001",
  54624=>"010101101",
  54625=>"111100111",
  54626=>"110001010",
  54627=>"011100101",
  54628=>"001011001",
  54629=>"001001011",
  54630=>"011110011",
  54631=>"000000011",
  54632=>"010101101",
  54633=>"111100011",
  54634=>"111011111",
  54635=>"100101000",
  54636=>"101100010",
  54637=>"001011100",
  54638=>"100001010",
  54639=>"001100010",
  54640=>"000100110",
  54641=>"011111011",
  54642=>"101011111",
  54643=>"111000011",
  54644=>"100000101",
  54645=>"100101101",
  54646=>"101100100",
  54647=>"110101101",
  54648=>"000100010",
  54649=>"001011111",
  54650=>"001101111",
  54651=>"000010011",
  54652=>"110000111",
  54653=>"100000000",
  54654=>"101111010",
  54655=>"001011001",
  54656=>"110000010",
  54657=>"101010011",
  54658=>"101111111",
  54659=>"001011100",
  54660=>"000100010",
  54661=>"111110001",
  54662=>"001111010",
  54663=>"011000000",
  54664=>"000001000",
  54665=>"111010111",
  54666=>"111110011",
  54667=>"000111110",
  54668=>"100000010",
  54669=>"111000001",
  54670=>"101011111",
  54671=>"111100000",
  54672=>"011011101",
  54673=>"111000010",
  54674=>"111110110",
  54675=>"011100010",
  54676=>"100111001",
  54677=>"000001001",
  54678=>"010100000",
  54679=>"100010000",
  54680=>"000101110",
  54681=>"101000101",
  54682=>"111010011",
  54683=>"110000100",
  54684=>"110000111",
  54685=>"101111000",
  54686=>"111001000",
  54687=>"100110010",
  54688=>"000000010",
  54689=>"111101110",
  54690=>"100111000",
  54691=>"011110011",
  54692=>"010000101",
  54693=>"100100011",
  54694=>"010101100",
  54695=>"110011101",
  54696=>"011110000",
  54697=>"000010111",
  54698=>"001110101",
  54699=>"100001001",
  54700=>"110011001",
  54701=>"100110010",
  54702=>"110100111",
  54703=>"101010011",
  54704=>"100101111",
  54705=>"100111000",
  54706=>"000010111",
  54707=>"101100010",
  54708=>"110011110",
  54709=>"011101101",
  54710=>"001011110",
  54711=>"010111000",
  54712=>"011100101",
  54713=>"100000100",
  54714=>"111111101",
  54715=>"110000101",
  54716=>"011011011",
  54717=>"001011011",
  54718=>"010100010",
  54719=>"011111000",
  54720=>"101110001",
  54721=>"111110111",
  54722=>"110010101",
  54723=>"110100010",
  54724=>"000000011",
  54725=>"011011100",
  54726=>"101100100",
  54727=>"011100110",
  54728=>"111111010",
  54729=>"110010010",
  54730=>"110111110",
  54731=>"100011011",
  54732=>"111010100",
  54733=>"010011001",
  54734=>"000100100",
  54735=>"111001110",
  54736=>"001110011",
  54737=>"000110001",
  54738=>"011001110",
  54739=>"001110001",
  54740=>"000011010",
  54741=>"010100101",
  54742=>"000010000",
  54743=>"110001100",
  54744=>"010100110",
  54745=>"011100111",
  54746=>"010000101",
  54747=>"000111001",
  54748=>"101011101",
  54749=>"100100011",
  54750=>"000111011",
  54751=>"100111110",
  54752=>"011001100",
  54753=>"000111001",
  54754=>"000111001",
  54755=>"010100001",
  54756=>"011011110",
  54757=>"011110011",
  54758=>"110011110",
  54759=>"110001101",
  54760=>"100101000",
  54761=>"100100111",
  54762=>"111110100",
  54763=>"101011110",
  54764=>"000011000",
  54765=>"100011100",
  54766=>"001101110",
  54767=>"110110000",
  54768=>"111101111",
  54769=>"110011111",
  54770=>"001111101",
  54771=>"001001001",
  54772=>"101110100",
  54773=>"011001101",
  54774=>"111000001",
  54775=>"101101001",
  54776=>"101111000",
  54777=>"010110110",
  54778=>"000101110",
  54779=>"000010101",
  54780=>"111111110",
  54781=>"110000001",
  54782=>"010001000",
  54783=>"000011001",
  54784=>"011010110",
  54785=>"001110011",
  54786=>"101101100",
  54787=>"111001010",
  54788=>"100011100",
  54789=>"100011011",
  54790=>"100000010",
  54791=>"100010001",
  54792=>"000101101",
  54793=>"111001110",
  54794=>"000010110",
  54795=>"001010100",
  54796=>"001111100",
  54797=>"110000111",
  54798=>"101001110",
  54799=>"111010010",
  54800=>"100100110",
  54801=>"100000000",
  54802=>"001100000",
  54803=>"000101000",
  54804=>"011110110",
  54805=>"011001011",
  54806=>"110001000",
  54807=>"000011011",
  54808=>"010100010",
  54809=>"011101011",
  54810=>"010011000",
  54811=>"000101000",
  54812=>"011011100",
  54813=>"111111110",
  54814=>"010111110",
  54815=>"110011100",
  54816=>"111100010",
  54817=>"101111111",
  54818=>"101000001",
  54819=>"001111000",
  54820=>"110111101",
  54821=>"000001000",
  54822=>"111111111",
  54823=>"101011010",
  54824=>"000111011",
  54825=>"100001111",
  54826=>"110100000",
  54827=>"111101001",
  54828=>"001001000",
  54829=>"111110111",
  54830=>"001011111",
  54831=>"111001101",
  54832=>"000000001",
  54833=>"100011011",
  54834=>"100010000",
  54835=>"110101111",
  54836=>"010001010",
  54837=>"001111101",
  54838=>"010011000",
  54839=>"100001101",
  54840=>"111111001",
  54841=>"010111010",
  54842=>"101000010",
  54843=>"101101111",
  54844=>"000000110",
  54845=>"110010110",
  54846=>"000101101",
  54847=>"010111011",
  54848=>"111110111",
  54849=>"101011110",
  54850=>"000100000",
  54851=>"000100001",
  54852=>"011000110",
  54853=>"111101100",
  54854=>"100001101",
  54855=>"011000101",
  54856=>"010010000",
  54857=>"100011100",
  54858=>"001111111",
  54859=>"001011100",
  54860=>"100000100",
  54861=>"111111111",
  54862=>"010101100",
  54863=>"000010100",
  54864=>"011100000",
  54865=>"010100100",
  54866=>"001001100",
  54867=>"000110100",
  54868=>"111010100",
  54869=>"101010111",
  54870=>"111011111",
  54871=>"000100010",
  54872=>"101011001",
  54873=>"010001110",
  54874=>"110000100",
  54875=>"111110000",
  54876=>"000011001",
  54877=>"110000010",
  54878=>"100100101",
  54879=>"111100100",
  54880=>"100000000",
  54881=>"010101010",
  54882=>"010010100",
  54883=>"100100001",
  54884=>"010101101",
  54885=>"001001100",
  54886=>"111011001",
  54887=>"100000101",
  54888=>"001000110",
  54889=>"111111011",
  54890=>"110100000",
  54891=>"000110110",
  54892=>"011101010",
  54893=>"111111110",
  54894=>"110111111",
  54895=>"000010110",
  54896=>"011010101",
  54897=>"110101011",
  54898=>"101111011",
  54899=>"000001111",
  54900=>"001101010",
  54901=>"011111000",
  54902=>"110011011",
  54903=>"000111011",
  54904=>"110110010",
  54905=>"000000001",
  54906=>"110011000",
  54907=>"001000111",
  54908=>"110110001",
  54909=>"110110001",
  54910=>"010100101",
  54911=>"011100100",
  54912=>"011100001",
  54913=>"001011101",
  54914=>"101000010",
  54915=>"011110011",
  54916=>"111010111",
  54917=>"111011111",
  54918=>"101110001",
  54919=>"100011111",
  54920=>"101100001",
  54921=>"011011001",
  54922=>"011000101",
  54923=>"001000110",
  54924=>"000110101",
  54925=>"100011011",
  54926=>"000011111",
  54927=>"001001101",
  54928=>"111010001",
  54929=>"000011100",
  54930=>"001000000",
  54931=>"111000000",
  54932=>"110001110",
  54933=>"001101010",
  54934=>"011111011",
  54935=>"100110010",
  54936=>"100000101",
  54937=>"100000110",
  54938=>"001000011",
  54939=>"000010011",
  54940=>"110011011",
  54941=>"111101101",
  54942=>"111111111",
  54943=>"011000000",
  54944=>"111001001",
  54945=>"000000010",
  54946=>"101111011",
  54947=>"101110111",
  54948=>"110100100",
  54949=>"101000000",
  54950=>"101001111",
  54951=>"011100011",
  54952=>"110110101",
  54953=>"101100110",
  54954=>"100111010",
  54955=>"110011110",
  54956=>"110101000",
  54957=>"001110100",
  54958=>"111111001",
  54959=>"110011100",
  54960=>"101100011",
  54961=>"111101001",
  54962=>"001110101",
  54963=>"111001011",
  54964=>"000001111",
  54965=>"001000010",
  54966=>"110011010",
  54967=>"111011100",
  54968=>"010000001",
  54969=>"011001100",
  54970=>"111111011",
  54971=>"010000101",
  54972=>"010000010",
  54973=>"111001110",
  54974=>"010101100",
  54975=>"011111101",
  54976=>"111000000",
  54977=>"101101011",
  54978=>"111011101",
  54979=>"000011100",
  54980=>"001011001",
  54981=>"011010011",
  54982=>"000000000",
  54983=>"100000011",
  54984=>"100110011",
  54985=>"100100001",
  54986=>"010111110",
  54987=>"110111010",
  54988=>"001101011",
  54989=>"110101111",
  54990=>"000100110",
  54991=>"001010100",
  54992=>"001101011",
  54993=>"001011100",
  54994=>"010010001",
  54995=>"010011110",
  54996=>"001000101",
  54997=>"100101101",
  54998=>"011001011",
  54999=>"000011110",
  55000=>"100100110",
  55001=>"110110010",
  55002=>"110111011",
  55003=>"101100010",
  55004=>"011110000",
  55005=>"010101101",
  55006=>"000001100",
  55007=>"001101000",
  55008=>"000000111",
  55009=>"011001111",
  55010=>"010011000",
  55011=>"100010000",
  55012=>"000001000",
  55013=>"011100011",
  55014=>"010011000",
  55015=>"000000001",
  55016=>"001101001",
  55017=>"100110110",
  55018=>"000011110",
  55019=>"000101111",
  55020=>"111110001",
  55021=>"101110011",
  55022=>"111011010",
  55023=>"111101111",
  55024=>"100111100",
  55025=>"110101000",
  55026=>"001010100",
  55027=>"100000010",
  55028=>"011001010",
  55029=>"001101011",
  55030=>"010010110",
  55031=>"000000010",
  55032=>"010000110",
  55033=>"110000011",
  55034=>"111011100",
  55035=>"111011101",
  55036=>"111110110",
  55037=>"001001110",
  55038=>"101111100",
  55039=>"111000101",
  55040=>"111111101",
  55041=>"000010110",
  55042=>"000101010",
  55043=>"110101010",
  55044=>"011011000",
  55045=>"100001100",
  55046=>"011000000",
  55047=>"010011100",
  55048=>"111100001",
  55049=>"001010111",
  55050=>"011100010",
  55051=>"100001000",
  55052=>"001001100",
  55053=>"101011000",
  55054=>"011110010",
  55055=>"111101110",
  55056=>"101010011",
  55057=>"010000011",
  55058=>"011011111",
  55059=>"100010101",
  55060=>"111011100",
  55061=>"110110011",
  55062=>"011110111",
  55063=>"001111100",
  55064=>"101101101",
  55065=>"101100001",
  55066=>"101001001",
  55067=>"100010100",
  55068=>"111010001",
  55069=>"010000101",
  55070=>"100010001",
  55071=>"010100001",
  55072=>"110111101",
  55073=>"110000000",
  55074=>"000000110",
  55075=>"100010100",
  55076=>"110001001",
  55077=>"110100011",
  55078=>"011110111",
  55079=>"010011100",
  55080=>"001010011",
  55081=>"111000011",
  55082=>"000010001",
  55083=>"010010100",
  55084=>"001011100",
  55085=>"000001100",
  55086=>"101100100",
  55087=>"010101100",
  55088=>"000101111",
  55089=>"011110011",
  55090=>"110110010",
  55091=>"110000011",
  55092=>"101110110",
  55093=>"101110110",
  55094=>"110010011",
  55095=>"000001100",
  55096=>"000010010",
  55097=>"000000101",
  55098=>"011101111",
  55099=>"111011101",
  55100=>"010110100",
  55101=>"011100011",
  55102=>"010001111",
  55103=>"000111100",
  55104=>"000100100",
  55105=>"010100001",
  55106=>"010000011",
  55107=>"010000101",
  55108=>"011011001",
  55109=>"010011111",
  55110=>"101001111",
  55111=>"101010000",
  55112=>"011011011",
  55113=>"010101111",
  55114=>"001000111",
  55115=>"001101111",
  55116=>"011110011",
  55117=>"100111111",
  55118=>"011000000",
  55119=>"110000001",
  55120=>"111110011",
  55121=>"001110010",
  55122=>"111011101",
  55123=>"100101000",
  55124=>"110110010",
  55125=>"111100111",
  55126=>"010110101",
  55127=>"110011111",
  55128=>"000000000",
  55129=>"101101101",
  55130=>"100100101",
  55131=>"011000001",
  55132=>"000000010",
  55133=>"001100110",
  55134=>"111000000",
  55135=>"100101011",
  55136=>"111011000",
  55137=>"010101011",
  55138=>"101110000",
  55139=>"111111011",
  55140=>"110001010",
  55141=>"100110110",
  55142=>"100000001",
  55143=>"101101101",
  55144=>"111101110",
  55145=>"011000110",
  55146=>"010010111",
  55147=>"001100011",
  55148=>"111000011",
  55149=>"110110010",
  55150=>"011110111",
  55151=>"010010100",
  55152=>"000100001",
  55153=>"001110010",
  55154=>"011110100",
  55155=>"110101111",
  55156=>"000011010",
  55157=>"110011111",
  55158=>"001011111",
  55159=>"101111000",
  55160=>"001101000",
  55161=>"101101011",
  55162=>"010111010",
  55163=>"011100101",
  55164=>"011100000",
  55165=>"010111011",
  55166=>"110000100",
  55167=>"011100110",
  55168=>"101010000",
  55169=>"001100011",
  55170=>"000110010",
  55171=>"101011101",
  55172=>"011110011",
  55173=>"010100000",
  55174=>"001001101",
  55175=>"100010000",
  55176=>"111011001",
  55177=>"111000011",
  55178=>"010010000",
  55179=>"110001000",
  55180=>"000000011",
  55181=>"101101100",
  55182=>"001000001",
  55183=>"111111100",
  55184=>"101100000",
  55185=>"000011010",
  55186=>"111000001",
  55187=>"101110111",
  55188=>"101001000",
  55189=>"101011100",
  55190=>"001001101",
  55191=>"000010000",
  55192=>"110000100",
  55193=>"000101001",
  55194=>"001011101",
  55195=>"101100000",
  55196=>"001011100",
  55197=>"000011100",
  55198=>"110011011",
  55199=>"010100110",
  55200=>"011001101",
  55201=>"001001110",
  55202=>"011001110",
  55203=>"000001111",
  55204=>"000000110",
  55205=>"001011101",
  55206=>"001100101",
  55207=>"011000001",
  55208=>"100001001",
  55209=>"010010100",
  55210=>"000010000",
  55211=>"011100011",
  55212=>"001100100",
  55213=>"111011110",
  55214=>"000001101",
  55215=>"000111001",
  55216=>"100101000",
  55217=>"100010011",
  55218=>"010111011",
  55219=>"011110000",
  55220=>"110011111",
  55221=>"010100000",
  55222=>"100001000",
  55223=>"010010101",
  55224=>"110010111",
  55225=>"111010101",
  55226=>"000011100",
  55227=>"011010101",
  55228=>"010110011",
  55229=>"110011001",
  55230=>"001110110",
  55231=>"110110000",
  55232=>"010001010",
  55233=>"101001000",
  55234=>"110101110",
  55235=>"000100111",
  55236=>"011111000",
  55237=>"100100100",
  55238=>"100100011",
  55239=>"110100100",
  55240=>"111111010",
  55241=>"010100000",
  55242=>"110110010",
  55243=>"100011101",
  55244=>"110100101",
  55245=>"000100011",
  55246=>"000111110",
  55247=>"011000101",
  55248=>"111100010",
  55249=>"101000010",
  55250=>"111011110",
  55251=>"000010110",
  55252=>"001111111",
  55253=>"011000101",
  55254=>"101111011",
  55255=>"000101011",
  55256=>"000000011",
  55257=>"000000111",
  55258=>"100000001",
  55259=>"100111010",
  55260=>"000111101",
  55261=>"001111110",
  55262=>"010000101",
  55263=>"101100010",
  55264=>"101001011",
  55265=>"110000000",
  55266=>"111100101",
  55267=>"100101101",
  55268=>"111111011",
  55269=>"111110111",
  55270=>"101110010",
  55271=>"111100110",
  55272=>"011011001",
  55273=>"100010111",
  55274=>"110011110",
  55275=>"101101010",
  55276=>"101101111",
  55277=>"101011101",
  55278=>"111100110",
  55279=>"100101111",
  55280=>"101011001",
  55281=>"101011010",
  55282=>"010110110",
  55283=>"101011101",
  55284=>"101101001",
  55285=>"011010010",
  55286=>"111101000",
  55287=>"000100111",
  55288=>"000111111",
  55289=>"111111111",
  55290=>"000011111",
  55291=>"111011010",
  55292=>"000110000",
  55293=>"100001111",
  55294=>"111111111",
  55295=>"001101101",
  55296=>"000010111",
  55297=>"101001111",
  55298=>"110001110",
  55299=>"010101111",
  55300=>"000000110",
  55301=>"010001111",
  55302=>"101100000",
  55303=>"101001000",
  55304=>"101010110",
  55305=>"000000101",
  55306=>"001001000",
  55307=>"111010001",
  55308=>"101000011",
  55309=>"011010100",
  55310=>"011101001",
  55311=>"110110010",
  55312=>"100111110",
  55313=>"101000101",
  55314=>"100001001",
  55315=>"010111100",
  55316=>"111011111",
  55317=>"111101100",
  55318=>"110100010",
  55319=>"111101100",
  55320=>"100011110",
  55321=>"101100010",
  55322=>"110011110",
  55323=>"000111000",
  55324=>"110011110",
  55325=>"011111011",
  55326=>"010000100",
  55327=>"000000110",
  55328=>"111111110",
  55329=>"100001100",
  55330=>"110100100",
  55331=>"100111010",
  55332=>"110100111",
  55333=>"101001111",
  55334=>"101110101",
  55335=>"111000101",
  55336=>"000100000",
  55337=>"101000100",
  55338=>"110110100",
  55339=>"100001001",
  55340=>"001110100",
  55341=>"110110010",
  55342=>"000101010",
  55343=>"010111101",
  55344=>"101111111",
  55345=>"100011100",
  55346=>"010100000",
  55347=>"110011010",
  55348=>"101001000",
  55349=>"001011111",
  55350=>"011011000",
  55351=>"110001111",
  55352=>"011101111",
  55353=>"000010001",
  55354=>"100001110",
  55355=>"010101101",
  55356=>"010001000",
  55357=>"000000101",
  55358=>"010111011",
  55359=>"111111101",
  55360=>"110011100",
  55361=>"100000000",
  55362=>"011100110",
  55363=>"000101001",
  55364=>"100000100",
  55365=>"110111110",
  55366=>"101110010",
  55367=>"101100111",
  55368=>"101111010",
  55369=>"000010010",
  55370=>"011110101",
  55371=>"110011111",
  55372=>"000001011",
  55373=>"110100010",
  55374=>"100000000",
  55375=>"001111011",
  55376=>"101010010",
  55377=>"100101100",
  55378=>"000001110",
  55379=>"100110010",
  55380=>"001110100",
  55381=>"000001101",
  55382=>"011101111",
  55383=>"000000101",
  55384=>"010010001",
  55385=>"101110100",
  55386=>"100100101",
  55387=>"101101110",
  55388=>"011011010",
  55389=>"011000100",
  55390=>"011001100",
  55391=>"001101001",
  55392=>"001000000",
  55393=>"100111010",
  55394=>"011011110",
  55395=>"000000001",
  55396=>"000100101",
  55397=>"111111010",
  55398=>"110000011",
  55399=>"111000110",
  55400=>"111101001",
  55401=>"010110011",
  55402=>"100100000",
  55403=>"110110101",
  55404=>"101001101",
  55405=>"101011101",
  55406=>"100100001",
  55407=>"010110111",
  55408=>"101011101",
  55409=>"111100101",
  55410=>"000110111",
  55411=>"011101100",
  55412=>"001000000",
  55413=>"010010111",
  55414=>"011010100",
  55415=>"001110011",
  55416=>"001101011",
  55417=>"000001101",
  55418=>"110000111",
  55419=>"001001100",
  55420=>"000110010",
  55421=>"001100001",
  55422=>"101111111",
  55423=>"000111110",
  55424=>"110001111",
  55425=>"101010011",
  55426=>"000000001",
  55427=>"000110101",
  55428=>"010100111",
  55429=>"000001001",
  55430=>"001011101",
  55431=>"010111010",
  55432=>"100110110",
  55433=>"001001010",
  55434=>"110000100",
  55435=>"001000001",
  55436=>"111101000",
  55437=>"010000101",
  55438=>"001010001",
  55439=>"111110110",
  55440=>"011100001",
  55441=>"001101111",
  55442=>"001110001",
  55443=>"111011011",
  55444=>"111110010",
  55445=>"010110110",
  55446=>"000011001",
  55447=>"000101111",
  55448=>"111010011",
  55449=>"110101000",
  55450=>"000101001",
  55451=>"010000110",
  55452=>"110111100",
  55453=>"000001100",
  55454=>"110011100",
  55455=>"011110000",
  55456=>"100101010",
  55457=>"011100110",
  55458=>"110010001",
  55459=>"101110011",
  55460=>"010000011",
  55461=>"011110100",
  55462=>"001001111",
  55463=>"100000110",
  55464=>"110010100",
  55465=>"001011111",
  55466=>"100001010",
  55467=>"001101011",
  55468=>"000110010",
  55469=>"000111100",
  55470=>"001110000",
  55471=>"111001001",
  55472=>"101111001",
  55473=>"001000001",
  55474=>"110011110",
  55475=>"001000111",
  55476=>"100011000",
  55477=>"010010011",
  55478=>"001110000",
  55479=>"011000011",
  55480=>"100010101",
  55481=>"000001101",
  55482=>"101101100",
  55483=>"000010010",
  55484=>"011010011",
  55485=>"011010010",
  55486=>"100100110",
  55487=>"000101011",
  55488=>"001011100",
  55489=>"001100010",
  55490=>"111010001",
  55491=>"001011001",
  55492=>"100000101",
  55493=>"011000011",
  55494=>"100011110",
  55495=>"111000111",
  55496=>"011100011",
  55497=>"101111110",
  55498=>"110111000",
  55499=>"110101011",
  55500=>"110110000",
  55501=>"101000000",
  55502=>"011111111",
  55503=>"100110001",
  55504=>"110100101",
  55505=>"100000100",
  55506=>"010111000",
  55507=>"001010011",
  55508=>"100001001",
  55509=>"110001001",
  55510=>"101010011",
  55511=>"101011001",
  55512=>"001001001",
  55513=>"001100011",
  55514=>"011001101",
  55515=>"100001000",
  55516=>"100101110",
  55517=>"100100011",
  55518=>"001000100",
  55519=>"010011110",
  55520=>"100110001",
  55521=>"101010010",
  55522=>"001010100",
  55523=>"001011011",
  55524=>"101011010",
  55525=>"000101100",
  55526=>"110101001",
  55527=>"011111100",
  55528=>"000110100",
  55529=>"011011111",
  55530=>"000100001",
  55531=>"011100111",
  55532=>"010101000",
  55533=>"100100011",
  55534=>"010000000",
  55535=>"000000000",
  55536=>"001101011",
  55537=>"010000100",
  55538=>"110000101",
  55539=>"000010110",
  55540=>"010000011",
  55541=>"100101111",
  55542=>"000101111",
  55543=>"100011010",
  55544=>"011001001",
  55545=>"000000001",
  55546=>"111011010",
  55547=>"001011010",
  55548=>"000010111",
  55549=>"010110011",
  55550=>"001101101",
  55551=>"000000100",
  55552=>"001100110",
  55553=>"000110000",
  55554=>"111100011",
  55555=>"101001100",
  55556=>"001001000",
  55557=>"101010110",
  55558=>"001101101",
  55559=>"111101110",
  55560=>"000110110",
  55561=>"110000100",
  55562=>"110000100",
  55563=>"111110011",
  55564=>"011100101",
  55565=>"001000101",
  55566=>"001110111",
  55567=>"010001100",
  55568=>"011101110",
  55569=>"101111111",
  55570=>"110010110",
  55571=>"010100001",
  55572=>"010001101",
  55573=>"001101010",
  55574=>"000100111",
  55575=>"000101100",
  55576=>"010001010",
  55577=>"011001110",
  55578=>"101000000",
  55579=>"000110100",
  55580=>"000001010",
  55581=>"111100101",
  55582=>"110100010",
  55583=>"000010001",
  55584=>"011101010",
  55585=>"001100000",
  55586=>"001010100",
  55587=>"001000101",
  55588=>"000010011",
  55589=>"011100111",
  55590=>"100111111",
  55591=>"000111011",
  55592=>"111010111",
  55593=>"100011111",
  55594=>"001010000",
  55595=>"011100010",
  55596=>"101110111",
  55597=>"101000011",
  55598=>"000101001",
  55599=>"110001000",
  55600=>"010110100",
  55601=>"101110100",
  55602=>"111100011",
  55603=>"011011110",
  55604=>"101100101",
  55605=>"100011000",
  55606=>"011010010",
  55607=>"001010010",
  55608=>"011010000",
  55609=>"011010010",
  55610=>"101101111",
  55611=>"111001101",
  55612=>"001000111",
  55613=>"111100110",
  55614=>"101111101",
  55615=>"011100100",
  55616=>"101011001",
  55617=>"000010100",
  55618=>"000010100",
  55619=>"010011000",
  55620=>"101011111",
  55621=>"101110011",
  55622=>"011010100",
  55623=>"000001011",
  55624=>"111010110",
  55625=>"001001110",
  55626=>"011110101",
  55627=>"000000011",
  55628=>"010011011",
  55629=>"110011010",
  55630=>"110111001",
  55631=>"000100011",
  55632=>"100001110",
  55633=>"110001101",
  55634=>"001001100",
  55635=>"100001100",
  55636=>"111110111",
  55637=>"010110000",
  55638=>"110110101",
  55639=>"100100000",
  55640=>"010101111",
  55641=>"011011111",
  55642=>"111001101",
  55643=>"000110100",
  55644=>"101011011",
  55645=>"010111111",
  55646=>"010000010",
  55647=>"011001011",
  55648=>"111000101",
  55649=>"011101101",
  55650=>"011001111",
  55651=>"110110000",
  55652=>"000010010",
  55653=>"101100111",
  55654=>"001101011",
  55655=>"010100011",
  55656=>"011101111",
  55657=>"101101001",
  55658=>"001111001",
  55659=>"000111110",
  55660=>"000100101",
  55661=>"000001100",
  55662=>"001000101",
  55663=>"100011000",
  55664=>"100101100",
  55665=>"100110100",
  55666=>"100101001",
  55667=>"010000001",
  55668=>"101111111",
  55669=>"100010111",
  55670=>"001000011",
  55671=>"101000111",
  55672=>"100100100",
  55673=>"011000000",
  55674=>"011101110",
  55675=>"110000001",
  55676=>"110010111",
  55677=>"000000001",
  55678=>"011111101",
  55679=>"100011111",
  55680=>"010110100",
  55681=>"111110100",
  55682=>"011001001",
  55683=>"011101111",
  55684=>"011100010",
  55685=>"011101101",
  55686=>"001001101",
  55687=>"001001000",
  55688=>"101110000",
  55689=>"100110111",
  55690=>"101010011",
  55691=>"100110101",
  55692=>"010101000",
  55693=>"010100110",
  55694=>"100110011",
  55695=>"000000110",
  55696=>"011100100",
  55697=>"011000100",
  55698=>"001000010",
  55699=>"000111111",
  55700=>"110001111",
  55701=>"011110101",
  55702=>"100010010",
  55703=>"000001001",
  55704=>"101110000",
  55705=>"010011111",
  55706=>"111110011",
  55707=>"111111000",
  55708=>"111001110",
  55709=>"000001101",
  55710=>"001100000",
  55711=>"111000011",
  55712=>"000100100",
  55713=>"100011010",
  55714=>"100001000",
  55715=>"111011000",
  55716=>"111110011",
  55717=>"101111101",
  55718=>"100111101",
  55719=>"101110011",
  55720=>"101110001",
  55721=>"001010011",
  55722=>"001000011",
  55723=>"000011111",
  55724=>"101000011",
  55725=>"010000000",
  55726=>"110001111",
  55727=>"101011010",
  55728=>"001011001",
  55729=>"000001110",
  55730=>"001101100",
  55731=>"000011010",
  55732=>"100101011",
  55733=>"011001111",
  55734=>"110101011",
  55735=>"110111000",
  55736=>"100101011",
  55737=>"011001101",
  55738=>"000111110",
  55739=>"101000111",
  55740=>"100110010",
  55741=>"001010011",
  55742=>"011101011",
  55743=>"111010101",
  55744=>"111010011",
  55745=>"000001010",
  55746=>"101111100",
  55747=>"010110001",
  55748=>"011011101",
  55749=>"100101100",
  55750=>"011111011",
  55751=>"001000110",
  55752=>"110001110",
  55753=>"000110010",
  55754=>"101011110",
  55755=>"010011111",
  55756=>"000101110",
  55757=>"010010010",
  55758=>"010010101",
  55759=>"111011100",
  55760=>"000110011",
  55761=>"000100101",
  55762=>"100110000",
  55763=>"010011100",
  55764=>"110001111",
  55765=>"110110110",
  55766=>"010011101",
  55767=>"101011001",
  55768=>"011000100",
  55769=>"110110011",
  55770=>"100000000",
  55771=>"110010001",
  55772=>"110111010",
  55773=>"011010101",
  55774=>"001001101",
  55775=>"100100110",
  55776=>"100101000",
  55777=>"101000011",
  55778=>"000011101",
  55779=>"100010000",
  55780=>"010110101",
  55781=>"011010001",
  55782=>"111011010",
  55783=>"101001100",
  55784=>"011100100",
  55785=>"100111101",
  55786=>"101001010",
  55787=>"111111010",
  55788=>"000101001",
  55789=>"011110011",
  55790=>"010000001",
  55791=>"000110011",
  55792=>"011011000",
  55793=>"010000111",
  55794=>"110100110",
  55795=>"001010111",
  55796=>"110100101",
  55797=>"111110101",
  55798=>"100111110",
  55799=>"111111101",
  55800=>"010110101",
  55801=>"010111110",
  55802=>"100111100",
  55803=>"000010101",
  55804=>"101110000",
  55805=>"101011011",
  55806=>"000011000",
  55807=>"111010001",
  55808=>"101101001",
  55809=>"001110110",
  55810=>"000100011",
  55811=>"010111101",
  55812=>"001110100",
  55813=>"000001000",
  55814=>"000010011",
  55815=>"111000001",
  55816=>"010000011",
  55817=>"111100110",
  55818=>"111110011",
  55819=>"111101111",
  55820=>"110111010",
  55821=>"101100110",
  55822=>"001101000",
  55823=>"111111111",
  55824=>"001010011",
  55825=>"000110111",
  55826=>"011011001",
  55827=>"010010100",
  55828=>"001010001",
  55829=>"110001111",
  55830=>"100111111",
  55831=>"010010000",
  55832=>"010010001",
  55833=>"010001110",
  55834=>"001011001",
  55835=>"101101000",
  55836=>"011111000",
  55837=>"111110101",
  55838=>"001100001",
  55839=>"110110010",
  55840=>"111111000",
  55841=>"100111101",
  55842=>"011001110",
  55843=>"010000000",
  55844=>"110100101",
  55845=>"110011000",
  55846=>"100000101",
  55847=>"001111110",
  55848=>"000000011",
  55849=>"111110110",
  55850=>"000111100",
  55851=>"001000111",
  55852=>"010100101",
  55853=>"000100010",
  55854=>"101010000",
  55855=>"100001100",
  55856=>"100000010",
  55857=>"010111111",
  55858=>"111001010",
  55859=>"010010001",
  55860=>"100010101",
  55861=>"111010010",
  55862=>"000011111",
  55863=>"000111000",
  55864=>"111001110",
  55865=>"010111001",
  55866=>"101111001",
  55867=>"110100111",
  55868=>"000110110",
  55869=>"110101101",
  55870=>"110101100",
  55871=>"011100001",
  55872=>"110111110",
  55873=>"100000011",
  55874=>"011011011",
  55875=>"000010111",
  55876=>"001100000",
  55877=>"100011011",
  55878=>"001001111",
  55879=>"110101011",
  55880=>"001111010",
  55881=>"011111100",
  55882=>"000111010",
  55883=>"110100101",
  55884=>"001101100",
  55885=>"010101100",
  55886=>"101111110",
  55887=>"101110000",
  55888=>"111101111",
  55889=>"111000011",
  55890=>"000101000",
  55891=>"000100000",
  55892=>"111000010",
  55893=>"100000111",
  55894=>"010001111",
  55895=>"100001010",
  55896=>"010100000",
  55897=>"101101100",
  55898=>"000010000",
  55899=>"101011000",
  55900=>"001101011",
  55901=>"110110100",
  55902=>"100010001",
  55903=>"110001111",
  55904=>"011000010",
  55905=>"100001000",
  55906=>"111100010",
  55907=>"101000000",
  55908=>"010111011",
  55909=>"100101000",
  55910=>"101110100",
  55911=>"001111010",
  55912=>"101010011",
  55913=>"011011010",
  55914=>"110001000",
  55915=>"101111101",
  55916=>"010111001",
  55917=>"000100000",
  55918=>"100010110",
  55919=>"101110000",
  55920=>"100111010",
  55921=>"011011101",
  55922=>"001111001",
  55923=>"101101111",
  55924=>"000000000",
  55925=>"010100010",
  55926=>"000111000",
  55927=>"000011011",
  55928=>"101100000",
  55929=>"000100000",
  55930=>"011001100",
  55931=>"011100100",
  55932=>"001011101",
  55933=>"011011100",
  55934=>"111100111",
  55935=>"011111001",
  55936=>"000101110",
  55937=>"000010000",
  55938=>"001111011",
  55939=>"001000010",
  55940=>"000000100",
  55941=>"101000101",
  55942=>"111011011",
  55943=>"011011010",
  55944=>"110000111",
  55945=>"111111111",
  55946=>"010001100",
  55947=>"000101100",
  55948=>"001100100",
  55949=>"101011101",
  55950=>"101100010",
  55951=>"001000000",
  55952=>"100000010",
  55953=>"100001001",
  55954=>"000111001",
  55955=>"000000001",
  55956=>"100101111",
  55957=>"011010001",
  55958=>"011010000",
  55959=>"010011101",
  55960=>"010000010",
  55961=>"001111111",
  55962=>"110110111",
  55963=>"110011100",
  55964=>"100000001",
  55965=>"111110101",
  55966=>"110100101",
  55967=>"101000000",
  55968=>"010011001",
  55969=>"101101010",
  55970=>"011011000",
  55971=>"011001100",
  55972=>"001011001",
  55973=>"101110111",
  55974=>"010010000",
  55975=>"010100010",
  55976=>"011000000",
  55977=>"000100111",
  55978=>"100000011",
  55979=>"100001010",
  55980=>"111100100",
  55981=>"111110110",
  55982=>"000100101",
  55983=>"001110010",
  55984=>"000100110",
  55985=>"011110010",
  55986=>"101011011",
  55987=>"100101011",
  55988=>"101110100",
  55989=>"101001111",
  55990=>"111001101",
  55991=>"011101100",
  55992=>"001010000",
  55993=>"010001110",
  55994=>"101100101",
  55995=>"110010000",
  55996=>"010110110",
  55997=>"001001100",
  55998=>"001011010",
  55999=>"110100010",
  56000=>"010111110",
  56001=>"111111010",
  56002=>"011001001",
  56003=>"001100110",
  56004=>"001110001",
  56005=>"111001010",
  56006=>"110100011",
  56007=>"001110010",
  56008=>"101101001",
  56009=>"101101011",
  56010=>"010001000",
  56011=>"000100110",
  56012=>"011011111",
  56013=>"011100111",
  56014=>"000011001",
  56015=>"011110111",
  56016=>"111100010",
  56017=>"011010011",
  56018=>"111001110",
  56019=>"010001000",
  56020=>"111111110",
  56021=>"011000011",
  56022=>"100100111",
  56023=>"101110110",
  56024=>"111111001",
  56025=>"001100011",
  56026=>"011110011",
  56027=>"000001011",
  56028=>"101000000",
  56029=>"000100110",
  56030=>"101110000",
  56031=>"110111000",
  56032=>"010111001",
  56033=>"001001010",
  56034=>"011011000",
  56035=>"100100000",
  56036=>"101001010",
  56037=>"100011011",
  56038=>"000110111",
  56039=>"100011101",
  56040=>"100001011",
  56041=>"001111101",
  56042=>"111011011",
  56043=>"011110111",
  56044=>"010010011",
  56045=>"001111100",
  56046=>"000101000",
  56047=>"111010100",
  56048=>"010100100",
  56049=>"010011101",
  56050=>"010100000",
  56051=>"001001000",
  56052=>"100101000",
  56053=>"111100011",
  56054=>"010101101",
  56055=>"110010010",
  56056=>"110000100",
  56057=>"000111010",
  56058=>"101000000",
  56059=>"001100011",
  56060=>"011011110",
  56061=>"111100000",
  56062=>"111101010",
  56063=>"100011101",
  56064=>"111100011",
  56065=>"000111011",
  56066=>"001010010",
  56067=>"111110011",
  56068=>"011101011",
  56069=>"110110100",
  56070=>"100111001",
  56071=>"100000100",
  56072=>"000100100",
  56073=>"001101000",
  56074=>"010110011",
  56075=>"000111010",
  56076=>"000001001",
  56077=>"110011110",
  56078=>"110110001",
  56079=>"110111000",
  56080=>"110011011",
  56081=>"000101001",
  56082=>"001011010",
  56083=>"101010011",
  56084=>"001101111",
  56085=>"001100101",
  56086=>"111011110",
  56087=>"010011101",
  56088=>"001001010",
  56089=>"000001100",
  56090=>"101001111",
  56091=>"000110110",
  56092=>"001000110",
  56093=>"111011011",
  56094=>"100111111",
  56095=>"101111100",
  56096=>"101011100",
  56097=>"101011100",
  56098=>"110011111",
  56099=>"010111111",
  56100=>"111111111",
  56101=>"110100001",
  56102=>"010100111",
  56103=>"011101010",
  56104=>"000011010",
  56105=>"101100110",
  56106=>"100001000",
  56107=>"111001001",
  56108=>"100000011",
  56109=>"001111100",
  56110=>"101000100",
  56111=>"100110110",
  56112=>"000100010",
  56113=>"010011110",
  56114=>"100001111",
  56115=>"110010010",
  56116=>"101100000",
  56117=>"001000101",
  56118=>"000001001",
  56119=>"111101101",
  56120=>"000101111",
  56121=>"101010111",
  56122=>"100010001",
  56123=>"111100011",
  56124=>"101100111",
  56125=>"011011000",
  56126=>"101101001",
  56127=>"001101110",
  56128=>"101111010",
  56129=>"001100010",
  56130=>"100100001",
  56131=>"100001100",
  56132=>"101101011",
  56133=>"010110001",
  56134=>"000001100",
  56135=>"100011110",
  56136=>"011101011",
  56137=>"111111110",
  56138=>"100110100",
  56139=>"010101001",
  56140=>"000100011",
  56141=>"101000010",
  56142=>"110100000",
  56143=>"111111000",
  56144=>"101100100",
  56145=>"100100001",
  56146=>"001110011",
  56147=>"010110010",
  56148=>"011100000",
  56149=>"010000000",
  56150=>"011001011",
  56151=>"111011110",
  56152=>"011011101",
  56153=>"000010000",
  56154=>"100010001",
  56155=>"100001101",
  56156=>"010001011",
  56157=>"011101011",
  56158=>"101100000",
  56159=>"001101011",
  56160=>"100001010",
  56161=>"010100110",
  56162=>"110100011",
  56163=>"101010010",
  56164=>"010011111",
  56165=>"101001001",
  56166=>"010111111",
  56167=>"110001001",
  56168=>"100101000",
  56169=>"110111011",
  56170=>"110100010",
  56171=>"101111001",
  56172=>"000011000",
  56173=>"000011011",
  56174=>"100111110",
  56175=>"111010101",
  56176=>"010100000",
  56177=>"110100100",
  56178=>"011101001",
  56179=>"111101101",
  56180=>"001111011",
  56181=>"001111110",
  56182=>"000010010",
  56183=>"010000110",
  56184=>"011111100",
  56185=>"011101111",
  56186=>"011001101",
  56187=>"101001101",
  56188=>"000100011",
  56189=>"011010101",
  56190=>"011100011",
  56191=>"100110110",
  56192=>"111100100",
  56193=>"011101010",
  56194=>"001011110",
  56195=>"101001111",
  56196=>"011101001",
  56197=>"111101111",
  56198=>"010101010",
  56199=>"010100100",
  56200=>"101101100",
  56201=>"000111100",
  56202=>"110100110",
  56203=>"010010100",
  56204=>"011001011",
  56205=>"001001011",
  56206=>"111011010",
  56207=>"110100100",
  56208=>"010110101",
  56209=>"110000100",
  56210=>"000101101",
  56211=>"100010011",
  56212=>"101010100",
  56213=>"010001010",
  56214=>"000001001",
  56215=>"111111011",
  56216=>"011111001",
  56217=>"010111100",
  56218=>"011001010",
  56219=>"001011110",
  56220=>"010001101",
  56221=>"101100001",
  56222=>"001001000",
  56223=>"101011101",
  56224=>"010111110",
  56225=>"001101011",
  56226=>"011011011",
  56227=>"101110010",
  56228=>"101011011",
  56229=>"000101000",
  56230=>"010101010",
  56231=>"101111000",
  56232=>"101001111",
  56233=>"110011000",
  56234=>"010010000",
  56235=>"000000011",
  56236=>"100000100",
  56237=>"111111100",
  56238=>"100001011",
  56239=>"111110000",
  56240=>"111101101",
  56241=>"011010110",
  56242=>"101011101",
  56243=>"000110011",
  56244=>"111011111",
  56245=>"010010000",
  56246=>"000101101",
  56247=>"000010111",
  56248=>"011101111",
  56249=>"001000101",
  56250=>"001110110",
  56251=>"010000010",
  56252=>"111011000",
  56253=>"010101011",
  56254=>"111111111",
  56255=>"100010110",
  56256=>"110010110",
  56257=>"101010001",
  56258=>"100000101",
  56259=>"100110010",
  56260=>"111101010",
  56261=>"101110000",
  56262=>"011011011",
  56263=>"111100111",
  56264=>"001110101",
  56265=>"100111110",
  56266=>"001101110",
  56267=>"100110110",
  56268=>"100100110",
  56269=>"001110101",
  56270=>"110111110",
  56271=>"001010101",
  56272=>"110001110",
  56273=>"001101011",
  56274=>"111111110",
  56275=>"011110110",
  56276=>"010101111",
  56277=>"001110101",
  56278=>"101000100",
  56279=>"101111111",
  56280=>"001011110",
  56281=>"111100000",
  56282=>"110111100",
  56283=>"011000101",
  56284=>"110111101",
  56285=>"000001000",
  56286=>"101100011",
  56287=>"000001010",
  56288=>"001010111",
  56289=>"001010001",
  56290=>"110001001",
  56291=>"001111000",
  56292=>"110000001",
  56293=>"010101011",
  56294=>"010001001",
  56295=>"111110010",
  56296=>"000011010",
  56297=>"010011001",
  56298=>"100000000",
  56299=>"110010100",
  56300=>"001001010",
  56301=>"111111100",
  56302=>"110111101",
  56303=>"011110011",
  56304=>"000100000",
  56305=>"011111101",
  56306=>"101111100",
  56307=>"110011101",
  56308=>"110110110",
  56309=>"100001010",
  56310=>"100000001",
  56311=>"100101011",
  56312=>"000100010",
  56313=>"110111011",
  56314=>"000000101",
  56315=>"011001011",
  56316=>"110001001",
  56317=>"101010100",
  56318=>"011100000",
  56319=>"011000000",
  56320=>"010001011",
  56321=>"010011011",
  56322=>"010001001",
  56323=>"010000011",
  56324=>"011000010",
  56325=>"101101011",
  56326=>"100100111",
  56327=>"011000100",
  56328=>"000000110",
  56329=>"010011000",
  56330=>"001111010",
  56331=>"110011111",
  56332=>"011000100",
  56333=>"101011000",
  56334=>"010001100",
  56335=>"011010110",
  56336=>"010011100",
  56337=>"001100011",
  56338=>"000001110",
  56339=>"100010111",
  56340=>"101000110",
  56341=>"000100011",
  56342=>"110011010",
  56343=>"100001011",
  56344=>"001111100",
  56345=>"001101000",
  56346=>"010001110",
  56347=>"011101100",
  56348=>"011010010",
  56349=>"001100011",
  56350=>"000010111",
  56351=>"101011101",
  56352=>"010011001",
  56353=>"111011011",
  56354=>"110000100",
  56355=>"000011101",
  56356=>"000111010",
  56357=>"000011100",
  56358=>"011001111",
  56359=>"001101011",
  56360=>"100001010",
  56361=>"000000111",
  56362=>"101011111",
  56363=>"101001101",
  56364=>"010111000",
  56365=>"111110011",
  56366=>"110101111",
  56367=>"000111011",
  56368=>"100001010",
  56369=>"000101110",
  56370=>"001010111",
  56371=>"001011000",
  56372=>"001000100",
  56373=>"001100000",
  56374=>"010100010",
  56375=>"010000010",
  56376=>"010100100",
  56377=>"110001011",
  56378=>"101111111",
  56379=>"100000100",
  56380=>"011000010",
  56381=>"010010111",
  56382=>"011111010",
  56383=>"010111000",
  56384=>"110010000",
  56385=>"110100011",
  56386=>"001000000",
  56387=>"010101101",
  56388=>"110010100",
  56389=>"110110010",
  56390=>"101101001",
  56391=>"000010001",
  56392=>"011010001",
  56393=>"111111110",
  56394=>"010000000",
  56395=>"101001000",
  56396=>"010001001",
  56397=>"100000010",
  56398=>"100011101",
  56399=>"010100110",
  56400=>"111011110",
  56401=>"100110010",
  56402=>"101010100",
  56403=>"101010010",
  56404=>"001101111",
  56405=>"000000111",
  56406=>"100000110",
  56407=>"001000101",
  56408=>"101101010",
  56409=>"000000001",
  56410=>"101101110",
  56411=>"001100000",
  56412=>"000001010",
  56413=>"101100010",
  56414=>"001111111",
  56415=>"111000001",
  56416=>"101100110",
  56417=>"101010000",
  56418=>"011011011",
  56419=>"010010011",
  56420=>"000011001",
  56421=>"100100111",
  56422=>"011001010",
  56423=>"110011111",
  56424=>"001011010",
  56425=>"100110000",
  56426=>"101100000",
  56427=>"010100100",
  56428=>"001100011",
  56429=>"010110110",
  56430=>"011001111",
  56431=>"111111010",
  56432=>"100110101",
  56433=>"010100000",
  56434=>"000111111",
  56435=>"011101100",
  56436=>"110111111",
  56437=>"110100000",
  56438=>"110000011",
  56439=>"011010000",
  56440=>"110000000",
  56441=>"100100110",
  56442=>"010000111",
  56443=>"010100100",
  56444=>"110000001",
  56445=>"010110101",
  56446=>"110101001",
  56447=>"000101101",
  56448=>"111011000",
  56449=>"100000001",
  56450=>"001100010",
  56451=>"100110110",
  56452=>"101010100",
  56453=>"001011001",
  56454=>"011011011",
  56455=>"100000010",
  56456=>"010011110",
  56457=>"000000101",
  56458=>"101000111",
  56459=>"010101101",
  56460=>"101001011",
  56461=>"111110111",
  56462=>"000101010",
  56463=>"011111111",
  56464=>"001001010",
  56465=>"110011110",
  56466=>"110111010",
  56467=>"100110000",
  56468=>"000000111",
  56469=>"001111111",
  56470=>"010101110",
  56471=>"001100100",
  56472=>"110110100",
  56473=>"111000000",
  56474=>"111001011",
  56475=>"010111001",
  56476=>"111111001",
  56477=>"111111100",
  56478=>"001011010",
  56479=>"111000000",
  56480=>"010100101",
  56481=>"101110111",
  56482=>"010011100",
  56483=>"110010110",
  56484=>"110101000",
  56485=>"010010000",
  56486=>"011011111",
  56487=>"111010000",
  56488=>"011110010",
  56489=>"100100011",
  56490=>"001101000",
  56491=>"100011100",
  56492=>"011101011",
  56493=>"111001010",
  56494=>"100011111",
  56495=>"110001101",
  56496=>"000010100",
  56497=>"100100000",
  56498=>"010111010",
  56499=>"110100000",
  56500=>"100111110",
  56501=>"000000001",
  56502=>"001000110",
  56503=>"010001111",
  56504=>"011001110",
  56505=>"010100011",
  56506=>"111110000",
  56507=>"000110011",
  56508=>"010010100",
  56509=>"010100000",
  56510=>"000101000",
  56511=>"110010001",
  56512=>"011110011",
  56513=>"001010111",
  56514=>"011011110",
  56515=>"110101001",
  56516=>"001011101",
  56517=>"010100111",
  56518=>"010100111",
  56519=>"101100110",
  56520=>"100000000",
  56521=>"110000111",
  56522=>"111111110",
  56523=>"011010000",
  56524=>"111100101",
  56525=>"110010000",
  56526=>"001100111",
  56527=>"001110000",
  56528=>"011111001",
  56529=>"010011011",
  56530=>"001010010",
  56531=>"001000010",
  56532=>"010100011",
  56533=>"111101001",
  56534=>"100011111",
  56535=>"011011011",
  56536=>"000101111",
  56537=>"100000010",
  56538=>"101111000",
  56539=>"100100001",
  56540=>"111101100",
  56541=>"011010001",
  56542=>"111000111",
  56543=>"001101000",
  56544=>"011000110",
  56545=>"011100111",
  56546=>"100001000",
  56547=>"010010100",
  56548=>"010010010",
  56549=>"001101010",
  56550=>"110001000",
  56551=>"000000100",
  56552=>"100111101",
  56553=>"100000000",
  56554=>"011111000",
  56555=>"110001110",
  56556=>"010001110",
  56557=>"001111010",
  56558=>"010110011",
  56559=>"101010111",
  56560=>"101101110",
  56561=>"001000110",
  56562=>"001101101",
  56563=>"110101001",
  56564=>"001011001",
  56565=>"101001100",
  56566=>"110011010",
  56567=>"000001110",
  56568=>"111011010",
  56569=>"011010011",
  56570=>"001011100",
  56571=>"001001010",
  56572=>"111010010",
  56573=>"100100000",
  56574=>"100100111",
  56575=>"111110001",
  56576=>"011101011",
  56577=>"110110011",
  56578=>"010010001",
  56579=>"100011001",
  56580=>"011011111",
  56581=>"110110111",
  56582=>"101111101",
  56583=>"111010010",
  56584=>"101000110",
  56585=>"100100000",
  56586=>"001110001",
  56587=>"111100111",
  56588=>"000001001",
  56589=>"100000101",
  56590=>"111100100",
  56591=>"010100100",
  56592=>"001010100",
  56593=>"010111010",
  56594=>"001010001",
  56595=>"110010000",
  56596=>"110110001",
  56597=>"110000001",
  56598=>"111000000",
  56599=>"100000111",
  56600=>"110111000",
  56601=>"001111010",
  56602=>"100001101",
  56603=>"110110001",
  56604=>"001010111",
  56605=>"101111001",
  56606=>"011111000",
  56607=>"100101001",
  56608=>"100010010",
  56609=>"110011010",
  56610=>"001011110",
  56611=>"111001001",
  56612=>"111111001",
  56613=>"100001110",
  56614=>"111101010",
  56615=>"000010111",
  56616=>"011110001",
  56617=>"101101010",
  56618=>"001010110",
  56619=>"111011011",
  56620=>"000110000",
  56621=>"011111000",
  56622=>"001110000",
  56623=>"000110100",
  56624=>"000000101",
  56625=>"110010100",
  56626=>"010111101",
  56627=>"101101010",
  56628=>"001000000",
  56629=>"101110101",
  56630=>"010010010",
  56631=>"011000110",
  56632=>"110001100",
  56633=>"100100100",
  56634=>"111111111",
  56635=>"000000011",
  56636=>"110100000",
  56637=>"111101100",
  56638=>"010001100",
  56639=>"001011011",
  56640=>"001011010",
  56641=>"000010111",
  56642=>"011011001",
  56643=>"101001011",
  56644=>"001010011",
  56645=>"101000110",
  56646=>"110000001",
  56647=>"000111111",
  56648=>"101011010",
  56649=>"010101010",
  56650=>"101100001",
  56651=>"010100010",
  56652=>"010100101",
  56653=>"011101101",
  56654=>"000011000",
  56655=>"110010000",
  56656=>"011110010",
  56657=>"000011010",
  56658=>"101000000",
  56659=>"010101001",
  56660=>"011001001",
  56661=>"000011001",
  56662=>"100010111",
  56663=>"000000110",
  56664=>"110000100",
  56665=>"010011101",
  56666=>"010001100",
  56667=>"101111001",
  56668=>"111101110",
  56669=>"010000110",
  56670=>"111111111",
  56671=>"111101001",
  56672=>"111000011",
  56673=>"111101101",
  56674=>"011111001",
  56675=>"000101010",
  56676=>"101100110",
  56677=>"000100100",
  56678=>"111011110",
  56679=>"000101111",
  56680=>"101010101",
  56681=>"111111000",
  56682=>"011100101",
  56683=>"111010001",
  56684=>"110000000",
  56685=>"111011000",
  56686=>"001111010",
  56687=>"101010001",
  56688=>"100001101",
  56689=>"001100010",
  56690=>"001111001",
  56691=>"111110110",
  56692=>"110000011",
  56693=>"011100000",
  56694=>"100000000",
  56695=>"000011011",
  56696=>"001110110",
  56697=>"100011000",
  56698=>"100011111",
  56699=>"000011110",
  56700=>"000100001",
  56701=>"010001100",
  56702=>"110001110",
  56703=>"001011001",
  56704=>"010101101",
  56705=>"000110110",
  56706=>"100111011",
  56707=>"010101010",
  56708=>"111111010",
  56709=>"100010001",
  56710=>"011110111",
  56711=>"111010000",
  56712=>"001111101",
  56713=>"010111011",
  56714=>"101100000",
  56715=>"110111001",
  56716=>"001100000",
  56717=>"101010000",
  56718=>"011101101",
  56719=>"110010011",
  56720=>"111111101",
  56721=>"100010000",
  56722=>"101111101",
  56723=>"000110010",
  56724=>"000011001",
  56725=>"101101011",
  56726=>"100011111",
  56727=>"101001111",
  56728=>"000110100",
  56729=>"101001101",
  56730=>"100110001",
  56731=>"110100101",
  56732=>"011010010",
  56733=>"101001001",
  56734=>"011111101",
  56735=>"000100110",
  56736=>"011111101",
  56737=>"000001010",
  56738=>"101111110",
  56739=>"111111111",
  56740=>"101111101",
  56741=>"100001001",
  56742=>"100001111",
  56743=>"100001111",
  56744=>"101000110",
  56745=>"010101011",
  56746=>"010111010",
  56747=>"001100001",
  56748=>"101110011",
  56749=>"011111010",
  56750=>"001000001",
  56751=>"110111110",
  56752=>"011011111",
  56753=>"010111001",
  56754=>"001110011",
  56755=>"010100101",
  56756=>"101010100",
  56757=>"001101111",
  56758=>"010100000",
  56759=>"010001110",
  56760=>"001101100",
  56761=>"011011111",
  56762=>"110011110",
  56763=>"100010111",
  56764=>"100111111",
  56765=>"000000001",
  56766=>"101100100",
  56767=>"001000010",
  56768=>"111000100",
  56769=>"001100100",
  56770=>"000011011",
  56771=>"111110100",
  56772=>"111011010",
  56773=>"011110001",
  56774=>"101000101",
  56775=>"111011001",
  56776=>"001111100",
  56777=>"011010101",
  56778=>"111110111",
  56779=>"111000011",
  56780=>"110001111",
  56781=>"001100011",
  56782=>"000001011",
  56783=>"000011000",
  56784=>"000100110",
  56785=>"100100010",
  56786=>"100010110",
  56787=>"000100101",
  56788=>"011111000",
  56789=>"010100111",
  56790=>"101111000",
  56791=>"101100000",
  56792=>"001000011",
  56793=>"100000100",
  56794=>"101001110",
  56795=>"100100011",
  56796=>"101110100",
  56797=>"100001101",
  56798=>"101111010",
  56799=>"100000010",
  56800=>"111010010",
  56801=>"010001101",
  56802=>"111101110",
  56803=>"000101000",
  56804=>"010110011",
  56805=>"110001100",
  56806=>"100011001",
  56807=>"111100101",
  56808=>"011011110",
  56809=>"110111110",
  56810=>"010100010",
  56811=>"011001010",
  56812=>"000000011",
  56813=>"111010000",
  56814=>"100010101",
  56815=>"110111011",
  56816=>"001100101",
  56817=>"111011010",
  56818=>"110000101",
  56819=>"001100000",
  56820=>"011011110",
  56821=>"010101010",
  56822=>"000010001",
  56823=>"001110111",
  56824=>"100110001",
  56825=>"111100010",
  56826=>"101000011",
  56827=>"100011110",
  56828=>"011011100",
  56829=>"011001000",
  56830=>"000111010",
  56831=>"110000011",
  56832=>"110011101",
  56833=>"100000100",
  56834=>"000011110",
  56835=>"110011110",
  56836=>"010010001",
  56837=>"011111101",
  56838=>"000110100",
  56839=>"010101000",
  56840=>"101011101",
  56841=>"100010001",
  56842=>"100111110",
  56843=>"100001100",
  56844=>"001010011",
  56845=>"010011001",
  56846=>"000011101",
  56847=>"001111111",
  56848=>"100100001",
  56849=>"110010000",
  56850=>"010111111",
  56851=>"101001001",
  56852=>"000100010",
  56853=>"000111011",
  56854=>"111101001",
  56855=>"101110011",
  56856=>"000111110",
  56857=>"111100010",
  56858=>"100101110",
  56859=>"101010100",
  56860=>"011111101",
  56861=>"101001111",
  56862=>"011110001",
  56863=>"110100011",
  56864=>"100100001",
  56865=>"011000111",
  56866=>"001011001",
  56867=>"111111101",
  56868=>"110110010",
  56869=>"010111110",
  56870=>"001010100",
  56871=>"010110101",
  56872=>"001101101",
  56873=>"001111010",
  56874=>"111100011",
  56875=>"011010001",
  56876=>"111001101",
  56877=>"110011100",
  56878=>"101010101",
  56879=>"101001110",
  56880=>"100000000",
  56881=>"001010000",
  56882=>"100000011",
  56883=>"010011110",
  56884=>"101011000",
  56885=>"010000110",
  56886=>"001111000",
  56887=>"100010000",
  56888=>"000111100",
  56889=>"111110111",
  56890=>"111011011",
  56891=>"100101010",
  56892=>"111010010",
  56893=>"001000101",
  56894=>"110000101",
  56895=>"000100001",
  56896=>"100111010",
  56897=>"111010000",
  56898=>"100010110",
  56899=>"001110011",
  56900=>"001110010",
  56901=>"100100010",
  56902=>"001100111",
  56903=>"101111000",
  56904=>"101101000",
  56905=>"001110101",
  56906=>"100111011",
  56907=>"000101101",
  56908=>"101100000",
  56909=>"110011111",
  56910=>"000000000",
  56911=>"011000001",
  56912=>"001101010",
  56913=>"010000001",
  56914=>"100010000",
  56915=>"111100011",
  56916=>"111110110",
  56917=>"100000100",
  56918=>"000001000",
  56919=>"001001011",
  56920=>"100101100",
  56921=>"111110001",
  56922=>"011000100",
  56923=>"100001010",
  56924=>"010110010",
  56925=>"101000011",
  56926=>"000001110",
  56927=>"101111001",
  56928=>"010111100",
  56929=>"010011010",
  56930=>"011000101",
  56931=>"001001110",
  56932=>"011110100",
  56933=>"111111111",
  56934=>"110111001",
  56935=>"000110010",
  56936=>"100111101",
  56937=>"010111111",
  56938=>"011100000",
  56939=>"111110101",
  56940=>"100011000",
  56941=>"111111110",
  56942=>"110000111",
  56943=>"000100000",
  56944=>"000101101",
  56945=>"010010011",
  56946=>"011010000",
  56947=>"111110110",
  56948=>"101010101",
  56949=>"000111010",
  56950=>"100011111",
  56951=>"100000010",
  56952=>"000000101",
  56953=>"101011001",
  56954=>"110111101",
  56955=>"100010011",
  56956=>"100000000",
  56957=>"100010011",
  56958=>"100000010",
  56959=>"111110001",
  56960=>"101100001",
  56961=>"011010011",
  56962=>"001001010",
  56963=>"110001001",
  56964=>"100100101",
  56965=>"011011101",
  56966=>"011010101",
  56967=>"011001000",
  56968=>"110011111",
  56969=>"010010111",
  56970=>"001100111",
  56971=>"000011001",
  56972=>"011000011",
  56973=>"111010000",
  56974=>"011101101",
  56975=>"111100001",
  56976=>"101110110",
  56977=>"111110111",
  56978=>"111011001",
  56979=>"110101010",
  56980=>"100100010",
  56981=>"101100010",
  56982=>"000111010",
  56983=>"111110001",
  56984=>"000001010",
  56985=>"000100101",
  56986=>"111100110",
  56987=>"000111010",
  56988=>"001011001",
  56989=>"100100001",
  56990=>"110110010",
  56991=>"001000011",
  56992=>"110101101",
  56993=>"010101001",
  56994=>"110111101",
  56995=>"101110011",
  56996=>"011100101",
  56997=>"111101010",
  56998=>"111111111",
  56999=>"010110110",
  57000=>"010111001",
  57001=>"100000000",
  57002=>"101001110",
  57003=>"110010011",
  57004=>"110001000",
  57005=>"101101101",
  57006=>"001100000",
  57007=>"011001000",
  57008=>"001100100",
  57009=>"111100110",
  57010=>"111100101",
  57011=>"000110011",
  57012=>"111100100",
  57013=>"110001001",
  57014=>"010001010",
  57015=>"100011110",
  57016=>"000001000",
  57017=>"001011001",
  57018=>"101001001",
  57019=>"000000111",
  57020=>"101000101",
  57021=>"001001101",
  57022=>"111101010",
  57023=>"111011010",
  57024=>"011011000",
  57025=>"110110100",
  57026=>"110001100",
  57027=>"110011101",
  57028=>"101110100",
  57029=>"001010111",
  57030=>"010110100",
  57031=>"110010100",
  57032=>"000111101",
  57033=>"000010010",
  57034=>"111100101",
  57035=>"110100011",
  57036=>"100001100",
  57037=>"000001111",
  57038=>"111001001",
  57039=>"100101111",
  57040=>"000100001",
  57041=>"101110000",
  57042=>"111100000",
  57043=>"111001100",
  57044=>"100010010",
  57045=>"011110001",
  57046=>"101001111",
  57047=>"100000110",
  57048=>"101001000",
  57049=>"011100100",
  57050=>"000000101",
  57051=>"111001010",
  57052=>"111011110",
  57053=>"100011001",
  57054=>"111110001",
  57055=>"001010111",
  57056=>"110001010",
  57057=>"101101011",
  57058=>"101011110",
  57059=>"010111010",
  57060=>"001100010",
  57061=>"110000111",
  57062=>"001110110",
  57063=>"011001011",
  57064=>"010110101",
  57065=>"000011100",
  57066=>"100110010",
  57067=>"101011111",
  57068=>"000111010",
  57069=>"011111110",
  57070=>"010011001",
  57071=>"000001000",
  57072=>"110011101",
  57073=>"110001110",
  57074=>"001001001",
  57075=>"010111110",
  57076=>"110111010",
  57077=>"010000000",
  57078=>"101110101",
  57079=>"001011110",
  57080=>"010111101",
  57081=>"100011100",
  57082=>"001101101",
  57083=>"011100100",
  57084=>"110111111",
  57085=>"110110111",
  57086=>"001001100",
  57087=>"110010000",
  57088=>"000010011",
  57089=>"100010011",
  57090=>"101001000",
  57091=>"010000000",
  57092=>"101001011",
  57093=>"110001011",
  57094=>"011000101",
  57095=>"111000111",
  57096=>"100110101",
  57097=>"010010110",
  57098=>"101001000",
  57099=>"100110001",
  57100=>"001111010",
  57101=>"001100101",
  57102=>"111001000",
  57103=>"001101100",
  57104=>"000000000",
  57105=>"111010010",
  57106=>"010011010",
  57107=>"001110100",
  57108=>"010000001",
  57109=>"111110000",
  57110=>"101010101",
  57111=>"110011001",
  57112=>"000000101",
  57113=>"000000001",
  57114=>"011111111",
  57115=>"010001110",
  57116=>"110110111",
  57117=>"001101110",
  57118=>"100000110",
  57119=>"110111100",
  57120=>"000100101",
  57121=>"000110111",
  57122=>"100000001",
  57123=>"010101101",
  57124=>"011101100",
  57125=>"000000011",
  57126=>"101001011",
  57127=>"111011101",
  57128=>"110110110",
  57129=>"011010110",
  57130=>"000110011",
  57131=>"110110001",
  57132=>"010100100",
  57133=>"100010110",
  57134=>"100001001",
  57135=>"100110000",
  57136=>"000110101",
  57137=>"011010101",
  57138=>"011001001",
  57139=>"001001101",
  57140=>"010011000",
  57141=>"011100001",
  57142=>"111000111",
  57143=>"101101111",
  57144=>"111011111",
  57145=>"000110110",
  57146=>"111000000",
  57147=>"110101010",
  57148=>"010110010",
  57149=>"101101101",
  57150=>"111001110",
  57151=>"000101000",
  57152=>"010100100",
  57153=>"001100010",
  57154=>"010011010",
  57155=>"011101000",
  57156=>"011010010",
  57157=>"000101011",
  57158=>"001111100",
  57159=>"000111001",
  57160=>"001111100",
  57161=>"101010001",
  57162=>"110110110",
  57163=>"110110001",
  57164=>"100011100",
  57165=>"000011011",
  57166=>"110010001",
  57167=>"100101100",
  57168=>"000111011",
  57169=>"111100000",
  57170=>"010000001",
  57171=>"001111010",
  57172=>"100100001",
  57173=>"010010101",
  57174=>"010110100",
  57175=>"011000000",
  57176=>"101000101",
  57177=>"100110100",
  57178=>"011010111",
  57179=>"000100110",
  57180=>"110100011",
  57181=>"000111010",
  57182=>"010000011",
  57183=>"000110100",
  57184=>"100111100",
  57185=>"000110010",
  57186=>"100101011",
  57187=>"011010101",
  57188=>"000111011",
  57189=>"011001110",
  57190=>"011110000",
  57191=>"010000010",
  57192=>"011000111",
  57193=>"001100010",
  57194=>"111100001",
  57195=>"111111011",
  57196=>"110000100",
  57197=>"000111011",
  57198=>"100001111",
  57199=>"001010101",
  57200=>"100010000",
  57201=>"000000001",
  57202=>"000011111",
  57203=>"000100000",
  57204=>"010101101",
  57205=>"010100101",
  57206=>"000001000",
  57207=>"000010100",
  57208=>"111011001",
  57209=>"100010111",
  57210=>"111100010",
  57211=>"110001110",
  57212=>"000011000",
  57213=>"100000000",
  57214=>"000001000",
  57215=>"001111101",
  57216=>"011101001",
  57217=>"001110101",
  57218=>"110100100",
  57219=>"111000000",
  57220=>"101111101",
  57221=>"000001000",
  57222=>"011101111",
  57223=>"110011111",
  57224=>"100011011",
  57225=>"010100001",
  57226=>"000001110",
  57227=>"111010111",
  57228=>"000110111",
  57229=>"000111010",
  57230=>"000011000",
  57231=>"000100000",
  57232=>"110010010",
  57233=>"010111101",
  57234=>"100110010",
  57235=>"001111101",
  57236=>"110110110",
  57237=>"011010101",
  57238=>"111111010",
  57239=>"100000100",
  57240=>"011100000",
  57241=>"010110001",
  57242=>"101100111",
  57243=>"001011011",
  57244=>"110111001",
  57245=>"001011010",
  57246=>"001100111",
  57247=>"000010001",
  57248=>"010000110",
  57249=>"111111010",
  57250=>"010000011",
  57251=>"101110111",
  57252=>"110101001",
  57253=>"101110111",
  57254=>"000111101",
  57255=>"111010111",
  57256=>"101010101",
  57257=>"001101001",
  57258=>"110111001",
  57259=>"010000110",
  57260=>"111111000",
  57261=>"010110001",
  57262=>"100111110",
  57263=>"010111011",
  57264=>"000001100",
  57265=>"001001011",
  57266=>"011100110",
  57267=>"111001110",
  57268=>"010011101",
  57269=>"111010011",
  57270=>"100000100",
  57271=>"110011001",
  57272=>"001110000",
  57273=>"111100100",
  57274=>"001101001",
  57275=>"110110000",
  57276=>"110011111",
  57277=>"100010011",
  57278=>"100100111",
  57279=>"100100000",
  57280=>"101111011",
  57281=>"101000111",
  57282=>"010101000",
  57283=>"100100000",
  57284=>"000011011",
  57285=>"110010110",
  57286=>"101110010",
  57287=>"011110000",
  57288=>"010001111",
  57289=>"000111110",
  57290=>"011111011",
  57291=>"000111100",
  57292=>"111001011",
  57293=>"010001001",
  57294=>"101011000",
  57295=>"011000101",
  57296=>"110110101",
  57297=>"001000100",
  57298=>"011111000",
  57299=>"111110010",
  57300=>"000111111",
  57301=>"000111011",
  57302=>"111111001",
  57303=>"101110011",
  57304=>"101110100",
  57305=>"110111010",
  57306=>"111000001",
  57307=>"010001001",
  57308=>"001100010",
  57309=>"111011110",
  57310=>"110000101",
  57311=>"000001111",
  57312=>"010100011",
  57313=>"100110001",
  57314=>"000011101",
  57315=>"000100001",
  57316=>"100010100",
  57317=>"011000011",
  57318=>"000100001",
  57319=>"100011000",
  57320=>"101001101",
  57321=>"110110111",
  57322=>"101010000",
  57323=>"100001001",
  57324=>"100100011",
  57325=>"011010001",
  57326=>"001010001",
  57327=>"000110000",
  57328=>"010001001",
  57329=>"001111101",
  57330=>"001000011",
  57331=>"111000000",
  57332=>"011110111",
  57333=>"000010000",
  57334=>"000000100",
  57335=>"001011000",
  57336=>"001010000",
  57337=>"000010000",
  57338=>"101000011",
  57339=>"110100101",
  57340=>"001010011",
  57341=>"101011000",
  57342=>"001101101",
  57343=>"111111001",
  57344=>"000000001",
  57345=>"011110000",
  57346=>"100100001",
  57347=>"010010000",
  57348=>"111010101",
  57349=>"110111000",
  57350=>"010011011",
  57351=>"000111101",
  57352=>"011010010",
  57353=>"010011011",
  57354=>"010100000",
  57355=>"101000000",
  57356=>"111000000",
  57357=>"011001010",
  57358=>"101011111",
  57359=>"011111011",
  57360=>"100111011",
  57361=>"001101001",
  57362=>"010111001",
  57363=>"110001100",
  57364=>"000010011",
  57365=>"010100110",
  57366=>"111011100",
  57367=>"110111001",
  57368=>"000100101",
  57369=>"100110101",
  57370=>"001010110",
  57371=>"100101011",
  57372=>"010010010",
  57373=>"001111111",
  57374=>"100101001",
  57375=>"101010100",
  57376=>"100010101",
  57377=>"110011101",
  57378=>"100101011",
  57379=>"101010011",
  57380=>"100000001",
  57381=>"110001011",
  57382=>"010001110",
  57383=>"001110111",
  57384=>"100000010",
  57385=>"000101011",
  57386=>"100010001",
  57387=>"011110101",
  57388=>"010110010",
  57389=>"111110111",
  57390=>"010000101",
  57391=>"110100100",
  57392=>"101000010",
  57393=>"111111111",
  57394=>"111111100",
  57395=>"111010100",
  57396=>"110110111",
  57397=>"001011011",
  57398=>"101001101",
  57399=>"110110110",
  57400=>"001001001",
  57401=>"110011100",
  57402=>"111110110",
  57403=>"011010011",
  57404=>"011010110",
  57405=>"110110100",
  57406=>"111000111",
  57407=>"010100001",
  57408=>"010000001",
  57409=>"000101001",
  57410=>"001101011",
  57411=>"011001000",
  57412=>"011110100",
  57413=>"011010111",
  57414=>"101011011",
  57415=>"111001011",
  57416=>"001110010",
  57417=>"111000100",
  57418=>"000111101",
  57419=>"001000110",
  57420=>"001011101",
  57421=>"011001010",
  57422=>"001011001",
  57423=>"011011000",
  57424=>"110010110",
  57425=>"101000010",
  57426=>"110100000",
  57427=>"110010110",
  57428=>"111011110",
  57429=>"011010101",
  57430=>"101101110",
  57431=>"000000101",
  57432=>"000000110",
  57433=>"001101110",
  57434=>"010010111",
  57435=>"000111001",
  57436=>"101101010",
  57437=>"000101001",
  57438=>"101110110",
  57439=>"010010001",
  57440=>"101010000",
  57441=>"010100111",
  57442=>"000110001",
  57443=>"100101000",
  57444=>"100001100",
  57445=>"101100001",
  57446=>"110000010",
  57447=>"101011010",
  57448=>"001001000",
  57449=>"001010011",
  57450=>"000011111",
  57451=>"100001110",
  57452=>"100011000",
  57453=>"000000011",
  57454=>"001000110",
  57455=>"000100100",
  57456=>"010111110",
  57457=>"101110010",
  57458=>"111110010",
  57459=>"101110100",
  57460=>"010111011",
  57461=>"000111111",
  57462=>"010111100",
  57463=>"100100110",
  57464=>"001111000",
  57465=>"100101010",
  57466=>"101111010",
  57467=>"100110100",
  57468=>"001101100",
  57469=>"100010010",
  57470=>"000111110",
  57471=>"001000011",
  57472=>"010110110",
  57473=>"000100010",
  57474=>"100011101",
  57475=>"001000010",
  57476=>"110100100",
  57477=>"001010011",
  57478=>"011100101",
  57479=>"100010010",
  57480=>"011111101",
  57481=>"010010000",
  57482=>"010111001",
  57483=>"000110000",
  57484=>"010100011",
  57485=>"110100011",
  57486=>"011100101",
  57487=>"110010101",
  57488=>"001011001",
  57489=>"001011011",
  57490=>"100101101",
  57491=>"100110100",
  57492=>"000001110",
  57493=>"100110100",
  57494=>"010011011",
  57495=>"101100001",
  57496=>"101011000",
  57497=>"100100001",
  57498=>"010100111",
  57499=>"110011110",
  57500=>"101110100",
  57501=>"110111011",
  57502=>"101100110",
  57503=>"011110101",
  57504=>"100000001",
  57505=>"001100111",
  57506=>"100011111",
  57507=>"001000110",
  57508=>"110101011",
  57509=>"110011001",
  57510=>"110011000",
  57511=>"101101000",
  57512=>"111100011",
  57513=>"101110010",
  57514=>"011000000",
  57515=>"000001000",
  57516=>"110100000",
  57517=>"001101111",
  57518=>"001110000",
  57519=>"001001111",
  57520=>"001001100",
  57521=>"111000101",
  57522=>"001100010",
  57523=>"100110011",
  57524=>"001101110",
  57525=>"110010000",
  57526=>"011110101",
  57527=>"000011000",
  57528=>"111101010",
  57529=>"010011100",
  57530=>"101000101",
  57531=>"110101100",
  57532=>"101110010",
  57533=>"001101010",
  57534=>"101010001",
  57535=>"011011011",
  57536=>"010000011",
  57537=>"000011010",
  57538=>"101111101",
  57539=>"001011101",
  57540=>"100011110",
  57541=>"000101110",
  57542=>"000011010",
  57543=>"100111101",
  57544=>"111111100",
  57545=>"111110001",
  57546=>"101101101",
  57547=>"011001110",
  57548=>"111100110",
  57549=>"001110010",
  57550=>"010101001",
  57551=>"101000100",
  57552=>"000000000",
  57553=>"010101010",
  57554=>"010111101",
  57555=>"111011101",
  57556=>"011100101",
  57557=>"000000101",
  57558=>"110011001",
  57559=>"110101101",
  57560=>"101010000",
  57561=>"001011011",
  57562=>"011111011",
  57563=>"100111000",
  57564=>"101011110",
  57565=>"100011001",
  57566=>"000001101",
  57567=>"011100111",
  57568=>"101101100",
  57569=>"101010111",
  57570=>"101000001",
  57571=>"010001111",
  57572=>"110111010",
  57573=>"011101011",
  57574=>"101111000",
  57575=>"010011010",
  57576=>"110110100",
  57577=>"110011001",
  57578=>"011011010",
  57579=>"011111100",
  57580=>"101010111",
  57581=>"010111111",
  57582=>"000000011",
  57583=>"000100001",
  57584=>"010000100",
  57585=>"010010000",
  57586=>"100100110",
  57587=>"011111001",
  57588=>"111110110",
  57589=>"111000010",
  57590=>"110111001",
  57591=>"111001011",
  57592=>"000111000",
  57593=>"100011111",
  57594=>"010111101",
  57595=>"100001000",
  57596=>"001010011",
  57597=>"010000100",
  57598=>"000011111",
  57599=>"001100110",
  57600=>"110110111",
  57601=>"001101101",
  57602=>"001001100",
  57603=>"111111011",
  57604=>"011001110",
  57605=>"111011110",
  57606=>"010100110",
  57607=>"010100000",
  57608=>"000111111",
  57609=>"001101010",
  57610=>"101111001",
  57611=>"010100111",
  57612=>"001010100",
  57613=>"000100000",
  57614=>"100101010",
  57615=>"000001110",
  57616=>"001000011",
  57617=>"001000011",
  57618=>"001100110",
  57619=>"111111001",
  57620=>"111011011",
  57621=>"011001110",
  57622=>"000011100",
  57623=>"010001000",
  57624=>"100110100",
  57625=>"100101110",
  57626=>"011100010",
  57627=>"111010010",
  57628=>"000101110",
  57629=>"011011101",
  57630=>"001101001",
  57631=>"110001111",
  57632=>"111111100",
  57633=>"010001111",
  57634=>"000000110",
  57635=>"000011001",
  57636=>"101111011",
  57637=>"111101101",
  57638=>"110000001",
  57639=>"000101000",
  57640=>"001101001",
  57641=>"011011001",
  57642=>"001010110",
  57643=>"000001100",
  57644=>"110011011",
  57645=>"100000011",
  57646=>"000100011",
  57647=>"111100100",
  57648=>"101100011",
  57649=>"111110001",
  57650=>"100101010",
  57651=>"110111110",
  57652=>"101010101",
  57653=>"000100010",
  57654=>"000000110",
  57655=>"111111011",
  57656=>"111110100",
  57657=>"010011101",
  57658=>"011001111",
  57659=>"101000110",
  57660=>"000110000",
  57661=>"000100111",
  57662=>"010001101",
  57663=>"101100000",
  57664=>"100000000",
  57665=>"100000000",
  57666=>"001100110",
  57667=>"101100000",
  57668=>"111011011",
  57669=>"101000100",
  57670=>"110011011",
  57671=>"010100001",
  57672=>"000111110",
  57673=>"010010000",
  57674=>"101101010",
  57675=>"000001111",
  57676=>"111101001",
  57677=>"011101100",
  57678=>"011000100",
  57679=>"101001010",
  57680=>"001000001",
  57681=>"010001011",
  57682=>"010101011",
  57683=>"001101010",
  57684=>"111101111",
  57685=>"011000011",
  57686=>"100100010",
  57687=>"010000010",
  57688=>"000000111",
  57689=>"010011101",
  57690=>"100000000",
  57691=>"110100101",
  57692=>"000000110",
  57693=>"111101110",
  57694=>"011101101",
  57695=>"000001110",
  57696=>"001010011",
  57697=>"001010001",
  57698=>"101111110",
  57699=>"001110010",
  57700=>"101000001",
  57701=>"000100110",
  57702=>"110100111",
  57703=>"111010111",
  57704=>"111000010",
  57705=>"010011011",
  57706=>"100101010",
  57707=>"010011000",
  57708=>"001001000",
  57709=>"001111001",
  57710=>"100010011",
  57711=>"011000000",
  57712=>"000001100",
  57713=>"100101110",
  57714=>"010101111",
  57715=>"011111100",
  57716=>"010011101",
  57717=>"101101101",
  57718=>"100110000",
  57719=>"000010111",
  57720=>"010000001",
  57721=>"000000011",
  57722=>"100100011",
  57723=>"011001010",
  57724=>"110001001",
  57725=>"100111000",
  57726=>"000011110",
  57727=>"101101010",
  57728=>"101001110",
  57729=>"011110110",
  57730=>"110110111",
  57731=>"010101011",
  57732=>"101000000",
  57733=>"010100111",
  57734=>"100011100",
  57735=>"011001110",
  57736=>"101110100",
  57737=>"110111100",
  57738=>"111100101",
  57739=>"101101010",
  57740=>"111100111",
  57741=>"111101001",
  57742=>"101101100",
  57743=>"000111111",
  57744=>"101010010",
  57745=>"001010000",
  57746=>"000101111",
  57747=>"010001010",
  57748=>"100010000",
  57749=>"111111100",
  57750=>"011000011",
  57751=>"110001010",
  57752=>"010110011",
  57753=>"011000001",
  57754=>"100000111",
  57755=>"010100010",
  57756=>"101001001",
  57757=>"100100011",
  57758=>"000100010",
  57759=>"000110000",
  57760=>"001001000",
  57761=>"111010110",
  57762=>"101000111",
  57763=>"101010110",
  57764=>"111100110",
  57765=>"111111010",
  57766=>"001000001",
  57767=>"000100000",
  57768=>"110000000",
  57769=>"010101011",
  57770=>"111101100",
  57771=>"000101010",
  57772=>"000110000",
  57773=>"111001110",
  57774=>"110111111",
  57775=>"010101000",
  57776=>"000011011",
  57777=>"011000111",
  57778=>"011001101",
  57779=>"010111100",
  57780=>"110101010",
  57781=>"000001110",
  57782=>"000011101",
  57783=>"110011100",
  57784=>"000110101",
  57785=>"000111110",
  57786=>"000010001",
  57787=>"011111110",
  57788=>"111101100",
  57789=>"101101001",
  57790=>"111001010",
  57791=>"010101111",
  57792=>"110101010",
  57793=>"001111101",
  57794=>"100110110",
  57795=>"110011001",
  57796=>"110111111",
  57797=>"001001110",
  57798=>"111010001",
  57799=>"100100011",
  57800=>"000111011",
  57801=>"001000100",
  57802=>"010011111",
  57803=>"101101110",
  57804=>"110111100",
  57805=>"100111110",
  57806=>"000000011",
  57807=>"110000100",
  57808=>"110101001",
  57809=>"010000010",
  57810=>"111011110",
  57811=>"110000101",
  57812=>"000100011",
  57813=>"001111101",
  57814=>"010010011",
  57815=>"101110001",
  57816=>"000110000",
  57817=>"111110110",
  57818=>"010100111",
  57819=>"110101110",
  57820=>"101100011",
  57821=>"111110100",
  57822=>"000000011",
  57823=>"010001111",
  57824=>"100111010",
  57825=>"011110010",
  57826=>"000100100",
  57827=>"000100111",
  57828=>"000101101",
  57829=>"101001110",
  57830=>"011111100",
  57831=>"100100001",
  57832=>"011110000",
  57833=>"010000111",
  57834=>"000100000",
  57835=>"100010000",
  57836=>"010011111",
  57837=>"110111010",
  57838=>"100101110",
  57839=>"010011000",
  57840=>"110011101",
  57841=>"000101011",
  57842=>"000100011",
  57843=>"011011101",
  57844=>"110011001",
  57845=>"100101010",
  57846=>"010111111",
  57847=>"101111110",
  57848=>"001110010",
  57849=>"110000000",
  57850=>"101010100",
  57851=>"101000000",
  57852=>"111110001",
  57853=>"000010011",
  57854=>"011111001",
  57855=>"101000000",
  57856=>"100001100",
  57857=>"000010000",
  57858=>"000101110",
  57859=>"010110111",
  57860=>"111010111",
  57861=>"001000101",
  57862=>"110101110",
  57863=>"010001010",
  57864=>"000011000",
  57865=>"110111111",
  57866=>"111010111",
  57867=>"000001110",
  57868=>"010001100",
  57869=>"001111000",
  57870=>"110110001",
  57871=>"000100010",
  57872=>"100000110",
  57873=>"111100011",
  57874=>"010010111",
  57875=>"110011011",
  57876=>"111000100",
  57877=>"101110000",
  57878=>"110000111",
  57879=>"000101110",
  57880=>"100100100",
  57881=>"000010101",
  57882=>"111011111",
  57883=>"101101101",
  57884=>"011110000",
  57885=>"010000011",
  57886=>"111110011",
  57887=>"001110101",
  57888=>"000010101",
  57889=>"100111011",
  57890=>"000100000",
  57891=>"110111100",
  57892=>"111111101",
  57893=>"011111111",
  57894=>"001111011",
  57895=>"111010110",
  57896=>"110010111",
  57897=>"011001111",
  57898=>"011110011",
  57899=>"001010100",
  57900=>"111100100",
  57901=>"000001000",
  57902=>"011000110",
  57903=>"000000100",
  57904=>"011101100",
  57905=>"101110010",
  57906=>"111110011",
  57907=>"110001111",
  57908=>"110101111",
  57909=>"111000110",
  57910=>"101111111",
  57911=>"111000101",
  57912=>"111010000",
  57913=>"110110100",
  57914=>"011000011",
  57915=>"101111011",
  57916=>"001001110",
  57917=>"100110111",
  57918=>"010100110",
  57919=>"101000010",
  57920=>"101010111",
  57921=>"001111000",
  57922=>"011111010",
  57923=>"111100101",
  57924=>"101010011",
  57925=>"110101111",
  57926=>"100101111",
  57927=>"111101111",
  57928=>"100110110",
  57929=>"111001101",
  57930=>"101010011",
  57931=>"101001001",
  57932=>"010111010",
  57933=>"000010100",
  57934=>"000111010",
  57935=>"000111010",
  57936=>"111100000",
  57937=>"010110110",
  57938=>"101000111",
  57939=>"010111110",
  57940=>"010000110",
  57941=>"011001010",
  57942=>"000110011",
  57943=>"001010100",
  57944=>"010001001",
  57945=>"111001001",
  57946=>"000001100",
  57947=>"010100100",
  57948=>"101111011",
  57949=>"110011111",
  57950=>"000100010",
  57951=>"110111000",
  57952=>"100111001",
  57953=>"000100000",
  57954=>"000000100",
  57955=>"111011001",
  57956=>"100000001",
  57957=>"011011011",
  57958=>"110000111",
  57959=>"100100111",
  57960=>"010000110",
  57961=>"010111110",
  57962=>"010100000",
  57963=>"111001101",
  57964=>"000110101",
  57965=>"100000000",
  57966=>"100100111",
  57967=>"110000110",
  57968=>"001100001",
  57969=>"011100000",
  57970=>"010000010",
  57971=>"101110000",
  57972=>"111000010",
  57973=>"110000111",
  57974=>"100111111",
  57975=>"001011001",
  57976=>"000010001",
  57977=>"110000110",
  57978=>"001111100",
  57979=>"000001100",
  57980=>"001110010",
  57981=>"100110110",
  57982=>"100010101",
  57983=>"010110011",
  57984=>"011000101",
  57985=>"111111011",
  57986=>"101011101",
  57987=>"101000011",
  57988=>"101000100",
  57989=>"100011000",
  57990=>"110110010",
  57991=>"110010000",
  57992=>"101010001",
  57993=>"100100111",
  57994=>"010100111",
  57995=>"011110011",
  57996=>"011010000",
  57997=>"100000011",
  57998=>"000000010",
  57999=>"001001010",
  58000=>"001111110",
  58001=>"001110011",
  58002=>"110100101",
  58003=>"001111101",
  58004=>"000001001",
  58005=>"110100011",
  58006=>"111001010",
  58007=>"000101010",
  58008=>"000001001",
  58009=>"111000010",
  58010=>"000101001",
  58011=>"011001100",
  58012=>"011000011",
  58013=>"101101110",
  58014=>"011111010",
  58015=>"000011000",
  58016=>"000010010",
  58017=>"110001001",
  58018=>"111010111",
  58019=>"110000111",
  58020=>"011111111",
  58021=>"101010101",
  58022=>"110110111",
  58023=>"110110001",
  58024=>"001111000",
  58025=>"010010101",
  58026=>"101100000",
  58027=>"111111001",
  58028=>"011011101",
  58029=>"000110100",
  58030=>"011000101",
  58031=>"100001011",
  58032=>"100010111",
  58033=>"110011110",
  58034=>"110101110",
  58035=>"111111000",
  58036=>"000011000",
  58037=>"000100011",
  58038=>"110110100",
  58039=>"001011011",
  58040=>"001011110",
  58041=>"111001100",
  58042=>"111111010",
  58043=>"000101111",
  58044=>"100101010",
  58045=>"000101001",
  58046=>"100011010",
  58047=>"000111001",
  58048=>"110001100",
  58049=>"100000110",
  58050=>"101001101",
  58051=>"000101110",
  58052=>"000011101",
  58053=>"101101101",
  58054=>"010010010",
  58055=>"001000111",
  58056=>"110100000",
  58057=>"111100110",
  58058=>"110000011",
  58059=>"000001010",
  58060=>"010100011",
  58061=>"100000011",
  58062=>"010111011",
  58063=>"000101010",
  58064=>"101010011",
  58065=>"010101111",
  58066=>"101011100",
  58067=>"100110110",
  58068=>"001101100",
  58069=>"100110011",
  58070=>"011000001",
  58071=>"111011010",
  58072=>"111000010",
  58073=>"000001111",
  58074=>"001001101",
  58075=>"110110000",
  58076=>"100010011",
  58077=>"110101100",
  58078=>"011110101",
  58079=>"010111010",
  58080=>"010110000",
  58081=>"010000101",
  58082=>"100110110",
  58083=>"011111111",
  58084=>"001001110",
  58085=>"111000101",
  58086=>"100111101",
  58087=>"111010001",
  58088=>"010101000",
  58089=>"011010111",
  58090=>"001001011",
  58091=>"000101000",
  58092=>"000100101",
  58093=>"110001011",
  58094=>"010000011",
  58095=>"001100101",
  58096=>"110101100",
  58097=>"110000100",
  58098=>"010110101",
  58099=>"001000010",
  58100=>"011101100",
  58101=>"001100110",
  58102=>"011111101",
  58103=>"010010000",
  58104=>"110100100",
  58105=>"110000100",
  58106=>"111000110",
  58107=>"000110110",
  58108=>"101001001",
  58109=>"001111111",
  58110=>"111011011",
  58111=>"000101001",
  58112=>"101001010",
  58113=>"000101101",
  58114=>"010011110",
  58115=>"011010000",
  58116=>"010110111",
  58117=>"101111000",
  58118=>"001011011",
  58119=>"011110101",
  58120=>"000110100",
  58121=>"111011100",
  58122=>"101010001",
  58123=>"100110000",
  58124=>"111010110",
  58125=>"011001100",
  58126=>"110100011",
  58127=>"010010011",
  58128=>"000001001",
  58129=>"100000000",
  58130=>"100100111",
  58131=>"010101111",
  58132=>"110010101",
  58133=>"110001000",
  58134=>"000101010",
  58135=>"110101001",
  58136=>"101010111",
  58137=>"101100100",
  58138=>"100111100",
  58139=>"001101001",
  58140=>"111101110",
  58141=>"110011011",
  58142=>"111010110",
  58143=>"101100000",
  58144=>"010010011",
  58145=>"000010110",
  58146=>"010111001",
  58147=>"000111010",
  58148=>"000010101",
  58149=>"010110101",
  58150=>"111010011",
  58151=>"011101111",
  58152=>"000111000",
  58153=>"100011001",
  58154=>"010000111",
  58155=>"100110101",
  58156=>"100001110",
  58157=>"010100010",
  58158=>"100000011",
  58159=>"100101101",
  58160=>"110100010",
  58161=>"100011000",
  58162=>"100101100",
  58163=>"111100110",
  58164=>"100011000",
  58165=>"001110000",
  58166=>"101110111",
  58167=>"101001000",
  58168=>"100111001",
  58169=>"100101101",
  58170=>"111000000",
  58171=>"001101010",
  58172=>"010101011",
  58173=>"100111100",
  58174=>"111101001",
  58175=>"010010100",
  58176=>"110110100",
  58177=>"011101111",
  58178=>"001101100",
  58179=>"000011001",
  58180=>"111100000",
  58181=>"100000000",
  58182=>"001100001",
  58183=>"110001101",
  58184=>"011101111",
  58185=>"100100110",
  58186=>"101011000",
  58187=>"000000100",
  58188=>"001000000",
  58189=>"111100110",
  58190=>"000111001",
  58191=>"000000010",
  58192=>"101100101",
  58193=>"100111001",
  58194=>"100100111",
  58195=>"100000101",
  58196=>"010101000",
  58197=>"010001000",
  58198=>"000100010",
  58199=>"001000101",
  58200=>"010001100",
  58201=>"011110010",
  58202=>"011100001",
  58203=>"010011101",
  58204=>"010101001",
  58205=>"000110011",
  58206=>"110100110",
  58207=>"000010110",
  58208=>"000100010",
  58209=>"001000010",
  58210=>"001010001",
  58211=>"011111010",
  58212=>"110000100",
  58213=>"000001100",
  58214=>"110100011",
  58215=>"101000000",
  58216=>"110000111",
  58217=>"111011101",
  58218=>"100101001",
  58219=>"001000001",
  58220=>"110010011",
  58221=>"111001100",
  58222=>"001100110",
  58223=>"011111110",
  58224=>"110101010",
  58225=>"001011110",
  58226=>"001111000",
  58227=>"101011010",
  58228=>"011100001",
  58229=>"101011100",
  58230=>"000000100",
  58231=>"111111111",
  58232=>"110111010",
  58233=>"000011111",
  58234=>"011100100",
  58235=>"111000001",
  58236=>"000000000",
  58237=>"101011000",
  58238=>"100111010",
  58239=>"000001011",
  58240=>"110111100",
  58241=>"011000101",
  58242=>"011101000",
  58243=>"101000110",
  58244=>"010011000",
  58245=>"010011101",
  58246=>"110111101",
  58247=>"010000110",
  58248=>"101010110",
  58249=>"010010001",
  58250=>"101101011",
  58251=>"101110111",
  58252=>"001100001",
  58253=>"010010000",
  58254=>"111100101",
  58255=>"111000000",
  58256=>"101110111",
  58257=>"010101100",
  58258=>"100000010",
  58259=>"010101000",
  58260=>"100110111",
  58261=>"100010111",
  58262=>"101110000",
  58263=>"010111100",
  58264=>"001011000",
  58265=>"110000100",
  58266=>"011110100",
  58267=>"000100000",
  58268=>"110010011",
  58269=>"110001110",
  58270=>"111101010",
  58271=>"011110111",
  58272=>"000100100",
  58273=>"101001111",
  58274=>"010100111",
  58275=>"010111010",
  58276=>"001011011",
  58277=>"011111001",
  58278=>"011010111",
  58279=>"111101011",
  58280=>"000000100",
  58281=>"001001100",
  58282=>"000110011",
  58283=>"010110001",
  58284=>"011000011",
  58285=>"110010000",
  58286=>"111011101",
  58287=>"001111111",
  58288=>"101010101",
  58289=>"111111111",
  58290=>"011000110",
  58291=>"000000111",
  58292=>"100011010",
  58293=>"000110110",
  58294=>"010010001",
  58295=>"011011000",
  58296=>"111010010",
  58297=>"101101010",
  58298=>"011000110",
  58299=>"010011001",
  58300=>"010100101",
  58301=>"001100001",
  58302=>"110010110",
  58303=>"110001011",
  58304=>"111101111",
  58305=>"101101001",
  58306=>"001110101",
  58307=>"111110000",
  58308=>"010010010",
  58309=>"111000010",
  58310=>"010001110",
  58311=>"001101111",
  58312=>"010110010",
  58313=>"010001001",
  58314=>"101001010",
  58315=>"111111111",
  58316=>"110011000",
  58317=>"111101010",
  58318=>"011011000",
  58319=>"101000000",
  58320=>"010110011",
  58321=>"010000000",
  58322=>"101101110",
  58323=>"000010111",
  58324=>"000000110",
  58325=>"111110001",
  58326=>"000000110",
  58327=>"110111101",
  58328=>"010101100",
  58329=>"001101011",
  58330=>"100111001",
  58331=>"011101000",
  58332=>"101001110",
  58333=>"111110111",
  58334=>"110101111",
  58335=>"010110000",
  58336=>"010000011",
  58337=>"010011000",
  58338=>"100110000",
  58339=>"110100011",
  58340=>"010100000",
  58341=>"011011110",
  58342=>"000110111",
  58343=>"000010110",
  58344=>"111111011",
  58345=>"100110101",
  58346=>"100001001",
  58347=>"110101101",
  58348=>"000101010",
  58349=>"001000110",
  58350=>"011100001",
  58351=>"011100000",
  58352=>"000010111",
  58353=>"000010011",
  58354=>"111011110",
  58355=>"010010000",
  58356=>"100001111",
  58357=>"000110110",
  58358=>"111111110",
  58359=>"001110011",
  58360=>"101001100",
  58361=>"000110001",
  58362=>"001110101",
  58363=>"110111110",
  58364=>"111110001",
  58365=>"010010011",
  58366=>"001010001",
  58367=>"101011011",
  58368=>"110101111",
  58369=>"100001001",
  58370=>"111010111",
  58371=>"101111101",
  58372=>"100000101",
  58373=>"011010001",
  58374=>"011011111",
  58375=>"110000010",
  58376=>"111111110",
  58377=>"100110000",
  58378=>"001110111",
  58379=>"000000011",
  58380=>"110010100",
  58381=>"100010100",
  58382=>"010100001",
  58383=>"110111010",
  58384=>"000000011",
  58385=>"111011001",
  58386=>"110111100",
  58387=>"100110111",
  58388=>"000001110",
  58389=>"111111101",
  58390=>"110001100",
  58391=>"110000000",
  58392=>"000001011",
  58393=>"011011101",
  58394=>"001101101",
  58395=>"110010101",
  58396=>"011001111",
  58397=>"111001110",
  58398=>"100100110",
  58399=>"001011111",
  58400=>"111011011",
  58401=>"110001001",
  58402=>"111100001",
  58403=>"001011110",
  58404=>"110011110",
  58405=>"101101011",
  58406=>"011110011",
  58407=>"011101111",
  58408=>"101110000",
  58409=>"110111000",
  58410=>"100000010",
  58411=>"010010000",
  58412=>"001101111",
  58413=>"011101010",
  58414=>"000101110",
  58415=>"011100010",
  58416=>"001111110",
  58417=>"011110011",
  58418=>"000110000",
  58419=>"001010000",
  58420=>"110101101",
  58421=>"100100111",
  58422=>"110011100",
  58423=>"001111110",
  58424=>"110011000",
  58425=>"101101101",
  58426=>"001000101",
  58427=>"111100111",
  58428=>"000111111",
  58429=>"011100111",
  58430=>"101101100",
  58431=>"111100110",
  58432=>"001100101",
  58433=>"100000011",
  58434=>"101100110",
  58435=>"111100101",
  58436=>"000011000",
  58437=>"101000010",
  58438=>"110100100",
  58439=>"001111011",
  58440=>"000000011",
  58441=>"010101000",
  58442=>"010011011",
  58443=>"000111001",
  58444=>"111001101",
  58445=>"110101101",
  58446=>"101100000",
  58447=>"100100000",
  58448=>"111100100",
  58449=>"001011010",
  58450=>"110101011",
  58451=>"001111000",
  58452=>"001110011",
  58453=>"111101010",
  58454=>"110100110",
  58455=>"100011100",
  58456=>"110111000",
  58457=>"110100100",
  58458=>"010000000",
  58459=>"001000011",
  58460=>"011001110",
  58461=>"110110000",
  58462=>"011110110",
  58463=>"011100011",
  58464=>"011010110",
  58465=>"110000011",
  58466=>"010110000",
  58467=>"010110100",
  58468=>"110111100",
  58469=>"111011110",
  58470=>"101110101",
  58471=>"110101001",
  58472=>"010001001",
  58473=>"111111110",
  58474=>"011100101",
  58475=>"100001111",
  58476=>"110101001",
  58477=>"001100010",
  58478=>"011011000",
  58479=>"001001001",
  58480=>"000000000",
  58481=>"000011000",
  58482=>"011010001",
  58483=>"011000100",
  58484=>"100001111",
  58485=>"001100110",
  58486=>"010111100",
  58487=>"110011011",
  58488=>"111001000",
  58489=>"101100010",
  58490=>"100011100",
  58491=>"111101010",
  58492=>"011001001",
  58493=>"111011111",
  58494=>"001110111",
  58495=>"000100001",
  58496=>"110101000",
  58497=>"011001111",
  58498=>"000010101",
  58499=>"111110101",
  58500=>"110111000",
  58501=>"011101001",
  58502=>"110011000",
  58503=>"001010000",
  58504=>"000010011",
  58505=>"111001100",
  58506=>"100111100",
  58507=>"111111001",
  58508=>"001000101",
  58509=>"100111111",
  58510=>"001101010",
  58511=>"010000000",
  58512=>"011010111",
  58513=>"000011001",
  58514=>"111101011",
  58515=>"010101101",
  58516=>"100011110",
  58517=>"000010110",
  58518=>"011101100",
  58519=>"010110000",
  58520=>"000110110",
  58521=>"010010001",
  58522=>"011011111",
  58523=>"010000010",
  58524=>"111010000",
  58525=>"010110010",
  58526=>"001111101",
  58527=>"001001001",
  58528=>"110011100",
  58529=>"001000101",
  58530=>"110100000",
  58531=>"011110100",
  58532=>"011011010",
  58533=>"110010001",
  58534=>"011111001",
  58535=>"101110010",
  58536=>"010100111",
  58537=>"010100110",
  58538=>"001011101",
  58539=>"011010100",
  58540=>"001011011",
  58541=>"000110000",
  58542=>"111001111",
  58543=>"011010011",
  58544=>"111101101",
  58545=>"110100010",
  58546=>"110010010",
  58547=>"001010101",
  58548=>"001011101",
  58549=>"001001001",
  58550=>"100111111",
  58551=>"001101100",
  58552=>"011111001",
  58553=>"110010110",
  58554=>"000101001",
  58555=>"111011010",
  58556=>"011011000",
  58557=>"111011000",
  58558=>"110011001",
  58559=>"101001101",
  58560=>"011011011",
  58561=>"011011101",
  58562=>"101101010",
  58563=>"101000001",
  58564=>"111011010",
  58565=>"110101111",
  58566=>"000001001",
  58567=>"000001110",
  58568=>"100111111",
  58569=>"100011101",
  58570=>"000010000",
  58571=>"011011000",
  58572=>"110100101",
  58573=>"010100001",
  58574=>"111011000",
  58575=>"110000001",
  58576=>"111111110",
  58577=>"011111100",
  58578=>"101011100",
  58579=>"100000010",
  58580=>"011011010",
  58581=>"110010011",
  58582=>"001100011",
  58583=>"001000010",
  58584=>"111110110",
  58585=>"101110100",
  58586=>"010110101",
  58587=>"100100110",
  58588=>"010000001",
  58589=>"000101111",
  58590=>"000101101",
  58591=>"101001011",
  58592=>"010000100",
  58593=>"001001000",
  58594=>"110010011",
  58595=>"111001101",
  58596=>"011101110",
  58597=>"101111000",
  58598=>"010001011",
  58599=>"111111001",
  58600=>"100101100",
  58601=>"001100110",
  58602=>"010101000",
  58603=>"100101101",
  58604=>"111110111",
  58605=>"110000001",
  58606=>"101101011",
  58607=>"001011011",
  58608=>"001101010",
  58609=>"000111101",
  58610=>"010011010",
  58611=>"110001000",
  58612=>"101001000",
  58613=>"010000001",
  58614=>"001001100",
  58615=>"100001010",
  58616=>"001111011",
  58617=>"110101001",
  58618=>"010001100",
  58619=>"111100011",
  58620=>"110101110",
  58621=>"000000011",
  58622=>"110101111",
  58623=>"100110110",
  58624=>"000100001",
  58625=>"000001101",
  58626=>"001000111",
  58627=>"001111110",
  58628=>"110101010",
  58629=>"101111110",
  58630=>"100100011",
  58631=>"100100001",
  58632=>"000101100",
  58633=>"111010111",
  58634=>"111110011",
  58635=>"110100110",
  58636=>"111001111",
  58637=>"011011100",
  58638=>"011001001",
  58639=>"111010111",
  58640=>"100001000",
  58641=>"101010110",
  58642=>"110101010",
  58643=>"111000001",
  58644=>"000011010",
  58645=>"011111100",
  58646=>"011100111",
  58647=>"111001111",
  58648=>"011001110",
  58649=>"101010001",
  58650=>"100110100",
  58651=>"111010000",
  58652=>"100000111",
  58653=>"100100110",
  58654=>"111000100",
  58655=>"110100111",
  58656=>"100111001",
  58657=>"101100001",
  58658=>"111100111",
  58659=>"010010110",
  58660=>"111001001",
  58661=>"100011000",
  58662=>"011011011",
  58663=>"001000111",
  58664=>"011010011",
  58665=>"111101110",
  58666=>"001111110",
  58667=>"010000011",
  58668=>"001010001",
  58669=>"111100000",
  58670=>"111000011",
  58671=>"011001101",
  58672=>"101101011",
  58673=>"111111001",
  58674=>"000010110",
  58675=>"111101010",
  58676=>"000000111",
  58677=>"110110010",
  58678=>"111111000",
  58679=>"111010010",
  58680=>"110111101",
  58681=>"001110110",
  58682=>"000000110",
  58683=>"101001000",
  58684=>"001010110",
  58685=>"010001011",
  58686=>"000001010",
  58687=>"001101101",
  58688=>"101011001",
  58689=>"001000110",
  58690=>"010111111",
  58691=>"011010111",
  58692=>"100001001",
  58693=>"000110000",
  58694=>"110010010",
  58695=>"110101110",
  58696=>"011101011",
  58697=>"101110000",
  58698=>"111001111",
  58699=>"011110010",
  58700=>"011111110",
  58701=>"110110101",
  58702=>"010101000",
  58703=>"001111000",
  58704=>"111101100",
  58705=>"101010000",
  58706=>"111001100",
  58707=>"100101101",
  58708=>"001010010",
  58709=>"010110101",
  58710=>"010111101",
  58711=>"110100100",
  58712=>"010110110",
  58713=>"010100111",
  58714=>"110111110",
  58715=>"100010111",
  58716=>"111110110",
  58717=>"011100111",
  58718=>"111101000",
  58719=>"111101011",
  58720=>"010110111",
  58721=>"101101001",
  58722=>"011000011",
  58723=>"110101011",
  58724=>"000111110",
  58725=>"001001110",
  58726=>"111100000",
  58727=>"100010110",
  58728=>"111001111",
  58729=>"100110011",
  58730=>"111010000",
  58731=>"110110110",
  58732=>"101010111",
  58733=>"001100000",
  58734=>"000010001",
  58735=>"000010000",
  58736=>"001000111",
  58737=>"001011010",
  58738=>"110100011",
  58739=>"000110110",
  58740=>"101010011",
  58741=>"001111111",
  58742=>"010100101",
  58743=>"110011101",
  58744=>"111110011",
  58745=>"101001000",
  58746=>"100000101",
  58747=>"100101010",
  58748=>"001010101",
  58749=>"001000100",
  58750=>"101111101",
  58751=>"001110111",
  58752=>"100000000",
  58753=>"001100010",
  58754=>"100110001",
  58755=>"101000011",
  58756=>"010100110",
  58757=>"110110000",
  58758=>"011001110",
  58759=>"011001001",
  58760=>"011011111",
  58761=>"011000000",
  58762=>"001011101",
  58763=>"011000010",
  58764=>"001001001",
  58765=>"010100101",
  58766=>"110001111",
  58767=>"010110001",
  58768=>"100011111",
  58769=>"100100100",
  58770=>"101100000",
  58771=>"001101011",
  58772=>"001100010",
  58773=>"110110001",
  58774=>"011010110",
  58775=>"101001101",
  58776=>"111100010",
  58777=>"110110010",
  58778=>"001001010",
  58779=>"111110101",
  58780=>"100001100",
  58781=>"001011011",
  58782=>"011110011",
  58783=>"011011011",
  58784=>"100110100",
  58785=>"000000101",
  58786=>"001100100",
  58787=>"001001000",
  58788=>"111001000",
  58789=>"000001110",
  58790=>"110100100",
  58791=>"010110011",
  58792=>"001101010",
  58793=>"101101101",
  58794=>"001111000",
  58795=>"010010001",
  58796=>"000001010",
  58797=>"000011010",
  58798=>"011101110",
  58799=>"011110100",
  58800=>"000011111",
  58801=>"010110001",
  58802=>"001101111",
  58803=>"100110100",
  58804=>"000111100",
  58805=>"001101101",
  58806=>"010111011",
  58807=>"111001010",
  58808=>"110010110",
  58809=>"100110111",
  58810=>"010100110",
  58811=>"110011011",
  58812=>"000100010",
  58813=>"110000101",
  58814=>"111011110",
  58815=>"010100101",
  58816=>"000100000",
  58817=>"001101101",
  58818=>"100110010",
  58819=>"000011110",
  58820=>"011001001",
  58821=>"000001000",
  58822=>"000111001",
  58823=>"010000110",
  58824=>"110101110",
  58825=>"011100011",
  58826=>"101001000",
  58827=>"001000111",
  58828=>"111011100",
  58829=>"100110100",
  58830=>"100111100",
  58831=>"100101100",
  58832=>"111101101",
  58833=>"010011010",
  58834=>"111111011",
  58835=>"101011100",
  58836=>"110110110",
  58837=>"111001001",
  58838=>"001000101",
  58839=>"010111101",
  58840=>"010011011",
  58841=>"000100100",
  58842=>"101111100",
  58843=>"100000000",
  58844=>"000010010",
  58845=>"101101101",
  58846=>"111110011",
  58847=>"101100101",
  58848=>"100101111",
  58849=>"100011011",
  58850=>"000011011",
  58851=>"001000010",
  58852=>"111101101",
  58853=>"110110101",
  58854=>"001011011",
  58855=>"111010010",
  58856=>"111110101",
  58857=>"101000011",
  58858=>"100110100",
  58859=>"000101011",
  58860=>"100000011",
  58861=>"110010111",
  58862=>"000010010",
  58863=>"100011001",
  58864=>"110000011",
  58865=>"001001110",
  58866=>"001000111",
  58867=>"100111101",
  58868=>"110111000",
  58869=>"001000011",
  58870=>"000001010",
  58871=>"100101110",
  58872=>"100101111",
  58873=>"000110000",
  58874=>"110110011",
  58875=>"111001100",
  58876=>"000000001",
  58877=>"000000011",
  58878=>"011011001",
  58879=>"010100001",
  58880=>"010001001",
  58881=>"000110110",
  58882=>"000010000",
  58883=>"111111100",
  58884=>"010110110",
  58885=>"001010011",
  58886=>"000101011",
  58887=>"001010000",
  58888=>"100111101",
  58889=>"000101111",
  58890=>"101101110",
  58891=>"011011111",
  58892=>"010010000",
  58893=>"010010001",
  58894=>"011110111",
  58895=>"110010101",
  58896=>"001011111",
  58897=>"011001001",
  58898=>"101111101",
  58899=>"010111101",
  58900=>"100001000",
  58901=>"011101111",
  58902=>"110001001",
  58903=>"010110011",
  58904=>"011011110",
  58905=>"110111111",
  58906=>"100111110",
  58907=>"111010000",
  58908=>"011010001",
  58909=>"001010010",
  58910=>"001100110",
  58911=>"101001000",
  58912=>"111001011",
  58913=>"010011001",
  58914=>"100000001",
  58915=>"101010011",
  58916=>"111001001",
  58917=>"000010100",
  58918=>"001101011",
  58919=>"001001101",
  58920=>"111100100",
  58921=>"111011100",
  58922=>"110111100",
  58923=>"111010000",
  58924=>"001100001",
  58925=>"000001111",
  58926=>"110100000",
  58927=>"111111011",
  58928=>"010011000",
  58929=>"011001101",
  58930=>"000101011",
  58931=>"000000110",
  58932=>"110110100",
  58933=>"111010001",
  58934=>"011111011",
  58935=>"101110010",
  58936=>"011101010",
  58937=>"011100010",
  58938=>"000011110",
  58939=>"111011100",
  58940=>"110010111",
  58941=>"000001000",
  58942=>"111010010",
  58943=>"110001111",
  58944=>"001111100",
  58945=>"010100110",
  58946=>"110111010",
  58947=>"001110111",
  58948=>"101100110",
  58949=>"001001100",
  58950=>"000110010",
  58951=>"001010011",
  58952=>"111101000",
  58953=>"110001000",
  58954=>"111100100",
  58955=>"000000010",
  58956=>"000000111",
  58957=>"010111111",
  58958=>"100001001",
  58959=>"011100110",
  58960=>"001111100",
  58961=>"101111010",
  58962=>"111101001",
  58963=>"010111110",
  58964=>"011111001",
  58965=>"010000110",
  58966=>"100100100",
  58967=>"111101111",
  58968=>"100001110",
  58969=>"000000011",
  58970=>"000110010",
  58971=>"110100111",
  58972=>"100001011",
  58973=>"000100111",
  58974=>"111010111",
  58975=>"101001001",
  58976=>"000100011",
  58977=>"101100010",
  58978=>"111100011",
  58979=>"010111011",
  58980=>"101101111",
  58981=>"101100111",
  58982=>"100100100",
  58983=>"011001001",
  58984=>"101111110",
  58985=>"001000111",
  58986=>"101000111",
  58987=>"110110000",
  58988=>"011010001",
  58989=>"010111111",
  58990=>"011011100",
  58991=>"000010011",
  58992=>"010101001",
  58993=>"101101010",
  58994=>"101000111",
  58995=>"111000111",
  58996=>"011010011",
  58997=>"010010101",
  58998=>"100111000",
  58999=>"101011001",
  59000=>"110011000",
  59001=>"010010010",
  59002=>"011011000",
  59003=>"011101000",
  59004=>"001110110",
  59005=>"101111010",
  59006=>"000010000",
  59007=>"111010101",
  59008=>"001110111",
  59009=>"001101010",
  59010=>"001101010",
  59011=>"111110111",
  59012=>"000111000",
  59013=>"011000000",
  59014=>"101110110",
  59015=>"011111010",
  59016=>"101111101",
  59017=>"101111101",
  59018=>"011111011",
  59019=>"111111100",
  59020=>"010100000",
  59021=>"001000111",
  59022=>"000011000",
  59023=>"000010101",
  59024=>"001101011",
  59025=>"011001011",
  59026=>"001001111",
  59027=>"011110011",
  59028=>"001010110",
  59029=>"101101010",
  59030=>"000111111",
  59031=>"100100101",
  59032=>"101010111",
  59033=>"101100011",
  59034=>"111001111",
  59035=>"100101100",
  59036=>"100010010",
  59037=>"010011010",
  59038=>"001100011",
  59039=>"111000011",
  59040=>"011111000",
  59041=>"110011111",
  59042=>"001110101",
  59043=>"111100010",
  59044=>"101011001",
  59045=>"010000011",
  59046=>"100010100",
  59047=>"100010010",
  59048=>"100010000",
  59049=>"000000010",
  59050=>"100000101",
  59051=>"001100001",
  59052=>"111010000",
  59053=>"001000100",
  59054=>"001000000",
  59055=>"001100100",
  59056=>"000101011",
  59057=>"110010001",
  59058=>"000100101",
  59059=>"101001011",
  59060=>"000101000",
  59061=>"101011001",
  59062=>"100100001",
  59063=>"110010110",
  59064=>"001111001",
  59065=>"000000000",
  59066=>"001000110",
  59067=>"100010110",
  59068=>"000101100",
  59069=>"011101101",
  59070=>"100100100",
  59071=>"100000111",
  59072=>"110001111",
  59073=>"000110000",
  59074=>"111011011",
  59075=>"100000001",
  59076=>"011111101",
  59077=>"000111011",
  59078=>"000110010",
  59079=>"000000001",
  59080=>"000100001",
  59081=>"101101011",
  59082=>"110101100",
  59083=>"000110101",
  59084=>"000000000",
  59085=>"101010101",
  59086=>"101100101",
  59087=>"000111111",
  59088=>"011110000",
  59089=>"000011010",
  59090=>"000001000",
  59091=>"100100001",
  59092=>"100000000",
  59093=>"000001110",
  59094=>"010001001",
  59095=>"111010011",
  59096=>"001101011",
  59097=>"101100111",
  59098=>"001010000",
  59099=>"001010000",
  59100=>"110110001",
  59101=>"000000010",
  59102=>"101110000",
  59103=>"011100110",
  59104=>"000110001",
  59105=>"001110000",
  59106=>"010001011",
  59107=>"001111111",
  59108=>"110000010",
  59109=>"001000100",
  59110=>"100110001",
  59111=>"000010010",
  59112=>"100010101",
  59113=>"011101001",
  59114=>"110010110",
  59115=>"000110111",
  59116=>"111101001",
  59117=>"000111100",
  59118=>"010010001",
  59119=>"011000001",
  59120=>"101100110",
  59121=>"011000100",
  59122=>"010101110",
  59123=>"000000110",
  59124=>"000110100",
  59125=>"101001101",
  59126=>"010001101",
  59127=>"001011101",
  59128=>"001101001",
  59129=>"101101111",
  59130=>"110110101",
  59131=>"001101110",
  59132=>"100000110",
  59133=>"011011010",
  59134=>"110101101",
  59135=>"011010101",
  59136=>"000000011",
  59137=>"000010101",
  59138=>"000010000",
  59139=>"000110001",
  59140=>"011011010",
  59141=>"111001111",
  59142=>"011100111",
  59143=>"010001100",
  59144=>"110010010",
  59145=>"011100110",
  59146=>"110110100",
  59147=>"101010110",
  59148=>"100010110",
  59149=>"001110110",
  59150=>"110000110",
  59151=>"001000101",
  59152=>"101101001",
  59153=>"111011010",
  59154=>"111101110",
  59155=>"110100001",
  59156=>"111011010",
  59157=>"000010000",
  59158=>"000101110",
  59159=>"000010000",
  59160=>"101101101",
  59161=>"001100111",
  59162=>"110111110",
  59163=>"000011010",
  59164=>"101111000",
  59165=>"110000010",
  59166=>"010110000",
  59167=>"100000010",
  59168=>"100000001",
  59169=>"101000000",
  59170=>"100111111",
  59171=>"001000100",
  59172=>"100000000",
  59173=>"010110111",
  59174=>"110011100",
  59175=>"111010001",
  59176=>"100010001",
  59177=>"010101111",
  59178=>"011111110",
  59179=>"010111110",
  59180=>"110100011",
  59181=>"100100001",
  59182=>"101100000",
  59183=>"100001111",
  59184=>"110110000",
  59185=>"001101001",
  59186=>"100101000",
  59187=>"001100110",
  59188=>"111011111",
  59189=>"101000010",
  59190=>"010011011",
  59191=>"100110010",
  59192=>"110111111",
  59193=>"010101000",
  59194=>"000010100",
  59195=>"000000110",
  59196=>"110101100",
  59197=>"001010100",
  59198=>"001100110",
  59199=>"001101110",
  59200=>"101101001",
  59201=>"011001000",
  59202=>"000001001",
  59203=>"110100110",
  59204=>"000110101",
  59205=>"010111101",
  59206=>"000011111",
  59207=>"101110011",
  59208=>"000011100",
  59209=>"010000000",
  59210=>"111111111",
  59211=>"010000001",
  59212=>"001001000",
  59213=>"111100100",
  59214=>"110000000",
  59215=>"101001000",
  59216=>"010010111",
  59217=>"000011110",
  59218=>"001111011",
  59219=>"011111000",
  59220=>"110110100",
  59221=>"110110011",
  59222=>"111000000",
  59223=>"001101111",
  59224=>"011001001",
  59225=>"110010111",
  59226=>"010101110",
  59227=>"011111011",
  59228=>"101101111",
  59229=>"100000100",
  59230=>"111011011",
  59231=>"010010110",
  59232=>"111100100",
  59233=>"001110000",
  59234=>"100010010",
  59235=>"100110011",
  59236=>"100010110",
  59237=>"010011001",
  59238=>"010100010",
  59239=>"111000100",
  59240=>"001001101",
  59241=>"010001110",
  59242=>"010000000",
  59243=>"001101100",
  59244=>"010000110",
  59245=>"100101111",
  59246=>"100010000",
  59247=>"011001110",
  59248=>"110011000",
  59249=>"111100011",
  59250=>"010111011",
  59251=>"101000001",
  59252=>"100100101",
  59253=>"101111100",
  59254=>"100001101",
  59255=>"001100011",
  59256=>"111111000",
  59257=>"101000110",
  59258=>"000011011",
  59259=>"001101000",
  59260=>"000011011",
  59261=>"000001110",
  59262=>"010000001",
  59263=>"111010001",
  59264=>"100101111",
  59265=>"100010000",
  59266=>"110111100",
  59267=>"110101011",
  59268=>"011100000",
  59269=>"010100010",
  59270=>"110001110",
  59271=>"000001111",
  59272=>"111100111",
  59273=>"111110010",
  59274=>"110110100",
  59275=>"001001001",
  59276=>"100100000",
  59277=>"000111111",
  59278=>"101101110",
  59279=>"100010010",
  59280=>"011001010",
  59281=>"001100101",
  59282=>"010110100",
  59283=>"001011100",
  59284=>"111110111",
  59285=>"011111100",
  59286=>"001111110",
  59287=>"110111110",
  59288=>"110111010",
  59289=>"000001110",
  59290=>"000011000",
  59291=>"010110000",
  59292=>"100000110",
  59293=>"010101110",
  59294=>"111111010",
  59295=>"010011011",
  59296=>"000100100",
  59297=>"000111100",
  59298=>"010110001",
  59299=>"000110100",
  59300=>"100110110",
  59301=>"011100100",
  59302=>"101011100",
  59303=>"001000111",
  59304=>"011000110",
  59305=>"011111101",
  59306=>"101110100",
  59307=>"110111011",
  59308=>"111110011",
  59309=>"011101100",
  59310=>"010110101",
  59311=>"111100000",
  59312=>"010111110",
  59313=>"110100011",
  59314=>"010000000",
  59315=>"100010010",
  59316=>"010011010",
  59317=>"101110001",
  59318=>"011000111",
  59319=>"001011001",
  59320=>"010011001",
  59321=>"100110000",
  59322=>"110111000",
  59323=>"000100011",
  59324=>"010101000",
  59325=>"010010100",
  59326=>"011111010",
  59327=>"011100011",
  59328=>"110010111",
  59329=>"000110011",
  59330=>"110110110",
  59331=>"000011001",
  59332=>"001000110",
  59333=>"101110010",
  59334=>"110010010",
  59335=>"111100001",
  59336=>"100010110",
  59337=>"010101100",
  59338=>"111001101",
  59339=>"110100000",
  59340=>"100001110",
  59341=>"010110010",
  59342=>"000100011",
  59343=>"010111111",
  59344=>"111111010",
  59345=>"000101001",
  59346=>"100110101",
  59347=>"001010111",
  59348=>"111110100",
  59349=>"101111101",
  59350=>"101100100",
  59351=>"100001011",
  59352=>"010100101",
  59353=>"010100101",
  59354=>"001000110",
  59355=>"011110111",
  59356=>"101110111",
  59357=>"001110110",
  59358=>"000000111",
  59359=>"101010011",
  59360=>"101010101",
  59361=>"001100011",
  59362=>"001000110",
  59363=>"011100011",
  59364=>"000000100",
  59365=>"001000010",
  59366=>"010110001",
  59367=>"110000101",
  59368=>"001000001",
  59369=>"100010100",
  59370=>"110100011",
  59371=>"111111100",
  59372=>"110111010",
  59373=>"101110101",
  59374=>"001100110",
  59375=>"000010101",
  59376=>"000100101",
  59377=>"010011101",
  59378=>"000110101",
  59379=>"010000100",
  59380=>"010110011",
  59381=>"110001011",
  59382=>"001011111",
  59383=>"111110110",
  59384=>"010001000",
  59385=>"011100000",
  59386=>"110001011",
  59387=>"110101010",
  59388=>"101111111",
  59389=>"100011100",
  59390=>"100100101",
  59391=>"000100001",
  59392=>"101100000",
  59393=>"101100100",
  59394=>"100010101",
  59395=>"111111111",
  59396=>"110010111",
  59397=>"100110000",
  59398=>"001001011",
  59399=>"010110011",
  59400=>"110101100",
  59401=>"111100000",
  59402=>"110111110",
  59403=>"111010111",
  59404=>"010010001",
  59405=>"000011001",
  59406=>"110100011",
  59407=>"100101010",
  59408=>"000001010",
  59409=>"000100110",
  59410=>"010111000",
  59411=>"100100101",
  59412=>"011011001",
  59413=>"001100100",
  59414=>"100110001",
  59415=>"000000110",
  59416=>"111010101",
  59417=>"000011110",
  59418=>"000111011",
  59419=>"111001010",
  59420=>"111111101",
  59421=>"101100001",
  59422=>"001000101",
  59423=>"001110001",
  59424=>"000010011",
  59425=>"000101111",
  59426=>"010111010",
  59427=>"001001110",
  59428=>"000000001",
  59429=>"010001011",
  59430=>"000010111",
  59431=>"011111000",
  59432=>"101011111",
  59433=>"101011111",
  59434=>"110100100",
  59435=>"100001111",
  59436=>"100101000",
  59437=>"010111010",
  59438=>"000011011",
  59439=>"010101011",
  59440=>"100101101",
  59441=>"100111111",
  59442=>"101000011",
  59443=>"011101100",
  59444=>"110000101",
  59445=>"111101001",
  59446=>"100000101",
  59447=>"100110001",
  59448=>"000011111",
  59449=>"011100010",
  59450=>"110101100",
  59451=>"101011010",
  59452=>"101001000",
  59453=>"110101010",
  59454=>"110101110",
  59455=>"000111111",
  59456=>"100111111",
  59457=>"111101100",
  59458=>"110000101",
  59459=>"001010011",
  59460=>"111100100",
  59461=>"010000001",
  59462=>"111100101",
  59463=>"100110000",
  59464=>"101101011",
  59465=>"100000010",
  59466=>"010001101",
  59467=>"010100101",
  59468=>"010000111",
  59469=>"000100011",
  59470=>"110011000",
  59471=>"100000011",
  59472=>"100011101",
  59473=>"100110101",
  59474=>"100100001",
  59475=>"001100101",
  59476=>"111111011",
  59477=>"011000100",
  59478=>"011111110",
  59479=>"110110110",
  59480=>"011100101",
  59481=>"111001110",
  59482=>"011101101",
  59483=>"000011101",
  59484=>"010100110",
  59485=>"000110011",
  59486=>"100001100",
  59487=>"000000111",
  59488=>"000000011",
  59489=>"001100010",
  59490=>"001110001",
  59491=>"010001010",
  59492=>"100000010",
  59493=>"001101011",
  59494=>"011011001",
  59495=>"101011000",
  59496=>"101101111",
  59497=>"101010111",
  59498=>"000000000",
  59499=>"010001101",
  59500=>"111100011",
  59501=>"100100101",
  59502=>"011010111",
  59503=>"011000001",
  59504=>"010110001",
  59505=>"100001010",
  59506=>"110010000",
  59507=>"010111010",
  59508=>"111011000",
  59509=>"001010000",
  59510=>"100010001",
  59511=>"011100000",
  59512=>"110111101",
  59513=>"101001001",
  59514=>"110011011",
  59515=>"110111001",
  59516=>"101010101",
  59517=>"100000000",
  59518=>"011100001",
  59519=>"000110100",
  59520=>"001101010",
  59521=>"001000101",
  59522=>"000101001",
  59523=>"001001001",
  59524=>"010010001",
  59525=>"000100011",
  59526=>"100111111",
  59527=>"001010100",
  59528=>"001111111",
  59529=>"011011001",
  59530=>"100010000",
  59531=>"100011110",
  59532=>"001110010",
  59533=>"001110101",
  59534=>"011111010",
  59535=>"101001110",
  59536=>"100001011",
  59537=>"000010011",
  59538=>"110000011",
  59539=>"101001001",
  59540=>"001110010",
  59541=>"101110001",
  59542=>"101011011",
  59543=>"000111111",
  59544=>"101101111",
  59545=>"111111001",
  59546=>"001001101",
  59547=>"111011101",
  59548=>"011001100",
  59549=>"010011101",
  59550=>"110000111",
  59551=>"010001000",
  59552=>"111101001",
  59553=>"111101010",
  59554=>"011010001",
  59555=>"000100100",
  59556=>"001100100",
  59557=>"000011101",
  59558=>"000011011",
  59559=>"111100101",
  59560=>"011010110",
  59561=>"010101011",
  59562=>"000010110",
  59563=>"000110101",
  59564=>"010110100",
  59565=>"000000101",
  59566=>"001110111",
  59567=>"110111001",
  59568=>"001110101",
  59569=>"110101011",
  59570=>"100101101",
  59571=>"100010001",
  59572=>"111011110",
  59573=>"101010010",
  59574=>"100101100",
  59575=>"110100110",
  59576=>"011011001",
  59577=>"000101011",
  59578=>"010011100",
  59579=>"101111110",
  59580=>"010001000",
  59581=>"010011010",
  59582=>"001101001",
  59583=>"110011110",
  59584=>"100111111",
  59585=>"100011000",
  59586=>"110111110",
  59587=>"000000000",
  59588=>"011110010",
  59589=>"010011101",
  59590=>"110001100",
  59591=>"100010101",
  59592=>"011011110",
  59593=>"000100110",
  59594=>"101001001",
  59595=>"001000011",
  59596=>"001111000",
  59597=>"001111101",
  59598=>"101011100",
  59599=>"101111010",
  59600=>"110110000",
  59601=>"001001001",
  59602=>"000010110",
  59603=>"011010110",
  59604=>"001000010",
  59605=>"000101000",
  59606=>"011101001",
  59607=>"100101001",
  59608=>"000000000",
  59609=>"001010010",
  59610=>"111001100",
  59611=>"010000111",
  59612=>"000010010",
  59613=>"011111000",
  59614=>"011000011",
  59615=>"110110101",
  59616=>"001000100",
  59617=>"000101011",
  59618=>"110111100",
  59619=>"010011100",
  59620=>"001011001",
  59621=>"100000111",
  59622=>"110100000",
  59623=>"010001110",
  59624=>"001110001",
  59625=>"010010010",
  59626=>"110100011",
  59627=>"100110110",
  59628=>"011101100",
  59629=>"111001111",
  59630=>"110000010",
  59631=>"100100010",
  59632=>"010011110",
  59633=>"101001010",
  59634=>"010000101",
  59635=>"111111010",
  59636=>"010001011",
  59637=>"110001000",
  59638=>"100111111",
  59639=>"001100111",
  59640=>"010110010",
  59641=>"001011011",
  59642=>"000101101",
  59643=>"010100000",
  59644=>"001101000",
  59645=>"010001111",
  59646=>"001001100",
  59647=>"100001000",
  59648=>"101111111",
  59649=>"001110111",
  59650=>"010011101",
  59651=>"000101100",
  59652=>"111110010",
  59653=>"111000000",
  59654=>"100000001",
  59655=>"101111100",
  59656=>"000011010",
  59657=>"110010100",
  59658=>"111101001",
  59659=>"101000111",
  59660=>"010010110",
  59661=>"011100010",
  59662=>"011011111",
  59663=>"000100010",
  59664=>"110011110",
  59665=>"010100001",
  59666=>"100100001",
  59667=>"110010010",
  59668=>"010011111",
  59669=>"110100001",
  59670=>"110000001",
  59671=>"111111001",
  59672=>"111111100",
  59673=>"111000111",
  59674=>"110101110",
  59675=>"100000111",
  59676=>"111110000",
  59677=>"111000000",
  59678=>"011001111",
  59679=>"101111011",
  59680=>"001110101",
  59681=>"010111010",
  59682=>"011111000",
  59683=>"011001101",
  59684=>"001100101",
  59685=>"011011010",
  59686=>"110000001",
  59687=>"101111100",
  59688=>"010000000",
  59689=>"101001110",
  59690=>"110001010",
  59691=>"001110000",
  59692=>"001100101",
  59693=>"100100001",
  59694=>"111010001",
  59695=>"100001110",
  59696=>"011101100",
  59697=>"100010011",
  59698=>"110000110",
  59699=>"000001000",
  59700=>"000010100",
  59701=>"100111100",
  59702=>"111000001",
  59703=>"011010001",
  59704=>"111000100",
  59705=>"101100100",
  59706=>"111110110",
  59707=>"101000011",
  59708=>"100010100",
  59709=>"101100011",
  59710=>"001101000",
  59711=>"010001000",
  59712=>"101010111",
  59713=>"110101101",
  59714=>"000011101",
  59715=>"110110110",
  59716=>"001100001",
  59717=>"111001111",
  59718=>"110001000",
  59719=>"111100010",
  59720=>"101010000",
  59721=>"001111111",
  59722=>"101101110",
  59723=>"100000111",
  59724=>"110110111",
  59725=>"111110000",
  59726=>"001110110",
  59727=>"100101001",
  59728=>"101110001",
  59729=>"000110111",
  59730=>"101000010",
  59731=>"000010101",
  59732=>"010111001",
  59733=>"010010011",
  59734=>"001111110",
  59735=>"001000000",
  59736=>"101111110",
  59737=>"011000111",
  59738=>"111100001",
  59739=>"111010001",
  59740=>"111111101",
  59741=>"101110110",
  59742=>"111001011",
  59743=>"101111101",
  59744=>"010010110",
  59745=>"011101111",
  59746=>"001101110",
  59747=>"001001011",
  59748=>"001110111",
  59749=>"000000000",
  59750=>"000101000",
  59751=>"111000100",
  59752=>"011100111",
  59753=>"010010011",
  59754=>"101000101",
  59755=>"101001111",
  59756=>"110000000",
  59757=>"010111101",
  59758=>"010110011",
  59759=>"010110010",
  59760=>"001101100",
  59761=>"010000010",
  59762=>"110101100",
  59763=>"010101011",
  59764=>"101011111",
  59765=>"101010001",
  59766=>"001000111",
  59767=>"001000001",
  59768=>"000110001",
  59769=>"000000011",
  59770=>"101011011",
  59771=>"000111111",
  59772=>"111110111",
  59773=>"010000110",
  59774=>"010010010",
  59775=>"101111000",
  59776=>"001111010",
  59777=>"001110000",
  59778=>"100100110",
  59779=>"001010011",
  59780=>"111100110",
  59781=>"000110000",
  59782=>"010011010",
  59783=>"011110000",
  59784=>"110100000",
  59785=>"001100010",
  59786=>"100100101",
  59787=>"110010010",
  59788=>"010101000",
  59789=>"100100101",
  59790=>"101101111",
  59791=>"110010110",
  59792=>"011110110",
  59793=>"110001100",
  59794=>"111000010",
  59795=>"001111011",
  59796=>"000011111",
  59797=>"001000110",
  59798=>"001110011",
  59799=>"001101001",
  59800=>"011010011",
  59801=>"001001111",
  59802=>"100100001",
  59803=>"011011010",
  59804=>"110111000",
  59805=>"001000001",
  59806=>"101111110",
  59807=>"100000111",
  59808=>"100100111",
  59809=>"111000111",
  59810=>"011010010",
  59811=>"110000001",
  59812=>"010111111",
  59813=>"111110001",
  59814=>"111100001",
  59815=>"111001010",
  59816=>"000000101",
  59817=>"100101000",
  59818=>"100110110",
  59819=>"000111110",
  59820=>"000101001",
  59821=>"010000001",
  59822=>"111000101",
  59823=>"100101000",
  59824=>"100101100",
  59825=>"011111101",
  59826=>"100110000",
  59827=>"100000101",
  59828=>"101101111",
  59829=>"010010001",
  59830=>"000001100",
  59831=>"111001010",
  59832=>"001110111",
  59833=>"100111101",
  59834=>"100001111",
  59835=>"011000111",
  59836=>"111111000",
  59837=>"101000100",
  59838=>"000010000",
  59839=>"100101011",
  59840=>"010101111",
  59841=>"000011010",
  59842=>"010110100",
  59843=>"110010011",
  59844=>"111100010",
  59845=>"111001000",
  59846=>"000111001",
  59847=>"111000001",
  59848=>"110000000",
  59849=>"101010101",
  59850=>"110101100",
  59851=>"010111000",
  59852=>"000000010",
  59853=>"101010000",
  59854=>"111010010",
  59855=>"010001110",
  59856=>"011000111",
  59857=>"000001001",
  59858=>"010100000",
  59859=>"111011000",
  59860=>"011110100",
  59861=>"110000110",
  59862=>"110010110",
  59863=>"110100100",
  59864=>"100110000",
  59865=>"010110011",
  59866=>"011101101",
  59867=>"001011111",
  59868=>"001011100",
  59869=>"100111100",
  59870=>"101111011",
  59871=>"010000011",
  59872=>"100001001",
  59873=>"000111010",
  59874=>"101011011",
  59875=>"001010101",
  59876=>"000110101",
  59877=>"001000010",
  59878=>"010000100",
  59879=>"110111110",
  59880=>"001011101",
  59881=>"000000001",
  59882=>"011010011",
  59883=>"010111011",
  59884=>"110111101",
  59885=>"100010000",
  59886=>"111000010",
  59887=>"011101011",
  59888=>"111100101",
  59889=>"001001111",
  59890=>"010000011",
  59891=>"011101101",
  59892=>"110011001",
  59893=>"010100000",
  59894=>"110010110",
  59895=>"100110100",
  59896=>"100110000",
  59897=>"111001001",
  59898=>"000110001",
  59899=>"100111010",
  59900=>"001000001",
  59901=>"110011010",
  59902=>"101101111",
  59903=>"100001011",
  59904=>"101111101",
  59905=>"110001101",
  59906=>"101011000",
  59907=>"110100101",
  59908=>"000011110",
  59909=>"110000001",
  59910=>"010001000",
  59911=>"110110100",
  59912=>"000011111",
  59913=>"110101010",
  59914=>"100111011",
  59915=>"101000010",
  59916=>"101100001",
  59917=>"101001000",
  59918=>"010100100",
  59919=>"001000001",
  59920=>"100110111",
  59921=>"101100100",
  59922=>"001000011",
  59923=>"011101111",
  59924=>"011100110",
  59925=>"111110010",
  59926=>"010001000",
  59927=>"010101100",
  59928=>"101000011",
  59929=>"011111111",
  59930=>"100000111",
  59931=>"110100110",
  59932=>"011100100",
  59933=>"010100000",
  59934=>"100101110",
  59935=>"110110010",
  59936=>"111010001",
  59937=>"001101111",
  59938=>"011100000",
  59939=>"011010011",
  59940=>"001010100",
  59941=>"011001111",
  59942=>"001011001",
  59943=>"000011010",
  59944=>"110100000",
  59945=>"101110101",
  59946=>"001101010",
  59947=>"010001001",
  59948=>"110001100",
  59949=>"010100101",
  59950=>"011111111",
  59951=>"101100101",
  59952=>"001001011",
  59953=>"110111011",
  59954=>"111000010",
  59955=>"010101111",
  59956=>"011000101",
  59957=>"111000110",
  59958=>"100010110",
  59959=>"001111001",
  59960=>"111000100",
  59961=>"000101100",
  59962=>"000101011",
  59963=>"000100011",
  59964=>"010100111",
  59965=>"100110000",
  59966=>"010110001",
  59967=>"111111101",
  59968=>"001110100",
  59969=>"010110100",
  59970=>"011010101",
  59971=>"111010011",
  59972=>"010011110",
  59973=>"100110111",
  59974=>"000100110",
  59975=>"111000100",
  59976=>"010110110",
  59977=>"101101101",
  59978=>"011010100",
  59979=>"011001110",
  59980=>"010111111",
  59981=>"001101100",
  59982=>"001111001",
  59983=>"010110011",
  59984=>"110111011",
  59985=>"000000011",
  59986=>"111010110",
  59987=>"011010000",
  59988=>"111110001",
  59989=>"000010101",
  59990=>"010010011",
  59991=>"100001001",
  59992=>"001110010",
  59993=>"110010100",
  59994=>"110110110",
  59995=>"110001000",
  59996=>"110100000",
  59997=>"001000000",
  59998=>"000001110",
  59999=>"110010000",
  60000=>"111011000",
  60001=>"001100101",
  60002=>"100110011",
  60003=>"000011001",
  60004=>"101000000",
  60005=>"101010011",
  60006=>"111001111",
  60007=>"111011010",
  60008=>"101111001",
  60009=>"010000111",
  60010=>"100010101",
  60011=>"101101111",
  60012=>"010000111",
  60013=>"000111000",
  60014=>"011000101",
  60015=>"100010010",
  60016=>"001100001",
  60017=>"001111110",
  60018=>"110001000",
  60019=>"110001110",
  60020=>"100111110",
  60021=>"100101110",
  60022=>"101110010",
  60023=>"110110011",
  60024=>"110001001",
  60025=>"000000110",
  60026=>"011111110",
  60027=>"110010001",
  60028=>"100010101",
  60029=>"100100101",
  60030=>"110110101",
  60031=>"001110110",
  60032=>"100100100",
  60033=>"011101100",
  60034=>"111111011",
  60035=>"110100110",
  60036=>"010010010",
  60037=>"111000101",
  60038=>"011010000",
  60039=>"000000110",
  60040=>"101000101",
  60041=>"010000001",
  60042=>"000110101",
  60043=>"011010110",
  60044=>"010100010",
  60045=>"011100111",
  60046=>"011011010",
  60047=>"010010111",
  60048=>"000100010",
  60049=>"011101100",
  60050=>"010110011",
  60051=>"001111010",
  60052=>"001001001",
  60053=>"110001101",
  60054=>"100101100",
  60055=>"100100110",
  60056=>"000000011",
  60057=>"111001100",
  60058=>"010000011",
  60059=>"001011110",
  60060=>"011110110",
  60061=>"101110011",
  60062=>"101110010",
  60063=>"011011100",
  60064=>"100011100",
  60065=>"011010110",
  60066=>"011010001",
  60067=>"100000001",
  60068=>"000011010",
  60069=>"000011001",
  60070=>"100100000",
  60071=>"011010001",
  60072=>"011110000",
  60073=>"110110101",
  60074=>"001111000",
  60075=>"111100000",
  60076=>"000100111",
  60077=>"010100100",
  60078=>"100010111",
  60079=>"011010100",
  60080=>"110100100",
  60081=>"001110000",
  60082=>"111001000",
  60083=>"010111100",
  60084=>"000010000",
  60085=>"010000010",
  60086=>"110100111",
  60087=>"110111000",
  60088=>"001110101",
  60089=>"000011101",
  60090=>"001110000",
  60091=>"100010100",
  60092=>"000101110",
  60093=>"111011110",
  60094=>"011010000",
  60095=>"001000101",
  60096=>"010100110",
  60097=>"011111101",
  60098=>"111010101",
  60099=>"001111010",
  60100=>"001100001",
  60101=>"011111110",
  60102=>"011110100",
  60103=>"011000010",
  60104=>"111010101",
  60105=>"000100101",
  60106=>"000011001",
  60107=>"001011001",
  60108=>"011100001",
  60109=>"001000010",
  60110=>"110101011",
  60111=>"011111111",
  60112=>"110100001",
  60113=>"111101011",
  60114=>"100001101",
  60115=>"110000101",
  60116=>"010100001",
  60117=>"001101110",
  60118=>"110100010",
  60119=>"000000001",
  60120=>"000011010",
  60121=>"010110001",
  60122=>"010110101",
  60123=>"010101011",
  60124=>"100001110",
  60125=>"101000010",
  60126=>"000110111",
  60127=>"110100111",
  60128=>"111100011",
  60129=>"100101001",
  60130=>"100001110",
  60131=>"111110111",
  60132=>"001000010",
  60133=>"111011101",
  60134=>"010000110",
  60135=>"000011011",
  60136=>"001001100",
  60137=>"011010100",
  60138=>"000111011",
  60139=>"111000011",
  60140=>"001100010",
  60141=>"000111010",
  60142=>"000100110",
  60143=>"101000111",
  60144=>"010110100",
  60145=>"101100000",
  60146=>"010000011",
  60147=>"011010101",
  60148=>"000011111",
  60149=>"111011100",
  60150=>"111100110",
  60151=>"011011010",
  60152=>"101100000",
  60153=>"011011010",
  60154=>"101000111",
  60155=>"010100001",
  60156=>"011111101",
  60157=>"010001110",
  60158=>"001110101",
  60159=>"000101100",
  60160=>"110010101",
  60161=>"100101011",
  60162=>"110011111",
  60163=>"011000011",
  60164=>"011000011",
  60165=>"011000010",
  60166=>"000001110",
  60167=>"000001110",
  60168=>"011101000",
  60169=>"110110011",
  60170=>"111001010",
  60171=>"111110100",
  60172=>"111100000",
  60173=>"101001101",
  60174=>"100101000",
  60175=>"101111011",
  60176=>"010100000",
  60177=>"101001111",
  60178=>"101001101",
  60179=>"110010111",
  60180=>"111001111",
  60181=>"010001001",
  60182=>"100101001",
  60183=>"000101100",
  60184=>"110101000",
  60185=>"100101111",
  60186=>"000000001",
  60187=>"011001000",
  60188=>"000000111",
  60189=>"111101010",
  60190=>"110010010",
  60191=>"000011110",
  60192=>"010111000",
  60193=>"000000001",
  60194=>"111010111",
  60195=>"011000111",
  60196=>"000101000",
  60197=>"000000100",
  60198=>"110000010",
  60199=>"001011110",
  60200=>"010111101",
  60201=>"110111101",
  60202=>"111101011",
  60203=>"000011001",
  60204=>"001011001",
  60205=>"001100001",
  60206=>"010110100",
  60207=>"000010100",
  60208=>"000000010",
  60209=>"111001111",
  60210=>"011100000",
  60211=>"000011110",
  60212=>"011011000",
  60213=>"111101001",
  60214=>"100001011",
  60215=>"011011000",
  60216=>"110111101",
  60217=>"000001011",
  60218=>"001101101",
  60219=>"111001011",
  60220=>"001000101",
  60221=>"010000110",
  60222=>"101000000",
  60223=>"011110101",
  60224=>"010010000",
  60225=>"111010110",
  60226=>"000110100",
  60227=>"100011011",
  60228=>"101111000",
  60229=>"110110100",
  60230=>"110100100",
  60231=>"110100110",
  60232=>"000101001",
  60233=>"010101100",
  60234=>"010010001",
  60235=>"110101100",
  60236=>"000001010",
  60237=>"010010101",
  60238=>"010100011",
  60239=>"011000110",
  60240=>"010001011",
  60241=>"001000011",
  60242=>"101000110",
  60243=>"001001011",
  60244=>"110001001",
  60245=>"110000101",
  60246=>"000000011",
  60247=>"111111001",
  60248=>"011100101",
  60249=>"000001111",
  60250=>"110000100",
  60251=>"100001000",
  60252=>"100101100",
  60253=>"000001110",
  60254=>"111110001",
  60255=>"000000101",
  60256=>"100110110",
  60257=>"110001100",
  60258=>"000101010",
  60259=>"000011110",
  60260=>"110000011",
  60261=>"011000001",
  60262=>"010111011",
  60263=>"110001000",
  60264=>"111010000",
  60265=>"010101011",
  60266=>"011110110",
  60267=>"110001101",
  60268=>"000001001",
  60269=>"011111000",
  60270=>"101110010",
  60271=>"010001001",
  60272=>"010001101",
  60273=>"011000100",
  60274=>"000010010",
  60275=>"000010110",
  60276=>"000010000",
  60277=>"000011101",
  60278=>"001111000",
  60279=>"010101101",
  60280=>"101000111",
  60281=>"100011000",
  60282=>"000111000",
  60283=>"000110100",
  60284=>"010010101",
  60285=>"100100010",
  60286=>"000000000",
  60287=>"110010011",
  60288=>"111110000",
  60289=>"100110011",
  60290=>"001010101",
  60291=>"100011000",
  60292=>"010111111",
  60293=>"001011101",
  60294=>"011000010",
  60295=>"000001100",
  60296=>"111000101",
  60297=>"001001100",
  60298=>"101100010",
  60299=>"010100010",
  60300=>"101111110",
  60301=>"111110110",
  60302=>"111000011",
  60303=>"101001101",
  60304=>"111111000",
  60305=>"000010010",
  60306=>"100111011",
  60307=>"000011100",
  60308=>"000110101",
  60309=>"101101001",
  60310=>"110110111",
  60311=>"101010001",
  60312=>"101010011",
  60313=>"101100100",
  60314=>"101110101",
  60315=>"100000011",
  60316=>"110111100",
  60317=>"001001111",
  60318=>"110101001",
  60319=>"110001101",
  60320=>"111100000",
  60321=>"001111010",
  60322=>"111010111",
  60323=>"011101111",
  60324=>"111001001",
  60325=>"001111001",
  60326=>"010100100",
  60327=>"011111111",
  60328=>"101000011",
  60329=>"101001101",
  60330=>"110110111",
  60331=>"111101101",
  60332=>"111100001",
  60333=>"001101001",
  60334=>"010011101",
  60335=>"000111001",
  60336=>"110011010",
  60337=>"010001101",
  60338=>"001111011",
  60339=>"110101111",
  60340=>"111101001",
  60341=>"011110111",
  60342=>"010011111",
  60343=>"011000101",
  60344=>"100001011",
  60345=>"001000000",
  60346=>"011100101",
  60347=>"001110000",
  60348=>"110101001",
  60349=>"111011101",
  60350=>"010111111",
  60351=>"111010010",
  60352=>"010011000",
  60353=>"001010000",
  60354=>"111001010",
  60355=>"101111110",
  60356=>"000000011",
  60357=>"010010001",
  60358=>"111111010",
  60359=>"011010001",
  60360=>"100010101",
  60361=>"010011111",
  60362=>"000100010",
  60363=>"110111100",
  60364=>"110101111",
  60365=>"100000100",
  60366=>"001101010",
  60367=>"111110111",
  60368=>"101000111",
  60369=>"100110110",
  60370=>"111000110",
  60371=>"111110101",
  60372=>"000010010",
  60373=>"100001000",
  60374=>"000101011",
  60375=>"100010100",
  60376=>"111000010",
  60377=>"011001011",
  60378=>"111111000",
  60379=>"011110000",
  60380=>"000010100",
  60381=>"110110100",
  60382=>"001111110",
  60383=>"110011000",
  60384=>"000100100",
  60385=>"000001011",
  60386=>"100110000",
  60387=>"110001011",
  60388=>"000000011",
  60389=>"110000111",
  60390=>"000010001",
  60391=>"011110110",
  60392=>"011101111",
  60393=>"101101101",
  60394=>"110101100",
  60395=>"100001010",
  60396=>"100101010",
  60397=>"110110111",
  60398=>"001000100",
  60399=>"101010000",
  60400=>"011000000",
  60401=>"111000110",
  60402=>"000110100",
  60403=>"101101101",
  60404=>"010001011",
  60405=>"000010100",
  60406=>"001110010",
  60407=>"010001010",
  60408=>"010000110",
  60409=>"101101111",
  60410=>"000001001",
  60411=>"110010000",
  60412=>"011111001",
  60413=>"110001000",
  60414=>"001000101",
  60415=>"101111001",
  60416=>"010111000",
  60417=>"000011101",
  60418=>"011010110",
  60419=>"101101101",
  60420=>"111110010",
  60421=>"100010010",
  60422=>"110000111",
  60423=>"111000110",
  60424=>"101011101",
  60425=>"111011011",
  60426=>"111000100",
  60427=>"110110101",
  60428=>"010111111",
  60429=>"010011001",
  60430=>"100100001",
  60431=>"100001000",
  60432=>"011111110",
  60433=>"010001000",
  60434=>"000000001",
  60435=>"100010100",
  60436=>"000001011",
  60437=>"000000111",
  60438=>"101000100",
  60439=>"100100011",
  60440=>"101111101",
  60441=>"111001110",
  60442=>"110110010",
  60443=>"001000111",
  60444=>"000011100",
  60445=>"110101100",
  60446=>"001011111",
  60447=>"000000000",
  60448=>"101011001",
  60449=>"001100101",
  60450=>"000100011",
  60451=>"111000011",
  60452=>"000011001",
  60453=>"000000000",
  60454=>"110000110",
  60455=>"011001011",
  60456=>"011001000",
  60457=>"010000011",
  60458=>"101110010",
  60459=>"101111110",
  60460=>"110000101",
  60461=>"001100011",
  60462=>"101111101",
  60463=>"000010111",
  60464=>"110111110",
  60465=>"100110011",
  60466=>"010101000",
  60467=>"000100111",
  60468=>"111000011",
  60469=>"000000010",
  60470=>"111101011",
  60471=>"001010001",
  60472=>"000000111",
  60473=>"100000010",
  60474=>"100100000",
  60475=>"000111101",
  60476=>"011001111",
  60477=>"111110010",
  60478=>"110001101",
  60479=>"001010101",
  60480=>"111110000",
  60481=>"000001010",
  60482=>"100111101",
  60483=>"101111100",
  60484=>"010001101",
  60485=>"000101111",
  60486=>"101001000",
  60487=>"111011001",
  60488=>"010111011",
  60489=>"001110101",
  60490=>"000001000",
  60491=>"101000110",
  60492=>"101001010",
  60493=>"010111101",
  60494=>"100110011",
  60495=>"001111000",
  60496=>"001010001",
  60497=>"010011000",
  60498=>"111010111",
  60499=>"010111110",
  60500=>"110000111",
  60501=>"010101101",
  60502=>"101101110",
  60503=>"000100100",
  60504=>"111111110",
  60505=>"011111100",
  60506=>"000110100",
  60507=>"111100101",
  60508=>"011000101",
  60509=>"000000111",
  60510=>"111001100",
  60511=>"111101100",
  60512=>"100100001",
  60513=>"110010011",
  60514=>"000101011",
  60515=>"110100001",
  60516=>"101100001",
  60517=>"110101111",
  60518=>"101101101",
  60519=>"001101111",
  60520=>"010110010",
  60521=>"100110000",
  60522=>"001101001",
  60523=>"011011110",
  60524=>"111000000",
  60525=>"011100010",
  60526=>"000010111",
  60527=>"111100101",
  60528=>"111001101",
  60529=>"011001101",
  60530=>"000011010",
  60531=>"111111011",
  60532=>"000011100",
  60533=>"100101100",
  60534=>"110111101",
  60535=>"100111011",
  60536=>"011011000",
  60537=>"100010010",
  60538=>"100101110",
  60539=>"000000101",
  60540=>"000100010",
  60541=>"100110000",
  60542=>"001110111",
  60543=>"111000000",
  60544=>"010110110",
  60545=>"011111101",
  60546=>"011100110",
  60547=>"111011111",
  60548=>"100000101",
  60549=>"100100001",
  60550=>"010110011",
  60551=>"001100111",
  60552=>"100100101",
  60553=>"100000110",
  60554=>"100111001",
  60555=>"000111011",
  60556=>"011010001",
  60557=>"011111010",
  60558=>"011101001",
  60559=>"111110110",
  60560=>"100110000",
  60561=>"110010011",
  60562=>"011000100",
  60563=>"010110101",
  60564=>"001001110",
  60565=>"011101100",
  60566=>"010100111",
  60567=>"101001101",
  60568=>"000100100",
  60569=>"011000111",
  60570=>"100011011",
  60571=>"010000111",
  60572=>"001111001",
  60573=>"111111000",
  60574=>"010100100",
  60575=>"001000011",
  60576=>"100101001",
  60577=>"000111001",
  60578=>"000100010",
  60579=>"110111110",
  60580=>"100000000",
  60581=>"111111100",
  60582=>"001111010",
  60583=>"010000110",
  60584=>"001110000",
  60585=>"011011001",
  60586=>"010011000",
  60587=>"111101011",
  60588=>"000100000",
  60589=>"010010110",
  60590=>"101100011",
  60591=>"000110000",
  60592=>"001001101",
  60593=>"000110011",
  60594=>"101011100",
  60595=>"000010011",
  60596=>"111010000",
  60597=>"101010000",
  60598=>"011011000",
  60599=>"000001001",
  60600=>"010000000",
  60601=>"110110001",
  60602=>"000111001",
  60603=>"000111100",
  60604=>"010101001",
  60605=>"000001001",
  60606=>"000111001",
  60607=>"001101011",
  60608=>"110000100",
  60609=>"110111110",
  60610=>"101011111",
  60611=>"111110100",
  60612=>"011000010",
  60613=>"011001100",
  60614=>"000010100",
  60615=>"010011010",
  60616=>"100101110",
  60617=>"011111100",
  60618=>"111001110",
  60619=>"010101100",
  60620=>"111100010",
  60621=>"110010010",
  60622=>"101011100",
  60623=>"000011011",
  60624=>"001010101",
  60625=>"101101100",
  60626=>"010000100",
  60627=>"110010100",
  60628=>"011011100",
  60629=>"000110001",
  60630=>"010001011",
  60631=>"010110001",
  60632=>"010010101",
  60633=>"001101100",
  60634=>"101100110",
  60635=>"001000110",
  60636=>"111110100",
  60637=>"111111011",
  60638=>"100011110",
  60639=>"100101100",
  60640=>"000100000",
  60641=>"100111010",
  60642=>"000101000",
  60643=>"010001100",
  60644=>"001101011",
  60645=>"100011100",
  60646=>"100101010",
  60647=>"100010110",
  60648=>"010011101",
  60649=>"000100011",
  60650=>"110011011",
  60651=>"110010110",
  60652=>"000101111",
  60653=>"011011011",
  60654=>"001001100",
  60655=>"111010110",
  60656=>"100011010",
  60657=>"001101100",
  60658=>"010010011",
  60659=>"010101110",
  60660=>"011100000",
  60661=>"011011101",
  60662=>"101110100",
  60663=>"110100100",
  60664=>"110101011",
  60665=>"010010100",
  60666=>"100010010",
  60667=>"010001010",
  60668=>"001010010",
  60669=>"101101000",
  60670=>"011010100",
  60671=>"010111010",
  60672=>"001100101",
  60673=>"101001000",
  60674=>"101111101",
  60675=>"011010010",
  60676=>"100001111",
  60677=>"110100011",
  60678=>"001000101",
  60679=>"100010010",
  60680=>"111101001",
  60681=>"011010010",
  60682=>"110111010",
  60683=>"101111101",
  60684=>"000111011",
  60685=>"111111110",
  60686=>"000000000",
  60687=>"110101110",
  60688=>"100011010",
  60689=>"111010001",
  60690=>"100100010",
  60691=>"101110100",
  60692=>"101001101",
  60693=>"011100110",
  60694=>"001010010",
  60695=>"000001011",
  60696=>"011110110",
  60697=>"100100110",
  60698=>"111100011",
  60699=>"101100000",
  60700=>"111100101",
  60701=>"110110010",
  60702=>"011010101",
  60703=>"111010001",
  60704=>"001111010",
  60705=>"000101101",
  60706=>"101101011",
  60707=>"110101101",
  60708=>"000110101",
  60709=>"101011000",
  60710=>"011101011",
  60711=>"101110101",
  60712=>"000110000",
  60713=>"101101001",
  60714=>"011110101",
  60715=>"010000110",
  60716=>"100010001",
  60717=>"110111111",
  60718=>"000000000",
  60719=>"000011100",
  60720=>"101100011",
  60721=>"000111010",
  60722=>"100010101",
  60723=>"010111111",
  60724=>"110110000",
  60725=>"000110110",
  60726=>"110111111",
  60727=>"101000001",
  60728=>"111010001",
  60729=>"001101100",
  60730=>"110110111",
  60731=>"110101011",
  60732=>"110001001",
  60733=>"100100111",
  60734=>"001001001",
  60735=>"110100111",
  60736=>"101111111",
  60737=>"000010011",
  60738=>"001010101",
  60739=>"001111000",
  60740=>"011000100",
  60741=>"000100110",
  60742=>"101101001",
  60743=>"111000011",
  60744=>"010110100",
  60745=>"000001111",
  60746=>"111010111",
  60747=>"101011001",
  60748=>"100100010",
  60749=>"000100001",
  60750=>"101101100",
  60751=>"001111111",
  60752=>"101001011",
  60753=>"000010010",
  60754=>"001010000",
  60755=>"110111010",
  60756=>"001011001",
  60757=>"111110111",
  60758=>"111010110",
  60759=>"100100111",
  60760=>"111000000",
  60761=>"010110111",
  60762=>"011001101",
  60763=>"110101110",
  60764=>"110001101",
  60765=>"111100011",
  60766=>"001100001",
  60767=>"010010001",
  60768=>"001011010",
  60769=>"101000001",
  60770=>"001011111",
  60771=>"011101101",
  60772=>"110110101",
  60773=>"001110011",
  60774=>"100010110",
  60775=>"111000000",
  60776=>"110000010",
  60777=>"101000000",
  60778=>"000101001",
  60779=>"101111001",
  60780=>"010101001",
  60781=>"111011111",
  60782=>"110110000",
  60783=>"101010100",
  60784=>"001010000",
  60785=>"101101110",
  60786=>"111110100",
  60787=>"100010011",
  60788=>"111010000",
  60789=>"100010010",
  60790=>"101111001",
  60791=>"011001001",
  60792=>"001110111",
  60793=>"001111101",
  60794=>"100011101",
  60795=>"000111100",
  60796=>"101101010",
  60797=>"010001111",
  60798=>"000011010",
  60799=>"100100101",
  60800=>"011000000",
  60801=>"111000101",
  60802=>"000000000",
  60803=>"111100000",
  60804=>"111001011",
  60805=>"000010111",
  60806=>"101001110",
  60807=>"000100101",
  60808=>"110111100",
  60809=>"011110111",
  60810=>"010011111",
  60811=>"000111001",
  60812=>"101000110",
  60813=>"001111111",
  60814=>"110110110",
  60815=>"011011110",
  60816=>"010010001",
  60817=>"101010101",
  60818=>"101010100",
  60819=>"111010000",
  60820=>"000011100",
  60821=>"001001001",
  60822=>"110101101",
  60823=>"001110001",
  60824=>"101000101",
  60825=>"110100101",
  60826=>"101001011",
  60827=>"001011001",
  60828=>"110011110",
  60829=>"101001111",
  60830=>"101111001",
  60831=>"101101111",
  60832=>"100110000",
  60833=>"110110000",
  60834=>"000001100",
  60835=>"101111011",
  60836=>"011111000",
  60837=>"011000101",
  60838=>"110100001",
  60839=>"111110011",
  60840=>"110000010",
  60841=>"110110001",
  60842=>"010001111",
  60843=>"110110010",
  60844=>"011000111",
  60845=>"111111110",
  60846=>"000000100",
  60847=>"000100011",
  60848=>"000110100",
  60849=>"010001011",
  60850=>"111011000",
  60851=>"101001111",
  60852=>"101001111",
  60853=>"001010011",
  60854=>"000000111",
  60855=>"111011001",
  60856=>"110101111",
  60857=>"111110111",
  60858=>"011100111",
  60859=>"111101000",
  60860=>"010110111",
  60861=>"111011110",
  60862=>"001100101",
  60863=>"101101101",
  60864=>"011001001",
  60865=>"011110010",
  60866=>"010001010",
  60867=>"001110011",
  60868=>"011000000",
  60869=>"000101000",
  60870=>"000000011",
  60871=>"001110000",
  60872=>"101100100",
  60873=>"100111101",
  60874=>"001010001",
  60875=>"111010100",
  60876=>"001010001",
  60877=>"001010010",
  60878=>"001011001",
  60879=>"001100011",
  60880=>"000001100",
  60881=>"010111101",
  60882=>"001111111",
  60883=>"110100101",
  60884=>"100011111",
  60885=>"001000011",
  60886=>"100100010",
  60887=>"111111110",
  60888=>"010011101",
  60889=>"111110101",
  60890=>"000000111",
  60891=>"111000000",
  60892=>"110111100",
  60893=>"101000111",
  60894=>"111100100",
  60895=>"100011001",
  60896=>"001010110",
  60897=>"011110011",
  60898=>"001000100",
  60899=>"111111000",
  60900=>"111101100",
  60901=>"011111111",
  60902=>"011100011",
  60903=>"101011010",
  60904=>"010111010",
  60905=>"000111100",
  60906=>"110100100",
  60907=>"100100011",
  60908=>"000001000",
  60909=>"011010001",
  60910=>"100001000",
  60911=>"001010010",
  60912=>"100001111",
  60913=>"011010111",
  60914=>"000011000",
  60915=>"100101111",
  60916=>"100000000",
  60917=>"010000001",
  60918=>"010000110",
  60919=>"011111010",
  60920=>"001110001",
  60921=>"110011000",
  60922=>"001100001",
  60923=>"001110000",
  60924=>"100001111",
  60925=>"111101110",
  60926=>"100111101",
  60927=>"110100000",
  60928=>"000100000",
  60929=>"010010111",
  60930=>"000001001",
  60931=>"000100101",
  60932=>"011001111",
  60933=>"101100111",
  60934=>"101000101",
  60935=>"101110111",
  60936=>"100110001",
  60937=>"101100010",
  60938=>"000001110",
  60939=>"001111101",
  60940=>"000010001",
  60941=>"010101011",
  60942=>"110110111",
  60943=>"001000001",
  60944=>"110000101",
  60945=>"010011011",
  60946=>"000110011",
  60947=>"111111100",
  60948=>"010100001",
  60949=>"010000011",
  60950=>"000100100",
  60951=>"010000010",
  60952=>"001111010",
  60953=>"101101000",
  60954=>"100100100",
  60955=>"100000000",
  60956=>"000000011",
  60957=>"110000001",
  60958=>"000110101",
  60959=>"101110110",
  60960=>"011101110",
  60961=>"101001101",
  60962=>"001100101",
  60963=>"110110111",
  60964=>"111001100",
  60965=>"100101011",
  60966=>"010110001",
  60967=>"001010100",
  60968=>"001011100",
  60969=>"001001101",
  60970=>"100111010",
  60971=>"010110000",
  60972=>"001001010",
  60973=>"101111001",
  60974=>"100010101",
  60975=>"010001100",
  60976=>"110110010",
  60977=>"010111110",
  60978=>"101110011",
  60979=>"110001001",
  60980=>"001000100",
  60981=>"000111010",
  60982=>"100000000",
  60983=>"000000111",
  60984=>"011101111",
  60985=>"001110100",
  60986=>"110010001",
  60987=>"011000011",
  60988=>"110100100",
  60989=>"110110001",
  60990=>"100111110",
  60991=>"010111010",
  60992=>"000000100",
  60993=>"100101010",
  60994=>"101001000",
  60995=>"111110100",
  60996=>"011001001",
  60997=>"100001100",
  60998=>"111100110",
  60999=>"111011011",
  61000=>"000100010",
  61001=>"101110010",
  61002=>"100000101",
  61003=>"001100101",
  61004=>"100111011",
  61005=>"100001101",
  61006=>"101110101",
  61007=>"111110110",
  61008=>"100010001",
  61009=>"111001000",
  61010=>"011011101",
  61011=>"000000010",
  61012=>"110110101",
  61013=>"000110111",
  61014=>"111000111",
  61015=>"110000100",
  61016=>"111100000",
  61017=>"010101110",
  61018=>"110010011",
  61019=>"000110000",
  61020=>"011010000",
  61021=>"011001101",
  61022=>"000100110",
  61023=>"011011100",
  61024=>"101100111",
  61025=>"011110010",
  61026=>"100101011",
  61027=>"001100011",
  61028=>"100011100",
  61029=>"010111100",
  61030=>"011001100",
  61031=>"100101100",
  61032=>"101000111",
  61033=>"000010000",
  61034=>"111111011",
  61035=>"110110101",
  61036=>"000111001",
  61037=>"001111111",
  61038=>"110111100",
  61039=>"010111111",
  61040=>"111000010",
  61041=>"111011000",
  61042=>"000010000",
  61043=>"101011100",
  61044=>"101011100",
  61045=>"111000101",
  61046=>"010010010",
  61047=>"110000000",
  61048=>"011100000",
  61049=>"011001001",
  61050=>"111101100",
  61051=>"011010100",
  61052=>"010010000",
  61053=>"111111011",
  61054=>"010011001",
  61055=>"001000110",
  61056=>"010001000",
  61057=>"000001000",
  61058=>"011111111",
  61059=>"000000011",
  61060=>"111001011",
  61061=>"011010000",
  61062=>"101110011",
  61063=>"110010111",
  61064=>"110110000",
  61065=>"101110000",
  61066=>"010100010",
  61067=>"000000011",
  61068=>"011000010",
  61069=>"001001110",
  61070=>"111010110",
  61071=>"101101110",
  61072=>"111000101",
  61073=>"111010010",
  61074=>"010010001",
  61075=>"101100100",
  61076=>"100000110",
  61077=>"010001111",
  61078=>"111100100",
  61079=>"000001110",
  61080=>"001111111",
  61081=>"110001010",
  61082=>"010011001",
  61083=>"001100101",
  61084=>"010000000",
  61085=>"000100001",
  61086=>"101100100",
  61087=>"111101011",
  61088=>"010101010",
  61089=>"011011010",
  61090=>"000100010",
  61091=>"011101011",
  61092=>"101101000",
  61093=>"010111001",
  61094=>"010000110",
  61095=>"010000000",
  61096=>"010101010",
  61097=>"111111001",
  61098=>"001010101",
  61099=>"001010010",
  61100=>"110011111",
  61101=>"011101111",
  61102=>"111000100",
  61103=>"001101100",
  61104=>"010010110",
  61105=>"100001001",
  61106=>"101000111",
  61107=>"110010110",
  61108=>"011110000",
  61109=>"100001001",
  61110=>"101110000",
  61111=>"000110111",
  61112=>"111011110",
  61113=>"000000010",
  61114=>"010101111",
  61115=>"100000000",
  61116=>"000000111",
  61117=>"111101011",
  61118=>"111000000",
  61119=>"101111100",
  61120=>"001001111",
  61121=>"111011100",
  61122=>"001000011",
  61123=>"111000101",
  61124=>"110101000",
  61125=>"000001100",
  61126=>"111110110",
  61127=>"011100101",
  61128=>"111110010",
  61129=>"110001000",
  61130=>"110111010",
  61131=>"110001000",
  61132=>"000011010",
  61133=>"011110010",
  61134=>"111011111",
  61135=>"000110111",
  61136=>"011001111",
  61137=>"010010011",
  61138=>"101110101",
  61139=>"010100110",
  61140=>"000001000",
  61141=>"111100101",
  61142=>"100101100",
  61143=>"111000000",
  61144=>"000101010",
  61145=>"011011001",
  61146=>"110111101",
  61147=>"100000000",
  61148=>"000100011",
  61149=>"011010000",
  61150=>"000101010",
  61151=>"100110001",
  61152=>"110011011",
  61153=>"001000001",
  61154=>"001010010",
  61155=>"101110001",
  61156=>"101010010",
  61157=>"000001111",
  61158=>"110011101",
  61159=>"101100111",
  61160=>"111100000",
  61161=>"000000111",
  61162=>"110010001",
  61163=>"010000101",
  61164=>"010000101",
  61165=>"110000111",
  61166=>"111111000",
  61167=>"010010000",
  61168=>"101110101",
  61169=>"111010000",
  61170=>"100000000",
  61171=>"010110000",
  61172=>"101111010",
  61173=>"101100100",
  61174=>"111111110",
  61175=>"011111000",
  61176=>"000010000",
  61177=>"100111110",
  61178=>"100011101",
  61179=>"011110101",
  61180=>"100000011",
  61181=>"111010010",
  61182=>"000110100",
  61183=>"101010010",
  61184=>"000010010",
  61185=>"101100100",
  61186=>"010000010",
  61187=>"010000010",
  61188=>"110000111",
  61189=>"010001110",
  61190=>"000010111",
  61191=>"000000101",
  61192=>"101001001",
  61193=>"001000000",
  61194=>"000000110",
  61195=>"000011111",
  61196=>"100000111",
  61197=>"011101110",
  61198=>"010100000",
  61199=>"111101101",
  61200=>"101011101",
  61201=>"111110100",
  61202=>"011001111",
  61203=>"000011010",
  61204=>"000010110",
  61205=>"100001111",
  61206=>"011111001",
  61207=>"101010110",
  61208=>"101001100",
  61209=>"101100000",
  61210=>"000000110",
  61211=>"101010000",
  61212=>"101111110",
  61213=>"001000101",
  61214=>"000000101",
  61215=>"110000110",
  61216=>"011111000",
  61217=>"111111101",
  61218=>"000101101",
  61219=>"010001011",
  61220=>"101011101",
  61221=>"110111011",
  61222=>"111011101",
  61223=>"101000000",
  61224=>"101111001",
  61225=>"010100111",
  61226=>"110000010",
  61227=>"110111000",
  61228=>"111010011",
  61229=>"111000011",
  61230=>"011001101",
  61231=>"111111011",
  61232=>"010001101",
  61233=>"000010001",
  61234=>"100110000",
  61235=>"011111101",
  61236=>"101001000",
  61237=>"011111000",
  61238=>"111110110",
  61239=>"111010011",
  61240=>"101000101",
  61241=>"110011011",
  61242=>"011100111",
  61243=>"011100110",
  61244=>"001111111",
  61245=>"010011000",
  61246=>"101010110",
  61247=>"101000110",
  61248=>"010101100",
  61249=>"111000101",
  61250=>"000001000",
  61251=>"000101100",
  61252=>"000100101",
  61253=>"101110011",
  61254=>"001000101",
  61255=>"100110100",
  61256=>"001110111",
  61257=>"111101111",
  61258=>"111111000",
  61259=>"101001001",
  61260=>"010000100",
  61261=>"001101010",
  61262=>"100000111",
  61263=>"111010111",
  61264=>"000001010",
  61265=>"000100101",
  61266=>"000011001",
  61267=>"110000110",
  61268=>"000101111",
  61269=>"010100111",
  61270=>"010000110",
  61271=>"101011100",
  61272=>"010101111",
  61273=>"000001001",
  61274=>"010111110",
  61275=>"111110101",
  61276=>"001000100",
  61277=>"011101110",
  61278=>"100010111",
  61279=>"000000101",
  61280=>"010101010",
  61281=>"110000000",
  61282=>"001000011",
  61283=>"101000001",
  61284=>"001100111",
  61285=>"010010001",
  61286=>"000101110",
  61287=>"000011000",
  61288=>"111011010",
  61289=>"101100000",
  61290=>"111101111",
  61291=>"111110001",
  61292=>"111011100",
  61293=>"110001011",
  61294=>"010101011",
  61295=>"010011111",
  61296=>"110101110",
  61297=>"111101111",
  61298=>"100011010",
  61299=>"010000101",
  61300=>"000010111",
  61301=>"000101011",
  61302=>"011100011",
  61303=>"000110010",
  61304=>"101101101",
  61305=>"100110001",
  61306=>"101110111",
  61307=>"000001110",
  61308=>"100101011",
  61309=>"101000000",
  61310=>"001011111",
  61311=>"001000101",
  61312=>"101001011",
  61313=>"110101000",
  61314=>"001011111",
  61315=>"101000100",
  61316=>"001001111",
  61317=>"111111110",
  61318=>"001000100",
  61319=>"101000100",
  61320=>"101011111",
  61321=>"000010010",
  61322=>"110011111",
  61323=>"010000010",
  61324=>"010001111",
  61325=>"000100101",
  61326=>"101011101",
  61327=>"101011010",
  61328=>"110011111",
  61329=>"110101100",
  61330=>"010000010",
  61331=>"110111011",
  61332=>"110011101",
  61333=>"001101010",
  61334=>"001101010",
  61335=>"010101010",
  61336=>"101000010",
  61337=>"000001010",
  61338=>"101100101",
  61339=>"000101111",
  61340=>"111010000",
  61341=>"100010111",
  61342=>"011100111",
  61343=>"110110110",
  61344=>"100011000",
  61345=>"110011001",
  61346=>"101000000",
  61347=>"011101111",
  61348=>"000101101",
  61349=>"010001100",
  61350=>"000011000",
  61351=>"001010000",
  61352=>"101111011",
  61353=>"010011101",
  61354=>"110111010",
  61355=>"011101000",
  61356=>"010011011",
  61357=>"000111000",
  61358=>"101110011",
  61359=>"100001000",
  61360=>"100000100",
  61361=>"010001101",
  61362=>"010000001",
  61363=>"001100111",
  61364=>"011111110",
  61365=>"110111110",
  61366=>"001000000",
  61367=>"011100111",
  61368=>"010000101",
  61369=>"111100111",
  61370=>"110101100",
  61371=>"111100000",
  61372=>"001111111",
  61373=>"001101001",
  61374=>"101000101",
  61375=>"101101000",
  61376=>"110000000",
  61377=>"101000001",
  61378=>"111111101",
  61379=>"101001011",
  61380=>"111011011",
  61381=>"011101100",
  61382=>"000011001",
  61383=>"110110101",
  61384=>"100000100",
  61385=>"011001000",
  61386=>"001101000",
  61387=>"011011000",
  61388=>"010110000",
  61389=>"010101010",
  61390=>"001001000",
  61391=>"110100000",
  61392=>"011011001",
  61393=>"000000101",
  61394=>"100111010",
  61395=>"110111001",
  61396=>"101000111",
  61397=>"111001011",
  61398=>"000011111",
  61399=>"101011110",
  61400=>"000110110",
  61401=>"000001010",
  61402=>"010110010",
  61403=>"000000001",
  61404=>"011101001",
  61405=>"111000001",
  61406=>"111100101",
  61407=>"000011110",
  61408=>"111111011",
  61409=>"110110001",
  61410=>"111000011",
  61411=>"001000011",
  61412=>"010010001",
  61413=>"100010100",
  61414=>"110101001",
  61415=>"111101010",
  61416=>"110100000",
  61417=>"100000000",
  61418=>"011100001",
  61419=>"001110110",
  61420=>"101110010",
  61421=>"000100001",
  61422=>"001110100",
  61423=>"111100100",
  61424=>"110001111",
  61425=>"111011000",
  61426=>"000000111",
  61427=>"100101000",
  61428=>"110101110",
  61429=>"101001010",
  61430=>"110000101",
  61431=>"000110101",
  61432=>"111011110",
  61433=>"101001000",
  61434=>"101010011",
  61435=>"001000101",
  61436=>"010110100",
  61437=>"101101011",
  61438=>"010001111",
  61439=>"001001110",
  61440=>"100000111",
  61441=>"100010111",
  61442=>"110011001",
  61443=>"101000000",
  61444=>"100110001",
  61445=>"010011001",
  61446=>"100110010",
  61447=>"101111110",
  61448=>"101011110",
  61449=>"100111011",
  61450=>"001111011",
  61451=>"000101110",
  61452=>"010010100",
  61453=>"001111111",
  61454=>"100101000",
  61455=>"110111100",
  61456=>"011010100",
  61457=>"101001111",
  61458=>"010111111",
  61459=>"001101101",
  61460=>"000000011",
  61461=>"111100110",
  61462=>"110001000",
  61463=>"011000101",
  61464=>"001000111",
  61465=>"000001100",
  61466=>"110010000",
  61467=>"101110110",
  61468=>"000101011",
  61469=>"000011010",
  61470=>"101111010",
  61471=>"011100111",
  61472=>"100110110",
  61473=>"100010111",
  61474=>"111010100",
  61475=>"000001011",
  61476=>"101011011",
  61477=>"010010111",
  61478=>"111010100",
  61479=>"011010110",
  61480=>"110101101",
  61481=>"001100100",
  61482=>"001111010",
  61483=>"001000001",
  61484=>"000000100",
  61485=>"001100100",
  61486=>"011000001",
  61487=>"110100100",
  61488=>"001001001",
  61489=>"010100110",
  61490=>"011011001",
  61491=>"010111001",
  61492=>"111111011",
  61493=>"101100001",
  61494=>"100111101",
  61495=>"010101101",
  61496=>"000001010",
  61497=>"011011101",
  61498=>"111011010",
  61499=>"001010100",
  61500=>"001011100",
  61501=>"111000000",
  61502=>"101100000",
  61503=>"000001000",
  61504=>"100100010",
  61505=>"001101010",
  61506=>"101100110",
  61507=>"011010110",
  61508=>"010110100",
  61509=>"110101110",
  61510=>"110010011",
  61511=>"010100011",
  61512=>"100011010",
  61513=>"010011011",
  61514=>"011000000",
  61515=>"101010011",
  61516=>"001000011",
  61517=>"010100011",
  61518=>"110111101",
  61519=>"110101010",
  61520=>"011001000",
  61521=>"111101110",
  61522=>"010101001",
  61523=>"100010101",
  61524=>"111100000",
  61525=>"110000010",
  61526=>"000011111",
  61527=>"010110100",
  61528=>"001100101",
  61529=>"110101110",
  61530=>"000100010",
  61531=>"010000111",
  61532=>"000111011",
  61533=>"110110101",
  61534=>"100000110",
  61535=>"010001000",
  61536=>"111111111",
  61537=>"000001000",
  61538=>"011101101",
  61539=>"101111111",
  61540=>"111101001",
  61541=>"010010110",
  61542=>"000010011",
  61543=>"010100001",
  61544=>"010011111",
  61545=>"110001111",
  61546=>"010100011",
  61547=>"111011100",
  61548=>"010011100",
  61549=>"011011111",
  61550=>"101010100",
  61551=>"111100100",
  61552=>"010010000",
  61553=>"010000011",
  61554=>"101110011",
  61555=>"000110010",
  61556=>"000001011",
  61557=>"110001011",
  61558=>"000101001",
  61559=>"100110101",
  61560=>"001001101",
  61561=>"001111100",
  61562=>"011101000",
  61563=>"101110010",
  61564=>"101100001",
  61565=>"010100000",
  61566=>"001010000",
  61567=>"010110001",
  61568=>"001011001",
  61569=>"101010000",
  61570=>"000110111",
  61571=>"001000001",
  61572=>"001010101",
  61573=>"000000101",
  61574=>"001100110",
  61575=>"111101101",
  61576=>"101100111",
  61577=>"001011111",
  61578=>"101000001",
  61579=>"111110001",
  61580=>"100001111",
  61581=>"100100011",
  61582=>"010011001",
  61583=>"110100001",
  61584=>"000011110",
  61585=>"011001000",
  61586=>"011111010",
  61587=>"111011101",
  61588=>"101000000",
  61589=>"111000000",
  61590=>"110010100",
  61591=>"000001101",
  61592=>"000000010",
  61593=>"000110110",
  61594=>"111100010",
  61595=>"000101000",
  61596=>"000110010",
  61597=>"100001101",
  61598=>"110011011",
  61599=>"011100101",
  61600=>"100101100",
  61601=>"100001100",
  61602=>"111001111",
  61603=>"110101001",
  61604=>"000011001",
  61605=>"110001100",
  61606=>"100001100",
  61607=>"000001000",
  61608=>"101101100",
  61609=>"100011001",
  61610=>"111111000",
  61611=>"101001000",
  61612=>"100111000",
  61613=>"100010101",
  61614=>"111010000",
  61615=>"101111001",
  61616=>"111001001",
  61617=>"000000001",
  61618=>"111001010",
  61619=>"110111011",
  61620=>"001110011",
  61621=>"000000101",
  61622=>"100000010",
  61623=>"011110111",
  61624=>"111001100",
  61625=>"110011000",
  61626=>"111111101",
  61627=>"100010010",
  61628=>"010010101",
  61629=>"000111011",
  61630=>"100000111",
  61631=>"111110111",
  61632=>"001001011",
  61633=>"010011011",
  61634=>"100011010",
  61635=>"000100110",
  61636=>"100010011",
  61637=>"110011011",
  61638=>"010001001",
  61639=>"010101001",
  61640=>"010100001",
  61641=>"110010000",
  61642=>"001111110",
  61643=>"000111000",
  61644=>"000100100",
  61645=>"010111111",
  61646=>"001111010",
  61647=>"001010110",
  61648=>"110101011",
  61649=>"101010110",
  61650=>"110010111",
  61651=>"111110000",
  61652=>"100101011",
  61653=>"001101110",
  61654=>"100101000",
  61655=>"101100110",
  61656=>"101111101",
  61657=>"101100010",
  61658=>"111001101",
  61659=>"001110110",
  61660=>"001000101",
  61661=>"101001100",
  61662=>"000010000",
  61663=>"111101001",
  61664=>"111110010",
  61665=>"000001110",
  61666=>"101111101",
  61667=>"011111111",
  61668=>"011110111",
  61669=>"101111111",
  61670=>"011101010",
  61671=>"011010000",
  61672=>"101010101",
  61673=>"101000001",
  61674=>"111011000",
  61675=>"101101111",
  61676=>"100100100",
  61677=>"000000110",
  61678=>"000110011",
  61679=>"010111101",
  61680=>"100011110",
  61681=>"010000111",
  61682=>"000100001",
  61683=>"010110001",
  61684=>"111110100",
  61685=>"110100011",
  61686=>"101101000",
  61687=>"010010111",
  61688=>"001111111",
  61689=>"001101101",
  61690=>"001100000",
  61691=>"101001001",
  61692=>"111001110",
  61693=>"000010001",
  61694=>"010100101",
  61695=>"101111010",
  61696=>"111011011",
  61697=>"010101100",
  61698=>"010111110",
  61699=>"011110000",
  61700=>"000100101",
  61701=>"010110010",
  61702=>"101101100",
  61703=>"000101100",
  61704=>"010000011",
  61705=>"000100000",
  61706=>"010101010",
  61707=>"000111100",
  61708=>"110110111",
  61709=>"110000000",
  61710=>"101110010",
  61711=>"000011101",
  61712=>"110010101",
  61713=>"101100011",
  61714=>"101101001",
  61715=>"110101111",
  61716=>"010100111",
  61717=>"100111011",
  61718=>"010101010",
  61719=>"011110101",
  61720=>"011101111",
  61721=>"010000010",
  61722=>"100101111",
  61723=>"011111111",
  61724=>"001011101",
  61725=>"101111011",
  61726=>"001110110",
  61727=>"001011000",
  61728=>"111001001",
  61729=>"100101001",
  61730=>"101010010",
  61731=>"100011101",
  61732=>"001100001",
  61733=>"100100101",
  61734=>"101111011",
  61735=>"111010001",
  61736=>"001000000",
  61737=>"011010011",
  61738=>"111110100",
  61739=>"001110111",
  61740=>"000100111",
  61741=>"011111110",
  61742=>"101000101",
  61743=>"001111100",
  61744=>"010010100",
  61745=>"101001100",
  61746=>"100101000",
  61747=>"001101100",
  61748=>"100110101",
  61749=>"000110001",
  61750=>"111000110",
  61751=>"001101111",
  61752=>"111101101",
  61753=>"000011101",
  61754=>"010001111",
  61755=>"100111010",
  61756=>"010010110",
  61757=>"110010000",
  61758=>"001101111",
  61759=>"101110010",
  61760=>"110110000",
  61761=>"000111101",
  61762=>"100111010",
  61763=>"010101100",
  61764=>"110011011",
  61765=>"001100011",
  61766=>"011101100",
  61767=>"110011011",
  61768=>"000001000",
  61769=>"001011110",
  61770=>"100100000",
  61771=>"110101001",
  61772=>"101001111",
  61773=>"000111111",
  61774=>"110111110",
  61775=>"000011110",
  61776=>"111100110",
  61777=>"101100101",
  61778=>"101111011",
  61779=>"111000101",
  61780=>"001011010",
  61781=>"000010100",
  61782=>"001010111",
  61783=>"001111101",
  61784=>"000000101",
  61785=>"100111011",
  61786=>"111010010",
  61787=>"000110101",
  61788=>"110100111",
  61789=>"001010110",
  61790=>"011010011",
  61791=>"001001110",
  61792=>"110111010",
  61793=>"110111101",
  61794=>"000101100",
  61795=>"010111001",
  61796=>"010000101",
  61797=>"101000100",
  61798=>"111101011",
  61799=>"111111100",
  61800=>"111100110",
  61801=>"000001000",
  61802=>"101001010",
  61803=>"000001000",
  61804=>"001101011",
  61805=>"010011100",
  61806=>"101100110",
  61807=>"100011101",
  61808=>"000000110",
  61809=>"000000011",
  61810=>"110110000",
  61811=>"110001110",
  61812=>"001110000",
  61813=>"110010111",
  61814=>"010011000",
  61815=>"001001001",
  61816=>"011001110",
  61817=>"101001100",
  61818=>"111101000",
  61819=>"001010111",
  61820=>"000011001",
  61821=>"110011101",
  61822=>"000011011",
  61823=>"110111010",
  61824=>"111110111",
  61825=>"011000010",
  61826=>"100011100",
  61827=>"001001111",
  61828=>"000110100",
  61829=>"111001011",
  61830=>"010011001",
  61831=>"011100011",
  61832=>"001001111",
  61833=>"011010101",
  61834=>"000011100",
  61835=>"100000000",
  61836=>"011111110",
  61837=>"101111100",
  61838=>"100101110",
  61839=>"100101101",
  61840=>"110011110",
  61841=>"011100000",
  61842=>"110110010",
  61843=>"100010100",
  61844=>"001100101",
  61845=>"000100100",
  61846=>"001111001",
  61847=>"110110011",
  61848=>"100011001",
  61849=>"110010010",
  61850=>"110110101",
  61851=>"000101100",
  61852=>"011010010",
  61853=>"010011010",
  61854=>"000011101",
  61855=>"000110011",
  61856=>"101101001",
  61857=>"000111100",
  61858=>"111100101",
  61859=>"011101101",
  61860=>"010111000",
  61861=>"001101011",
  61862=>"110011110",
  61863=>"100111111",
  61864=>"011110101",
  61865=>"011111110",
  61866=>"010000001",
  61867=>"100111101",
  61868=>"110011111",
  61869=>"100000011",
  61870=>"000100111",
  61871=>"110011000",
  61872=>"111110010",
  61873=>"000001011",
  61874=>"001011111",
  61875=>"101111110",
  61876=>"011000100",
  61877=>"011100111",
  61878=>"100001000",
  61879=>"011101011",
  61880=>"010101100",
  61881=>"100011001",
  61882=>"001111101",
  61883=>"111101100",
  61884=>"110100101",
  61885=>"100010110",
  61886=>"101100011",
  61887=>"111001100",
  61888=>"110111110",
  61889=>"010101001",
  61890=>"100111101",
  61891=>"000000101",
  61892=>"010000010",
  61893=>"101000011",
  61894=>"000011010",
  61895=>"010101000",
  61896=>"000100010",
  61897=>"001001110",
  61898=>"010000000",
  61899=>"000111100",
  61900=>"011001110",
  61901=>"000110110",
  61902=>"000111100",
  61903=>"001000011",
  61904=>"000110100",
  61905=>"100001000",
  61906=>"011101010",
  61907=>"001111010",
  61908=>"111010011",
  61909=>"101100101",
  61910=>"001011111",
  61911=>"111010011",
  61912=>"110001100",
  61913=>"110101000",
  61914=>"001100100",
  61915=>"111001001",
  61916=>"010010000",
  61917=>"101001101",
  61918=>"000010010",
  61919=>"000000100",
  61920=>"010011010",
  61921=>"011000101",
  61922=>"100011001",
  61923=>"101000010",
  61924=>"000101111",
  61925=>"100011101",
  61926=>"010010111",
  61927=>"101000011",
  61928=>"010000010",
  61929=>"000010001",
  61930=>"010110111",
  61931=>"101000001",
  61932=>"010101101",
  61933=>"101101011",
  61934=>"011001101",
  61935=>"000101100",
  61936=>"101001010",
  61937=>"110101001",
  61938=>"101100111",
  61939=>"011101011",
  61940=>"001011011",
  61941=>"100000010",
  61942=>"000111100",
  61943=>"000000110",
  61944=>"011000010",
  61945=>"000100000",
  61946=>"010001010",
  61947=>"110101101",
  61948=>"000110111",
  61949=>"001101110",
  61950=>"100011011",
  61951=>"000111110",
  61952=>"010100011",
  61953=>"000100100",
  61954=>"010001010",
  61955=>"110010100",
  61956=>"011000010",
  61957=>"101010000",
  61958=>"100101010",
  61959=>"011001001",
  61960=>"011100000",
  61961=>"010111111",
  61962=>"110011001",
  61963=>"100111100",
  61964=>"111101010",
  61965=>"111000000",
  61966=>"011001111",
  61967=>"110101011",
  61968=>"001000101",
  61969=>"101110000",
  61970=>"010001010",
  61971=>"000000000",
  61972=>"010111111",
  61973=>"001001001",
  61974=>"001111011",
  61975=>"000010011",
  61976=>"011110111",
  61977=>"010110001",
  61978=>"100100000",
  61979=>"011011100",
  61980=>"000101100",
  61981=>"001100000",
  61982=>"000001111",
  61983=>"100011001",
  61984=>"100001111",
  61985=>"100010111",
  61986=>"010010111",
  61987=>"100100000",
  61988=>"100101111",
  61989=>"000000111",
  61990=>"011000010",
  61991=>"111111111",
  61992=>"000111010",
  61993=>"111101000",
  61994=>"000001100",
  61995=>"100011110",
  61996=>"010000010",
  61997=>"110001011",
  61998=>"011000110",
  61999=>"000010110",
  62000=>"010010101",
  62001=>"100100010",
  62002=>"111100001",
  62003=>"111000110",
  62004=>"110001010",
  62005=>"101101111",
  62006=>"001111001",
  62007=>"111000001",
  62008=>"000011111",
  62009=>"111011011",
  62010=>"100100000",
  62011=>"111010100",
  62012=>"011101000",
  62013=>"000001011",
  62014=>"100010101",
  62015=>"011011011",
  62016=>"100001111",
  62017=>"010001010",
  62018=>"011010010",
  62019=>"101111100",
  62020=>"010110111",
  62021=>"000111101",
  62022=>"101111111",
  62023=>"001001110",
  62024=>"010101001",
  62025=>"111101000",
  62026=>"011100111",
  62027=>"011110110",
  62028=>"000001100",
  62029=>"000101111",
  62030=>"111000011",
  62031=>"110001110",
  62032=>"000001011",
  62033=>"001000101",
  62034=>"011111011",
  62035=>"101001011",
  62036=>"100011001",
  62037=>"100000101",
  62038=>"000100101",
  62039=>"000101001",
  62040=>"000010011",
  62041=>"111000110",
  62042=>"010101001",
  62043=>"000011011",
  62044=>"000010111",
  62045=>"110110010",
  62046=>"010101001",
  62047=>"100011111",
  62048=>"000001100",
  62049=>"111011001",
  62050=>"110011100",
  62051=>"000111111",
  62052=>"000111100",
  62053=>"110101111",
  62054=>"001000111",
  62055=>"010000001",
  62056=>"011100101",
  62057=>"010010001",
  62058=>"011100010",
  62059=>"000100011",
  62060=>"011001011",
  62061=>"001111000",
  62062=>"011101110",
  62063=>"100111011",
  62064=>"000111101",
  62065=>"110101111",
  62066=>"001101111",
  62067=>"010010001",
  62068=>"000010010",
  62069=>"101010000",
  62070=>"101000000",
  62071=>"000110110",
  62072=>"010011100",
  62073=>"010000111",
  62074=>"000110110",
  62075=>"001111110",
  62076=>"111011010",
  62077=>"010110110",
  62078=>"011010111",
  62079=>"100100001",
  62080=>"001111100",
  62081=>"101101110",
  62082=>"001000110",
  62083=>"100011001",
  62084=>"110110110",
  62085=>"001010010",
  62086=>"100101010",
  62087=>"111111010",
  62088=>"001000011",
  62089=>"001001111",
  62090=>"010100101",
  62091=>"001000001",
  62092=>"000001001",
  62093=>"111000101",
  62094=>"111011000",
  62095=>"010101011",
  62096=>"000101100",
  62097=>"010011011",
  62098=>"001001111",
  62099=>"110111110",
  62100=>"110110100",
  62101=>"100010001",
  62102=>"100110100",
  62103=>"101101000",
  62104=>"111010011",
  62105=>"011011101",
  62106=>"000011011",
  62107=>"101001000",
  62108=>"010110111",
  62109=>"110111110",
  62110=>"010010000",
  62111=>"001100100",
  62112=>"001111011",
  62113=>"110100011",
  62114=>"111111110",
  62115=>"100001101",
  62116=>"110001000",
  62117=>"000011110",
  62118=>"111110001",
  62119=>"110111110",
  62120=>"110101000",
  62121=>"000001001",
  62122=>"000000001",
  62123=>"111100001",
  62124=>"101010000",
  62125=>"101100001",
  62126=>"000000101",
  62127=>"000100100",
  62128=>"010111011",
  62129=>"010101011",
  62130=>"111010011",
  62131=>"110110001",
  62132=>"110100000",
  62133=>"001000000",
  62134=>"111111011",
  62135=>"011000001",
  62136=>"100100111",
  62137=>"001001010",
  62138=>"111001110",
  62139=>"000111001",
  62140=>"001011111",
  62141=>"101011100",
  62142=>"110111010",
  62143=>"011001111",
  62144=>"100000001",
  62145=>"001000100",
  62146=>"110110111",
  62147=>"100001110",
  62148=>"001100010",
  62149=>"010011110",
  62150=>"000111000",
  62151=>"000010111",
  62152=>"101001000",
  62153=>"001001101",
  62154=>"000110111",
  62155=>"110110110",
  62156=>"001100010",
  62157=>"000011110",
  62158=>"101001110",
  62159=>"110001011",
  62160=>"111111010",
  62161=>"100000011",
  62162=>"101000000",
  62163=>"100000101",
  62164=>"001110100",
  62165=>"001110010",
  62166=>"101101000",
  62167=>"000001011",
  62168=>"001101100",
  62169=>"110101101",
  62170=>"110110001",
  62171=>"111111001",
  62172=>"111010011",
  62173=>"100111100",
  62174=>"111111000",
  62175=>"000100000",
  62176=>"111110000",
  62177=>"110111001",
  62178=>"100100001",
  62179=>"111010101",
  62180=>"100001011",
  62181=>"101111110",
  62182=>"000101000",
  62183=>"111110100",
  62184=>"000000010",
  62185=>"101101001",
  62186=>"110011000",
  62187=>"000000001",
  62188=>"110100101",
  62189=>"101101110",
  62190=>"111010110",
  62191=>"001110111",
  62192=>"001100110",
  62193=>"011001000",
  62194=>"010010010",
  62195=>"000000000",
  62196=>"000101011",
  62197=>"000000110",
  62198=>"001000111",
  62199=>"100111101",
  62200=>"011011000",
  62201=>"111101110",
  62202=>"100010111",
  62203=>"001110110",
  62204=>"101111101",
  62205=>"110010110",
  62206=>"101101001",
  62207=>"100010111",
  62208=>"000100101",
  62209=>"010111000",
  62210=>"010111000",
  62211=>"001000010",
  62212=>"101110100",
  62213=>"110100000",
  62214=>"100000010",
  62215=>"111100011",
  62216=>"110100000",
  62217=>"011111101",
  62218=>"100110111",
  62219=>"101110011",
  62220=>"010100011",
  62221=>"011110110",
  62222=>"101001001",
  62223=>"101010110",
  62224=>"100000001",
  62225=>"011011011",
  62226=>"111100010",
  62227=>"001101010",
  62228=>"010100000",
  62229=>"110100101",
  62230=>"100111100",
  62231=>"001000001",
  62232=>"110011001",
  62233=>"000101001",
  62234=>"111000111",
  62235=>"100000000",
  62236=>"011110011",
  62237=>"011111110",
  62238=>"011000000",
  62239=>"111000111",
  62240=>"101101001",
  62241=>"001000011",
  62242=>"101011111",
  62243=>"110111101",
  62244=>"011000111",
  62245=>"101101101",
  62246=>"000000000",
  62247=>"110110110",
  62248=>"110000010",
  62249=>"111101000",
  62250=>"110110001",
  62251=>"101010000",
  62252=>"100100010",
  62253=>"011111100",
  62254=>"011111101",
  62255=>"001011111",
  62256=>"111000111",
  62257=>"001100000",
  62258=>"100100110",
  62259=>"000110010",
  62260=>"110001011",
  62261=>"010010001",
  62262=>"110110111",
  62263=>"100010000",
  62264=>"100101111",
  62265=>"000111011",
  62266=>"001000100",
  62267=>"010111111",
  62268=>"011001001",
  62269=>"000111111",
  62270=>"100111000",
  62271=>"110001101",
  62272=>"100000100",
  62273=>"000001010",
  62274=>"100010000",
  62275=>"100111110",
  62276=>"011111010",
  62277=>"101010111",
  62278=>"111111010",
  62279=>"110101011",
  62280=>"001010000",
  62281=>"010110100",
  62282=>"001101011",
  62283=>"101111011",
  62284=>"100101001",
  62285=>"110101101",
  62286=>"000001010",
  62287=>"010100101",
  62288=>"110101110",
  62289=>"010000101",
  62290=>"011010000",
  62291=>"000000010",
  62292=>"000011010",
  62293=>"100010101",
  62294=>"110001111",
  62295=>"111100011",
  62296=>"111100011",
  62297=>"111000000",
  62298=>"110101101",
  62299=>"101100101",
  62300=>"111100000",
  62301=>"000000000",
  62302=>"110111000",
  62303=>"111110010",
  62304=>"000111010",
  62305=>"111011110",
  62306=>"110110101",
  62307=>"101100001",
  62308=>"011110010",
  62309=>"100110011",
  62310=>"101110010",
  62311=>"111010111",
  62312=>"010011100",
  62313=>"010110100",
  62314=>"111001100",
  62315=>"001101010",
  62316=>"010010011",
  62317=>"101101111",
  62318=>"011110101",
  62319=>"000011101",
  62320=>"100100110",
  62321=>"000100100",
  62322=>"111011101",
  62323=>"011011101",
  62324=>"011100111",
  62325=>"000001101",
  62326=>"011101000",
  62327=>"010100100",
  62328=>"110101111",
  62329=>"011001111",
  62330=>"001001101",
  62331=>"001011111",
  62332=>"000110100",
  62333=>"100111010",
  62334=>"100011010",
  62335=>"100010000",
  62336=>"101011110",
  62337=>"011010101",
  62338=>"001010111",
  62339=>"010110010",
  62340=>"001011111",
  62341=>"011101001",
  62342=>"110101101",
  62343=>"000010111",
  62344=>"111010111",
  62345=>"101101111",
  62346=>"111101111",
  62347=>"101110000",
  62348=>"111010100",
  62349=>"011001101",
  62350=>"000011010",
  62351=>"011100000",
  62352=>"100101001",
  62353=>"010110000",
  62354=>"001001000",
  62355=>"101111100",
  62356=>"111110100",
  62357=>"010000011",
  62358=>"011000001",
  62359=>"100011110",
  62360=>"111111000",
  62361=>"001010000",
  62362=>"000010010",
  62363=>"110011011",
  62364=>"011000010",
  62365=>"100110000",
  62366=>"100000011",
  62367=>"010100100",
  62368=>"001000110",
  62369=>"010000101",
  62370=>"110110010",
  62371=>"101000011",
  62372=>"110110001",
  62373=>"110011101",
  62374=>"010101000",
  62375=>"000001101",
  62376=>"101000100",
  62377=>"000000001",
  62378=>"010011100",
  62379=>"101001110",
  62380=>"000001110",
  62381=>"001101111",
  62382=>"110010100",
  62383=>"101100010",
  62384=>"010010010",
  62385=>"110011111",
  62386=>"011000001",
  62387=>"111111001",
  62388=>"000100111",
  62389=>"011110001",
  62390=>"001010010",
  62391=>"111001100",
  62392=>"001100000",
  62393=>"000011011",
  62394=>"100010100",
  62395=>"001010000",
  62396=>"111000011",
  62397=>"111001001",
  62398=>"010001010",
  62399=>"111010100",
  62400=>"100100001",
  62401=>"010111010",
  62402=>"111100100",
  62403=>"001001010",
  62404=>"010000011",
  62405=>"001010111",
  62406=>"100000000",
  62407=>"010000000",
  62408=>"000000110",
  62409=>"011000011",
  62410=>"110011011",
  62411=>"100111100",
  62412=>"111101100",
  62413=>"010011101",
  62414=>"111100111",
  62415=>"001001000",
  62416=>"111001011",
  62417=>"001000110",
  62418=>"001110100",
  62419=>"100000001",
  62420=>"111111101",
  62421=>"001101101",
  62422=>"101011100",
  62423=>"000100010",
  62424=>"110100010",
  62425=>"000100010",
  62426=>"111111101",
  62427=>"000000101",
  62428=>"100111000",
  62429=>"111000110",
  62430=>"011010001",
  62431=>"011101000",
  62432=>"011111011",
  62433=>"000101111",
  62434=>"111100101",
  62435=>"111000111",
  62436=>"011101101",
  62437=>"111010001",
  62438=>"010011110",
  62439=>"011010101",
  62440=>"100100010",
  62441=>"110100100",
  62442=>"100111010",
  62443=>"101100010",
  62444=>"001011111",
  62445=>"100000011",
  62446=>"101000001",
  62447=>"000111010",
  62448=>"011010010",
  62449=>"010011111",
  62450=>"100110100",
  62451=>"110101100",
  62452=>"010011111",
  62453=>"000110000",
  62454=>"100110111",
  62455=>"110010010",
  62456=>"100001101",
  62457=>"111100001",
  62458=>"001010001",
  62459=>"101000011",
  62460=>"010101110",
  62461=>"100110100",
  62462=>"000000000",
  62463=>"111111111",
  62464=>"111100000",
  62465=>"100011011",
  62466=>"000001011",
  62467=>"111010110",
  62468=>"011100000",
  62469=>"011000000",
  62470=>"000000101",
  62471=>"011000101",
  62472=>"110100101",
  62473=>"011110010",
  62474=>"011010011",
  62475=>"000101011",
  62476=>"000111110",
  62477=>"010101111",
  62478=>"100101100",
  62479=>"101101001",
  62480=>"100000000",
  62481=>"011111001",
  62482=>"101000100",
  62483=>"001100101",
  62484=>"000001100",
  62485=>"001000011",
  62486=>"000101111",
  62487=>"110010111",
  62488=>"000111111",
  62489=>"100100111",
  62490=>"001111000",
  62491=>"010111110",
  62492=>"000000111",
  62493=>"010110010",
  62494=>"011001001",
  62495=>"100010000",
  62496=>"110011111",
  62497=>"101000011",
  62498=>"111011000",
  62499=>"110110000",
  62500=>"101111010",
  62501=>"011100010",
  62502=>"011000100",
  62503=>"000001110",
  62504=>"111101100",
  62505=>"001011100",
  62506=>"111110101",
  62507=>"110110101",
  62508=>"011000011",
  62509=>"011101111",
  62510=>"001000100",
  62511=>"011100011",
  62512=>"010011001",
  62513=>"101110111",
  62514=>"011111101",
  62515=>"000001101",
  62516=>"001000101",
  62517=>"111010100",
  62518=>"101000010",
  62519=>"001111101",
  62520=>"110111001",
  62521=>"001110000",
  62522=>"000110000",
  62523=>"010110000",
  62524=>"100000001",
  62525=>"000101011",
  62526=>"000110011",
  62527=>"111110101",
  62528=>"010101001",
  62529=>"001110100",
  62530=>"011001100",
  62531=>"111000110",
  62532=>"110011110",
  62533=>"011010011",
  62534=>"110000010",
  62535=>"111101001",
  62536=>"100111111",
  62537=>"000110001",
  62538=>"011001001",
  62539=>"101100101",
  62540=>"110110010",
  62541=>"111110001",
  62542=>"101100111",
  62543=>"011011011",
  62544=>"110010100",
  62545=>"111101101",
  62546=>"101111111",
  62547=>"000001000",
  62548=>"010011000",
  62549=>"010111101",
  62550=>"110001010",
  62551=>"011000011",
  62552=>"110010010",
  62553=>"000100011",
  62554=>"001001111",
  62555=>"010010100",
  62556=>"111111110",
  62557=>"110001000",
  62558=>"000100011",
  62559=>"001000000",
  62560=>"000001100",
  62561=>"111110111",
  62562=>"110111100",
  62563=>"000000101",
  62564=>"111011010",
  62565=>"011101101",
  62566=>"101100100",
  62567=>"000000000",
  62568=>"001100100",
  62569=>"101010010",
  62570=>"001000000",
  62571=>"100111010",
  62572=>"111001000",
  62573=>"000010111",
  62574=>"111000010",
  62575=>"000110100",
  62576=>"101100010",
  62577=>"000001000",
  62578=>"010010000",
  62579=>"000100001",
  62580=>"100011000",
  62581=>"101101111",
  62582=>"011111110",
  62583=>"011010110",
  62584=>"010110101",
  62585=>"010010010",
  62586=>"001111000",
  62587=>"010001100",
  62588=>"010101001",
  62589=>"000001111",
  62590=>"010110110",
  62591=>"111000000",
  62592=>"101000000",
  62593=>"001111110",
  62594=>"100011000",
  62595=>"101001100",
  62596=>"110000011",
  62597=>"000001111",
  62598=>"001001011",
  62599=>"010010110",
  62600=>"011000101",
  62601=>"000100000",
  62602=>"011101010",
  62603=>"111011000",
  62604=>"111011101",
  62605=>"010100010",
  62606=>"001001000",
  62607=>"010000111",
  62608=>"111000000",
  62609=>"101101101",
  62610=>"010111100",
  62611=>"110101111",
  62612=>"010101001",
  62613=>"110000010",
  62614=>"011100101",
  62615=>"110011000",
  62616=>"101101001",
  62617=>"110101110",
  62618=>"010100110",
  62619=>"110011010",
  62620=>"111101111",
  62621=>"111101011",
  62622=>"011011111",
  62623=>"111101111",
  62624=>"001101011",
  62625=>"101000011",
  62626=>"010111111",
  62627=>"000001110",
  62628=>"100010101",
  62629=>"101110101",
  62630=>"110110000",
  62631=>"100000011",
  62632=>"010011110",
  62633=>"000101011",
  62634=>"111010111",
  62635=>"111100111",
  62636=>"101100100",
  62637=>"110101001",
  62638=>"111110001",
  62639=>"011011010",
  62640=>"010111100",
  62641=>"010001110",
  62642=>"001000110",
  62643=>"111100011",
  62644=>"001000111",
  62645=>"000110000",
  62646=>"101111101",
  62647=>"001010110",
  62648=>"110001000",
  62649=>"101101100",
  62650=>"001000100",
  62651=>"010111110",
  62652=>"010101010",
  62653=>"010010001",
  62654=>"001111101",
  62655=>"110001001",
  62656=>"011010000",
  62657=>"110011101",
  62658=>"001001000",
  62659=>"010011011",
  62660=>"010111010",
  62661=>"101100110",
  62662=>"110100101",
  62663=>"101010111",
  62664=>"000111101",
  62665=>"000110000",
  62666=>"011001111",
  62667=>"111111011",
  62668=>"100101011",
  62669=>"100011110",
  62670=>"000001001",
  62671=>"001100100",
  62672=>"110101100",
  62673=>"110001100",
  62674=>"000000000",
  62675=>"000100010",
  62676=>"101001000",
  62677=>"110101011",
  62678=>"010001101",
  62679=>"001101101",
  62680=>"010111100",
  62681=>"011001011",
  62682=>"101100001",
  62683=>"011011001",
  62684=>"010011101",
  62685=>"111000001",
  62686=>"001101101",
  62687=>"011011011",
  62688=>"011110011",
  62689=>"111101010",
  62690=>"101100001",
  62691=>"111111111",
  62692=>"111110001",
  62693=>"011010101",
  62694=>"101100111",
  62695=>"101110001",
  62696=>"111101010",
  62697=>"000110010",
  62698=>"110010111",
  62699=>"000110110",
  62700=>"011001011",
  62701=>"100111001",
  62702=>"000100100",
  62703=>"011010110",
  62704=>"000110010",
  62705=>"000111010",
  62706=>"000111110",
  62707=>"001111100",
  62708=>"011111010",
  62709=>"111100001",
  62710=>"111111011",
  62711=>"011111110",
  62712=>"100000100",
  62713=>"001100010",
  62714=>"101001011",
  62715=>"100011010",
  62716=>"011010110",
  62717=>"000110000",
  62718=>"010100100",
  62719=>"000011001",
  62720=>"010101011",
  62721=>"101001000",
  62722=>"010000110",
  62723=>"010001111",
  62724=>"010101000",
  62725=>"000010100",
  62726=>"010001011",
  62727=>"101100000",
  62728=>"001100001",
  62729=>"000110111",
  62730=>"110110111",
  62731=>"111000110",
  62732=>"010101010",
  62733=>"011110100",
  62734=>"011101111",
  62735=>"001001001",
  62736=>"101111100",
  62737=>"100100000",
  62738=>"000110111",
  62739=>"000011010",
  62740=>"101101110",
  62741=>"100101110",
  62742=>"000110111",
  62743=>"010100001",
  62744=>"111010001",
  62745=>"000000001",
  62746=>"010000111",
  62747=>"100000101",
  62748=>"010110101",
  62749=>"010101000",
  62750=>"000110011",
  62751=>"011111010",
  62752=>"000111111",
  62753=>"110110010",
  62754=>"010011111",
  62755=>"110111101",
  62756=>"101111110",
  62757=>"010000001",
  62758=>"000000010",
  62759=>"111011011",
  62760=>"100011001",
  62761=>"010000101",
  62762=>"111111010",
  62763=>"011111111",
  62764=>"000000010",
  62765=>"111001100",
  62766=>"010010111",
  62767=>"001111010",
  62768=>"100011100",
  62769=>"010110101",
  62770=>"110100111",
  62771=>"001001001",
  62772=>"001111001",
  62773=>"001000111",
  62774=>"100101011",
  62775=>"000000000",
  62776=>"111010001",
  62777=>"011101000",
  62778=>"101110101",
  62779=>"100001001",
  62780=>"100001100",
  62781=>"011110100",
  62782=>"101101011",
  62783=>"100111101",
  62784=>"010100011",
  62785=>"000101111",
  62786=>"111111111",
  62787=>"001100001",
  62788=>"010011100",
  62789=>"000010100",
  62790=>"101000101",
  62791=>"000100010",
  62792=>"101001001",
  62793=>"000010001",
  62794=>"011011110",
  62795=>"001001010",
  62796=>"011000011",
  62797=>"011101101",
  62798=>"000101100",
  62799=>"101011111",
  62800=>"111100101",
  62801=>"111011010",
  62802=>"101100001",
  62803=>"000010111",
  62804=>"000000001",
  62805=>"100011111",
  62806=>"100010000",
  62807=>"111110100",
  62808=>"110111110",
  62809=>"010111100",
  62810=>"100000111",
  62811=>"000000111",
  62812=>"010110101",
  62813=>"001000100",
  62814=>"100101010",
  62815=>"001110000",
  62816=>"011011101",
  62817=>"000100110",
  62818=>"000001000",
  62819=>"011110010",
  62820=>"111101011",
  62821=>"101011010",
  62822=>"100110110",
  62823=>"110100000",
  62824=>"011010111",
  62825=>"111010011",
  62826=>"000000101",
  62827=>"000101101",
  62828=>"011001011",
  62829=>"001001110",
  62830=>"001011111",
  62831=>"011010111",
  62832=>"000100111",
  62833=>"010100010",
  62834=>"110111011",
  62835=>"101011011",
  62836=>"110001011",
  62837=>"110111101",
  62838=>"000001101",
  62839=>"100001001",
  62840=>"000000111",
  62841=>"010111011",
  62842=>"110000101",
  62843=>"010100001",
  62844=>"001011101",
  62845=>"011100100",
  62846=>"110000010",
  62847=>"001100111",
  62848=>"101111001",
  62849=>"101011001",
  62850=>"101001100",
  62851=>"011101100",
  62852=>"011111111",
  62853=>"001000001",
  62854=>"100001110",
  62855=>"100010101",
  62856=>"101000110",
  62857=>"111111110",
  62858=>"011111010",
  62859=>"010011100",
  62860=>"101001110",
  62861=>"100111110",
  62862=>"010000000",
  62863=>"100101100",
  62864=>"100001011",
  62865=>"010110000",
  62866=>"101001001",
  62867=>"100011011",
  62868=>"101000000",
  62869=>"000101010",
  62870=>"000100100",
  62871=>"101111000",
  62872=>"110101011",
  62873=>"101101001",
  62874=>"111110000",
  62875=>"010001111",
  62876=>"111011010",
  62877=>"101011111",
  62878=>"100111010",
  62879=>"101111101",
  62880=>"111101100",
  62881=>"000011010",
  62882=>"100100111",
  62883=>"110001110",
  62884=>"001000110",
  62885=>"010000011",
  62886=>"111100100",
  62887=>"010110000",
  62888=>"000100000",
  62889=>"111111001",
  62890=>"011011000",
  62891=>"111011011",
  62892=>"100110111",
  62893=>"000010111",
  62894=>"001010100",
  62895=>"111010111",
  62896=>"110011000",
  62897=>"010000000",
  62898=>"001010001",
  62899=>"010001101",
  62900=>"011111110",
  62901=>"011111001",
  62902=>"110100000",
  62903=>"001111100",
  62904=>"111000110",
  62905=>"001000111",
  62906=>"101011110",
  62907=>"000000100",
  62908=>"000011111",
  62909=>"010011011",
  62910=>"100111001",
  62911=>"010100000",
  62912=>"101101100",
  62913=>"111010110",
  62914=>"010000010",
  62915=>"100110101",
  62916=>"000000010",
  62917=>"100111001",
  62918=>"000001001",
  62919=>"100011010",
  62920=>"010111111",
  62921=>"010010111",
  62922=>"101000011",
  62923=>"010000011",
  62924=>"001110001",
  62925=>"011100110",
  62926=>"000000010",
  62927=>"110100010",
  62928=>"001110011",
  62929=>"010110011",
  62930=>"000110110",
  62931=>"010000101",
  62932=>"100111000",
  62933=>"110010000",
  62934=>"100101001",
  62935=>"000000110",
  62936=>"101010000",
  62937=>"111001100",
  62938=>"001011001",
  62939=>"101001000",
  62940=>"111110110",
  62941=>"110100000",
  62942=>"111011011",
  62943=>"110110010",
  62944=>"000000101",
  62945=>"110001100",
  62946=>"010011111",
  62947=>"111110000",
  62948=>"110111100",
  62949=>"111101100",
  62950=>"100000000",
  62951=>"010111110",
  62952=>"111101001",
  62953=>"000011101",
  62954=>"101100010",
  62955=>"100000111",
  62956=>"100000110",
  62957=>"000010101",
  62958=>"110001001",
  62959=>"001011000",
  62960=>"010101101",
  62961=>"100001110",
  62962=>"001101001",
  62963=>"111101110",
  62964=>"001000110",
  62965=>"001001100",
  62966=>"111100110",
  62967=>"001110000",
  62968=>"010101101",
  62969=>"101110011",
  62970=>"000111111",
  62971=>"000111001",
  62972=>"110110110",
  62973=>"001110001",
  62974=>"011011010",
  62975=>"110000100",
  62976=>"010010011",
  62977=>"000010110",
  62978=>"111011110",
  62979=>"000010001",
  62980=>"001011001",
  62981=>"100110100",
  62982=>"010111110",
  62983=>"000001111",
  62984=>"001111000",
  62985=>"101101110",
  62986=>"001110011",
  62987=>"010101101",
  62988=>"000111011",
  62989=>"111101001",
  62990=>"000110000",
  62991=>"010101111",
  62992=>"100100010",
  62993=>"101101100",
  62994=>"111011001",
  62995=>"001111000",
  62996=>"000100111",
  62997=>"111001100",
  62998=>"111010011",
  62999=>"010000110",
  63000=>"110111010",
  63001=>"000000010",
  63002=>"100000000",
  63003=>"000101110",
  63004=>"111100011",
  63005=>"010100111",
  63006=>"110001001",
  63007=>"110010100",
  63008=>"001101010",
  63009=>"111100111",
  63010=>"011011110",
  63011=>"111001000",
  63012=>"111001110",
  63013=>"001101100",
  63014=>"000111111",
  63015=>"000000001",
  63016=>"111100101",
  63017=>"010000111",
  63018=>"011011110",
  63019=>"110000000",
  63020=>"000100100",
  63021=>"000100100",
  63022=>"110110001",
  63023=>"000000000",
  63024=>"110110101",
  63025=>"000100001",
  63026=>"101100101",
  63027=>"010100001",
  63028=>"110000111",
  63029=>"000111011",
  63030=>"100010011",
  63031=>"001011110",
  63032=>"001010010",
  63033=>"111010110",
  63034=>"101101011",
  63035=>"000001011",
  63036=>"000110001",
  63037=>"001101001",
  63038=>"000101000",
  63039=>"110000101",
  63040=>"101111101",
  63041=>"110010011",
  63042=>"110010001",
  63043=>"011000011",
  63044=>"110101101",
  63045=>"000100000",
  63046=>"000101100",
  63047=>"110111010",
  63048=>"110111011",
  63049=>"111111010",
  63050=>"111010111",
  63051=>"001100010",
  63052=>"101001010",
  63053=>"100101010",
  63054=>"001011100",
  63055=>"100011101",
  63056=>"000000010",
  63057=>"101110011",
  63058=>"001000100",
  63059=>"000011001",
  63060=>"110110100",
  63061=>"111100111",
  63062=>"110001000",
  63063=>"111111000",
  63064=>"110010010",
  63065=>"000010111",
  63066=>"010101001",
  63067=>"001000100",
  63068=>"000101000",
  63069=>"111010011",
  63070=>"000101110",
  63071=>"000100100",
  63072=>"101010100",
  63073=>"011011011",
  63074=>"000011100",
  63075=>"110001100",
  63076=>"101010100",
  63077=>"100110010",
  63078=>"111000011",
  63079=>"000001100",
  63080=>"000000010",
  63081=>"111010101",
  63082=>"011011010",
  63083=>"110111011",
  63084=>"100110110",
  63085=>"110001100",
  63086=>"000000101",
  63087=>"111011111",
  63088=>"000110110",
  63089=>"000010000",
  63090=>"001011001",
  63091=>"011100011",
  63092=>"010011010",
  63093=>"000110011",
  63094=>"011011111",
  63095=>"010000011",
  63096=>"111001111",
  63097=>"100110110",
  63098=>"111111001",
  63099=>"001011011",
  63100=>"000010111",
  63101=>"001010000",
  63102=>"000100011",
  63103=>"001100111",
  63104=>"110011000",
  63105=>"110110001",
  63106=>"101101110",
  63107=>"001000100",
  63108=>"001010010",
  63109=>"101011100",
  63110=>"111101110",
  63111=>"000000010",
  63112=>"110100100",
  63113=>"000000101",
  63114=>"011000110",
  63115=>"111010010",
  63116=>"111101011",
  63117=>"000110100",
  63118=>"111111111",
  63119=>"100011111",
  63120=>"001010001",
  63121=>"010001000",
  63122=>"010100000",
  63123=>"010010111",
  63124=>"111111011",
  63125=>"111010110",
  63126=>"001101110",
  63127=>"001101111",
  63128=>"010111101",
  63129=>"010110011",
  63130=>"010011101",
  63131=>"001001001",
  63132=>"001101000",
  63133=>"111110000",
  63134=>"010001100",
  63135=>"111011110",
  63136=>"010110111",
  63137=>"001000101",
  63138=>"100111000",
  63139=>"000000110",
  63140=>"010010001",
  63141=>"100000010",
  63142=>"000100001",
  63143=>"110001110",
  63144=>"000111101",
  63145=>"111110111",
  63146=>"011001110",
  63147=>"010010110",
  63148=>"111111100",
  63149=>"101100010",
  63150=>"000111011",
  63151=>"110110110",
  63152=>"000100000",
  63153=>"100010001",
  63154=>"011100110",
  63155=>"000110111",
  63156=>"000010000",
  63157=>"111110111",
  63158=>"110100010",
  63159=>"000110010",
  63160=>"100101010",
  63161=>"100111010",
  63162=>"111110111",
  63163=>"001010010",
  63164=>"100010010",
  63165=>"011000000",
  63166=>"100100100",
  63167=>"001111001",
  63168=>"101111011",
  63169=>"110000010",
  63170=>"100100000",
  63171=>"111001010",
  63172=>"100011110",
  63173=>"101101010",
  63174=>"101110011",
  63175=>"000101110",
  63176=>"100111011",
  63177=>"010011001",
  63178=>"111010110",
  63179=>"101100111",
  63180=>"010100011",
  63181=>"110010000",
  63182=>"101010000",
  63183=>"000100010",
  63184=>"011011101",
  63185=>"111101111",
  63186=>"111001000",
  63187=>"001001010",
  63188=>"000001100",
  63189=>"111011111",
  63190=>"111110101",
  63191=>"000101000",
  63192=>"000111000",
  63193=>"100111011",
  63194=>"000000100",
  63195=>"000110100",
  63196=>"010000010",
  63197=>"000011111",
  63198=>"001110010",
  63199=>"000101111",
  63200=>"001111111",
  63201=>"000010000",
  63202=>"101110101",
  63203=>"101111001",
  63204=>"101010101",
  63205=>"010011000",
  63206=>"101110000",
  63207=>"000101011",
  63208=>"101000110",
  63209=>"001110111",
  63210=>"110000001",
  63211=>"011111100",
  63212=>"010101011",
  63213=>"010010111",
  63214=>"101000100",
  63215=>"000011001",
  63216=>"011011100",
  63217=>"111011000",
  63218=>"111101000",
  63219=>"010111111",
  63220=>"101001111",
  63221=>"111110000",
  63222=>"011000111",
  63223=>"101100000",
  63224=>"000110011",
  63225=>"010111000",
  63226=>"000011001",
  63227=>"010010100",
  63228=>"011001011",
  63229=>"000000110",
  63230=>"010111001",
  63231=>"000111010",
  63232=>"111011100",
  63233=>"011000110",
  63234=>"110101100",
  63235=>"000000000",
  63236=>"000000010",
  63237=>"000101100",
  63238=>"010000000",
  63239=>"111011111",
  63240=>"010001010",
  63241=>"010110001",
  63242=>"001100000",
  63243=>"010110000",
  63244=>"011100100",
  63245=>"001101100",
  63246=>"011110000",
  63247=>"000010101",
  63248=>"111101010",
  63249=>"111001110",
  63250=>"011010101",
  63251=>"001101011",
  63252=>"011111011",
  63253=>"110110000",
  63254=>"100000011",
  63255=>"011011011",
  63256=>"011010110",
  63257=>"011101011",
  63258=>"000001000",
  63259=>"000100000",
  63260=>"101001110",
  63261=>"010010100",
  63262=>"111011111",
  63263=>"000100111",
  63264=>"101101100",
  63265=>"000100101",
  63266=>"111100100",
  63267=>"111101000",
  63268=>"011000110",
  63269=>"100111010",
  63270=>"000001010",
  63271=>"100000110",
  63272=>"001001101",
  63273=>"110110110",
  63274=>"010111110",
  63275=>"111110101",
  63276=>"111000110",
  63277=>"000000110",
  63278=>"110111111",
  63279=>"001011001",
  63280=>"011110111",
  63281=>"010100001",
  63282=>"010000000",
  63283=>"001101111",
  63284=>"010101000",
  63285=>"100000110",
  63286=>"000001001",
  63287=>"101101111",
  63288=>"111101010",
  63289=>"011000110",
  63290=>"001001010",
  63291=>"111100101",
  63292=>"101110000",
  63293=>"000000100",
  63294=>"100000110",
  63295=>"011010011",
  63296=>"011111011",
  63297=>"001001000",
  63298=>"101100110",
  63299=>"111011110",
  63300=>"111001111",
  63301=>"110101100",
  63302=>"100011111",
  63303=>"001010000",
  63304=>"100101100",
  63305=>"110011011",
  63306=>"111111001",
  63307=>"010100110",
  63308=>"111110010",
  63309=>"111110010",
  63310=>"011100001",
  63311=>"010110010",
  63312=>"101011011",
  63313=>"010010110",
  63314=>"000000001",
  63315=>"101111100",
  63316=>"000101001",
  63317=>"001001010",
  63318=>"111101111",
  63319=>"001111110",
  63320=>"000000111",
  63321=>"100110001",
  63322=>"110011100",
  63323=>"100001111",
  63324=>"011111010",
  63325=>"111000110",
  63326=>"100100001",
  63327=>"110100010",
  63328=>"001000111",
  63329=>"011011101",
  63330=>"101101001",
  63331=>"011011010",
  63332=>"111110100",
  63333=>"000101101",
  63334=>"010101101",
  63335=>"000010010",
  63336=>"010001000",
  63337=>"011010010",
  63338=>"001110011",
  63339=>"111110110",
  63340=>"101110100",
  63341=>"100111011",
  63342=>"000001100",
  63343=>"100011100",
  63344=>"010110110",
  63345=>"101000110",
  63346=>"011101000",
  63347=>"101001100",
  63348=>"100110101",
  63349=>"101111111",
  63350=>"101000101",
  63351=>"101110111",
  63352=>"110010110",
  63353=>"001001000",
  63354=>"000110100",
  63355=>"100110000",
  63356=>"101111010",
  63357=>"110001110",
  63358=>"000100000",
  63359=>"000010011",
  63360=>"100000010",
  63361=>"110000111",
  63362=>"101001101",
  63363=>"111111011",
  63364=>"010110010",
  63365=>"010100010",
  63366=>"111000011",
  63367=>"101100000",
  63368=>"110110111",
  63369=>"100011110",
  63370=>"100000001",
  63371=>"111111011",
  63372=>"000100000",
  63373=>"010001010",
  63374=>"011000001",
  63375=>"100011011",
  63376=>"101011010",
  63377=>"001111010",
  63378=>"010111000",
  63379=>"010111111",
  63380=>"001101111",
  63381=>"010000101",
  63382=>"100110111",
  63383=>"011001010",
  63384=>"100110000",
  63385=>"000111111",
  63386=>"000111111",
  63387=>"000101110",
  63388=>"111001010",
  63389=>"011110110",
  63390=>"100011101",
  63391=>"010110010",
  63392=>"000011000",
  63393=>"110100011",
  63394=>"100011100",
  63395=>"111111111",
  63396=>"110100001",
  63397=>"000000010",
  63398=>"011110000",
  63399=>"011100101",
  63400=>"100110011",
  63401=>"001101000",
  63402=>"010000000",
  63403=>"110110110",
  63404=>"001100110",
  63405=>"101101010",
  63406=>"010010100",
  63407=>"000001011",
  63408=>"001111000",
  63409=>"010011101",
  63410=>"110101000",
  63411=>"001011101",
  63412=>"110001001",
  63413=>"011111010",
  63414=>"100011110",
  63415=>"111010010",
  63416=>"101101101",
  63417=>"101101011",
  63418=>"100010001",
  63419=>"101011001",
  63420=>"100111011",
  63421=>"000100000",
  63422=>"111001000",
  63423=>"001000101",
  63424=>"100111010",
  63425=>"000011110",
  63426=>"011110100",
  63427=>"111111011",
  63428=>"000100101",
  63429=>"011001001",
  63430=>"101111011",
  63431=>"010111000",
  63432=>"111000011",
  63433=>"001011010",
  63434=>"110100000",
  63435=>"010000111",
  63436=>"111001111",
  63437=>"000000101",
  63438=>"100101010",
  63439=>"101001001",
  63440=>"000000011",
  63441=>"000010111",
  63442=>"010011011",
  63443=>"011100000",
  63444=>"011011000",
  63445=>"011000010",
  63446=>"000100101",
  63447=>"101010110",
  63448=>"110100101",
  63449=>"000100011",
  63450=>"010100010",
  63451=>"000101001",
  63452=>"010100001",
  63453=>"000100001",
  63454=>"011100000",
  63455=>"101110011",
  63456=>"001010111",
  63457=>"100101000",
  63458=>"100011110",
  63459=>"011101101",
  63460=>"010111111",
  63461=>"111001111",
  63462=>"000101001",
  63463=>"000100111",
  63464=>"010111011",
  63465=>"111111111",
  63466=>"001001110",
  63467=>"010011000",
  63468=>"011000010",
  63469=>"000111111",
  63470=>"100111101",
  63471=>"111010100",
  63472=>"010111010",
  63473=>"100001110",
  63474=>"011010110",
  63475=>"010110101",
  63476=>"001000000",
  63477=>"110000101",
  63478=>"100111000",
  63479=>"011000111",
  63480=>"111010000",
  63481=>"011000100",
  63482=>"110010010",
  63483=>"001101001",
  63484=>"101001000",
  63485=>"110101010",
  63486=>"000100110",
  63487=>"111110110",
  63488=>"001010100",
  63489=>"101010010",
  63490=>"110001100",
  63491=>"011110101",
  63492=>"010000001",
  63493=>"111110011",
  63494=>"001011000",
  63495=>"101100000",
  63496=>"001011110",
  63497=>"001001000",
  63498=>"111011100",
  63499=>"010100000",
  63500=>"101000010",
  63501=>"101010001",
  63502=>"100110100",
  63503=>"001001011",
  63504=>"000110000",
  63505=>"100110001",
  63506=>"001100010",
  63507=>"111000001",
  63508=>"110110110",
  63509=>"110100100",
  63510=>"101100001",
  63511=>"001001100",
  63512=>"111001100",
  63513=>"010000101",
  63514=>"100101110",
  63515=>"001000011",
  63516=>"011000100",
  63517=>"001010000",
  63518=>"010011001",
  63519=>"000100010",
  63520=>"001000111",
  63521=>"001110111",
  63522=>"000001110",
  63523=>"101010111",
  63524=>"100101001",
  63525=>"110001001",
  63526=>"100010100",
  63527=>"010111110",
  63528=>"101000111",
  63529=>"000100000",
  63530=>"110000001",
  63531=>"011101000",
  63532=>"010010010",
  63533=>"010010100",
  63534=>"100001000",
  63535=>"111100011",
  63536=>"100111101",
  63537=>"001110110",
  63538=>"101010110",
  63539=>"111001010",
  63540=>"011011101",
  63541=>"100110111",
  63542=>"111010110",
  63543=>"100011111",
  63544=>"101011101",
  63545=>"001000101",
  63546=>"000001110",
  63547=>"001000100",
  63548=>"101001110",
  63549=>"000110001",
  63550=>"101110111",
  63551=>"110010010",
  63552=>"011010001",
  63553=>"000000110",
  63554=>"000000010",
  63555=>"110110111",
  63556=>"000011011",
  63557=>"111100001",
  63558=>"011100000",
  63559=>"000100001",
  63560=>"111110001",
  63561=>"110001110",
  63562=>"000000001",
  63563=>"100001010",
  63564=>"001001011",
  63565=>"100110001",
  63566=>"011010000",
  63567=>"000000001",
  63568=>"010001101",
  63569=>"000010101",
  63570=>"101001010",
  63571=>"101011110",
  63572=>"110101101",
  63573=>"111010010",
  63574=>"110011010",
  63575=>"101101101",
  63576=>"001101110",
  63577=>"111000010",
  63578=>"100011010",
  63579=>"111010010",
  63580=>"010001100",
  63581=>"101001011",
  63582=>"111010110",
  63583=>"100101111",
  63584=>"011110011",
  63585=>"010010011",
  63586=>"101001000",
  63587=>"011000100",
  63588=>"011111000",
  63589=>"010101110",
  63590=>"011000001",
  63591=>"100101111",
  63592=>"001111001",
  63593=>"010000011",
  63594=>"010000001",
  63595=>"100101100",
  63596=>"001101111",
  63597=>"100101111",
  63598=>"111010111",
  63599=>"000000101",
  63600=>"011011011",
  63601=>"111110101",
  63602=>"001111100",
  63603=>"011010001",
  63604=>"011111110",
  63605=>"111110010",
  63606=>"000011101",
  63607=>"101010100",
  63608=>"010111111",
  63609=>"100001001",
  63610=>"000100001",
  63611=>"111001001",
  63612=>"011111111",
  63613=>"110001011",
  63614=>"101010011",
  63615=>"101100001",
  63616=>"111111101",
  63617=>"101111011",
  63618=>"101111111",
  63619=>"010001111",
  63620=>"101000111",
  63621=>"001111001",
  63622=>"000000001",
  63623=>"001001000",
  63624=>"001010001",
  63625=>"011111111",
  63626=>"101100010",
  63627=>"011001010",
  63628=>"011010110",
  63629=>"101000110",
  63630=>"001001100",
  63631=>"111010010",
  63632=>"011010100",
  63633=>"010100011",
  63634=>"111001111",
  63635=>"010010000",
  63636=>"000010100",
  63637=>"111001000",
  63638=>"001000010",
  63639=>"100111100",
  63640=>"011001011",
  63641=>"010000100",
  63642=>"110011100",
  63643=>"001100111",
  63644=>"010011010",
  63645=>"110110100",
  63646=>"001001000",
  63647=>"011001001",
  63648=>"111110000",
  63649=>"011110011",
  63650=>"011000110",
  63651=>"001111000",
  63652=>"111110100",
  63653=>"011101011",
  63654=>"011101011",
  63655=>"010000000",
  63656=>"001010110",
  63657=>"001011001",
  63658=>"010100111",
  63659=>"001010000",
  63660=>"001111000",
  63661=>"001100001",
  63662=>"110100111",
  63663=>"110000111",
  63664=>"101011100",
  63665=>"010010101",
  63666=>"110110101",
  63667=>"111101011",
  63668=>"000011110",
  63669=>"000100010",
  63670=>"101000110",
  63671=>"001000000",
  63672=>"010101011",
  63673=>"101011001",
  63674=>"101111110",
  63675=>"000010110",
  63676=>"010110000",
  63677=>"101011010",
  63678=>"000000110",
  63679=>"101000000",
  63680=>"010100000",
  63681=>"010111100",
  63682=>"110111110",
  63683=>"111100001",
  63684=>"110111010",
  63685=>"000100111",
  63686=>"001100001",
  63687=>"101100110",
  63688=>"000111011",
  63689=>"111111011",
  63690=>"010000001",
  63691=>"011011010",
  63692=>"011010100",
  63693=>"001101011",
  63694=>"111000111",
  63695=>"010111110",
  63696=>"110001000",
  63697=>"101011111",
  63698=>"100100011",
  63699=>"100100000",
  63700=>"010000011",
  63701=>"111010100",
  63702=>"111010111",
  63703=>"010100110",
  63704=>"110101101",
  63705=>"111111101",
  63706=>"110100111",
  63707=>"011010010",
  63708=>"001111000",
  63709=>"000110100",
  63710=>"110011101",
  63711=>"001101111",
  63712=>"000100000",
  63713=>"010011111",
  63714=>"011001000",
  63715=>"010100111",
  63716=>"011001100",
  63717=>"010101011",
  63718=>"001101101",
  63719=>"000100100",
  63720=>"001111110",
  63721=>"100010010",
  63722=>"100101101",
  63723=>"001101001",
  63724=>"100110100",
  63725=>"001000101",
  63726=>"101001011",
  63727=>"111110111",
  63728=>"000000000",
  63729=>"111000001",
  63730=>"010111111",
  63731=>"100100110",
  63732=>"110001100",
  63733=>"100001000",
  63734=>"011101110",
  63735=>"101101111",
  63736=>"110111010",
  63737=>"010011010",
  63738=>"011000011",
  63739=>"100101100",
  63740=>"000101011",
  63741=>"100101100",
  63742=>"011100011",
  63743=>"111001101",
  63744=>"100010110",
  63745=>"010111010",
  63746=>"111011011",
  63747=>"001100011",
  63748=>"101111001",
  63749=>"010010001",
  63750=>"011011100",
  63751=>"001111100",
  63752=>"110000001",
  63753=>"110011111",
  63754=>"111010110",
  63755=>"111000001",
  63756=>"011001100",
  63757=>"100000000",
  63758=>"000011010",
  63759=>"111010010",
  63760=>"111001100",
  63761=>"000010101",
  63762=>"111100011",
  63763=>"101000110",
  63764=>"000111111",
  63765=>"001000011",
  63766=>"000100000",
  63767=>"111100011",
  63768=>"111010010",
  63769=>"110000111",
  63770=>"101101111",
  63771=>"111010101",
  63772=>"111101001",
  63773=>"110001000",
  63774=>"001011101",
  63775=>"111100000",
  63776=>"000100001",
  63777=>"010011000",
  63778=>"011100100",
  63779=>"011111011",
  63780=>"101100010",
  63781=>"111010000",
  63782=>"101000011",
  63783=>"101011010",
  63784=>"010101001",
  63785=>"000011101",
  63786=>"001011101",
  63787=>"110010111",
  63788=>"100000100",
  63789=>"110010010",
  63790=>"011101011",
  63791=>"011111110",
  63792=>"100101000",
  63793=>"000010000",
  63794=>"010100101",
  63795=>"010011010",
  63796=>"001100001",
  63797=>"000000000",
  63798=>"110110100",
  63799=>"110100111",
  63800=>"111111110",
  63801=>"100011111",
  63802=>"100001111",
  63803=>"001001111",
  63804=>"111110010",
  63805=>"111101011",
  63806=>"001010001",
  63807=>"111010011",
  63808=>"011010111",
  63809=>"001001011",
  63810=>"001001100",
  63811=>"101000001",
  63812=>"101100000",
  63813=>"001110000",
  63814=>"010111001",
  63815=>"110010001",
  63816=>"011110110",
  63817=>"110000001",
  63818=>"111100101",
  63819=>"100111111",
  63820=>"110111010",
  63821=>"000100110",
  63822=>"011011001",
  63823=>"110000011",
  63824=>"000001101",
  63825=>"111111111",
  63826=>"000011000",
  63827=>"110100011",
  63828=>"100100001",
  63829=>"011101101",
  63830=>"110001011",
  63831=>"110101001",
  63832=>"000001011",
  63833=>"111110100",
  63834=>"000010101",
  63835=>"110011101",
  63836=>"001011011",
  63837=>"000101010",
  63838=>"001110000",
  63839=>"110110110",
  63840=>"001110101",
  63841=>"001010110",
  63842=>"000000101",
  63843=>"111001000",
  63844=>"010101100",
  63845=>"101110000",
  63846=>"001000011",
  63847=>"001010101",
  63848=>"010010010",
  63849=>"110101001",
  63850=>"111111110",
  63851=>"101111100",
  63852=>"011001111",
  63853=>"000001111",
  63854=>"101100111",
  63855=>"000011001",
  63856=>"001001011",
  63857=>"001101000",
  63858=>"010001101",
  63859=>"110100000",
  63860=>"010101011",
  63861=>"001110100",
  63862=>"010001010",
  63863=>"001101101",
  63864=>"011001011",
  63865=>"101110011",
  63866=>"101111100",
  63867=>"000110000",
  63868=>"001111010",
  63869=>"110000101",
  63870=>"110011111",
  63871=>"111101101",
  63872=>"000101100",
  63873=>"000001001",
  63874=>"010011110",
  63875=>"101111001",
  63876=>"100000011",
  63877=>"110000001",
  63878=>"100101000",
  63879=>"000010011",
  63880=>"100100110",
  63881=>"111101010",
  63882=>"111101011",
  63883=>"010100000",
  63884=>"011011001",
  63885=>"000000100",
  63886=>"111111110",
  63887=>"010100111",
  63888=>"010011100",
  63889=>"001001010",
  63890=>"011001011",
  63891=>"110101011",
  63892=>"000110011",
  63893=>"000100110",
  63894=>"000101101",
  63895=>"110111000",
  63896=>"110001100",
  63897=>"100111001",
  63898=>"000111011",
  63899=>"000110100",
  63900=>"110101000",
  63901=>"001101101",
  63902=>"110101010",
  63903=>"010110010",
  63904=>"101101111",
  63905=>"110010100",
  63906=>"011010110",
  63907=>"001100000",
  63908=>"110000101",
  63909=>"100101111",
  63910=>"111111101",
  63911=>"001001011",
  63912=>"000010010",
  63913=>"011000111",
  63914=>"001000001",
  63915=>"100110111",
  63916=>"011100000",
  63917=>"101010001",
  63918=>"101100111",
  63919=>"011100110",
  63920=>"100101110",
  63921=>"101110000",
  63922=>"110001011",
  63923=>"001100010",
  63924=>"000110111",
  63925=>"100110000",
  63926=>"101100111",
  63927=>"000000011",
  63928=>"000010111",
  63929=>"111111110",
  63930=>"001111110",
  63931=>"001110110",
  63932=>"100011000",
  63933=>"010001000",
  63934=>"000000001",
  63935=>"111111001",
  63936=>"110111110",
  63937=>"101111110",
  63938=>"010000111",
  63939=>"011001010",
  63940=>"000010100",
  63941=>"110110101",
  63942=>"110001100",
  63943=>"110101101",
  63944=>"100111101",
  63945=>"101110001",
  63946=>"110000110",
  63947=>"001101110",
  63948=>"000101101",
  63949=>"000001001",
  63950=>"111101010",
  63951=>"001010010",
  63952=>"010111111",
  63953=>"000010100",
  63954=>"111110100",
  63955=>"111111111",
  63956=>"100110111",
  63957=>"110101011",
  63958=>"101100101",
  63959=>"010100101",
  63960=>"111110001",
  63961=>"011101100",
  63962=>"001001000",
  63963=>"110111100",
  63964=>"011100000",
  63965=>"000101000",
  63966=>"010010011",
  63967=>"100101001",
  63968=>"101111000",
  63969=>"111111000",
  63970=>"001100001",
  63971=>"011100101",
  63972=>"000100000",
  63973=>"100000001",
  63974=>"110011110",
  63975=>"000111001",
  63976=>"011010100",
  63977=>"101100111",
  63978=>"100101110",
  63979=>"001001000",
  63980=>"001100110",
  63981=>"001111101",
  63982=>"101111101",
  63983=>"101100000",
  63984=>"011110000",
  63985=>"100111100",
  63986=>"000111101",
  63987=>"101110100",
  63988=>"001010101",
  63989=>"000111000",
  63990=>"100111111",
  63991=>"101000111",
  63992=>"000110100",
  63993=>"110010100",
  63994=>"001001110",
  63995=>"010111011",
  63996=>"010100001",
  63997=>"101111000",
  63998=>"000110110",
  63999=>"110001110",
  64000=>"011001001",
  64001=>"110011110",
  64002=>"101011011",
  64003=>"001001111",
  64004=>"110011011",
  64005=>"000000010",
  64006=>"110011000",
  64007=>"101101100",
  64008=>"110011000",
  64009=>"101011101",
  64010=>"010100000",
  64011=>"011111111",
  64012=>"111110100",
  64013=>"100010000",
  64014=>"110110101",
  64015=>"000100100",
  64016=>"111101111",
  64017=>"101011111",
  64018=>"100110111",
  64019=>"001001101",
  64020=>"111001011",
  64021=>"000101011",
  64022=>"100011100",
  64023=>"000100111",
  64024=>"010000111",
  64025=>"010011010",
  64026=>"001001101",
  64027=>"010100000",
  64028=>"110000001",
  64029=>"010111011",
  64030=>"001000000",
  64031=>"100000010",
  64032=>"110111110",
  64033=>"110011010",
  64034=>"001100101",
  64035=>"111001111",
  64036=>"010000010",
  64037=>"011000010",
  64038=>"011101000",
  64039=>"010010000",
  64040=>"010011001",
  64041=>"101000101",
  64042=>"101110010",
  64043=>"001111100",
  64044=>"111011010",
  64045=>"000101101",
  64046=>"000100000",
  64047=>"011111000",
  64048=>"100111111",
  64049=>"111010010",
  64050=>"011001010",
  64051=>"110101101",
  64052=>"100011001",
  64053=>"010110110",
  64054=>"101000010",
  64055=>"010101001",
  64056=>"101000100",
  64057=>"001000000",
  64058=>"100101000",
  64059=>"100111000",
  64060=>"100101110",
  64061=>"101101010",
  64062=>"110010100",
  64063=>"001101101",
  64064=>"110101001",
  64065=>"101001000",
  64066=>"111101011",
  64067=>"011001101",
  64068=>"100001101",
  64069=>"000100000",
  64070=>"000111100",
  64071=>"010011001",
  64072=>"100111011",
  64073=>"010111010",
  64074=>"101110110",
  64075=>"000001010",
  64076=>"011011000",
  64077=>"101000000",
  64078=>"110000000",
  64079=>"010110010",
  64080=>"110000011",
  64081=>"011101001",
  64082=>"100111001",
  64083=>"001100001",
  64084=>"000000010",
  64085=>"100100001",
  64086=>"001100000",
  64087=>"101010010",
  64088=>"101001110",
  64089=>"001100100",
  64090=>"111101101",
  64091=>"111010100",
  64092=>"010010111",
  64093=>"110001111",
  64094=>"100101100",
  64095=>"010110110",
  64096=>"010111111",
  64097=>"001010000",
  64098=>"010010100",
  64099=>"010011010",
  64100=>"110100111",
  64101=>"110010001",
  64102=>"111111101",
  64103=>"111111110",
  64104=>"011000100",
  64105=>"110100000",
  64106=>"000011101",
  64107=>"101010000",
  64108=>"001110101",
  64109=>"111111011",
  64110=>"001101110",
  64111=>"111001111",
  64112=>"011110010",
  64113=>"011101110",
  64114=>"011011011",
  64115=>"110011000",
  64116=>"111101011",
  64117=>"011000011",
  64118=>"111001111",
  64119=>"101011111",
  64120=>"010011101",
  64121=>"000110100",
  64122=>"110011010",
  64123=>"101101111",
  64124=>"111100000",
  64125=>"000110011",
  64126=>"110011100",
  64127=>"101111101",
  64128=>"100110000",
  64129=>"010010011",
  64130=>"011001010",
  64131=>"001000101",
  64132=>"000010111",
  64133=>"110101101",
  64134=>"011100100",
  64135=>"110110000",
  64136=>"011100011",
  64137=>"101101000",
  64138=>"111111101",
  64139=>"001010111",
  64140=>"010111010",
  64141=>"110001100",
  64142=>"010001100",
  64143=>"000111000",
  64144=>"110100001",
  64145=>"001010000",
  64146=>"111101101",
  64147=>"101011010",
  64148=>"101111001",
  64149=>"001101001",
  64150=>"000110110",
  64151=>"001010111",
  64152=>"100000110",
  64153=>"010000000",
  64154=>"100010101",
  64155=>"010010011",
  64156=>"010001010",
  64157=>"101000001",
  64158=>"111011100",
  64159=>"100011001",
  64160=>"001111111",
  64161=>"101000010",
  64162=>"001101110",
  64163=>"010000110",
  64164=>"010010101",
  64165=>"000001011",
  64166=>"000101100",
  64167=>"000101110",
  64168=>"011000101",
  64169=>"110100110",
  64170=>"101101100",
  64171=>"100100000",
  64172=>"111110000",
  64173=>"010101000",
  64174=>"000111010",
  64175=>"000110010",
  64176=>"111010101",
  64177=>"110100101",
  64178=>"001001111",
  64179=>"100111001",
  64180=>"100110111",
  64181=>"001111110",
  64182=>"010000001",
  64183=>"010111000",
  64184=>"000101100",
  64185=>"110101100",
  64186=>"000101000",
  64187=>"001100100",
  64188=>"101010110",
  64189=>"010011010",
  64190=>"101101101",
  64191=>"110001101",
  64192=>"110011100",
  64193=>"110111110",
  64194=>"101000001",
  64195=>"110010011",
  64196=>"010101100",
  64197=>"111000110",
  64198=>"100000001",
  64199=>"111000011",
  64200=>"110010100",
  64201=>"000010110",
  64202=>"101110011",
  64203=>"101100100",
  64204=>"001101101",
  64205=>"110011100",
  64206=>"011110000",
  64207=>"001011100",
  64208=>"011111110",
  64209=>"000000000",
  64210=>"110111110",
  64211=>"100001001",
  64212=>"101000110",
  64213=>"101111111",
  64214=>"000010001",
  64215=>"001011100",
  64216=>"000000110",
  64217=>"001001011",
  64218=>"001100101",
  64219=>"100000011",
  64220=>"101101100",
  64221=>"001101100",
  64222=>"100111110",
  64223=>"001011101",
  64224=>"010001010",
  64225=>"111011100",
  64226=>"100100011",
  64227=>"010110100",
  64228=>"100101001",
  64229=>"110010001",
  64230=>"111111010",
  64231=>"010110100",
  64232=>"110011010",
  64233=>"000010100",
  64234=>"101000011",
  64235=>"110101100",
  64236=>"111110101",
  64237=>"110111110",
  64238=>"000011011",
  64239=>"100001100",
  64240=>"011101000",
  64241=>"110101100",
  64242=>"100001001",
  64243=>"000101100",
  64244=>"101110011",
  64245=>"111000110",
  64246=>"101011111",
  64247=>"001010001",
  64248=>"001100110",
  64249=>"001010101",
  64250=>"110000010",
  64251=>"010001100",
  64252=>"100001001",
  64253=>"001011000",
  64254=>"100110001",
  64255=>"101100110",
  64256=>"011100100",
  64257=>"101110010",
  64258=>"011101101",
  64259=>"111000010",
  64260=>"110100000",
  64261=>"100111110",
  64262=>"001001011",
  64263=>"111000101",
  64264=>"011000101",
  64265=>"000111111",
  64266=>"110000110",
  64267=>"011111100",
  64268=>"010001010",
  64269=>"110110001",
  64270=>"011011111",
  64271=>"111010011",
  64272=>"000100110",
  64273=>"110001111",
  64274=>"101000001",
  64275=>"111001111",
  64276=>"011001011",
  64277=>"010011111",
  64278=>"000010100",
  64279=>"110101011",
  64280=>"101000001",
  64281=>"001101000",
  64282=>"011111111",
  64283=>"000011001",
  64284=>"010110010",
  64285=>"111001110",
  64286=>"010100101",
  64287=>"110011011",
  64288=>"100010101",
  64289=>"011011011",
  64290=>"000001001",
  64291=>"001101001",
  64292=>"101001010",
  64293=>"101000100",
  64294=>"100111010",
  64295=>"101001110",
  64296=>"010110110",
  64297=>"100100001",
  64298=>"101010101",
  64299=>"110000011",
  64300=>"111001000",
  64301=>"001011101",
  64302=>"101001101",
  64303=>"111100000",
  64304=>"111001111",
  64305=>"001111011",
  64306=>"111101110",
  64307=>"111110011",
  64308=>"011111000",
  64309=>"000101001",
  64310=>"110100111",
  64311=>"011110000",
  64312=>"001100100",
  64313=>"000011111",
  64314=>"001110101",
  64315=>"100100110",
  64316=>"111100000",
  64317=>"101101000",
  64318=>"001111100",
  64319=>"111001111",
  64320=>"100000011",
  64321=>"011110011",
  64322=>"110100111",
  64323=>"000101101",
  64324=>"000100110",
  64325=>"111110100",
  64326=>"101000001",
  64327=>"100100000",
  64328=>"011111110",
  64329=>"101000011",
  64330=>"101111110",
  64331=>"110110100",
  64332=>"011010010",
  64333=>"010100110",
  64334=>"101100000",
  64335=>"001100110",
  64336=>"101101101",
  64337=>"101011110",
  64338=>"011101000",
  64339=>"110010001",
  64340=>"101111101",
  64341=>"100001100",
  64342=>"111111111",
  64343=>"011001011",
  64344=>"010110100",
  64345=>"111100101",
  64346=>"111110111",
  64347=>"001111101",
  64348=>"111001100",
  64349=>"000001111",
  64350=>"000011000",
  64351=>"110111111",
  64352=>"110100011",
  64353=>"100000100",
  64354=>"000010100",
  64355=>"110111110",
  64356=>"011001010",
  64357=>"110001010",
  64358=>"001010011",
  64359=>"010011110",
  64360=>"110101000",
  64361=>"110110000",
  64362=>"011111010",
  64363=>"111101001",
  64364=>"100100100",
  64365=>"000111111",
  64366=>"111100101",
  64367=>"011000000",
  64368=>"011001110",
  64369=>"101101100",
  64370=>"101000111",
  64371=>"111001010",
  64372=>"101111111",
  64373=>"101101111",
  64374=>"101101110",
  64375=>"111101000",
  64376=>"001111100",
  64377=>"101000001",
  64378=>"010001110",
  64379=>"000101000",
  64380=>"111111100",
  64381=>"000100110",
  64382=>"100000101",
  64383=>"000000100",
  64384=>"111010111",
  64385=>"100010001",
  64386=>"100001111",
  64387=>"111101000",
  64388=>"100111110",
  64389=>"001011000",
  64390=>"110000100",
  64391=>"000100011",
  64392=>"101000101",
  64393=>"110101100",
  64394=>"010001000",
  64395=>"001001000",
  64396=>"000011010",
  64397=>"001111111",
  64398=>"110101111",
  64399=>"110110110",
  64400=>"101000111",
  64401=>"000100000",
  64402=>"111101100",
  64403=>"100011001",
  64404=>"001110010",
  64405=>"011101110",
  64406=>"000000111",
  64407=>"111010010",
  64408=>"010111011",
  64409=>"000001110",
  64410=>"010101011",
  64411=>"100111111",
  64412=>"110010101",
  64413=>"110010000",
  64414=>"011100100",
  64415=>"011011100",
  64416=>"101100000",
  64417=>"010110101",
  64418=>"001011110",
  64419=>"101001101",
  64420=>"010110111",
  64421=>"010111011",
  64422=>"010101000",
  64423=>"100001011",
  64424=>"000011110",
  64425=>"100000101",
  64426=>"110001111",
  64427=>"011011111",
  64428=>"110111000",
  64429=>"111010110",
  64430=>"111111011",
  64431=>"100110101",
  64432=>"111101001",
  64433=>"101010100",
  64434=>"100000110",
  64435=>"101010000",
  64436=>"110000101",
  64437=>"001000000",
  64438=>"110101101",
  64439=>"010001000",
  64440=>"000001010",
  64441=>"000110111",
  64442=>"001100111",
  64443=>"111111110",
  64444=>"110100011",
  64445=>"001001110",
  64446=>"011100101",
  64447=>"001111001",
  64448=>"001111101",
  64449=>"001110000",
  64450=>"000011001",
  64451=>"110101011",
  64452=>"001001010",
  64453=>"010001100",
  64454=>"111100111",
  64455=>"010010101",
  64456=>"100110110",
  64457=>"010101011",
  64458=>"001011101",
  64459=>"111001010",
  64460=>"111110011",
  64461=>"101000100",
  64462=>"110011110",
  64463=>"111100100",
  64464=>"101100000",
  64465=>"000010000",
  64466=>"011000011",
  64467=>"001100011",
  64468=>"001100010",
  64469=>"000101110",
  64470=>"000010000",
  64471=>"111101101",
  64472=>"101101101",
  64473=>"100010010",
  64474=>"101011111",
  64475=>"100100001",
  64476=>"101110001",
  64477=>"101010001",
  64478=>"100100100",
  64479=>"011111001",
  64480=>"101101101",
  64481=>"011000001",
  64482=>"100111101",
  64483=>"101110000",
  64484=>"111101010",
  64485=>"100111110",
  64486=>"100001001",
  64487=>"011101001",
  64488=>"100101011",
  64489=>"010000011",
  64490=>"100111100",
  64491=>"010011100",
  64492=>"110010011",
  64493=>"101001010",
  64494=>"011010101",
  64495=>"110111011",
  64496=>"000001110",
  64497=>"100001111",
  64498=>"101110110",
  64499=>"101110111",
  64500=>"110111110",
  64501=>"101000110",
  64502=>"011000011",
  64503=>"000010111",
  64504=>"111101111",
  64505=>"111110111",
  64506=>"100010110",
  64507=>"011010111",
  64508=>"010001001",
  64509=>"011101110",
  64510=>"011011011",
  64511=>"110000011",
  64512=>"101010111",
  64513=>"000111001",
  64514=>"001001001",
  64515=>"111001100",
  64516=>"000001000",
  64517=>"101000110",
  64518=>"011011011",
  64519=>"111001001",
  64520=>"110011001",
  64521=>"100100011",
  64522=>"101100000",
  64523=>"111111110",
  64524=>"001010010",
  64525=>"100111001",
  64526=>"110001110",
  64527=>"111110010",
  64528=>"001100101",
  64529=>"110000111",
  64530=>"110111011",
  64531=>"111111100",
  64532=>"000010100",
  64533=>"111010100",
  64534=>"110100111",
  64535=>"100100000",
  64536=>"010110100",
  64537=>"011010101",
  64538=>"000110111",
  64539=>"001101001",
  64540=>"111101000",
  64541=>"101011001",
  64542=>"111110111",
  64543=>"111011110",
  64544=>"101000111",
  64545=>"100001110",
  64546=>"010000001",
  64547=>"110011111",
  64548=>"101101111",
  64549=>"111010010",
  64550=>"110010011",
  64551=>"010010100",
  64552=>"100110000",
  64553=>"100111111",
  64554=>"011010101",
  64555=>"110111101",
  64556=>"000101111",
  64557=>"011100101",
  64558=>"111001111",
  64559=>"011001011",
  64560=>"101110010",
  64561=>"101110100",
  64562=>"010110100",
  64563=>"000001111",
  64564=>"011110011",
  64565=>"110101000",
  64566=>"011110010",
  64567=>"010111011",
  64568=>"100110111",
  64569=>"100010001",
  64570=>"011011100",
  64571=>"100110100",
  64572=>"110010011",
  64573=>"111110011",
  64574=>"110101110",
  64575=>"110100001",
  64576=>"010000100",
  64577=>"101000100",
  64578=>"000011111",
  64579=>"110001100",
  64580=>"100100110",
  64581=>"110001010",
  64582=>"101110101",
  64583=>"110110000",
  64584=>"110101111",
  64585=>"110110100",
  64586=>"000110011",
  64587=>"011101110",
  64588=>"110000101",
  64589=>"011101101",
  64590=>"100011001",
  64591=>"001010100",
  64592=>"101100010",
  64593=>"011110101",
  64594=>"010001111",
  64595=>"001001111",
  64596=>"001000101",
  64597=>"010101111",
  64598=>"111110100",
  64599=>"000010110",
  64600=>"001100001",
  64601=>"111000001",
  64602=>"110110101",
  64603=>"101001110",
  64604=>"000110100",
  64605=>"110111101",
  64606=>"001010100",
  64607=>"111010111",
  64608=>"100111010",
  64609=>"111000001",
  64610=>"000111000",
  64611=>"110100111",
  64612=>"110101100",
  64613=>"111101111",
  64614=>"111011111",
  64615=>"100111111",
  64616=>"010011001",
  64617=>"001101110",
  64618=>"100011000",
  64619=>"010000110",
  64620=>"010010011",
  64621=>"111101001",
  64622=>"111110010",
  64623=>"110110001",
  64624=>"101000001",
  64625=>"100101001",
  64626=>"100001101",
  64627=>"110010001",
  64628=>"101100110",
  64629=>"011110010",
  64630=>"111101011",
  64631=>"011010101",
  64632=>"011011100",
  64633=>"110001111",
  64634=>"111110111",
  64635=>"101110110",
  64636=>"010011101",
  64637=>"001001010",
  64638=>"101010010",
  64639=>"001111101",
  64640=>"111101100",
  64641=>"011111101",
  64642=>"001110011",
  64643=>"011111001",
  64644=>"110110011",
  64645=>"000010110",
  64646=>"101101010",
  64647=>"000110000",
  64648=>"110100101",
  64649=>"100001111",
  64650=>"101100100",
  64651=>"111100110",
  64652=>"100101001",
  64653=>"111100100",
  64654=>"101100111",
  64655=>"001000011",
  64656=>"000001101",
  64657=>"000111010",
  64658=>"101100100",
  64659=>"010001101",
  64660=>"111111011",
  64661=>"101100110",
  64662=>"000010000",
  64663=>"100001010",
  64664=>"000010100",
  64665=>"101010100",
  64666=>"010111101",
  64667=>"111110111",
  64668=>"110110011",
  64669=>"110111101",
  64670=>"001010111",
  64671=>"101010011",
  64672=>"001010101",
  64673=>"100011110",
  64674=>"010101011",
  64675=>"100111000",
  64676=>"101111111",
  64677=>"011010111",
  64678=>"000010100",
  64679=>"100011100",
  64680=>"100010101",
  64681=>"001101111",
  64682=>"000000100",
  64683=>"101110011",
  64684=>"011011101",
  64685=>"100101001",
  64686=>"100010110",
  64687=>"111110001",
  64688=>"111011000",
  64689=>"100111110",
  64690=>"010111011",
  64691=>"011101110",
  64692=>"100101011",
  64693=>"110001000",
  64694=>"110111111",
  64695=>"010111111",
  64696=>"010010000",
  64697=>"111101110",
  64698=>"100001110",
  64699=>"001100010",
  64700=>"100111101",
  64701=>"001011000",
  64702=>"011100011",
  64703=>"101110101",
  64704=>"100000111",
  64705=>"101001011",
  64706=>"101011011",
  64707=>"101010000",
  64708=>"010000011",
  64709=>"100111001",
  64710=>"001110111",
  64711=>"101000110",
  64712=>"011010101",
  64713=>"000101101",
  64714=>"010111100",
  64715=>"001000000",
  64716=>"001001100",
  64717=>"000100001",
  64718=>"110100001",
  64719=>"111000110",
  64720=>"101110101",
  64721=>"101110100",
  64722=>"000100111",
  64723=>"100010000",
  64724=>"000101000",
  64725=>"101111101",
  64726=>"101000000",
  64727=>"111100011",
  64728=>"101011011",
  64729=>"111001010",
  64730=>"000010110",
  64731=>"101110001",
  64732=>"000100011",
  64733=>"001011111",
  64734=>"111111101",
  64735=>"010001011",
  64736=>"100100010",
  64737=>"011101100",
  64738=>"001001000",
  64739=>"110100000",
  64740=>"111010001",
  64741=>"011101111",
  64742=>"000001100",
  64743=>"100111000",
  64744=>"101001001",
  64745=>"100101110",
  64746=>"010111101",
  64747=>"001100011",
  64748=>"111100100",
  64749=>"100010001",
  64750=>"001100100",
  64751=>"101101110",
  64752=>"000101010",
  64753=>"111001000",
  64754=>"000000010",
  64755=>"110011110",
  64756=>"001111111",
  64757=>"001110101",
  64758=>"100001011",
  64759=>"001111111",
  64760=>"110101000",
  64761=>"010101010",
  64762=>"001000001",
  64763=>"110100110",
  64764=>"010100011",
  64765=>"000000001",
  64766=>"010111101",
  64767=>"011010110",
  64768=>"010011100",
  64769=>"001001000",
  64770=>"100101111",
  64771=>"111010000",
  64772=>"010000100",
  64773=>"001100100",
  64774=>"111110110",
  64775=>"100110010",
  64776=>"110110111",
  64777=>"111001100",
  64778=>"000011111",
  64779=>"111101001",
  64780=>"011110110",
  64781=>"111011011",
  64782=>"101110001",
  64783=>"011010110",
  64784=>"000111110",
  64785=>"000101010",
  64786=>"111100101",
  64787=>"011001001",
  64788=>"111010110",
  64789=>"001001111",
  64790=>"101100111",
  64791=>"111110011",
  64792=>"011000110",
  64793=>"101100000",
  64794=>"111100001",
  64795=>"111000001",
  64796=>"111111101",
  64797=>"111110000",
  64798=>"111001010",
  64799=>"010000110",
  64800=>"110101100",
  64801=>"101001011",
  64802=>"111001001",
  64803=>"111100101",
  64804=>"111011111",
  64805=>"010010111",
  64806=>"001001010",
  64807=>"110010000",
  64808=>"110010111",
  64809=>"001111100",
  64810=>"011001110",
  64811=>"101010100",
  64812=>"000001011",
  64813=>"111111101",
  64814=>"110010110",
  64815=>"001011011",
  64816=>"101000011",
  64817=>"100011000",
  64818=>"011110000",
  64819=>"001101110",
  64820=>"010100110",
  64821=>"100100100",
  64822=>"100001101",
  64823=>"000101010",
  64824=>"011111111",
  64825=>"010011011",
  64826=>"100000101",
  64827=>"000000010",
  64828=>"011010111",
  64829=>"100111100",
  64830=>"000110110",
  64831=>"111110100",
  64832=>"001110000",
  64833=>"000001010",
  64834=>"000100000",
  64835=>"111111111",
  64836=>"100010111",
  64837=>"100011011",
  64838=>"001111000",
  64839=>"101101101",
  64840=>"111011110",
  64841=>"000110001",
  64842=>"001101010",
  64843=>"001010001",
  64844=>"011111100",
  64845=>"011101011",
  64846=>"010000001",
  64847=>"001010110",
  64848=>"001001101",
  64849=>"011000011",
  64850=>"000011111",
  64851=>"000101000",
  64852=>"110100011",
  64853=>"001111111",
  64854=>"011100011",
  64855=>"101101010",
  64856=>"110000011",
  64857=>"111011010",
  64858=>"010100101",
  64859=>"111101111",
  64860=>"110111111",
  64861=>"010101110",
  64862=>"011111001",
  64863=>"010110101",
  64864=>"001111101",
  64865=>"011110000",
  64866=>"100100001",
  64867=>"111011101",
  64868=>"100010011",
  64869=>"100101110",
  64870=>"111101010",
  64871=>"111101001",
  64872=>"010100111",
  64873=>"110110111",
  64874=>"011100010",
  64875=>"110111000",
  64876=>"101011010",
  64877=>"011111101",
  64878=>"101100101",
  64879=>"100110100",
  64880=>"001100110",
  64881=>"001001000",
  64882=>"010001001",
  64883=>"111111111",
  64884=>"001000110",
  64885=>"000110011",
  64886=>"110101010",
  64887=>"010110111",
  64888=>"001110001",
  64889=>"101100110",
  64890=>"110001000",
  64891=>"000000001",
  64892=>"000001000",
  64893=>"011001101",
  64894=>"010110011",
  64895=>"110111110",
  64896=>"110101110",
  64897=>"011000100",
  64898=>"110101110",
  64899=>"110101100",
  64900=>"111001101",
  64901=>"010110011",
  64902=>"000101110",
  64903=>"110110110",
  64904=>"011101110",
  64905=>"001110011",
  64906=>"011101000",
  64907=>"001111000",
  64908=>"000010011",
  64909=>"100001100",
  64910=>"100110111",
  64911=>"000001011",
  64912=>"111010001",
  64913=>"001110010",
  64914=>"001000000",
  64915=>"000110011",
  64916=>"101001010",
  64917=>"010101000",
  64918=>"000111110",
  64919=>"110001010",
  64920=>"111011011",
  64921=>"111000110",
  64922=>"011101010",
  64923=>"011010100",
  64924=>"001000111",
  64925=>"110101110",
  64926=>"011011011",
  64927=>"111100011",
  64928=>"101011010",
  64929=>"001001111",
  64930=>"001000001",
  64931=>"011101101",
  64932=>"010000001",
  64933=>"101111001",
  64934=>"101100000",
  64935=>"111010000",
  64936=>"100100110",
  64937=>"001111000",
  64938=>"110101111",
  64939=>"111010011",
  64940=>"111101111",
  64941=>"001111111",
  64942=>"000010111",
  64943=>"010000101",
  64944=>"010101111",
  64945=>"010101111",
  64946=>"101110011",
  64947=>"000010110",
  64948=>"000001011",
  64949=>"010111101",
  64950=>"001111011",
  64951=>"001110101",
  64952=>"111111101",
  64953=>"010010111",
  64954=>"101101101",
  64955=>"111100101",
  64956=>"010011001",
  64957=>"111001010",
  64958=>"100001000",
  64959=>"100000100",
  64960=>"110001000",
  64961=>"111101110",
  64962=>"101001110",
  64963=>"000001101",
  64964=>"010111110",
  64965=>"101100100",
  64966=>"001000100",
  64967=>"111111110",
  64968=>"101110100",
  64969=>"111010001",
  64970=>"011110100",
  64971=>"001110011",
  64972=>"100000111",
  64973=>"000011110",
  64974=>"100111100",
  64975=>"111100111",
  64976=>"110111011",
  64977=>"110011110",
  64978=>"001100011",
  64979=>"100001011",
  64980=>"100110101",
  64981=>"110100111",
  64982=>"010101110",
  64983=>"111011111",
  64984=>"100111100",
  64985=>"000000001",
  64986=>"000010000",
  64987=>"011111000",
  64988=>"101011010",
  64989=>"110010100",
  64990=>"000101001",
  64991=>"001100001",
  64992=>"100111011",
  64993=>"101110100",
  64994=>"101001011",
  64995=>"000111110",
  64996=>"101100101",
  64997=>"111000111",
  64998=>"000001101",
  64999=>"001111010",
  65000=>"000001000",
  65001=>"000010101",
  65002=>"101001111",
  65003=>"101110110",
  65004=>"110000100",
  65005=>"100110111",
  65006=>"110001010",
  65007=>"010111110",
  65008=>"001001100",
  65009=>"011000000",
  65010=>"011000011",
  65011=>"011000011",
  65012=>"011100001",
  65013=>"011011111",
  65014=>"101101011",
  65015=>"101100110",
  65016=>"100110011",
  65017=>"111101000",
  65018=>"110110110",
  65019=>"100001100",
  65020=>"000101110",
  65021=>"000101101",
  65022=>"011110101",
  65023=>"001100001",
  65024=>"101001110",
  65025=>"011000011",
  65026=>"000110000",
  65027=>"100100010",
  65028=>"000010110",
  65029=>"011000110",
  65030=>"001100011",
  65031=>"011001100",
  65032=>"100001001",
  65033=>"000011101",
  65034=>"100011001",
  65035=>"110010001",
  65036=>"101110010",
  65037=>"011011111",
  65038=>"000111101",
  65039=>"001101100",
  65040=>"010010111",
  65041=>"101011001",
  65042=>"111010111",
  65043=>"111110011",
  65044=>"011101100",
  65045=>"001000100",
  65046=>"101110110",
  65047=>"010011111",
  65048=>"110110110",
  65049=>"010011000",
  65050=>"101110110",
  65051=>"000011111",
  65052=>"110010111",
  65053=>"011100011",
  65054=>"101011101",
  65055=>"010011010",
  65056=>"000011000",
  65057=>"011110000",
  65058=>"010110001",
  65059=>"101010011",
  65060=>"010010011",
  65061=>"100101010",
  65062=>"001011101",
  65063=>"000110001",
  65064=>"011011010",
  65065=>"110100001",
  65066=>"011111000",
  65067=>"000010111",
  65068=>"110111111",
  65069=>"110101100",
  65070=>"001001110",
  65071=>"100100111",
  65072=>"010010100",
  65073=>"011000000",
  65074=>"100011001",
  65075=>"110001110",
  65076=>"100000010",
  65077=>"001011111",
  65078=>"100011100",
  65079=>"010110001",
  65080=>"100000001",
  65081=>"111101111",
  65082=>"110101101",
  65083=>"000100101",
  65084=>"010011100",
  65085=>"011001010",
  65086=>"010011011",
  65087=>"100111110",
  65088=>"100010000",
  65089=>"111010111",
  65090=>"100101100",
  65091=>"100111000",
  65092=>"101110110",
  65093=>"110010101",
  65094=>"001011111",
  65095=>"110011011",
  65096=>"000000111",
  65097=>"111000001",
  65098=>"110100010",
  65099=>"110101011",
  65100=>"000101111",
  65101=>"110100101",
  65102=>"000100011",
  65103=>"001010011",
  65104=>"000010011",
  65105=>"011101000",
  65106=>"100111001",
  65107=>"100011010",
  65108=>"110001000",
  65109=>"101010001",
  65110=>"010101110",
  65111=>"010010100",
  65112=>"110011111",
  65113=>"110111110",
  65114=>"001100100",
  65115=>"100010111",
  65116=>"011101111",
  65117=>"110101010",
  65118=>"110010010",
  65119=>"100001111",
  65120=>"011001011",
  65121=>"001001100",
  65122=>"011001100",
  65123=>"101011011",
  65124=>"100001010",
  65125=>"100111100",
  65126=>"010100011",
  65127=>"111111001",
  65128=>"001011001",
  65129=>"001011100",
  65130=>"111111000",
  65131=>"111111010",
  65132=>"000110011",
  65133=>"000001010",
  65134=>"001110011",
  65135=>"100001010",
  65136=>"101101101",
  65137=>"111110001",
  65138=>"101001011",
  65139=>"111101111",
  65140=>"111111000",
  65141=>"000001110",
  65142=>"001011010",
  65143=>"101001010",
  65144=>"111000001",
  65145=>"011001001",
  65146=>"111011100",
  65147=>"010110010",
  65148=>"101100111",
  65149=>"000010101",
  65150=>"110100110",
  65151=>"001010101",
  65152=>"100001110",
  65153=>"010000100",
  65154=>"000000011",
  65155=>"001011100",
  65156=>"010001110",
  65157=>"011011001",
  65158=>"101011110",
  65159=>"001011100",
  65160=>"110101001",
  65161=>"011010111",
  65162=>"111111101",
  65163=>"010000000",
  65164=>"011111110",
  65165=>"100110101",
  65166=>"101000111",
  65167=>"011100100",
  65168=>"010101100",
  65169=>"000111101",
  65170=>"010101111",
  65171=>"001111100",
  65172=>"100100000",
  65173=>"101100010",
  65174=>"110000110",
  65175=>"011001000",
  65176=>"101010110",
  65177=>"010101101",
  65178=>"011011101",
  65179=>"110011011",
  65180=>"000011010",
  65181=>"001010110",
  65182=>"010010011",
  65183=>"111001001",
  65184=>"000001010",
  65185=>"110110111",
  65186=>"100110000",
  65187=>"111110101",
  65188=>"001101001",
  65189=>"000111110",
  65190=>"110111001",
  65191=>"100001111",
  65192=>"100001100",
  65193=>"000101101",
  65194=>"110000011",
  65195=>"111111010",
  65196=>"011101101",
  65197=>"110000111",
  65198=>"110011000",
  65199=>"101111001",
  65200=>"100101000",
  65201=>"011111100",
  65202=>"001010010",
  65203=>"101101110",
  65204=>"111111001",
  65205=>"111001101",
  65206=>"011101011",
  65207=>"010100001",
  65208=>"011111011",
  65209=>"010111000",
  65210=>"000001100",
  65211=>"001100101",
  65212=>"101110110",
  65213=>"000100100",
  65214=>"100001000",
  65215=>"100011001",
  65216=>"110111011",
  65217=>"000101010",
  65218=>"100000000",
  65219=>"010000111",
  65220=>"000101001",
  65221=>"100101011",
  65222=>"000100010",
  65223=>"000000101",
  65224=>"001100000",
  65225=>"000111011",
  65226=>"011101101",
  65227=>"100000101",
  65228=>"010111000",
  65229=>"110001011",
  65230=>"110100101",
  65231=>"011110011",
  65232=>"100010000",
  65233=>"000001001",
  65234=>"100001001",
  65235=>"001001110",
  65236=>"111000000",
  65237=>"011011010",
  65238=>"110001011",
  65239=>"000110100",
  65240=>"100000000",
  65241=>"000010111",
  65242=>"011001011",
  65243=>"001000101",
  65244=>"100101010",
  65245=>"101110010",
  65246=>"111101110",
  65247=>"100101111",
  65248=>"011101011",
  65249=>"110110111",
  65250=>"100110111",
  65251=>"000111000",
  65252=>"010010100",
  65253=>"101101010",
  65254=>"101010111",
  65255=>"110101001",
  65256=>"011010100",
  65257=>"110110110",
  65258=>"101000111",
  65259=>"101000010",
  65260=>"110100111",
  65261=>"000010100",
  65262=>"000010001",
  65263=>"101011110",
  65264=>"100000110",
  65265=>"011001000",
  65266=>"100001101",
  65267=>"110111110",
  65268=>"011010101",
  65269=>"111000111",
  65270=>"111011100",
  65271=>"010001011",
  65272=>"010001110",
  65273=>"111011011",
  65274=>"111011000",
  65275=>"101010110",
  65276=>"000001110",
  65277=>"110011001",
  65278=>"001010001",
  65279=>"101011101",
  65280=>"101011011",
  65281=>"101011001",
  65282=>"011000100",
  65283=>"110110110",
  65284=>"111011100",
  65285=>"100011011",
  65286=>"100111110",
  65287=>"111001100",
  65288=>"101111001",
  65289=>"100111001",
  65290=>"101000011",
  65291=>"100111010",
  65292=>"111110110",
  65293=>"111001110",
  65294=>"011111101",
  65295=>"101101010",
  65296=>"111100001",
  65297=>"001000001",
  65298=>"011111101",
  65299=>"110101100",
  65300=>"011000011",
  65301=>"010010110",
  65302=>"101010111",
  65303=>"100101101",
  65304=>"100100100",
  65305=>"000010100",
  65306=>"001010011",
  65307=>"010000111",
  65308=>"010111101",
  65309=>"010000100",
  65310=>"010101011",
  65311=>"001001100",
  65312=>"111110001",
  65313=>"000101111",
  65314=>"000000011",
  65315=>"101001010",
  65316=>"111101111",
  65317=>"011101100",
  65318=>"011110001",
  65319=>"100010100",
  65320=>"000011001",
  65321=>"000101010",
  65322=>"110011000",
  65323=>"100010011",
  65324=>"000100000",
  65325=>"010011100",
  65326=>"110110111",
  65327=>"111010111",
  65328=>"111011000",
  65329=>"001010101",
  65330=>"101100100",
  65331=>"101111001",
  65332=>"000001110",
  65333=>"001110111",
  65334=>"000000000",
  65335=>"100010101",
  65336=>"000000110",
  65337=>"000110001",
  65338=>"001001001",
  65339=>"101010110",
  65340=>"111011011",
  65341=>"001100111",
  65342=>"101100001",
  65343=>"010111011",
  65344=>"101110001",
  65345=>"010110100",
  65346=>"001101000",
  65347=>"000110011",
  65348=>"110001010",
  65349=>"110011111",
  65350=>"111101111",
  65351=>"101000000",
  65352=>"110000001",
  65353=>"111101101",
  65354=>"111000100",
  65355=>"000001000",
  65356=>"000010011",
  65357=>"100001011",
  65358=>"000011110",
  65359=>"001011111",
  65360=>"110111011",
  65361=>"100101110",
  65362=>"000100011",
  65363=>"000111101",
  65364=>"000000111",
  65365=>"110100111",
  65366=>"010111110",
  65367=>"001001100",
  65368=>"011001001",
  65369=>"010001011",
  65370=>"001111101",
  65371=>"000111010",
  65372=>"100010010",
  65373=>"000001100",
  65374=>"011000010",
  65375=>"010110111",
  65376=>"001001110",
  65377=>"000110111",
  65378=>"111010110",
  65379=>"001010000",
  65380=>"100000101",
  65381=>"011110011",
  65382=>"100111100",
  65383=>"101101101",
  65384=>"110100000",
  65385=>"101110001",
  65386=>"101000100",
  65387=>"010010110",
  65388=>"101100101",
  65389=>"100100111",
  65390=>"000100101",
  65391=>"101111111",
  65392=>"101100111",
  65393=>"101000000",
  65394=>"011011101",
  65395=>"100111111",
  65396=>"111101000",
  65397=>"100100100",
  65398=>"101010111",
  65399=>"001110000",
  65400=>"110001100",
  65401=>"011001011",
  65402=>"000001111",
  65403=>"111110001",
  65404=>"100100111",
  65405=>"000101011",
  65406=>"010010011",
  65407=>"111011011",
  65408=>"101110010",
  65409=>"101111111",
  65410=>"111111101",
  65411=>"000110111",
  65412=>"110001011",
  65413=>"110001000",
  65414=>"011111110",
  65415=>"011000111",
  65416=>"011010010",
  65417=>"001100001",
  65418=>"001111011",
  65419=>"000000111",
  65420=>"011001001",
  65421=>"010011000",
  65422=>"001001110",
  65423=>"110100001",
  65424=>"110101110",
  65425=>"111101100",
  65426=>"000010111",
  65427=>"000001000",
  65428=>"001110010",
  65429=>"000000001",
  65430=>"110001000",
  65431=>"011001111",
  65432=>"100000110",
  65433=>"110110010",
  65434=>"101000101",
  65435=>"110010001",
  65436=>"110111010",
  65437=>"000110010",
  65438=>"111001101",
  65439=>"011101011",
  65440=>"010001010",
  65441=>"001010000",
  65442=>"011111111",
  65443=>"010100010",
  65444=>"110100100",
  65445=>"010100111",
  65446=>"001110111",
  65447=>"011000100",
  65448=>"000010010",
  65449=>"010011001",
  65450=>"000000111",
  65451=>"110111011",
  65452=>"101101011",
  65453=>"111001100",
  65454=>"010111000",
  65455=>"010101000",
  65456=>"100000010",
  65457=>"101000001",
  65458=>"010110001",
  65459=>"010100010",
  65460=>"010011110",
  65461=>"000000101",
  65462=>"110111110",
  65463=>"010111101",
  65464=>"101101111",
  65465=>"001000110",
  65466=>"001110101",
  65467=>"100010000",
  65468=>"000100100",
  65469=>"010001100",
  65470=>"011101000",
  65471=>"010101111",
  65472=>"110010011",
  65473=>"111000001",
  65474=>"101101011",
  65475=>"111110010",
  65476=>"011001011",
  65477=>"101111100",
  65478=>"110111100",
  65479=>"101111101",
  65480=>"111111110",
  65481=>"010111100",
  65482=>"101110111",
  65483=>"110011101",
  65484=>"011011011",
  65485=>"101111011",
  65486=>"011001000",
  65487=>"001111110",
  65488=>"010110101",
  65489=>"000001000",
  65490=>"111011100",
  65491=>"010110110",
  65492=>"010000010",
  65493=>"001000101",
  65494=>"100011101",
  65495=>"100000001",
  65496=>"111111101",
  65497=>"100011000",
  65498=>"010010011",
  65499=>"000100000",
  65500=>"010100110",
  65501=>"000000110",
  65502=>"000000001",
  65503=>"111111110",
  65504=>"011001000",
  65505=>"100101000",
  65506=>"111111001",
  65507=>"010010100",
  65508=>"100010111",
  65509=>"010000111",
  65510=>"101101011",
  65511=>"001000000",
  65512=>"111111000",
  65513=>"001111111",
  65514=>"010001110",
  65515=>"110000100",
  65516=>"101111100",
  65517=>"001001101",
  65518=>"000001100",
  65519=>"010110011",
  65520=>"100111111",
  65521=>"000110000",
  65522=>"101011101",
  65523=>"001000100",
  65524=>"110110100",
  65525=>"010111010",
  65526=>"110011001",
  65527=>"110101101",
  65528=>"010011110",
  65529=>"010001111",
  65530=>"101111110",
  65531=>"100010010",
  65532=>"000110101",
  65533=>"001000111",
  65534=>"110100011",
  65535=>"001000111");

BEGIN
  weight <= ROM_content(to_integer(address));
END RTL;