LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L9_2_WROM IS
  PORT (
    weight : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    address : IN unsigned(weightsbitsAddress(9)-1 DOWNTO 0));
END L9_2_WROM;

ARCHITECTURE RTL OF L9_2_WROM IS

  TYPE ROM_mem IS ARRAY (0 TO 64511) OF STD_LOGIC_VECTOR(7 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem := (0=>"11111110",
  1=>"00000010",
  2=>"00000010",
  3=>"00000100",
  4=>"11111110",
  5=>"11111110",
  6=>"11111110",
  7=>"00000010",
  8=>"11111101",
  9=>"11111111",
  10=>"00000000",
  11=>"11111101",
  12=>"11111110",
  13=>"00000100",
  14=>"00000100",
  15=>"11111111",
  16=>"11111111",
  17=>"11111111",
  18=>"11111100",
  19=>"00000000",
  20=>"00000011",
  21=>"00000001",
  22=>"00000000",
  23=>"11111101",
  24=>"00000001",
  25=>"00000010",
  26=>"11111101",
  27=>"00000011",
  28=>"00000011",
  29=>"00000001",
  30=>"00000000",
  31=>"11111101",
  32=>"11111111",
  33=>"11111111",
  34=>"00000010",
  35=>"00000011",
  36=>"00000001",
  37=>"11111111",
  38=>"00000001",
  39=>"11111110",
  40=>"00000010",
  41=>"00000011",
  42=>"11111101",
  43=>"11111101",
  44=>"00000010",
  45=>"00000001",
  46=>"11111110",
  47=>"11111110",
  48=>"00000000",
  49=>"11111111",
  50=>"00000001",
  51=>"00000000",
  52=>"11111101",
  53=>"11111101",
  54=>"00000000",
  55=>"00000010",
  56=>"00000011",
  57=>"11111111",
  58=>"00000010",
  59=>"00000100",
  60=>"11111111",
  61=>"00000011",
  62=>"11111111",
  63=>"11111111",
  64=>"00000000",
  65=>"11111111",
  66=>"00000010",
  67=>"00000100",
  68=>"00000100",
  69=>"00000011",
  70=>"00000111",
  71=>"00000010",
  72=>"11111110",
  73=>"11111100",
  74=>"00000100",
  75=>"00000010",
  76=>"00000001",
  77=>"00000001",
  78=>"00000010",
  79=>"00000000",
  80=>"11111111",
  81=>"00000000",
  82=>"00000100",
  83=>"11111111",
  84=>"00000100",
  85=>"11111101",
  86=>"11111101",
  87=>"00000011",
  88=>"00000100",
  89=>"00000000",
  90=>"00000001",
  91=>"11111101",
  92=>"00000001",
  93=>"11111100",
  94=>"11111111",
  95=>"00000011",
  96=>"00000001",
  97=>"00000011",
  98=>"00001000",
  99=>"00000000",
  100=>"00000010",
  101=>"00000010",
  102=>"11111101",
  103=>"00000011",
  104=>"00000100",
  105=>"00000100",
  106=>"00000010",
  107=>"00000000",
  108=>"00000101",
  109=>"00000001",
  110=>"00000101",
  111=>"11111110",
  112=>"00000000",
  113=>"00000001",
  114=>"00000010",
  115=>"11111110",
  116=>"00000011",
  117=>"00000101",
  118=>"11111101",
  119=>"00000010",
  120=>"00000000",
  121=>"11111101",
  122=>"11111100",
  123=>"11111111",
  124=>"11111101",
  125=>"11111110",
  126=>"11111111",
  127=>"00000011",
  128=>"11111101",
  129=>"11111100",
  130=>"11111100",
  131=>"00000101",
  132=>"00000010",
  133=>"00000010",
  134=>"00000010",
  135=>"00000000",
  136=>"11111101",
  137=>"11111111",
  138=>"11111111",
  139=>"11111100",
  140=>"11111110",
  141=>"00000001",
  142=>"11111111",
  143=>"00000011",
  144=>"11111101",
  145=>"11111111",
  146=>"00000010",
  147=>"11111110",
  148=>"11111100",
  149=>"11111100",
  150=>"11111101",
  151=>"00000010",
  152=>"11111110",
  153=>"11111101",
  154=>"00000010",
  155=>"11111111",
  156=>"11111111",
  157=>"11111101",
  158=>"11111101",
  159=>"00000011",
  160=>"00000000",
  161=>"11111110",
  162=>"00000001",
  163=>"11111110",
  164=>"00000000",
  165=>"11111110",
  166=>"00000001",
  167=>"00000001",
  168=>"00000010",
  169=>"00000001",
  170=>"00000011",
  171=>"00000011",
  172=>"00000011",
  173=>"00000000",
  174=>"11111110",
  175=>"11111100",
  176=>"00000010",
  177=>"11111111",
  178=>"11111101",
  179=>"00000001",
  180=>"00000000",
  181=>"11111110",
  182=>"11111100",
  183=>"00000001",
  184=>"11111111",
  185=>"11111111",
  186=>"11111100",
  187=>"00000001",
  188=>"11111110",
  189=>"11111111",
  190=>"11111111",
  191=>"00000010",
  192=>"11111101",
  193=>"00000001",
  194=>"00000001",
  195=>"00000000",
  196=>"00000010",
  197=>"00000011",
  198=>"00000000",
  199=>"11111111",
  200=>"00000000",
  201=>"11111110",
  202=>"00000011",
  203=>"00000001",
  204=>"00000010",
  205=>"11111110",
  206=>"00000001",
  207=>"00000001",
  208=>"11111110",
  209=>"00000010",
  210=>"11111110",
  211=>"00000001",
  212=>"11111101",
  213=>"11111101",
  214=>"11111111",
  215=>"00000000",
  216=>"00000000",
  217=>"00000000",
  218=>"11111111",
  219=>"00000000",
  220=>"00000000",
  221=>"00000011",
  222=>"11111110",
  223=>"00000100",
  224=>"11111110",
  225=>"11111101",
  226=>"11111111",
  227=>"11111111",
  228=>"11111100",
  229=>"00000001",
  230=>"11111100",
  231=>"00000001",
  232=>"11111111",
  233=>"11111110",
  234=>"11111110",
  235=>"00000011",
  236=>"00000000",
  237=>"00000001",
  238=>"11111111",
  239=>"00000000",
  240=>"00000001",
  241=>"11111110",
  242=>"00000000",
  243=>"00000101",
  244=>"00000011",
  245=>"00000000",
  246=>"11111111",
  247=>"11111111",
  248=>"00000000",
  249=>"00000001",
  250=>"11111101",
  251=>"00000000",
  252=>"11111100",
  253=>"11111111",
  254=>"11111110",
  255=>"11111111",
  256=>"00000000",
  257=>"00000011",
  258=>"11111110",
  259=>"00000100",
  260=>"00000000",
  261=>"00000010",
  262=>"11111111",
  263=>"00000001",
  264=>"11111101",
  265=>"11111111",
  266=>"11111111",
  267=>"00000001",
  268=>"11111110",
  269=>"11111111",
  270=>"11111110",
  271=>"11111111",
  272=>"00000101",
  273=>"11111111",
  274=>"11111111",
  275=>"00000000",
  276=>"00000110",
  277=>"00000001",
  278=>"11111110",
  279=>"00000100",
  280=>"00000111",
  281=>"11111111",
  282=>"11111111",
  283=>"11111101",
  284=>"00000001",
  285=>"00000000",
  286=>"00000001",
  287=>"11111100",
  288=>"00000000",
  289=>"00001000",
  290=>"00000001",
  291=>"00000010",
  292=>"00000001",
  293=>"11111100",
  294=>"11111111",
  295=>"00000110",
  296=>"11111110",
  297=>"11111100",
  298=>"11111110",
  299=>"11111110",
  300=>"11111110",
  301=>"11111111",
  302=>"00000100",
  303=>"00000011",
  304=>"11111111",
  305=>"11111110",
  306=>"11111111",
  307=>"11111111",
  308=>"00000000",
  309=>"00000000",
  310=>"11111101",
  311=>"00000010",
  312=>"00000001",
  313=>"11111111",
  314=>"00000001",
  315=>"11111111",
  316=>"00000101",
  317=>"11111110",
  318=>"11111111",
  319=>"11111110",
  320=>"00000011",
  321=>"11111100",
  322=>"00000010",
  323=>"00000001",
  324=>"00000000",
  325=>"00000001",
  326=>"11111111",
  327=>"00000000",
  328=>"11111110",
  329=>"00000000",
  330=>"00000001",
  331=>"00000000",
  332=>"00000100",
  333=>"00000010",
  334=>"11111110",
  335=>"00000010",
  336=>"11111111",
  337=>"00000001",
  338=>"00000000",
  339=>"00000100",
  340=>"11111110",
  341=>"00000010",
  342=>"00000000",
  343=>"11111111",
  344=>"00000011",
  345=>"11111111",
  346=>"00000011",
  347=>"00000011",
  348=>"11111111",
  349=>"11111110",
  350=>"00000100",
  351=>"11111110",
  352=>"11111110",
  353=>"00000100",
  354=>"11111101",
  355=>"11111111",
  356=>"11111111",
  357=>"00000001",
  358=>"11111101",
  359=>"00000011",
  360=>"11111110",
  361=>"00000000",
  362=>"00000000",
  363=>"00000100",
  364=>"11111101",
  365=>"00000000",
  366=>"00000000",
  367=>"00000000",
  368=>"11111111",
  369=>"00000110",
  370=>"11111111",
  371=>"00000001",
  372=>"11111110",
  373=>"00000011",
  374=>"00000011",
  375=>"11111101",
  376=>"00000110",
  377=>"00000000",
  378=>"00000100",
  379=>"00000000",
  380=>"00000100",
  381=>"00000001",
  382=>"00000001",
  383=>"11111101",
  384=>"00000100",
  385=>"00000011",
  386=>"00000010",
  387=>"00000011",
  388=>"11111111",
  389=>"11111110",
  390=>"00000010",
  391=>"00000001",
  392=>"00000000",
  393=>"11111101",
  394=>"11111110",
  395=>"00000000",
  396=>"00000010",
  397=>"00000010",
  398=>"00000001",
  399=>"00000100",
  400=>"00000001",
  401=>"11111100",
  402=>"00000000",
  403=>"00000011",
  404=>"00000001",
  405=>"11111110",
  406=>"11111100",
  407=>"00000001",
  408=>"00000101",
  409=>"11111100",
  410=>"11111111",
  411=>"00000010",
  412=>"00000100",
  413=>"00000101",
  414=>"00000011",
  415=>"00000000",
  416=>"00000000",
  417=>"00000010",
  418=>"11111111",
  419=>"00000010",
  420=>"00000011",
  421=>"11111110",
  422=>"11111101",
  423=>"00000100",
  424=>"11111101",
  425=>"11111111",
  426=>"11111111",
  427=>"00000011",
  428=>"11111101",
  429=>"11111101",
  430=>"00000010",
  431=>"00000100",
  432=>"00000000",
  433=>"11111101",
  434=>"00000001",
  435=>"11111101",
  436=>"00000010",
  437=>"00000001",
  438=>"00000100",
  439=>"00000000",
  440=>"00000000",
  441=>"00000010",
  442=>"00000010",
  443=>"00000001",
  444=>"00000001",
  445=>"00000000",
  446=>"11111101",
  447=>"11111111",
  448=>"11111110",
  449=>"00000001",
  450=>"11111101",
  451=>"11111100",
  452=>"00000011",
  453=>"00000000",
  454=>"11111100",
  455=>"00000000",
  456=>"00000100",
  457=>"11111111",
  458=>"11111100",
  459=>"11111011",
  460=>"00000011",
  461=>"00000100",
  462=>"00000001",
  463=>"11111100",
  464=>"11111101",
  465=>"11111110",
  466=>"11111110",
  467=>"00000000",
  468=>"00000010",
  469=>"00000101",
  470=>"00000010",
  471=>"11111111",
  472=>"00000011",
  473=>"00000010",
  474=>"00000101",
  475=>"11111111",
  476=>"00000010",
  477=>"11111111",
  478=>"11111100",
  479=>"00000011",
  480=>"00000100",
  481=>"00000001",
  482=>"11111100",
  483=>"00000001",
  484=>"00000001",
  485=>"11111011",
  486=>"00000011",
  487=>"00000001",
  488=>"00000010",
  489=>"00000011",
  490=>"11111110",
  491=>"00000000",
  492=>"00000011",
  493=>"11111101",
  494=>"11111111",
  495=>"11111100",
  496=>"11111111",
  497=>"00000011",
  498=>"00000001",
  499=>"11111101",
  500=>"00000001",
  501=>"11111111",
  502=>"00000010",
  503=>"00000000",
  504=>"00000011",
  505=>"11111111",
  506=>"11111110",
  507=>"11111111",
  508=>"00000011",
  509=>"11111101",
  510=>"11111111",
  511=>"11111110",
  512=>"00000000",
  513=>"11111111",
  514=>"11111110",
  515=>"11111101",
  516=>"00000000",
  517=>"11111110",
  518=>"11111111",
  519=>"11111101",
  520=>"11111101",
  521=>"00000100",
  522=>"00000000",
  523=>"00000011",
  524=>"11111100",
  525=>"11111101",
  526=>"00000110",
  527=>"11111111",
  528=>"00000001",
  529=>"11111110",
  530=>"11111110",
  531=>"00000000",
  532=>"00000101",
  533=>"00000011",
  534=>"00000110",
  535=>"00000011",
  536=>"11111111",
  537=>"11111110",
  538=>"11111110",
  539=>"11111110",
  540=>"00000001",
  541=>"00000010",
  542=>"00000000",
  543=>"00000100",
  544=>"11111101",
  545=>"00000001",
  546=>"00000101",
  547=>"00000000",
  548=>"00000010",
  549=>"11111110",
  550=>"00000010",
  551=>"00000001",
  552=>"00000000",
  553=>"11111111",
  554=>"00000011",
  555=>"11111110",
  556=>"00000011",
  557=>"00000001",
  558=>"00000000",
  559=>"00000001",
  560=>"00000110",
  561=>"00000001",
  562=>"11111110",
  563=>"00000001",
  564=>"00000100",
  565=>"11111100",
  566=>"11111111",
  567=>"11111110",
  568=>"11111111",
  569=>"00000001",
  570=>"11111111",
  571=>"00000100",
  572=>"11111111",
  573=>"00000101",
  574=>"11111111",
  575=>"00000000",
  576=>"11111101",
  577=>"00000010",
  578=>"11111101",
  579=>"00000100",
  580=>"00000010",
  581=>"11111011",
  582=>"00000001",
  583=>"11111101",
  584=>"00000000",
  585=>"11111110",
  586=>"00000010",
  587=>"11111100",
  588=>"00000010",
  589=>"11111101",
  590=>"00000011",
  591=>"00000010",
  592=>"11111101",
  593=>"00000011",
  594=>"00000000",
  595=>"00000011",
  596=>"00000010",
  597=>"00000100",
  598=>"11111101",
  599=>"11111101",
  600=>"00000010",
  601=>"11111111",
  602=>"00000010",
  603=>"00000001",
  604=>"11111101",
  605=>"11111110",
  606=>"11111110",
  607=>"00000001",
  608=>"00000001",
  609=>"11111111",
  610=>"11111111",
  611=>"11111111",
  612=>"00000000",
  613=>"00000100",
  614=>"00000010",
  615=>"00000111",
  616=>"11111101",
  617=>"11111111",
  618=>"11111111",
  619=>"00000100",
  620=>"11111110",
  621=>"00000011",
  622=>"00000100",
  623=>"11111110",
  624=>"00000010",
  625=>"11111101",
  626=>"00000000",
  627=>"00000011",
  628=>"11111101",
  629=>"00000000",
  630=>"00000010",
  631=>"00000001",
  632=>"00000011",
  633=>"11111110",
  634=>"11111111",
  635=>"11111101",
  636=>"00000001",
  637=>"00000011",
  638=>"00000010",
  639=>"11111101",
  640=>"11111101",
  641=>"00000011",
  642=>"00000010",
  643=>"00000100",
  644=>"00000100",
  645=>"11111100",
  646=>"11111111",
  647=>"11111101",
  648=>"00000000",
  649=>"00000000",
  650=>"11111110",
  651=>"00000100",
  652=>"00000000",
  653=>"00000010",
  654=>"11111101",
  655=>"11111111",
  656=>"00000001",
  657=>"00000010",
  658=>"11111011",
  659=>"00000010",
  660=>"11111111",
  661=>"00000010",
  662=>"00000000",
  663=>"11111110",
  664=>"00000100",
  665=>"00000010",
  666=>"11111111",
  667=>"00000000",
  668=>"00000000",
  669=>"00000101",
  670=>"00000000",
  671=>"00000001",
  672=>"00000001",
  673=>"11111110",
  674=>"11111101",
  675=>"00000001",
  676=>"11111111",
  677=>"00000000",
  678=>"00000100",
  679=>"00000011",
  680=>"11111100",
  681=>"00000010",
  682=>"00000000",
  683=>"00000010",
  684=>"00000000",
  685=>"00000010",
  686=>"00000011",
  687=>"11111110",
  688=>"00000011",
  689=>"00000010",
  690=>"11111110",
  691=>"00000101",
  692=>"00000001",
  693=>"11111111",
  694=>"11111101",
  695=>"00000000",
  696=>"00000000",
  697=>"11111111",
  698=>"11111110",
  699=>"11111101",
  700=>"11111110",
  701=>"00000100",
  702=>"00000010",
  703=>"11111111",
  704=>"00000010",
  705=>"00000010",
  706=>"00000001",
  707=>"11111101",
  708=>"00000000",
  709=>"00000010",
  710=>"11111101",
  711=>"00000000",
  712=>"00000010",
  713=>"00000011",
  714=>"00000011",
  715=>"00000001",
  716=>"00000001",
  717=>"00000001",
  718=>"11111110",
  719=>"11111110",
  720=>"00000010",
  721=>"11111111",
  722=>"00000110",
  723=>"00000000",
  724=>"11111100",
  725=>"11111101",
  726=>"00000011",
  727=>"00000000",
  728=>"00000000",
  729=>"00000010",
  730=>"00000000",
  731=>"00000000",
  732=>"00000000",
  733=>"00000000",
  734=>"00000001",
  735=>"11111110",
  736=>"11111111",
  737=>"00000000",
  738=>"11111110",
  739=>"00000001",
  740=>"00000000",
  741=>"11111111",
  742=>"00000010",
  743=>"00000101",
  744=>"11111101",
  745=>"00000001",
  746=>"00000001",
  747=>"00000010",
  748=>"00000001",
  749=>"00000100",
  750=>"00000011",
  751=>"11111110",
  752=>"00000001",
  753=>"00000010",
  754=>"00000000",
  755=>"11111111",
  756=>"00000100",
  757=>"11111111",
  758=>"00000011",
  759=>"11111101",
  760=>"11111110",
  761=>"00000000",
  762=>"00000010",
  763=>"00000001",
  764=>"00000010",
  765=>"00000001",
  766=>"00000001",
  767=>"11111110",
  768=>"00000000",
  769=>"11111110",
  770=>"00000010",
  771=>"00000000",
  772=>"00000000",
  773=>"00000010",
  774=>"11111111",
  775=>"00000010",
  776=>"11111111",
  777=>"00000101",
  778=>"11111110",
  779=>"00001000",
  780=>"00000000",
  781=>"11111101",
  782=>"00000001",
  783=>"11111111",
  784=>"00000101",
  785=>"11111111",
  786=>"00000001",
  787=>"00000100",
  788=>"00000000",
  789=>"00000001",
  790=>"00000111",
  791=>"00000001",
  792=>"11111101",
  793=>"00000001",
  794=>"11111110",
  795=>"11111110",
  796=>"11111111",
  797=>"11111101",
  798=>"11111111",
  799=>"00000000",
  800=>"00000000",
  801=>"11111100",
  802=>"11111110",
  803=>"00000010",
  804=>"00000000",
  805=>"11111101",
  806=>"00000000",
  807=>"00000100",
  808=>"11111110",
  809=>"00000110",
  810=>"00000010",
  811=>"00000010",
  812=>"11111101",
  813=>"00000000",
  814=>"11111110",
  815=>"00000001",
  816=>"00000010",
  817=>"00000100",
  818=>"00000000",
  819=>"00000001",
  820=>"00000001",
  821=>"11111110",
  822=>"00000101",
  823=>"00000010",
  824=>"11111110",
  825=>"11111110",
  826=>"00000011",
  827=>"00000001",
  828=>"11111110",
  829=>"11111111",
  830=>"11111101",
  831=>"00000010",
  832=>"11111110",
  833=>"00000000",
  834=>"11111111",
  835=>"00000010",
  836=>"00000000",
  837=>"00000010",
  838=>"00000111",
  839=>"00000000",
  840=>"00000000",
  841=>"00000010",
  842=>"11111110",
  843=>"11111111",
  844=>"11111101",
  845=>"11111110",
  846=>"11111111",
  847=>"00000011",
  848=>"00000100",
  849=>"11111111",
  850=>"11111110",
  851=>"00000001",
  852=>"00000101",
  853=>"11111110",
  854=>"11111111",
  855=>"00000101",
  856=>"00000000",
  857=>"11111101",
  858=>"00000010",
  859=>"00000000",
  860=>"11111111",
  861=>"00000010",
  862=>"11111110",
  863=>"00000011",
  864=>"00000001",
  865=>"11111110",
  866=>"00000010",
  867=>"11111101",
  868=>"11111101",
  869=>"00000010",
  870=>"11111111",
  871=>"00000001",
  872=>"00000011",
  873=>"00000001",
  874=>"00000010",
  875=>"11111100",
  876=>"00000001",
  877=>"11111101",
  878=>"00000010",
  879=>"00000011",
  880=>"00000000",
  881=>"11111111",
  882=>"11111111",
  883=>"11111101",
  884=>"00000001",
  885=>"11111110",
  886=>"11111101",
  887=>"00000011",
  888=>"00000001",
  889=>"00000000",
  890=>"00000010",
  891=>"00000001",
  892=>"11111101",
  893=>"00000000",
  894=>"11111111",
  895=>"00000100",
  896=>"00000010",
  897=>"00000100",
  898=>"11111110",
  899=>"00000011",
  900=>"11111110",
  901=>"11111110",
  902=>"00000001",
  903=>"11111111",
  904=>"11111101",
  905=>"11111110",
  906=>"11111111",
  907=>"00000011",
  908=>"11111111",
  909=>"11111111",
  910=>"11111111",
  911=>"00000100",
  912=>"00000000",
  913=>"00000101",
  914=>"00000000",
  915=>"00000010",
  916=>"00000011",
  917=>"11111111",
  918=>"00000010",
  919=>"11111110",
  920=>"00000010",
  921=>"11111110",
  922=>"00000100",
  923=>"11111011",
  924=>"00000011",
  925=>"11111101",
  926=>"11111001",
  927=>"00000100",
  928=>"00000111",
  929=>"11111110",
  930=>"00000001",
  931=>"11111110",
  932=>"00000000",
  933=>"11111101",
  934=>"11111101",
  935=>"00000001",
  936=>"00000000",
  937=>"00000000",
  938=>"00000010",
  939=>"00000100",
  940=>"00000011",
  941=>"00000001",
  942=>"00000010",
  943=>"11111110",
  944=>"00000000",
  945=>"00000101",
  946=>"11111100",
  947=>"00000000",
  948=>"00000101",
  949=>"00000100",
  950=>"00000010",
  951=>"00000000",
  952=>"11111110",
  953=>"00000001",
  954=>"00000011",
  955=>"00000100",
  956=>"00000001",
  957=>"00000010",
  958=>"00000001",
  959=>"00000001",
  960=>"00000100",
  961=>"11111101",
  962=>"00000011",
  963=>"11111111",
  964=>"00000001",
  965=>"11111110",
  966=>"00000010",
  967=>"11111101",
  968=>"00000011",
  969=>"00000000",
  970=>"00000011",
  971=>"00000000",
  972=>"11111111",
  973=>"00000010",
  974=>"00000001",
  975=>"00000101",
  976=>"00000010",
  977=>"00000001",
  978=>"00000010",
  979=>"00000000",
  980=>"00000000",
  981=>"11111110",
  982=>"11111101",
  983=>"11111110",
  984=>"11111111",
  985=>"11111101",
  986=>"00000110",
  987=>"00000011",
  988=>"00000100",
  989=>"11111111",
  990=>"00000011",
  991=>"00000000",
  992=>"11111111",
  993=>"11111110",
  994=>"11111110",
  995=>"00000100",
  996=>"00000000",
  997=>"11111101",
  998=>"00000010",
  999=>"11111110",
  1000=>"00000010",
  1001=>"00000100",
  1002=>"00000100",
  1003=>"00000010",
  1004=>"00000010",
  1005=>"11111111",
  1006=>"11111110",
  1007=>"00000000",
  1008=>"00000000",
  1009=>"00000100",
  1010=>"00000001",
  1011=>"00000100",
  1012=>"00000001",
  1013=>"11111100",
  1014=>"00000000",
  1015=>"00000001",
  1016=>"11111110",
  1017=>"11111110",
  1018=>"11111110",
  1019=>"11111101",
  1020=>"11111111",
  1021=>"11111101",
  1022=>"00000010",
  1023=>"00000010",
  1024=>"11111111",
  1025=>"00000100",
  1026=>"00000001",
  1027=>"00000010",
  1028=>"11111100",
  1029=>"11111111",
  1030=>"11111110",
  1031=>"11111111",
  1032=>"11111110",
  1033=>"11111101",
  1034=>"00000001",
  1035=>"11111100",
  1036=>"00000000",
  1037=>"11111110",
  1038=>"00000000",
  1039=>"00000100",
  1040=>"00000000",
  1041=>"11111100",
  1042=>"00000010",
  1043=>"00000000",
  1044=>"11111110",
  1045=>"11111111",
  1046=>"00000000",
  1047=>"11111111",
  1048=>"00000000",
  1049=>"00000000",
  1050=>"11111111",
  1051=>"00000011",
  1052=>"00000011",
  1053=>"00000000",
  1054=>"00000000",
  1055=>"11111100",
  1056=>"11111110",
  1057=>"11111101",
  1058=>"00000110",
  1059=>"11111111",
  1060=>"00000001",
  1061=>"11111100",
  1062=>"00000010",
  1063=>"11111110",
  1064=>"11111110",
  1065=>"00000001",
  1066=>"11111101",
  1067=>"00000000",
  1068=>"00000100",
  1069=>"00000000",
  1070=>"00000010",
  1071=>"11111101",
  1072=>"00000000",
  1073=>"00000000",
  1074=>"00000010",
  1075=>"00000001",
  1076=>"00000010",
  1077=>"11111100",
  1078=>"11111110",
  1079=>"00000001",
  1080=>"00000000",
  1081=>"00000011",
  1082=>"11111111",
  1083=>"11111111",
  1084=>"11111110",
  1085=>"11111110",
  1086=>"11111111",
  1087=>"00000001",
  1088=>"00000000",
  1089=>"11111110",
  1090=>"11111101",
  1091=>"11111101",
  1092=>"00000000",
  1093=>"11111101",
  1094=>"11111110",
  1095=>"11111111",
  1096=>"00000000",
  1097=>"00000000",
  1098=>"11111101",
  1099=>"00000000",
  1100=>"11111101",
  1101=>"00000001",
  1102=>"00000001",
  1103=>"00000000",
  1104=>"00000000",
  1105=>"00000001",
  1106=>"00000001",
  1107=>"11111111",
  1108=>"11111111",
  1109=>"00000000",
  1110=>"00000010",
  1111=>"11111110",
  1112=>"11111111",
  1113=>"11111101",
  1114=>"00000000",
  1115=>"11111111",
  1116=>"11111110",
  1117=>"11111110",
  1118=>"11111111",
  1119=>"00000000",
  1120=>"11111111",
  1121=>"00000000",
  1122=>"00000001",
  1123=>"00000001",
  1124=>"00000000",
  1125=>"11111110",
  1126=>"11111111",
  1127=>"11111101",
  1128=>"00000010",
  1129=>"11111110",
  1130=>"00000001",
  1131=>"00000011",
  1132=>"11111100",
  1133=>"11111111",
  1134=>"11111111",
  1135=>"00000001",
  1136=>"11111111",
  1137=>"00000000",
  1138=>"00000010",
  1139=>"00000000",
  1140=>"11111110",
  1141=>"00000000",
  1142=>"00000111",
  1143=>"11111110",
  1144=>"11111010",
  1145=>"11111111",
  1146=>"11111101",
  1147=>"11111111",
  1148=>"00000011",
  1149=>"11111111",
  1150=>"11111110",
  1151=>"00000100",
  1152=>"00000100",
  1153=>"11111101",
  1154=>"00000000",
  1155=>"00000000",
  1156=>"11111111",
  1157=>"00000001",
  1158=>"00000001",
  1159=>"11111101",
  1160=>"11111101",
  1161=>"00000001",
  1162=>"11111101",
  1163=>"11111110",
  1164=>"11111101",
  1165=>"11111111",
  1166=>"00000011",
  1167=>"11111110",
  1168=>"11111110",
  1169=>"00000000",
  1170=>"00000011",
  1171=>"11111111",
  1172=>"00000001",
  1173=>"11111111",
  1174=>"00000011",
  1175=>"00000000",
  1176=>"11111101",
  1177=>"00000011",
  1178=>"00000101",
  1179=>"00000000",
  1180=>"11111110",
  1181=>"11111101",
  1182=>"00000010",
  1183=>"11111101",
  1184=>"11111110",
  1185=>"11111110",
  1186=>"11111111",
  1187=>"00000000",
  1188=>"11111110",
  1189=>"11111111",
  1190=>"00000001",
  1191=>"11111101",
  1192=>"00000010",
  1193=>"00000011",
  1194=>"00000001",
  1195=>"11111101",
  1196=>"00000011",
  1197=>"11111111",
  1198=>"11111110",
  1199=>"00000011",
  1200=>"11111111",
  1201=>"11111100",
  1202=>"11111100",
  1203=>"00000010",
  1204=>"00000000",
  1205=>"00000010",
  1206=>"11111111",
  1207=>"11111110",
  1208=>"00000101",
  1209=>"11111111",
  1210=>"00000110",
  1211=>"11111100",
  1212=>"00000001",
  1213=>"00000000",
  1214=>"11111110",
  1215=>"00000001",
  1216=>"00000100",
  1217=>"00000010",
  1218=>"11111111",
  1219=>"00000100",
  1220=>"11111111",
  1221=>"11111110",
  1222=>"11111101",
  1223=>"11111101",
  1224=>"11111100",
  1225=>"00000010",
  1226=>"11111110",
  1227=>"00000001",
  1228=>"11111110",
  1229=>"00000010",
  1230=>"00000000",
  1231=>"00000000",
  1232=>"00000001",
  1233=>"00000010",
  1234=>"11111111",
  1235=>"00000010",
  1236=>"11111111",
  1237=>"00000011",
  1238=>"00000011",
  1239=>"00000001",
  1240=>"11111111",
  1241=>"00000001",
  1242=>"11111111",
  1243=>"00000010",
  1244=>"11111111",
  1245=>"00000001",
  1246=>"00000101",
  1247=>"11111110",
  1248=>"00000000",
  1249=>"11111111",
  1250=>"11111111",
  1251=>"00000001",
  1252=>"11111111",
  1253=>"11111111",
  1254=>"11111101",
  1255=>"00000001",
  1256=>"11111110",
  1257=>"11111110",
  1258=>"00000001",
  1259=>"00000000",
  1260=>"00000010",
  1261=>"11111110",
  1262=>"11111101",
  1263=>"00000001",
  1264=>"00000011",
  1265=>"00000110",
  1266=>"11111111",
  1267=>"11111110",
  1268=>"00000000",
  1269=>"11111111",
  1270=>"11111111",
  1271=>"00000010",
  1272=>"00000100",
  1273=>"00000010",
  1274=>"00000110",
  1275=>"00000000",
  1276=>"00000000",
  1277=>"00000000",
  1278=>"00000010",
  1279=>"11111101",
  1280=>"00000010",
  1281=>"00000011",
  1282=>"00000011",
  1283=>"11111111",
  1284=>"00000000",
  1285=>"00000010",
  1286=>"00000000",
  1287=>"00000000",
  1288=>"11111111",
  1289=>"11111101",
  1290=>"00000000",
  1291=>"11111111",
  1292=>"11111110",
  1293=>"11111111",
  1294=>"11111110",
  1295=>"00000100",
  1296=>"00000100",
  1297=>"11111111",
  1298=>"11111110",
  1299=>"00000001",
  1300=>"00000000",
  1301=>"00000010",
  1302=>"11111111",
  1303=>"00000000",
  1304=>"00000000",
  1305=>"11111101",
  1306=>"11111110",
  1307=>"11111111",
  1308=>"00000000",
  1309=>"00000001",
  1310=>"11111111",
  1311=>"00000011",
  1312=>"00000000",
  1313=>"11111110",
  1314=>"11111111",
  1315=>"00000011",
  1316=>"11111101",
  1317=>"00000000",
  1318=>"00000000",
  1319=>"11111111",
  1320=>"00000010",
  1321=>"00000010",
  1322=>"00000010",
  1323=>"11111101",
  1324=>"11111110",
  1325=>"00000010",
  1326=>"11111100",
  1327=>"00000101",
  1328=>"00000000",
  1329=>"11111111",
  1330=>"11111111",
  1331=>"11111101",
  1332=>"00000010",
  1333=>"00000001",
  1334=>"00000010",
  1335=>"00000001",
  1336=>"11111101",
  1337=>"00000100",
  1338=>"11111101",
  1339=>"00000100",
  1340=>"11111111",
  1341=>"11111111",
  1342=>"00000000",
  1343=>"11111101",
  1344=>"00000010",
  1345=>"00000110",
  1346=>"00000010",
  1347=>"11111110",
  1348=>"00000000",
  1349=>"11111110",
  1350=>"00000110",
  1351=>"11111110",
  1352=>"00000100",
  1353=>"11111111",
  1354=>"11111110",
  1355=>"11111101",
  1356=>"11111111",
  1357=>"11111111",
  1358=>"11111100",
  1359=>"11111011",
  1360=>"00000010",
  1361=>"11111111",
  1362=>"11111110",
  1363=>"11111111",
  1364=>"11111111",
  1365=>"11111101",
  1366=>"00000000",
  1367=>"00000001",
  1368=>"00000010",
  1369=>"00000000",
  1370=>"11111110",
  1371=>"11111110",
  1372=>"00000010",
  1373=>"00000010",
  1374=>"11111111",
  1375=>"00000110",
  1376=>"00000000",
  1377=>"11111111",
  1378=>"00000001",
  1379=>"00000000",
  1380=>"00000000",
  1381=>"00000000",
  1382=>"00000010",
  1383=>"00000001",
  1384=>"11111110",
  1385=>"11111110",
  1386=>"00000001",
  1387=>"00000101",
  1388=>"11111110",
  1389=>"00000000",
  1390=>"00000000",
  1391=>"11111101",
  1392=>"11111110",
  1393=>"11111100",
  1394=>"00000001",
  1395=>"11111111",
  1396=>"11111101",
  1397=>"11111100",
  1398=>"00000010",
  1399=>"00000011",
  1400=>"11111111",
  1401=>"11111100",
  1402=>"11111111",
  1403=>"11111110",
  1404=>"00000001",
  1405=>"00000011",
  1406=>"11111101",
  1407=>"11111111",
  1408=>"11111111",
  1409=>"00000100",
  1410=>"00000011",
  1411=>"00000001",
  1412=>"00000001",
  1413=>"11111111",
  1414=>"11111111",
  1415=>"00000000",
  1416=>"00000000",
  1417=>"11111110",
  1418=>"00000101",
  1419=>"11111110",
  1420=>"00000010",
  1421=>"00000000",
  1422=>"11111110",
  1423=>"00000010",
  1424=>"11111111",
  1425=>"00000010",
  1426=>"00000001",
  1427=>"00000000",
  1428=>"00000001",
  1429=>"11111110",
  1430=>"00000000",
  1431=>"00000000",
  1432=>"11111101",
  1433=>"00000101",
  1434=>"11111111",
  1435=>"11111110",
  1436=>"00000010",
  1437=>"00000101",
  1438=>"00000001",
  1439=>"00001001",
  1440=>"00000001",
  1441=>"00000000",
  1442=>"00000110",
  1443=>"11111101",
  1444=>"11111111",
  1445=>"11111101",
  1446=>"11111111",
  1447=>"00000011",
  1448=>"11111110",
  1449=>"00000010",
  1450=>"11111110",
  1451=>"11111100",
  1452=>"11111110",
  1453=>"11111111",
  1454=>"11111101",
  1455=>"00000001",
  1456=>"11111101",
  1457=>"11111111",
  1458=>"11111111",
  1459=>"11111101",
  1460=>"00000000",
  1461=>"00000001",
  1462=>"00000001",
  1463=>"00000011",
  1464=>"00000001",
  1465=>"11111110",
  1466=>"11111110",
  1467=>"00000000",
  1468=>"11111110",
  1469=>"00000111",
  1470=>"00000010",
  1471=>"00000011",
  1472=>"00000000",
  1473=>"11111101",
  1474=>"11111101",
  1475=>"00000100",
  1476=>"11111111",
  1477=>"11111111",
  1478=>"00000001",
  1479=>"00000011",
  1480=>"11111101",
  1481=>"00000010",
  1482=>"00000001",
  1483=>"11111111",
  1484=>"11111101",
  1485=>"00000001",
  1486=>"11111110",
  1487=>"11111110",
  1488=>"11111111",
  1489=>"00000001",
  1490=>"11111110",
  1491=>"00000101",
  1492=>"00000000",
  1493=>"00000001",
  1494=>"00000011",
  1495=>"11111110",
  1496=>"11111111",
  1497=>"11111100",
  1498=>"00000001",
  1499=>"11111110",
  1500=>"00000001",
  1501=>"11111110",
  1502=>"11111101",
  1503=>"11111111",
  1504=>"11111111",
  1505=>"11111111",
  1506=>"11111111",
  1507=>"00000001",
  1508=>"00000001",
  1509=>"11111110",
  1510=>"11111111",
  1511=>"00000011",
  1512=>"11111100",
  1513=>"11111111",
  1514=>"11111111",
  1515=>"11111110",
  1516=>"00000001",
  1517=>"11111111",
  1518=>"11111111",
  1519=>"00000010",
  1520=>"11111110",
  1521=>"00000000",
  1522=>"00000000",
  1523=>"00000001",
  1524=>"00000011",
  1525=>"00000000",
  1526=>"00000010",
  1527=>"11111101",
  1528=>"11111111",
  1529=>"00000010",
  1530=>"11111111",
  1531=>"11111111",
  1532=>"11111101",
  1533=>"00000010",
  1534=>"11111100",
  1535=>"00000010",
  1536=>"11111101",
  1537=>"11111111",
  1538=>"11111110",
  1539=>"00000010",
  1540=>"00000000",
  1541=>"00000010",
  1542=>"00000000",
  1543=>"00000010",
  1544=>"11111111",
  1545=>"11111111",
  1546=>"00000010",
  1547=>"00000000",
  1548=>"11111111",
  1549=>"11111111",
  1550=>"11111101",
  1551=>"00000011",
  1552=>"11111111",
  1553=>"00000011",
  1554=>"11111111",
  1555=>"11111100",
  1556=>"11111101",
  1557=>"11111111",
  1558=>"11111111",
  1559=>"00000011",
  1560=>"11111100",
  1561=>"00000111",
  1562=>"00000001",
  1563=>"11111101",
  1564=>"00000000",
  1565=>"11111111",
  1566=>"00000000",
  1567=>"00000000",
  1568=>"00000000",
  1569=>"00000010",
  1570=>"00000000",
  1571=>"11111110",
  1572=>"00000001",
  1573=>"11111110",
  1574=>"11111110",
  1575=>"00000010",
  1576=>"11111110",
  1577=>"11111101",
  1578=>"00000010",
  1579=>"00000010",
  1580=>"11111111",
  1581=>"11111111",
  1582=>"11111111",
  1583=>"00000000",
  1584=>"11111111",
  1585=>"00000001",
  1586=>"11111101",
  1587=>"00000010",
  1588=>"11111110",
  1589=>"11111111",
  1590=>"00000010",
  1591=>"11111110",
  1592=>"11111111",
  1593=>"11111110",
  1594=>"11111111",
  1595=>"00000001",
  1596=>"00000011",
  1597=>"11111011",
  1598=>"00000000",
  1599=>"00000000",
  1600=>"00000010",
  1601=>"00000101",
  1602=>"11111101",
  1603=>"00000011",
  1604=>"11111101",
  1605=>"11111110",
  1606=>"00000000",
  1607=>"11111111",
  1608=>"11111111",
  1609=>"11111101",
  1610=>"11111101",
  1611=>"00000000",
  1612=>"00000011",
  1613=>"00000001",
  1614=>"00000000",
  1615=>"11111111",
  1616=>"00000000",
  1617=>"00000000",
  1618=>"00000000",
  1619=>"00000001",
  1620=>"11111110",
  1621=>"11111101",
  1622=>"11111111",
  1623=>"00000000",
  1624=>"11111110",
  1625=>"00000000",
  1626=>"11111111",
  1627=>"00000101",
  1628=>"00000101",
  1629=>"00000010",
  1630=>"11111111",
  1631=>"11111110",
  1632=>"00000001",
  1633=>"00000000",
  1634=>"11111101",
  1635=>"11111101",
  1636=>"00000001",
  1637=>"00000011",
  1638=>"00000000",
  1639=>"11111100",
  1640=>"00000111",
  1641=>"00000001",
  1642=>"00000010",
  1643=>"00000001",
  1644=>"11111110",
  1645=>"11111111",
  1646=>"11111101",
  1647=>"11111110",
  1648=>"11111101",
  1649=>"00000000",
  1650=>"00000001",
  1651=>"11111101",
  1652=>"00000000",
  1653=>"11111110",
  1654=>"00000000",
  1655=>"11111111",
  1656=>"00000001",
  1657=>"00000011",
  1658=>"00000000",
  1659=>"11111110",
  1660=>"00000001",
  1661=>"11111110",
  1662=>"11111111",
  1663=>"00000001",
  1664=>"00000001",
  1665=>"00000011",
  1666=>"00000000",
  1667=>"11111110",
  1668=>"00000001",
  1669=>"11111101",
  1670=>"11111111",
  1671=>"00000000",
  1672=>"00000010",
  1673=>"00000000",
  1674=>"11111110",
  1675=>"11111111",
  1676=>"00000010",
  1677=>"11111111",
  1678=>"11111110",
  1679=>"00000100",
  1680=>"00000001",
  1681=>"11111111",
  1682=>"11111101",
  1683=>"11111111",
  1684=>"11111111",
  1685=>"00000000",
  1686=>"11111111",
  1687=>"11111101",
  1688=>"00000001",
  1689=>"11111100",
  1690=>"00000000",
  1691=>"00000000",
  1692=>"11111110",
  1693=>"11111101",
  1694=>"11111110",
  1695=>"11111100",
  1696=>"11111110",
  1697=>"00000011",
  1698=>"00000000",
  1699=>"00000000",
  1700=>"11111110",
  1701=>"11111110",
  1702=>"11111101",
  1703=>"11111011",
  1704=>"00000000",
  1705=>"00000000",
  1706=>"00000000",
  1707=>"00000000",
  1708=>"11111111",
  1709=>"00000010",
  1710=>"00000000",
  1711=>"11111101",
  1712=>"11111101",
  1713=>"00000010",
  1714=>"00000000",
  1715=>"00000000",
  1716=>"11111110",
  1717=>"00000000",
  1718=>"00000001",
  1719=>"00000101",
  1720=>"00000001",
  1721=>"11111111",
  1722=>"11111111",
  1723=>"11111110",
  1724=>"00000000",
  1725=>"11111110",
  1726=>"00000000",
  1727=>"00000001",
  1728=>"11111111",
  1729=>"00000010",
  1730=>"00000010",
  1731=>"00000001",
  1732=>"11111110",
  1733=>"00000010",
  1734=>"00000001",
  1735=>"00000001",
  1736=>"11111111",
  1737=>"11111110",
  1738=>"11111110",
  1739=>"00000000",
  1740=>"11111101",
  1741=>"00000100",
  1742=>"00000000",
  1743=>"00000000",
  1744=>"11111111",
  1745=>"11111110",
  1746=>"11111100",
  1747=>"00000000",
  1748=>"00000010",
  1749=>"00000001",
  1750=>"11111111",
  1751=>"00000001",
  1752=>"11111101",
  1753=>"00000000",
  1754=>"11111110",
  1755=>"11111111",
  1756=>"11111101",
  1757=>"00000000",
  1758=>"11111111",
  1759=>"00000001",
  1760=>"00000000",
  1761=>"11111101",
  1762=>"00000001",
  1763=>"00000000",
  1764=>"00000010",
  1765=>"11111110",
  1766=>"11111111",
  1767=>"11111111",
  1768=>"11111110",
  1769=>"00000001",
  1770=>"11111100",
  1771=>"00000000",
  1772=>"00000000",
  1773=>"00000001",
  1774=>"00000001",
  1775=>"00000011",
  1776=>"00000001",
  1777=>"00000101",
  1778=>"11111111",
  1779=>"00000011",
  1780=>"00000010",
  1781=>"00000010",
  1782=>"00000000",
  1783=>"00000011",
  1784=>"11111111",
  1785=>"00000001",
  1786=>"00000000",
  1787=>"11111100",
  1788=>"11111111",
  1789=>"00000011",
  1790=>"00000011",
  1791=>"00000010",
  1792=>"00000001",
  1793=>"00000000",
  1794=>"11111111",
  1795=>"00000100",
  1796=>"00000000",
  1797=>"11111101",
  1798=>"11111110",
  1799=>"11111101",
  1800=>"11111100",
  1801=>"11111110",
  1802=>"00000000",
  1803=>"00000010",
  1804=>"11111111",
  1805=>"11111111",
  1806=>"00000000",
  1807=>"00000010",
  1808=>"11111101",
  1809=>"11111101",
  1810=>"00000000",
  1811=>"00000011",
  1812=>"00000010",
  1813=>"11111110",
  1814=>"00000010",
  1815=>"00000000",
  1816=>"11111110",
  1817=>"00000010",
  1818=>"00000000",
  1819=>"11111111",
  1820=>"11111111",
  1821=>"00000100",
  1822=>"11111110",
  1823=>"11111101",
  1824=>"11111110",
  1825=>"00000001",
  1826=>"00000010",
  1827=>"00000001",
  1828=>"11111101",
  1829=>"11111110",
  1830=>"00000011",
  1831=>"11111101",
  1832=>"00000000",
  1833=>"11111101",
  1834=>"00000010",
  1835=>"00000000",
  1836=>"00000001",
  1837=>"11111111",
  1838=>"11111111",
  1839=>"11111100",
  1840=>"00000001",
  1841=>"11111101",
  1842=>"00000110",
  1843=>"11111110",
  1844=>"11111111",
  1845=>"00000001",
  1846=>"11111101",
  1847=>"11111111",
  1848=>"00000101",
  1849=>"00000001",
  1850=>"11111101",
  1851=>"11111110",
  1852=>"11111111",
  1853=>"00000001",
  1854=>"11111101",
  1855=>"11111111",
  1856=>"11111111",
  1857=>"11111100",
  1858=>"11111110",
  1859=>"00000000",
  1860=>"11111110",
  1861=>"00000001",
  1862=>"00000001",
  1863=>"00000000",
  1864=>"11111110",
  1865=>"11111111",
  1866=>"00000000",
  1867=>"00000101",
  1868=>"00000001",
  1869=>"00000001",
  1870=>"00000010",
  1871=>"00000000",
  1872=>"00000010",
  1873=>"00000011",
  1874=>"00000001",
  1875=>"11111110",
  1876=>"00000000",
  1877=>"00000010",
  1878=>"00000010",
  1879=>"11111111",
  1880=>"11111111",
  1881=>"00000010",
  1882=>"11111111",
  1883=>"00000101",
  1884=>"00000000",
  1885=>"00000010",
  1886=>"11111101",
  1887=>"11111101",
  1888=>"00000010",
  1889=>"11111111",
  1890=>"00000001",
  1891=>"11111101",
  1892=>"00000011",
  1893=>"11111111",
  1894=>"00000010",
  1895=>"11111101",
  1896=>"00000011",
  1897=>"11111101",
  1898=>"11111110",
  1899=>"00000010",
  1900=>"11111101",
  1901=>"00000101",
  1902=>"00000000",
  1903=>"00000001",
  1904=>"00000001",
  1905=>"11111100",
  1906=>"11111110",
  1907=>"11111110",
  1908=>"00000001",
  1909=>"11111101",
  1910=>"00000010",
  1911=>"11111110",
  1912=>"11111100",
  1913=>"00000001",
  1914=>"11111101",
  1915=>"00000000",
  1916=>"00000010",
  1917=>"11111110",
  1918=>"00000011",
  1919=>"11111101",
  1920=>"11111111",
  1921=>"11111110",
  1922=>"11111110",
  1923=>"11111110",
  1924=>"00000010",
  1925=>"11111110",
  1926=>"00000001",
  1927=>"00000011",
  1928=>"11111111",
  1929=>"00000000",
  1930=>"00000001",
  1931=>"00000001",
  1932=>"11111110",
  1933=>"11111101",
  1934=>"00000011",
  1935=>"11111110",
  1936=>"11111101",
  1937=>"00000000",
  1938=>"00000100",
  1939=>"00000001",
  1940=>"00000001",
  1941=>"00000000",
  1942=>"11111110",
  1943=>"00000100",
  1944=>"11111110",
  1945=>"11111101",
  1946=>"11111110",
  1947=>"00000001",
  1948=>"11111110",
  1949=>"00000011",
  1950=>"00000100",
  1951=>"00000001",
  1952=>"11111110",
  1953=>"11111110",
  1954=>"11111110",
  1955=>"11111111",
  1956=>"00000000",
  1957=>"11111111",
  1958=>"11111100",
  1959=>"00000011",
  1960=>"00000010",
  1961=>"00000001",
  1962=>"11111111",
  1963=>"11111111",
  1964=>"00000001",
  1965=>"00000111",
  1966=>"00000001",
  1967=>"00000010",
  1968=>"11111111",
  1969=>"11111110",
  1970=>"00000011",
  1971=>"00000000",
  1972=>"11111110",
  1973=>"00000101",
  1974=>"11111110",
  1975=>"11111110",
  1976=>"11111101",
  1977=>"11111111",
  1978=>"11111110",
  1979=>"11111111",
  1980=>"11111111",
  1981=>"11111100",
  1982=>"11111110",
  1983=>"00000010",
  1984=>"00000000",
  1985=>"11111111",
  1986=>"11111101",
  1987=>"00000010",
  1988=>"00000001",
  1989=>"11111101",
  1990=>"00000000",
  1991=>"00000001",
  1992=>"11111101",
  1993=>"11111110",
  1994=>"11111110",
  1995=>"11111101",
  1996=>"11111110",
  1997=>"00000001",
  1998=>"11111101",
  1999=>"00000010",
  2000=>"11111110",
  2001=>"00000001",
  2002=>"11111111",
  2003=>"00000000",
  2004=>"00000001",
  2005=>"11111111",
  2006=>"11111100",
  2007=>"00000010",
  2008=>"00000010",
  2009=>"11111110",
  2010=>"11111101",
  2011=>"11111111",
  2012=>"00000000",
  2013=>"11111110",
  2014=>"11111101",
  2015=>"00000100",
  2016=>"11111111",
  2017=>"11111110",
  2018=>"00000000",
  2019=>"00000010",
  2020=>"11111111",
  2021=>"11111101",
  2022=>"00000011",
  2023=>"00000000",
  2024=>"11111111",
  2025=>"00000001",
  2026=>"11111111",
  2027=>"11111110",
  2028=>"00000000",
  2029=>"00000010",
  2030=>"00000000",
  2031=>"00000111",
  2032=>"11111110",
  2033=>"00000100",
  2034=>"11111111",
  2035=>"00000001",
  2036=>"11111110",
  2037=>"00000001",
  2038=>"00000001",
  2039=>"11111101",
  2040=>"00000000",
  2041=>"00000010",
  2042=>"00000000",
  2043=>"11111110",
  2044=>"11111110",
  2045=>"00000001",
  2046=>"00000001",
  2047=>"11111110",
  2048=>"00000010",
  2049=>"00000000",
  2050=>"00000010",
  2051=>"11111111",
  2052=>"00000000",
  2053=>"11111111",
  2054=>"00000010",
  2055=>"11111111",
  2056=>"11111101",
  2057=>"11111111",
  2058=>"00000010",
  2059=>"00000000",
  2060=>"00000010",
  2061=>"11111110",
  2062=>"00000011",
  2063=>"11111110",
  2064=>"11111110",
  2065=>"11111100",
  2066=>"11111110",
  2067=>"11111111",
  2068=>"00000010",
  2069=>"00000011",
  2070=>"00000001",
  2071=>"00000000",
  2072=>"00000010",
  2073=>"00000000",
  2074=>"00000010",
  2075=>"11111110",
  2076=>"11111110",
  2077=>"00000010",
  2078=>"00000010",
  2079=>"11111110",
  2080=>"11111100",
  2081=>"11111110",
  2082=>"00000000",
  2083=>"00000000",
  2084=>"00000001",
  2085=>"00000000",
  2086=>"00000001",
  2087=>"00000001",
  2088=>"00000001",
  2089=>"00000000",
  2090=>"11111111",
  2091=>"00000100",
  2092=>"00000100",
  2093=>"00000011",
  2094=>"00000011",
  2095=>"11111101",
  2096=>"00000000",
  2097=>"11111110",
  2098=>"11111111",
  2099=>"00000100",
  2100=>"11111110",
  2101=>"11111111",
  2102=>"11111111",
  2103=>"00000010",
  2104=>"00000010",
  2105=>"11111110",
  2106=>"11111101",
  2107=>"00000100",
  2108=>"00000010",
  2109=>"00000001",
  2110=>"11111101",
  2111=>"00000001",
  2112=>"00000001",
  2113=>"00000000",
  2114=>"11111111",
  2115=>"00000000",
  2116=>"11111110",
  2117=>"11111110",
  2118=>"11111100",
  2119=>"00000010",
  2120=>"00000001",
  2121=>"00000000",
  2122=>"00000011",
  2123=>"00000001",
  2124=>"00000000",
  2125=>"00000000",
  2126=>"00000001",
  2127=>"00000001",
  2128=>"00000010",
  2129=>"11111110",
  2130=>"11111110",
  2131=>"00000111",
  2132=>"00000001",
  2133=>"00000001",
  2134=>"00000100",
  2135=>"11111111",
  2136=>"00000011",
  2137=>"11111111",
  2138=>"11111110",
  2139=>"00000001",
  2140=>"00000010",
  2141=>"11111101",
  2142=>"00000000",
  2143=>"00000101",
  2144=>"00000001",
  2145=>"00000001",
  2146=>"11111100",
  2147=>"00000001",
  2148=>"00000011",
  2149=>"11111110",
  2150=>"00000000",
  2151=>"00000001",
  2152=>"00000011",
  2153=>"11111101",
  2154=>"11111110",
  2155=>"11111111",
  2156=>"00000010",
  2157=>"11111101",
  2158=>"00000010",
  2159=>"00000000",
  2160=>"11111110",
  2161=>"00000000",
  2162=>"00000001",
  2163=>"00000010",
  2164=>"11111111",
  2165=>"11111111",
  2166=>"00000010",
  2167=>"11111110",
  2168=>"11111110",
  2169=>"11111101",
  2170=>"00000010",
  2171=>"11111101",
  2172=>"11111101",
  2173=>"11111110",
  2174=>"00000001",
  2175=>"00000000",
  2176=>"11111100",
  2177=>"00000010",
  2178=>"00000000",
  2179=>"00000011",
  2180=>"11111101",
  2181=>"00000100",
  2182=>"00000001",
  2183=>"00000100",
  2184=>"11111111",
  2185=>"00000011",
  2186=>"11111110",
  2187=>"00000011",
  2188=>"11111100",
  2189=>"11111111",
  2190=>"11111111",
  2191=>"11111111",
  2192=>"00000001",
  2193=>"00000011",
  2194=>"11111110",
  2195=>"00000011",
  2196=>"00000010",
  2197=>"11111101",
  2198=>"11111111",
  2199=>"11111111",
  2200=>"11111101",
  2201=>"11111101",
  2202=>"11111110",
  2203=>"11111110",
  2204=>"00000000",
  2205=>"00000001",
  2206=>"00000011",
  2207=>"11111111",
  2208=>"00000001",
  2209=>"00000000",
  2210=>"00000000",
  2211=>"00000000",
  2212=>"11111110",
  2213=>"00000100",
  2214=>"11111110",
  2215=>"11111110",
  2216=>"00000011",
  2217=>"00000001",
  2218=>"11111101",
  2219=>"00000010",
  2220=>"00000010",
  2221=>"11111110",
  2222=>"11111110",
  2223=>"11111111",
  2224=>"00000010",
  2225=>"11111111",
  2226=>"00000000",
  2227=>"00000001",
  2228=>"11111110",
  2229=>"11111111",
  2230=>"00000100",
  2231=>"00000001",
  2232=>"11111111",
  2233=>"11111101",
  2234=>"00000001",
  2235=>"00000010",
  2236=>"00000011",
  2237=>"00000001",
  2238=>"11111111",
  2239=>"11111110",
  2240=>"00000011",
  2241=>"00000001",
  2242=>"00000011",
  2243=>"11111110",
  2244=>"00000001",
  2245=>"11111110",
  2246=>"00000000",
  2247=>"00000001",
  2248=>"00000011",
  2249=>"00000001",
  2250=>"11111111",
  2251=>"00000000",
  2252=>"00000101",
  2253=>"00000001",
  2254=>"11111110",
  2255=>"00000100",
  2256=>"00000001",
  2257=>"11111110",
  2258=>"00000000",
  2259=>"11111111",
  2260=>"00000001",
  2261=>"00000010",
  2262=>"00000011",
  2263=>"11111110",
  2264=>"00000001",
  2265=>"11111111",
  2266=>"11111110",
  2267=>"11111111",
  2268=>"11111101",
  2269=>"00000000",
  2270=>"00000010",
  2271=>"11111110",
  2272=>"11111101",
  2273=>"00000001",
  2274=>"11111110",
  2275=>"00000001",
  2276=>"00000001",
  2277=>"00000100",
  2278=>"11111100",
  2279=>"00000010",
  2280=>"00000001",
  2281=>"11111111",
  2282=>"00000000",
  2283=>"00000000",
  2284=>"11111101",
  2285=>"00000001",
  2286=>"11111111",
  2287=>"00000011",
  2288=>"00000111",
  2289=>"00000010",
  2290=>"00000001",
  2291=>"11111111",
  2292=>"11111111",
  2293=>"11111111",
  2294=>"00000011",
  2295=>"11111101",
  2296=>"00000001",
  2297=>"00000100",
  2298=>"11111111",
  2299=>"00000001",
  2300=>"11111110",
  2301=>"11111111",
  2302=>"00000000",
  2303=>"00000000",
  2304=>"11111110",
  2305=>"00000100",
  2306=>"11111100",
  2307=>"00000011",
  2308=>"00000010",
  2309=>"11111110",
  2310=>"00000010",
  2311=>"00000000",
  2312=>"11111111",
  2313=>"11111101",
  2314=>"00000010",
  2315=>"00000001",
  2316=>"00000010",
  2317=>"00000001",
  2318=>"00000000",
  2319=>"00000001",
  2320=>"11111110",
  2321=>"00000100",
  2322=>"11111111",
  2323=>"11111111",
  2324=>"00000110",
  2325=>"00000011",
  2326=>"00000010",
  2327=>"00000010",
  2328=>"00000011",
  2329=>"11111111",
  2330=>"11111110",
  2331=>"11111111",
  2332=>"00000001",
  2333=>"00000001",
  2334=>"00000001",
  2335=>"00000000",
  2336=>"00000010",
  2337=>"00000001",
  2338=>"00000001",
  2339=>"00000000",
  2340=>"00000101",
  2341=>"11111111",
  2342=>"11111101",
  2343=>"00000001",
  2344=>"00000000",
  2345=>"00000011",
  2346=>"11111110",
  2347=>"11111111",
  2348=>"11111110",
  2349=>"00000001",
  2350=>"11111110",
  2351=>"11111111",
  2352=>"00000000",
  2353=>"11111111",
  2354=>"11111111",
  2355=>"11111111",
  2356=>"11111111",
  2357=>"00000011",
  2358=>"00000011",
  2359=>"11111110",
  2360=>"11111110",
  2361=>"11111110",
  2362=>"00000000",
  2363=>"11111111",
  2364=>"00000011",
  2365=>"00000000",
  2366=>"11111111",
  2367=>"00000001",
  2368=>"11111111",
  2369=>"00000010",
  2370=>"11111111",
  2371=>"11111111",
  2372=>"11111111",
  2373=>"11111111",
  2374=>"00000011",
  2375=>"11111101",
  2376=>"11111110",
  2377=>"11111101",
  2378=>"00000011",
  2379=>"00000000",
  2380=>"00000011",
  2381=>"00000001",
  2382=>"00000010",
  2383=>"11111110",
  2384=>"11111101",
  2385=>"11111101",
  2386=>"00000001",
  2387=>"11111110",
  2388=>"11111110",
  2389=>"00000000",
  2390=>"11111111",
  2391=>"11111110",
  2392=>"00000000",
  2393=>"11111110",
  2394=>"00000010",
  2395=>"00000001",
  2396=>"00000001",
  2397=>"11111111",
  2398=>"11111110",
  2399=>"11111101",
  2400=>"11111110",
  2401=>"11111111",
  2402=>"00000000",
  2403=>"00000011",
  2404=>"00000010",
  2405=>"00000000",
  2406=>"00000011",
  2407=>"11111101",
  2408=>"00000000",
  2409=>"00000000",
  2410=>"00000000",
  2411=>"11111101",
  2412=>"11111101",
  2413=>"00000000",
  2414=>"11111110",
  2415=>"11111110",
  2416=>"00000001",
  2417=>"00000011",
  2418=>"00000000",
  2419=>"00000001",
  2420=>"00000000",
  2421=>"00000011",
  2422=>"00000010",
  2423=>"00000001",
  2424=>"00000010",
  2425=>"00000010",
  2426=>"11111111",
  2427=>"00000010",
  2428=>"11111111",
  2429=>"00000000",
  2430=>"00000000",
  2431=>"11111110",
  2432=>"11111110",
  2433=>"00000001",
  2434=>"00000010",
  2435=>"00000011",
  2436=>"11111111",
  2437=>"00000001",
  2438=>"00000101",
  2439=>"00000001",
  2440=>"11111110",
  2441=>"00000000",
  2442=>"00000001",
  2443=>"11111101",
  2444=>"00000011",
  2445=>"00000010",
  2446=>"11111110",
  2447=>"00000011",
  2448=>"00000001",
  2449=>"00000000",
  2450=>"11111110",
  2451=>"00000010",
  2452=>"11111111",
  2453=>"00000000",
  2454=>"00000010",
  2455=>"11111110",
  2456=>"00000100",
  2457=>"11111101",
  2458=>"00000010",
  2459=>"11111101",
  2460=>"00000010",
  2461=>"11111111",
  2462=>"11111110",
  2463=>"11111100",
  2464=>"11111110",
  2465=>"11111111",
  2466=>"11111100",
  2467=>"00000010",
  2468=>"11111110",
  2469=>"11111101",
  2470=>"00000000",
  2471=>"11111100",
  2472=>"00000000",
  2473=>"11111110",
  2474=>"11111111",
  2475=>"00000010",
  2476=>"11111101",
  2477=>"00000000",
  2478=>"11111101",
  2479=>"00000001",
  2480=>"00000010",
  2481=>"11111111",
  2482=>"00000011",
  2483=>"11111111",
  2484=>"00000001",
  2485=>"00000000",
  2486=>"00000001",
  2487=>"11111111",
  2488=>"00000010",
  2489=>"11111111",
  2490=>"00000000",
  2491=>"00000001",
  2492=>"00000001",
  2493=>"00000010",
  2494=>"00000001",
  2495=>"11111101",
  2496=>"11111110",
  2497=>"00000100",
  2498=>"00000001",
  2499=>"11111110",
  2500=>"00001000",
  2501=>"11111101",
  2502=>"00000001",
  2503=>"11111111",
  2504=>"11111110",
  2505=>"00000001",
  2506=>"00000001",
  2507=>"00000001",
  2508=>"11111110",
  2509=>"11111110",
  2510=>"11111111",
  2511=>"11111101",
  2512=>"00000000",
  2513=>"00000010",
  2514=>"00000001",
  2515=>"00001000",
  2516=>"00000000",
  2517=>"11111101",
  2518=>"00000000",
  2519=>"11111111",
  2520=>"11111111",
  2521=>"00000011",
  2522=>"11111101",
  2523=>"11111101",
  2524=>"00000001",
  2525=>"00000010",
  2526=>"11111110",
  2527=>"00000100",
  2528=>"00000101",
  2529=>"00000011",
  2530=>"11111101",
  2531=>"00000010",
  2532=>"00000011",
  2533=>"00000001",
  2534=>"11111110",
  2535=>"11111111",
  2536=>"11111110",
  2537=>"11111110",
  2538=>"00000001",
  2539=>"11111110",
  2540=>"11111111",
  2541=>"11111100",
  2542=>"00000000",
  2543=>"00000001",
  2544=>"00000010",
  2545=>"00000000",
  2546=>"00000011",
  2547=>"00000000",
  2548=>"00000010",
  2549=>"11111110",
  2550=>"00000010",
  2551=>"11111111",
  2552=>"11111101",
  2553=>"00000001",
  2554=>"11111110",
  2555=>"00000010",
  2556=>"11111111",
  2557=>"11111110",
  2558=>"00000000",
  2559=>"00000000",
  2560=>"11111111",
  2561=>"00000010",
  2562=>"00000010",
  2563=>"11111110",
  2564=>"11111111",
  2565=>"00000010",
  2566=>"11111110",
  2567=>"00000010",
  2568=>"11111101",
  2569=>"11111101",
  2570=>"11111110",
  2571=>"00000001",
  2572=>"11111110",
  2573=>"00000001",
  2574=>"00000000",
  2575=>"11111101",
  2576=>"11111111",
  2577=>"11111110",
  2578=>"00000000",
  2579=>"11111111",
  2580=>"11111111",
  2581=>"00000000",
  2582=>"00000001",
  2583=>"00000000",
  2584=>"11111111",
  2585=>"00000010",
  2586=>"00000000",
  2587=>"11111111",
  2588=>"11111111",
  2589=>"11111110",
  2590=>"00000010",
  2591=>"00000000",
  2592=>"00000010",
  2593=>"00000000",
  2594=>"00000010",
  2595=>"11111110",
  2596=>"11111111",
  2597=>"11111101",
  2598=>"11111101",
  2599=>"00000000",
  2600=>"11111110",
  2601=>"11111110",
  2602=>"00000011",
  2603=>"00000000",
  2604=>"00000001",
  2605=>"11111111",
  2606=>"00000000",
  2607=>"11111100",
  2608=>"00000011",
  2609=>"11111111",
  2610=>"11111111",
  2611=>"00000011",
  2612=>"00000000",
  2613=>"00000100",
  2614=>"00000001",
  2615=>"11111101",
  2616=>"00000010",
  2617=>"00000010",
  2618=>"00000000",
  2619=>"11111101",
  2620=>"11111110",
  2621=>"00000000",
  2622=>"00000010",
  2623=>"11111110",
  2624=>"00000010",
  2625=>"11111111",
  2626=>"11111111",
  2627=>"11111101",
  2628=>"00000000",
  2629=>"11111111",
  2630=>"00000000",
  2631=>"00000001",
  2632=>"00000001",
  2633=>"00000000",
  2634=>"11111111",
  2635=>"11111111",
  2636=>"00000100",
  2637=>"00000001",
  2638=>"11111110",
  2639=>"00000000",
  2640=>"00000100",
  2641=>"00000001",
  2642=>"11111111",
  2643=>"00000001",
  2644=>"00000001",
  2645=>"11111101",
  2646=>"00000001",
  2647=>"00000000",
  2648=>"00000101",
  2649=>"00000010",
  2650=>"00000001",
  2651=>"11111101",
  2652=>"11111110",
  2653=>"00000000",
  2654=>"11111110",
  2655=>"00000010",
  2656=>"00000011",
  2657=>"00000000",
  2658=>"11111101",
  2659=>"00000001",
  2660=>"11111101",
  2661=>"00000000",
  2662=>"11111111",
  2663=>"00000001",
  2664=>"11111111",
  2665=>"11111111",
  2666=>"00000010",
  2667=>"11111101",
  2668=>"11111110",
  2669=>"11111110",
  2670=>"00000011",
  2671=>"11111101",
  2672=>"00000001",
  2673=>"00000010",
  2674=>"00000011",
  2675=>"11111110",
  2676=>"00000011",
  2677=>"11111111",
  2678=>"00000001",
  2679=>"00000110",
  2680=>"11111111",
  2681=>"11111111",
  2682=>"11111100",
  2683=>"00000000",
  2684=>"00000010",
  2685=>"11111111",
  2686=>"00000100",
  2687=>"00000001",
  2688=>"00000000",
  2689=>"00000001",
  2690=>"11111111",
  2691=>"00000001",
  2692=>"11111110",
  2693=>"11111111",
  2694=>"11111111",
  2695=>"11111111",
  2696=>"00000101",
  2697=>"00000000",
  2698=>"00000000",
  2699=>"00000100",
  2700=>"00000001",
  2701=>"11111110",
  2702=>"11111101",
  2703=>"11111110",
  2704=>"00000000",
  2705=>"00000010",
  2706=>"00000001",
  2707=>"11111110",
  2708=>"11111110",
  2709=>"00000000",
  2710=>"11111101",
  2711=>"00000000",
  2712=>"11111111",
  2713=>"11111101",
  2714=>"11111110",
  2715=>"11111110",
  2716=>"11111110",
  2717=>"00000010",
  2718=>"00000001",
  2719=>"00000011",
  2720=>"00000001",
  2721=>"11111101",
  2722=>"00000001",
  2723=>"00000011",
  2724=>"00000000",
  2725=>"11111110",
  2726=>"11111110",
  2727=>"11111110",
  2728=>"00000011",
  2729=>"11111101",
  2730=>"11111110",
  2731=>"11111111",
  2732=>"11111110",
  2733=>"11111111",
  2734=>"00000010",
  2735=>"11111111",
  2736=>"11111110",
  2737=>"11111110",
  2738=>"00000000",
  2739=>"11111111",
  2740=>"11111111",
  2741=>"00000000",
  2742=>"11111110",
  2743=>"00000010",
  2744=>"00000001",
  2745=>"00000000",
  2746=>"11111101",
  2747=>"00000001",
  2748=>"00000010",
  2749=>"00000010",
  2750=>"00000101",
  2751=>"11111110",
  2752=>"00000010",
  2753=>"00000000",
  2754=>"11111110",
  2755=>"11111110",
  2756=>"11111101",
  2757=>"11111111",
  2758=>"11111111",
  2759=>"00000011",
  2760=>"00000001",
  2761=>"00000001",
  2762=>"11111110",
  2763=>"00000111",
  2764=>"11111101",
  2765=>"11111100",
  2766=>"00000010",
  2767=>"00000000",
  2768=>"11111111",
  2769=>"11111111",
  2770=>"00000011",
  2771=>"00000010",
  2772=>"00000001",
  2773=>"00000100",
  2774=>"00000000",
  2775=>"00000000",
  2776=>"11111111",
  2777=>"00000000",
  2778=>"11111111",
  2779=>"11111101",
  2780=>"11111111",
  2781=>"11111111",
  2782=>"11111110",
  2783=>"11111110",
  2784=>"00000011",
  2785=>"11111110",
  2786=>"00000000",
  2787=>"11111100",
  2788=>"00000000",
  2789=>"11111110",
  2790=>"00000100",
  2791=>"00000001",
  2792=>"11111110",
  2793=>"11111111",
  2794=>"11111111",
  2795=>"11111110",
  2796=>"11111111",
  2797=>"11111111",
  2798=>"11111111",
  2799=>"00000000",
  2800=>"00000001",
  2801=>"11111101",
  2802=>"11111111",
  2803=>"00000001",
  2804=>"11111101",
  2805=>"00000001",
  2806=>"11111101",
  2807=>"00000001",
  2808=>"11111111",
  2809=>"11111111",
  2810=>"00000001",
  2811=>"00000001",
  2812=>"00000010",
  2813=>"00000000",
  2814=>"11111111",
  2815=>"00000010",
  2816=>"00000010",
  2817=>"00000100",
  2818=>"00000001",
  2819=>"11111110",
  2820=>"11111110",
  2821=>"00000000",
  2822=>"11111110",
  2823=>"00000010",
  2824=>"00000010",
  2825=>"00000001",
  2826=>"11111111",
  2827=>"11111101",
  2828=>"11111110",
  2829=>"00000000",
  2830=>"00000010",
  2831=>"00000010",
  2832=>"00000010",
  2833=>"00000010",
  2834=>"00000001",
  2835=>"00000000",
  2836=>"00000010",
  2837=>"00000001",
  2838=>"11111110",
  2839=>"11111101",
  2840=>"11111100",
  2841=>"00000010",
  2842=>"11111100",
  2843=>"00000011",
  2844=>"00000001",
  2845=>"00000000",
  2846=>"11111111",
  2847=>"11111110",
  2848=>"11111111",
  2849=>"11111110",
  2850=>"11111111",
  2851=>"00000000",
  2852=>"00000001",
  2853=>"00000000",
  2854=>"00000010",
  2855=>"00000101",
  2856=>"00000000",
  2857=>"11111100",
  2858=>"00000000",
  2859=>"00000010",
  2860=>"00000010",
  2861=>"11111111",
  2862=>"00000010",
  2863=>"00000000",
  2864=>"11111110",
  2865=>"11111111",
  2866=>"11111110",
  2867=>"00000000",
  2868=>"00000011",
  2869=>"00000000",
  2870=>"11111111",
  2871=>"00000011",
  2872=>"11111110",
  2873=>"11111111",
  2874=>"00000010",
  2875=>"00000011",
  2876=>"00000001",
  2877=>"11111101",
  2878=>"11111101",
  2879=>"00000011",
  2880=>"11111110",
  2881=>"00000001",
  2882=>"11111111",
  2883=>"11111101",
  2884=>"00000000",
  2885=>"11111101",
  2886=>"00000010",
  2887=>"00000011",
  2888=>"11111110",
  2889=>"11111111",
  2890=>"00000000",
  2891=>"00000010",
  2892=>"00000010",
  2893=>"11111110",
  2894=>"11111111",
  2895=>"11111101",
  2896=>"00000000",
  2897=>"00000000",
  2898=>"11111110",
  2899=>"00000100",
  2900=>"00000011",
  2901=>"11111110",
  2902=>"00000000",
  2903=>"11111110",
  2904=>"11111111",
  2905=>"11111111",
  2906=>"11111101",
  2907=>"11111100",
  2908=>"11111111",
  2909=>"11111101",
  2910=>"00000001",
  2911=>"00000011",
  2912=>"00000000",
  2913=>"11111101",
  2914=>"00000011",
  2915=>"00000110",
  2916=>"11111101",
  2917=>"00000001",
  2918=>"11111111",
  2919=>"11111110",
  2920=>"00000001",
  2921=>"00000010",
  2922=>"11111110",
  2923=>"00000000",
  2924=>"11111110",
  2925=>"00000000",
  2926=>"00000000",
  2927=>"00000101",
  2928=>"00000010",
  2929=>"00000001",
  2930=>"11111111",
  2931=>"00000011",
  2932=>"11111101",
  2933=>"00000001",
  2934=>"11111101",
  2935=>"00000001",
  2936=>"00000001",
  2937=>"11111101",
  2938=>"00000010",
  2939=>"11111110",
  2940=>"11111101",
  2941=>"11111111",
  2942=>"00000010",
  2943=>"00000011",
  2944=>"00000000",
  2945=>"00000101",
  2946=>"11111111",
  2947=>"00000100",
  2948=>"11111110",
  2949=>"00000100",
  2950=>"00000010",
  2951=>"00000100",
  2952=>"00000011",
  2953=>"11111100",
  2954=>"00000001",
  2955=>"11111101",
  2956=>"11111110",
  2957=>"11111111",
  2958=>"00000001",
  2959=>"11111110",
  2960=>"11111110",
  2961=>"11111110",
  2962=>"11111100",
  2963=>"11111101",
  2964=>"00000001",
  2965=>"11111110",
  2966=>"00000000",
  2967=>"00000010",
  2968=>"11111110",
  2969=>"11111110",
  2970=>"11111110",
  2971=>"11111111",
  2972=>"11111111",
  2973=>"00000100",
  2974=>"11111101",
  2975=>"00000101",
  2976=>"00000010",
  2977=>"00000000",
  2978=>"11111111",
  2979=>"00000001",
  2980=>"00000000",
  2981=>"11111111",
  2982=>"00000010",
  2983=>"11111111",
  2984=>"00000000",
  2985=>"11111110",
  2986=>"11111111",
  2987=>"00000001",
  2988=>"00000001",
  2989=>"11111110",
  2990=>"11111101",
  2991=>"00000001",
  2992=>"11111101",
  2993=>"00000000",
  2994=>"00000001",
  2995=>"00000010",
  2996=>"11111111",
  2997=>"11111110",
  2998=>"00000001",
  2999=>"11111111",
  3000=>"00000000",
  3001=>"00000001",
  3002=>"00000100",
  3003=>"11111110",
  3004=>"00000000",
  3005=>"00000011",
  3006=>"00000100",
  3007=>"11111110",
  3008=>"11111111",
  3009=>"00000000",
  3010=>"00000010",
  3011=>"00000011",
  3012=>"00000010",
  3013=>"00000010",
  3014=>"11111110",
  3015=>"00000000",
  3016=>"00000100",
  3017=>"00000000",
  3018=>"11111111",
  3019=>"00000000",
  3020=>"00000001",
  3021=>"00000000",
  3022=>"11111110",
  3023=>"00000001",
  3024=>"00000000",
  3025=>"00000010",
  3026=>"00000000",
  3027=>"00000010",
  3028=>"11111111",
  3029=>"00000000",
  3030=>"11111110",
  3031=>"00000001",
  3032=>"11111110",
  3033=>"11111110",
  3034=>"00000011",
  3035=>"00000001",
  3036=>"11111101",
  3037=>"00000111",
  3038=>"00000100",
  3039=>"00000000",
  3040=>"00000000",
  3041=>"00000001",
  3042=>"00000000",
  3043=>"11111111",
  3044=>"00000000",
  3045=>"00000000",
  3046=>"00000001",
  3047=>"00000001",
  3048=>"11111110",
  3049=>"11111110",
  3050=>"00000100",
  3051=>"00000010",
  3052=>"00000001",
  3053=>"11111101",
  3054=>"11111110",
  3055=>"11111101",
  3056=>"11111101",
  3057=>"11111110",
  3058=>"00000010",
  3059=>"00000000",
  3060=>"00000000",
  3061=>"11111101",
  3062=>"11111110",
  3063=>"00000001",
  3064=>"11111110",
  3065=>"11111101",
  3066=>"11111101",
  3067=>"11111111",
  3068=>"00000010",
  3069=>"00000010",
  3070=>"00000010",
  3071=>"11111111",
  3072=>"00000001",
  3073=>"11111111",
  3074=>"00000001",
  3075=>"11111101",
  3076=>"11111100",
  3077=>"00000000",
  3078=>"00000000",
  3079=>"11111101",
  3080=>"00000010",
  3081=>"00000001",
  3082=>"00000001",
  3083=>"11111110",
  3084=>"00000001",
  3085=>"00000001",
  3086=>"00000000",
  3087=>"00000011",
  3088=>"11111111",
  3089=>"11111100",
  3090=>"00000010",
  3091=>"11111101",
  3092=>"11111111",
  3093=>"11111101",
  3094=>"00000000",
  3095=>"00000010",
  3096=>"11111110",
  3097=>"00000010",
  3098=>"11111101",
  3099=>"11111100",
  3100=>"00000011",
  3101=>"11111110",
  3102=>"11111111",
  3103=>"11111111",
  3104=>"11111111",
  3105=>"11111101",
  3106=>"00000010",
  3107=>"00000001",
  3108=>"11111111",
  3109=>"11111110",
  3110=>"00000010",
  3111=>"11111111",
  3112=>"00000101",
  3113=>"00000010",
  3114=>"11111111",
  3115=>"11111110",
  3116=>"00000101",
  3117=>"00000010",
  3118=>"00000011",
  3119=>"11111110",
  3120=>"11111101",
  3121=>"00000010",
  3122=>"11111111",
  3123=>"00000000",
  3124=>"00000000",
  3125=>"00000011",
  3126=>"11111111",
  3127=>"00000011",
  3128=>"00000000",
  3129=>"00000110",
  3130=>"00000010",
  3131=>"11111111",
  3132=>"00000001",
  3133=>"11111111",
  3134=>"11111101",
  3135=>"11111111",
  3136=>"11111101",
  3137=>"00000110",
  3138=>"00000110",
  3139=>"00000011",
  3140=>"11111100",
  3141=>"11111111",
  3142=>"11111111",
  3143=>"00000000",
  3144=>"11111110",
  3145=>"00000000",
  3146=>"00000001",
  3147=>"11111100",
  3148=>"00000001",
  3149=>"11111111",
  3150=>"11111111",
  3151=>"00000000",
  3152=>"11111110",
  3153=>"00000001",
  3154=>"11111111",
  3155=>"11111011",
  3156=>"00000010",
  3157=>"00000001",
  3158=>"00000100",
  3159=>"11111111",
  3160=>"00000010",
  3161=>"00000010",
  3162=>"00000010",
  3163=>"00000010",
  3164=>"00000011",
  3165=>"11111101",
  3166=>"00000010",
  3167=>"11111100",
  3168=>"00000011",
  3169=>"00000001",
  3170=>"11111101",
  3171=>"00000000",
  3172=>"00000000",
  3173=>"11111110",
  3174=>"00000000",
  3175=>"00000010",
  3176=>"00000011",
  3177=>"11111110",
  3178=>"00000100",
  3179=>"11111110",
  3180=>"00000010",
  3181=>"11111100",
  3182=>"11111111",
  3183=>"11111111",
  3184=>"00000000",
  3185=>"11111110",
  3186=>"11111110",
  3187=>"11111110",
  3188=>"00000001",
  3189=>"11111101",
  3190=>"00000010",
  3191=>"00000001",
  3192=>"00000011",
  3193=>"00000001",
  3194=>"11111101",
  3195=>"00000001",
  3196=>"00000001",
  3197=>"11111110",
  3198=>"00000100",
  3199=>"11111110",
  3200=>"00000110",
  3201=>"11111101",
  3202=>"11111110",
  3203=>"11111111",
  3204=>"11111101",
  3205=>"00000011",
  3206=>"11111110",
  3207=>"11111101",
  3208=>"11111100",
  3209=>"00000100",
  3210=>"11111110",
  3211=>"11111011",
  3212=>"00000010",
  3213=>"00000001",
  3214=>"00000000",
  3215=>"00000100",
  3216=>"00000001",
  3217=>"11111111",
  3218=>"00000011",
  3219=>"00000001",
  3220=>"00000000",
  3221=>"00000011",
  3222=>"11111101",
  3223=>"11111110",
  3224=>"11111111",
  3225=>"00000001",
  3226=>"00000110",
  3227=>"00000001",
  3228=>"11111111",
  3229=>"00000100",
  3230=>"00000000",
  3231=>"00000000",
  3232=>"00000010",
  3233=>"00000000",
  3234=>"00000010",
  3235=>"11111101",
  3236=>"11111111",
  3237=>"11111011",
  3238=>"11111101",
  3239=>"00000010",
  3240=>"11111101",
  3241=>"00000010",
  3242=>"00000010",
  3243=>"11111110",
  3244=>"11111101",
  3245=>"00000001",
  3246=>"00000001",
  3247=>"00000010",
  3248=>"11111100",
  3249=>"00000010",
  3250=>"11111111",
  3251=>"11111111",
  3252=>"11111110",
  3253=>"00000001",
  3254=>"11111111",
  3255=>"00000010",
  3256=>"00000110",
  3257=>"00000000",
  3258=>"00000010",
  3259=>"11111101",
  3260=>"00000000",
  3261=>"00000001",
  3262=>"00000000",
  3263=>"11111111",
  3264=>"00000001",
  3265=>"00000000",
  3266=>"11111110",
  3267=>"00000001",
  3268=>"00000010",
  3269=>"00000000",
  3270=>"11111101",
  3271=>"00000101",
  3272=>"11111111",
  3273=>"00000001",
  3274=>"00000010",
  3275=>"00000011",
  3276=>"00000001",
  3277=>"00000000",
  3278=>"11111111",
  3279=>"00000000",
  3280=>"00000001",
  3281=>"00000010",
  3282=>"00000010",
  3283=>"00000100",
  3284=>"11111111",
  3285=>"00000001",
  3286=>"00000000",
  3287=>"11111110",
  3288=>"11111100",
  3289=>"00000011",
  3290=>"11111111",
  3291=>"11111111",
  3292=>"00000001",
  3293=>"11111101",
  3294=>"00000001",
  3295=>"11111100",
  3296=>"00000000",
  3297=>"00000001",
  3298=>"11111100",
  3299=>"00000001",
  3300=>"00000011",
  3301=>"11111110",
  3302=>"00000000",
  3303=>"11111101",
  3304=>"11111101",
  3305=>"00000001",
  3306=>"11111111",
  3307=>"00000000",
  3308=>"11111101",
  3309=>"11111111",
  3310=>"11111110",
  3311=>"00000000",
  3312=>"00000001",
  3313=>"11111010",
  3314=>"11111111",
  3315=>"00000000",
  3316=>"00000010",
  3317=>"00000111",
  3318=>"00000100",
  3319=>"00000011",
  3320=>"00000010",
  3321=>"11111110",
  3322=>"00000110",
  3323=>"00000010",
  3324=>"11111110",
  3325=>"00000011",
  3326=>"00001000",
  3327=>"00000010",
  3328=>"00000011",
  3329=>"00000100",
  3330=>"00000010",
  3331=>"00000000",
  3332=>"11111110",
  3333=>"00000000",
  3334=>"00000010",
  3335=>"11111111",
  3336=>"11111110",
  3337=>"11111101",
  3338=>"00000010",
  3339=>"11111101",
  3340=>"11111110",
  3341=>"11111100",
  3342=>"00000001",
  3343=>"11111111",
  3344=>"11111101",
  3345=>"11111110",
  3346=>"00000000",
  3347=>"00000010",
  3348=>"11111101",
  3349=>"11111111",
  3350=>"11111110",
  3351=>"11111101",
  3352=>"00000001",
  3353=>"11111110",
  3354=>"00000001",
  3355=>"11111110",
  3356=>"00000000",
  3357=>"00000011",
  3358=>"11111100",
  3359=>"00000001",
  3360=>"00000010",
  3361=>"11111111",
  3362=>"00000001",
  3363=>"11111100",
  3364=>"00000001",
  3365=>"00000001",
  3366=>"11111110",
  3367=>"11111110",
  3368=>"00000001",
  3369=>"11111110",
  3370=>"00000000",
  3371=>"00000100",
  3372=>"00000000",
  3373=>"11111110",
  3374=>"11111110",
  3375=>"00000000",
  3376=>"00000000",
  3377=>"00000101",
  3378=>"11111110",
  3379=>"00000011",
  3380=>"11111111",
  3381=>"00000001",
  3382=>"00000000",
  3383=>"11111110",
  3384=>"11111111",
  3385=>"00000000",
  3386=>"11111111",
  3387=>"00000000",
  3388=>"00000001",
  3389=>"11111111",
  3390=>"11111110",
  3391=>"11111110",
  3392=>"00000010",
  3393=>"00000100",
  3394=>"11111110",
  3395=>"11111110",
  3396=>"11111111",
  3397=>"11111110",
  3398=>"00000010",
  3399=>"11111110",
  3400=>"00000011",
  3401=>"11111101",
  3402=>"11111101",
  3403=>"11111111",
  3404=>"11111110",
  3405=>"00000000",
  3406=>"00000001",
  3407=>"00000101",
  3408=>"11111111",
  3409=>"00000010",
  3410=>"11111111",
  3411=>"00000101",
  3412=>"11111111",
  3413=>"11111101",
  3414=>"11111100",
  3415=>"00000111",
  3416=>"11111111",
  3417=>"11111111",
  3418=>"11111110",
  3419=>"00000101",
  3420=>"00000001",
  3421=>"11111111",
  3422=>"00000100",
  3423=>"00000001",
  3424=>"11111111",
  3425=>"00000101",
  3426=>"00000010",
  3427=>"00000011",
  3428=>"00000000",
  3429=>"11111111",
  3430=>"00000011",
  3431=>"11111111",
  3432=>"11111111",
  3433=>"00000001",
  3434=>"00000000",
  3435=>"00000100",
  3436=>"00000001",
  3437=>"11111110",
  3438=>"00000010",
  3439=>"00000010",
  3440=>"11111110",
  3441=>"00000010",
  3442=>"00000000",
  3443=>"11111111",
  3444=>"00000100",
  3445=>"00000000",
  3446=>"00000010",
  3447=>"00000000",
  3448=>"11111110",
  3449=>"00000000",
  3450=>"11111100",
  3451=>"11111100",
  3452=>"00000101",
  3453=>"11111111",
  3454=>"00000001",
  3455=>"11111110",
  3456=>"11111011",
  3457=>"00000000",
  3458=>"00000100",
  3459=>"11111111",
  3460=>"00000010",
  3461=>"00000011",
  3462=>"00000000",
  3463=>"11111111",
  3464=>"00000001",
  3465=>"11111101",
  3466=>"11111101",
  3467=>"11111111",
  3468=>"11111111",
  3469=>"00000000",
  3470=>"11111101",
  3471=>"00000000",
  3472=>"00000001",
  3473=>"00000001",
  3474=>"11111100",
  3475=>"11111111",
  3476=>"00000110",
  3477=>"11111111",
  3478=>"00000001",
  3479=>"00000011",
  3480=>"00000101",
  3481=>"11111101",
  3482=>"00000100",
  3483=>"00000010",
  3484=>"11111101",
  3485=>"00000001",
  3486=>"11111111",
  3487=>"11111100",
  3488=>"11111100",
  3489=>"11111110",
  3490=>"00000000",
  3491=>"11111101",
  3492=>"11111101",
  3493=>"11111111",
  3494=>"00000011",
  3495=>"00000010",
  3496=>"11111110",
  3497=>"00000100",
  3498=>"11111110",
  3499=>"00000000",
  3500=>"00000001",
  3501=>"11111110",
  3502=>"11111010",
  3503=>"11111110",
  3504=>"11111111",
  3505=>"11111101",
  3506=>"00000001",
  3507=>"00000100",
  3508=>"11111111",
  3509=>"11111110",
  3510=>"00000101",
  3511=>"11111110",
  3512=>"11111101",
  3513=>"00000000",
  3514=>"11111111",
  3515=>"11111111",
  3516=>"11111111",
  3517=>"00000001",
  3518=>"00000011",
  3519=>"00000000",
  3520=>"00000010",
  3521=>"11111110",
  3522=>"00000101",
  3523=>"00000010",
  3524=>"11111111",
  3525=>"00000011",
  3526=>"00000001",
  3527=>"00000010",
  3528=>"11111111",
  3529=>"00000000",
  3530=>"11111111",
  3531=>"11111101",
  3532=>"11111100",
  3533=>"11111111",
  3534=>"11111101",
  3535=>"11111101",
  3536=>"00000000",
  3537=>"00000010",
  3538=>"00000011",
  3539=>"11111100",
  3540=>"11111111",
  3541=>"00000001",
  3542=>"11111111",
  3543=>"00000000",
  3544=>"11111111",
  3545=>"00000001",
  3546=>"11111110",
  3547=>"00000011",
  3548=>"11111111",
  3549=>"00000001",
  3550=>"00000010",
  3551=>"11111101",
  3552=>"11111100",
  3553=>"00000001",
  3554=>"00000000",
  3555=>"00000001",
  3556=>"11111110",
  3557=>"11111110",
  3558=>"11111111",
  3559=>"00000001",
  3560=>"00000011",
  3561=>"00000010",
  3562=>"00000011",
  3563=>"00000010",
  3564=>"00000000",
  3565=>"11111100",
  3566=>"11111101",
  3567=>"00000100",
  3568=>"11111101",
  3569=>"11111100",
  3570=>"00000011",
  3571=>"11111111",
  3572=>"00000010",
  3573=>"00000000",
  3574=>"00000101",
  3575=>"11111101",
  3576=>"11111101",
  3577=>"11111011",
  3578=>"11111101",
  3579=>"00000000",
  3580=>"00000011",
  3581=>"00000000",
  3582=>"00000010",
  3583=>"11111110",
  3584=>"11111111",
  3585=>"11111110",
  3586=>"00000100",
  3587=>"00000000",
  3588=>"11111101",
  3589=>"11111101",
  3590=>"11111101",
  3591=>"11111011",
  3592=>"00000011",
  3593=>"11111101",
  3594=>"11111101",
  3595=>"11111110",
  3596=>"00000000",
  3597=>"11111100",
  3598=>"00000010",
  3599=>"00000010",
  3600=>"11111101",
  3601=>"00000000",
  3602=>"00000010",
  3603=>"00000100",
  3604=>"11111101",
  3605=>"00000000",
  3606=>"00000010",
  3607=>"11111101",
  3608=>"00000001",
  3609=>"11111110",
  3610=>"00000010",
  3611=>"00000001",
  3612=>"00000010",
  3613=>"00000000",
  3614=>"00000000",
  3615=>"11111110",
  3616=>"00000011",
  3617=>"11111111",
  3618=>"00000010",
  3619=>"11111101",
  3620=>"11111111",
  3621=>"11111110",
  3622=>"11111111",
  3623=>"11111101",
  3624=>"00000000",
  3625=>"11111101",
  3626=>"11111110",
  3627=>"00000001",
  3628=>"11111111",
  3629=>"11111110",
  3630=>"11111110",
  3631=>"11111110",
  3632=>"00000010",
  3633=>"11111110",
  3634=>"11111110",
  3635=>"11111110",
  3636=>"00000000",
  3637=>"11111100",
  3638=>"11111111",
  3639=>"11111110",
  3640=>"11111110",
  3641=>"11111110",
  3642=>"00000001",
  3643=>"11111100",
  3644=>"00000010",
  3645=>"00000010",
  3646=>"11111110",
  3647=>"00000001",
  3648=>"00000101",
  3649=>"11111110",
  3650=>"11111110",
  3651=>"11111111",
  3652=>"00000010",
  3653=>"11111111",
  3654=>"00000000",
  3655=>"00000011",
  3656=>"11111111",
  3657=>"00000010",
  3658=>"00000010",
  3659=>"11111111",
  3660=>"11111101",
  3661=>"11111110",
  3662=>"00000010",
  3663=>"11111101",
  3664=>"11111110",
  3665=>"00000101",
  3666=>"11111101",
  3667=>"00000010",
  3668=>"11111110",
  3669=>"11111110",
  3670=>"11111101",
  3671=>"11111110",
  3672=>"00000000",
  3673=>"11111101",
  3674=>"11111110",
  3675=>"00000000",
  3676=>"00000100",
  3677=>"00000000",
  3678=>"00000010",
  3679=>"00000100",
  3680=>"00000000",
  3681=>"00000010",
  3682=>"00000100",
  3683=>"11111101",
  3684=>"00000001",
  3685=>"00000010",
  3686=>"11111101",
  3687=>"11111110",
  3688=>"11111101",
  3689=>"11111100",
  3690=>"00000001",
  3691=>"11111110",
  3692=>"11111110",
  3693=>"00000000",
  3694=>"11111101",
  3695=>"00000000",
  3696=>"00000001",
  3697=>"00000001",
  3698=>"11111110",
  3699=>"00000000",
  3700=>"00000001",
  3701=>"00000000",
  3702=>"00000010",
  3703=>"11111111",
  3704=>"00000001",
  3705=>"11111101",
  3706=>"00000100",
  3707=>"11111110",
  3708=>"00000011",
  3709=>"11111110",
  3710=>"00000010",
  3711=>"00000001",
  3712=>"00000011",
  3713=>"00000001",
  3714=>"00000101",
  3715=>"00000000",
  3716=>"11111011",
  3717=>"00000111",
  3718=>"00000001",
  3719=>"11111110",
  3720=>"00000010",
  3721=>"00000001",
  3722=>"00000000",
  3723=>"11111101",
  3724=>"11111101",
  3725=>"00000010",
  3726=>"00000100",
  3727=>"00000100",
  3728=>"11111110",
  3729=>"00000111",
  3730=>"00000000",
  3731=>"00000010",
  3732=>"00000000",
  3733=>"11111110",
  3734=>"00000000",
  3735=>"00000000",
  3736=>"11111111",
  3737=>"00000011",
  3738=>"11111101",
  3739=>"11111110",
  3740=>"11111101",
  3741=>"11111101",
  3742=>"00000100",
  3743=>"11111100",
  3744=>"00000010",
  3745=>"00000010",
  3746=>"11111111",
  3747=>"11111100",
  3748=>"00000001",
  3749=>"11111111",
  3750=>"11111101",
  3751=>"11111111",
  3752=>"00000011",
  3753=>"00000010",
  3754=>"00000010",
  3755=>"00000101",
  3756=>"11111111",
  3757=>"11111110",
  3758=>"11111111",
  3759=>"00000010",
  3760=>"11111101",
  3761=>"00000011",
  3762=>"11111111",
  3763=>"00000000",
  3764=>"11111101",
  3765=>"00000000",
  3766=>"11111111",
  3767=>"00000000",
  3768=>"00000000",
  3769=>"00000010",
  3770=>"00000010",
  3771=>"00000000",
  3772=>"00000001",
  3773=>"00000000",
  3774=>"00000100",
  3775=>"00000001",
  3776=>"11111111",
  3777=>"00000010",
  3778=>"00000010",
  3779=>"00000010",
  3780=>"00000011",
  3781=>"11111101",
  3782=>"11111111",
  3783=>"00000011",
  3784=>"00000010",
  3785=>"11111101",
  3786=>"00000011",
  3787=>"11111111",
  3788=>"11111100",
  3789=>"00000001",
  3790=>"11111110",
  3791=>"11111110",
  3792=>"11111111",
  3793=>"00000000",
  3794=>"00000001",
  3795=>"11111111",
  3796=>"11111110",
  3797=>"11111110",
  3798=>"11111101",
  3799=>"00000001",
  3800=>"00000110",
  3801=>"00000100",
  3802=>"11111111",
  3803=>"00000000",
  3804=>"00000000",
  3805=>"11111111",
  3806=>"00000000",
  3807=>"00000011",
  3808=>"00000010",
  3809=>"11111111",
  3810=>"00000010",
  3811=>"00000010",
  3812=>"11111111",
  3813=>"11111110",
  3814=>"00000010",
  3815=>"11111111",
  3816=>"11111110",
  3817=>"00000000",
  3818=>"00000001",
  3819=>"00000000",
  3820=>"11111101",
  3821=>"00000010",
  3822=>"00000001",
  3823=>"00000001",
  3824=>"00000000",
  3825=>"00000001",
  3826=>"00000011",
  3827=>"00000001",
  3828=>"00000011",
  3829=>"00000100",
  3830=>"00000011",
  3831=>"00000011",
  3832=>"00001000",
  3833=>"11111100",
  3834=>"00000001",
  3835=>"11111111",
  3836=>"00000000",
  3837=>"11111110",
  3838=>"11111111",
  3839=>"00000001",
  3840=>"11111111",
  3841=>"11111101",
  3842=>"11111110",
  3843=>"11111011",
  3844=>"11111111",
  3845=>"11111100",
  3846=>"11111111",
  3847=>"00000000",
  3848=>"11111111",
  3849=>"11111100",
  3850=>"00000100",
  3851=>"00000001",
  3852=>"11111110",
  3853=>"11111111",
  3854=>"11111101",
  3855=>"00000001",
  3856=>"11111110",
  3857=>"11111101",
  3858=>"00000000",
  3859=>"11111101",
  3860=>"11111101",
  3861=>"11111111",
  3862=>"00000011",
  3863=>"00000101",
  3864=>"00000010",
  3865=>"00000001",
  3866=>"11111111",
  3867=>"11111111",
  3868=>"00000100",
  3869=>"00000011",
  3870=>"11111110",
  3871=>"11111111",
  3872=>"00000011",
  3873=>"00000000",
  3874=>"11111111",
  3875=>"11111111",
  3876=>"00000001",
  3877=>"00000001",
  3878=>"00000000",
  3879=>"00000000",
  3880=>"00000101",
  3881=>"00000100",
  3882=>"11111100",
  3883=>"00000010",
  3884=>"00000001",
  3885=>"11111111",
  3886=>"00000000",
  3887=>"00000000",
  3888=>"11111101",
  3889=>"11111110",
  3890=>"00000001",
  3891=>"11111110",
  3892=>"11111111",
  3893=>"11111111",
  3894=>"11111110",
  3895=>"00000101",
  3896=>"00000101",
  3897=>"00000001",
  3898=>"11111101",
  3899=>"11111110",
  3900=>"11111111",
  3901=>"00000011",
  3902=>"00000100",
  3903=>"00000001",
  3904=>"11111100",
  3905=>"11111101",
  3906=>"00000100",
  3907=>"00000100",
  3908=>"11111101",
  3909=>"00000000",
  3910=>"00000000",
  3911=>"00000010",
  3912=>"11111111",
  3913=>"11111111",
  3914=>"00000101",
  3915=>"00000010",
  3916=>"00000001",
  3917=>"11111110",
  3918=>"11111101",
  3919=>"00000101",
  3920=>"11111110",
  3921=>"00000010",
  3922=>"11111110",
  3923=>"11111100",
  3924=>"11111101",
  3925=>"00000001",
  3926=>"11111101",
  3927=>"11111110",
  3928=>"11111101",
  3929=>"11111101",
  3930=>"00000010",
  3931=>"00000001",
  3932=>"11111111",
  3933=>"00000001",
  3934=>"11111101",
  3935=>"00000010",
  3936=>"00000010",
  3937=>"00000011",
  3938=>"00000010",
  3939=>"00000010",
  3940=>"11111101",
  3941=>"11111101",
  3942=>"00000010",
  3943=>"11111110",
  3944=>"11111111",
  3945=>"00000000",
  3946=>"00000010",
  3947=>"11111111",
  3948=>"00000011",
  3949=>"00000111",
  3950=>"11111101",
  3951=>"00000001",
  3952=>"00000100",
  3953=>"11111111",
  3954=>"00000000",
  3955=>"00000010",
  3956=>"00000011",
  3957=>"00000001",
  3958=>"00000001",
  3959=>"11111110",
  3960=>"00000001",
  3961=>"11111111",
  3962=>"11111111",
  3963=>"11111101",
  3964=>"11111101",
  3965=>"00000001",
  3966=>"00000010",
  3967=>"00000001",
  3968=>"00000000",
  3969=>"00000000",
  3970=>"00000100",
  3971=>"00000000",
  3972=>"00000001",
  3973=>"00000001",
  3974=>"00000011",
  3975=>"00000001",
  3976=>"11111101",
  3977=>"00000001",
  3978=>"00000000",
  3979=>"00000001",
  3980=>"00000010",
  3981=>"00000011",
  3982=>"11111111",
  3983=>"00000000",
  3984=>"11111110",
  3985=>"00000010",
  3986=>"11111111",
  3987=>"11111101",
  3988=>"11111111",
  3989=>"11111101",
  3990=>"11111111",
  3991=>"11111100",
  3992=>"00000000",
  3993=>"11111101",
  3994=>"11111101",
  3995=>"00000011",
  3996=>"00000100",
  3997=>"00000010",
  3998=>"00000011",
  3999=>"11111111",
  4000=>"00000010",
  4001=>"00000000",
  4002=>"00000101",
  4003=>"00000000",
  4004=>"11111110",
  4005=>"00000001",
  4006=>"00000001",
  4007=>"11111111",
  4008=>"00000000",
  4009=>"11111110",
  4010=>"11111110",
  4011=>"11111111",
  4012=>"00000110",
  4013=>"00000010",
  4014=>"00000011",
  4015=>"11111110",
  4016=>"00000000",
  4017=>"11111101",
  4018=>"00000000",
  4019=>"11111110",
  4020=>"11111111",
  4021=>"11111110",
  4022=>"11111111",
  4023=>"11111101",
  4024=>"00000000",
  4025=>"11111111",
  4026=>"00000010",
  4027=>"11111111",
  4028=>"11111111",
  4029=>"00000000",
  4030=>"00000010",
  4031=>"00000010",
  4032=>"11111100",
  4033=>"00000010",
  4034=>"00000000",
  4035=>"11111111",
  4036=>"00000001",
  4037=>"00000010",
  4038=>"00000001",
  4039=>"00000000",
  4040=>"11111100",
  4041=>"11111101",
  4042=>"00000010",
  4043=>"11111110",
  4044=>"00000010",
  4045=>"00000010",
  4046=>"11111111",
  4047=>"00000100",
  4048=>"11111101",
  4049=>"00000000",
  4050=>"11111110",
  4051=>"00000000",
  4052=>"11111111",
  4053=>"11111110",
  4054=>"11111111",
  4055=>"00000111",
  4056=>"00000010",
  4057=>"11111110",
  4058=>"00000000",
  4059=>"11111111",
  4060=>"00000010",
  4061=>"11111101",
  4062=>"11111110",
  4063=>"11111100",
  4064=>"00000000",
  4065=>"00000000",
  4066=>"00000010",
  4067=>"00000001",
  4068=>"00000001",
  4069=>"11111111",
  4070=>"11111101",
  4071=>"00000010",
  4072=>"11111110",
  4073=>"11111101",
  4074=>"11111100",
  4075=>"00000000",
  4076=>"00000001",
  4077=>"00000001",
  4078=>"11111110",
  4079=>"00000000",
  4080=>"11111100",
  4081=>"00000000",
  4082=>"11111110",
  4083=>"00000001",
  4084=>"11111101",
  4085=>"00000011",
  4086=>"00000000",
  4087=>"11111110",
  4088=>"11111101",
  4089=>"11111101",
  4090=>"00000010",
  4091=>"11111100",
  4092=>"11111100",
  4093=>"00000001",
  4094=>"11111110",
  4095=>"00000000",
  4096=>"00000001",
  4097=>"00000011",
  4098=>"00000000",
  4099=>"11111101",
  4100=>"11111110",
  4101=>"00000000",
  4102=>"00000011",
  4103=>"00000001",
  4104=>"00000000",
  4105=>"11111100",
  4106=>"11111111",
  4107=>"00000000",
  4108=>"11111111",
  4109=>"11111111",
  4110=>"11111111",
  4111=>"00000011",
  4112=>"00000010",
  4113=>"00000100",
  4114=>"11111111",
  4115=>"00000010",
  4116=>"11111110",
  4117=>"11111101",
  4118=>"00000011",
  4119=>"11111111",
  4120=>"11111101",
  4121=>"11111110",
  4122=>"00000000",
  4123=>"00000001",
  4124=>"11111101",
  4125=>"00000001",
  4126=>"11111110",
  4127=>"11111111",
  4128=>"00000011",
  4129=>"00000000",
  4130=>"11111111",
  4131=>"00000011",
  4132=>"11111110",
  4133=>"00000000",
  4134=>"11111111",
  4135=>"00000010",
  4136=>"00000011",
  4137=>"00000110",
  4138=>"11111101",
  4139=>"11111101",
  4140=>"11111110",
  4141=>"00000000",
  4142=>"00000010",
  4143=>"11111111",
  4144=>"11111110",
  4145=>"11111111",
  4146=>"11111111",
  4147=>"11111111",
  4148=>"11111111",
  4149=>"11111110",
  4150=>"00000001",
  4151=>"00000001",
  4152=>"00000001",
  4153=>"11111110",
  4154=>"11111101",
  4155=>"00000000",
  4156=>"11111101",
  4157=>"11111111",
  4158=>"11111110",
  4159=>"00000010",
  4160=>"00000110",
  4161=>"00000001",
  4162=>"00000010",
  4163=>"11111101",
  4164=>"11111111",
  4165=>"11111111",
  4166=>"00000011",
  4167=>"00000010",
  4168=>"00000000",
  4169=>"00000100",
  4170=>"00000011",
  4171=>"00000010",
  4172=>"00000001",
  4173=>"00000010",
  4174=>"11111111",
  4175=>"00000011",
  4176=>"11111111",
  4177=>"11111110",
  4178=>"11111101",
  4179=>"00000001",
  4180=>"00000010",
  4181=>"00000100",
  4182=>"00000001",
  4183=>"00000000",
  4184=>"11111110",
  4185=>"00000101",
  4186=>"11111110",
  4187=>"11111110",
  4188=>"11111101",
  4189=>"11111111",
  4190=>"11111101",
  4191=>"11111101",
  4192=>"11111111",
  4193=>"00000001",
  4194=>"11111101",
  4195=>"11111111",
  4196=>"11111110",
  4197=>"00000100",
  4198=>"11111111",
  4199=>"11111111",
  4200=>"00000011",
  4201=>"11111111",
  4202=>"00000001",
  4203=>"00000001",
  4204=>"11111110",
  4205=>"00000010",
  4206=>"11111110",
  4207=>"00000010",
  4208=>"11111111",
  4209=>"11111110",
  4210=>"00000001",
  4211=>"11111110",
  4212=>"11111111",
  4213=>"11111110",
  4214=>"00000011",
  4215=>"00000000",
  4216=>"11111100",
  4217=>"11111100",
  4218=>"00000000",
  4219=>"11111111",
  4220=>"00000000",
  4221=>"00000010",
  4222=>"00000001",
  4223=>"00000101",
  4224=>"00000010",
  4225=>"00000010",
  4226=>"11111111",
  4227=>"00000010",
  4228=>"00000010",
  4229=>"00000011",
  4230=>"00000000",
  4231=>"00000001",
  4232=>"11111111",
  4233=>"11111110",
  4234=>"11111101",
  4235=>"00000000",
  4236=>"00000010",
  4237=>"00000000",
  4238=>"00000001",
  4239=>"11111110",
  4240=>"00000001",
  4241=>"11111101",
  4242=>"00000000",
  4243=>"00000010",
  4244=>"00000010",
  4245=>"11111111",
  4246=>"11111110",
  4247=>"11111111",
  4248=>"11111101",
  4249=>"11111100",
  4250=>"11111101",
  4251=>"00000101",
  4252=>"00000010",
  4253=>"11111111",
  4254=>"00000010",
  4255=>"11111111",
  4256=>"00000000",
  4257=>"11111111",
  4258=>"11111100",
  4259=>"11111110",
  4260=>"00000000",
  4261=>"00000001",
  4262=>"11111101",
  4263=>"00000010",
  4264=>"00000001",
  4265=>"00000000",
  4266=>"00000011",
  4267=>"00000010",
  4268=>"00000011",
  4269=>"11111110",
  4270=>"11111101",
  4271=>"00000010",
  4272=>"11111111",
  4273=>"00000100",
  4274=>"00000001",
  4275=>"00000010",
  4276=>"11111110",
  4277=>"11111100",
  4278=>"11111111",
  4279=>"00000001",
  4280=>"11111101",
  4281=>"00000010",
  4282=>"11111111",
  4283=>"00000100",
  4284=>"11111101",
  4285=>"00000000",
  4286=>"11111110",
  4287=>"00000010",
  4288=>"00000110",
  4289=>"00000000",
  4290=>"11111110",
  4291=>"11111110",
  4292=>"11111110",
  4293=>"11111101",
  4294=>"11111110",
  4295=>"11111111",
  4296=>"00000010",
  4297=>"00000110",
  4298=>"11111101",
  4299=>"00000001",
  4300=>"11111100",
  4301=>"11111110",
  4302=>"11111110",
  4303=>"11111111",
  4304=>"00000011",
  4305=>"00000011",
  4306=>"11111111",
  4307=>"11111101",
  4308=>"00000001",
  4309=>"00000110",
  4310=>"00000010",
  4311=>"00000010",
  4312=>"00000000",
  4313=>"11111100",
  4314=>"00000010",
  4315=>"00000010",
  4316=>"11111111",
  4317=>"11111101",
  4318=>"00000001",
  4319=>"11111111",
  4320=>"00000000",
  4321=>"00000001",
  4322=>"00000000",
  4323=>"00000010",
  4324=>"00000010",
  4325=>"00000010",
  4326=>"11111110",
  4327=>"11111111",
  4328=>"00000001",
  4329=>"11111100",
  4330=>"00000001",
  4331=>"00000001",
  4332=>"11111111",
  4333=>"11111101",
  4334=>"11111111",
  4335=>"11111111",
  4336=>"00000010",
  4337=>"00000101",
  4338=>"11111111",
  4339=>"00000001",
  4340=>"00000000",
  4341=>"00000100",
  4342=>"00000010",
  4343=>"00000000",
  4344=>"00000100",
  4345=>"00000000",
  4346=>"11111010",
  4347=>"11111111",
  4348=>"00000001",
  4349=>"00000000",
  4350=>"00000010",
  4351=>"11111110",
  4352=>"11111111",
  4353=>"11111110",
  4354=>"00000000",
  4355=>"11111101",
  4356=>"11111111",
  4357=>"11111110",
  4358=>"11111111",
  4359=>"11111100",
  4360=>"11111111",
  4361=>"11111111",
  4362=>"00000001",
  4363=>"00000001",
  4364=>"00000001",
  4365=>"11111110",
  4366=>"11111101",
  4367=>"00000001",
  4368=>"00000010",
  4369=>"11111110",
  4370=>"11111110",
  4371=>"00000010",
  4372=>"11111110",
  4373=>"11111101",
  4374=>"00000001",
  4375=>"11111101",
  4376=>"11111111",
  4377=>"00000010",
  4378=>"00000000",
  4379=>"11111110",
  4380=>"11111111",
  4381=>"11111110",
  4382=>"11111111",
  4383=>"00000010",
  4384=>"00000001",
  4385=>"00000000",
  4386=>"00000010",
  4387=>"00000100",
  4388=>"11111011",
  4389=>"11111110",
  4390=>"00000011",
  4391=>"11111110",
  4392=>"00000001",
  4393=>"00000011",
  4394=>"11111110",
  4395=>"11111111",
  4396=>"00000010",
  4397=>"11111110",
  4398=>"00000001",
  4399=>"00000001",
  4400=>"11111111",
  4401=>"11111110",
  4402=>"11111101",
  4403=>"00000101",
  4404=>"11111101",
  4405=>"00000001",
  4406=>"00000010",
  4407=>"00000001",
  4408=>"00000000",
  4409=>"11111111",
  4410=>"00000010",
  4411=>"00000100",
  4412=>"00000001",
  4413=>"11111111",
  4414=>"00000000",
  4415=>"11111111",
  4416=>"11111110",
  4417=>"00000100",
  4418=>"11111110",
  4419=>"11111110",
  4420=>"00000010",
  4421=>"11111110",
  4422=>"00000110",
  4423=>"00000010",
  4424=>"00000011",
  4425=>"00000101",
  4426=>"11111101",
  4427=>"00000010",
  4428=>"00000011",
  4429=>"00000011",
  4430=>"00000000",
  4431=>"11111111",
  4432=>"11111101",
  4433=>"00000100",
  4434=>"11111110",
  4435=>"11111100",
  4436=>"11111111",
  4437=>"11111110",
  4438=>"00000011",
  4439=>"00000101",
  4440=>"11111111",
  4441=>"00000010",
  4442=>"00000100",
  4443=>"11111100",
  4444=>"11111111",
  4445=>"00000001",
  4446=>"11111110",
  4447=>"00000000",
  4448=>"11111101",
  4449=>"00000010",
  4450=>"00000001",
  4451=>"11111101",
  4452=>"00000001",
  4453=>"11111111",
  4454=>"00000101",
  4455=>"00000001",
  4456=>"11111110",
  4457=>"00000011",
  4458=>"11111111",
  4459=>"11111100",
  4460=>"00000011",
  4461=>"00000011",
  4462=>"00000000",
  4463=>"00000011",
  4464=>"00000001",
  4465=>"00000001",
  4466=>"11111101",
  4467=>"11111100",
  4468=>"00000011",
  4469=>"11111100",
  4470=>"11111101",
  4471=>"11111111",
  4472=>"11111100",
  4473=>"00000100",
  4474=>"00000000",
  4475=>"11111110",
  4476=>"00000010",
  4477=>"00000000",
  4478=>"11111101",
  4479=>"00000001",
  4480=>"11111111",
  4481=>"00000011",
  4482=>"00000011",
  4483=>"00000001",
  4484=>"11111110",
  4485=>"00000010",
  4486=>"00000000",
  4487=>"11111111",
  4488=>"00000000",
  4489=>"11111100",
  4490=>"11111111",
  4491=>"00000001",
  4492=>"00000011",
  4493=>"11111110",
  4494=>"00000000",
  4495=>"00000000",
  4496=>"11111101",
  4497=>"00000010",
  4498=>"00000011",
  4499=>"00000100",
  4500=>"00000010",
  4501=>"00000000",
  4502=>"11111110",
  4503=>"00000010",
  4504=>"11111111",
  4505=>"00000100",
  4506=>"11111110",
  4507=>"11111110",
  4508=>"00000000",
  4509=>"11111101",
  4510=>"11111101",
  4511=>"00000011",
  4512=>"11111110",
  4513=>"00000010",
  4514=>"00000000",
  4515=>"11111110",
  4516=>"00000001",
  4517=>"11111110",
  4518=>"00000011",
  4519=>"11111111",
  4520=>"00000000",
  4521=>"00000001",
  4522=>"11111100",
  4523=>"11111100",
  4524=>"00000001",
  4525=>"00000001",
  4526=>"00000011",
  4527=>"00000010",
  4528=>"11111110",
  4529=>"11111110",
  4530=>"00000001",
  4531=>"11111110",
  4532=>"00000010",
  4533=>"00000111",
  4534=>"11111101",
  4535=>"00000001",
  4536=>"00000000",
  4537=>"11111110",
  4538=>"00000010",
  4539=>"11111101",
  4540=>"00000001",
  4541=>"00000101",
  4542=>"00000010",
  4543=>"00000010",
  4544=>"00000010",
  4545=>"11111110",
  4546=>"11111111",
  4547=>"00000000",
  4548=>"11111111",
  4549=>"00000011",
  4550=>"00000111",
  4551=>"00000011",
  4552=>"11111110",
  4553=>"11111110",
  4554=>"00000010",
  4555=>"11111110",
  4556=>"11111111",
  4557=>"00000000",
  4558=>"00000010",
  4559=>"00000011",
  4560=>"00000011",
  4561=>"00000000",
  4562=>"11111101",
  4563=>"00000100",
  4564=>"11111111",
  4565=>"11111101",
  4566=>"11111111",
  4567=>"11111110",
  4568=>"00000000",
  4569=>"11111111",
  4570=>"11111110",
  4571=>"11111101",
  4572=>"11111101",
  4573=>"00000011",
  4574=>"00000011",
  4575=>"00000110",
  4576=>"11111110",
  4577=>"00000010",
  4578=>"11111111",
  4579=>"00000001",
  4580=>"00000010",
  4581=>"00000000",
  4582=>"11111111",
  4583=>"11111110",
  4584=>"11111111",
  4585=>"11111110",
  4586=>"00000000",
  4587=>"11111101",
  4588=>"00000100",
  4589=>"11111110",
  4590=>"11111101",
  4591=>"00000110",
  4592=>"00000011",
  4593=>"11111100",
  4594=>"00000010",
  4595=>"11111111",
  4596=>"11111110",
  4597=>"11111111",
  4598=>"00000000",
  4599=>"00000000",
  4600=>"00000000",
  4601=>"00000101",
  4602=>"00000011",
  4603=>"00000001",
  4604=>"00000010",
  4605=>"00000011",
  4606=>"00000000",
  4607=>"00000010",
  4608=>"00000001",
  4609=>"11111111",
  4610=>"00000001",
  4611=>"00000000",
  4612=>"00000001",
  4613=>"11111111",
  4614=>"11111101",
  4615=>"11111110",
  4616=>"00000000",
  4617=>"00000000",
  4618=>"11111111",
  4619=>"00000000",
  4620=>"00000011",
  4621=>"11111110",
  4622=>"11111111",
  4623=>"00000001",
  4624=>"11111110",
  4625=>"00000001",
  4626=>"11111111",
  4627=>"00000011",
  4628=>"00000010",
  4629=>"00000011",
  4630=>"11111110",
  4631=>"11111111",
  4632=>"00000010",
  4633=>"11111100",
  4634=>"11111101",
  4635=>"00000000",
  4636=>"00000010",
  4637=>"00000010",
  4638=>"00000000",
  4639=>"11111110",
  4640=>"11111100",
  4641=>"11111110",
  4642=>"11111100",
  4643=>"00000001",
  4644=>"00000000",
  4645=>"11111110",
  4646=>"00000011",
  4647=>"11111110",
  4648=>"00000000",
  4649=>"11111110",
  4650=>"00000011",
  4651=>"11111111",
  4652=>"11111111",
  4653=>"11111110",
  4654=>"11111111",
  4655=>"11111101",
  4656=>"00000000",
  4657=>"00000001",
  4658=>"00000010",
  4659=>"11111111",
  4660=>"00000010",
  4661=>"11111110",
  4662=>"11111111",
  4663=>"11111111",
  4664=>"11111101",
  4665=>"00000000",
  4666=>"11111110",
  4667=>"11111101",
  4668=>"00000000",
  4669=>"00000011",
  4670=>"00000000",
  4671=>"00000000",
  4672=>"00000011",
  4673=>"00000001",
  4674=>"11111101",
  4675=>"11111111",
  4676=>"00000001",
  4677=>"11111101",
  4678=>"11111111",
  4679=>"11111110",
  4680=>"11111111",
  4681=>"11111111",
  4682=>"11111101",
  4683=>"11111101",
  4684=>"11111111",
  4685=>"11111111",
  4686=>"11111101",
  4687=>"00000011",
  4688=>"11111110",
  4689=>"00000000",
  4690=>"11111110",
  4691=>"00000010",
  4692=>"00000010",
  4693=>"00000001",
  4694=>"11111110",
  4695=>"11111101",
  4696=>"11111110",
  4697=>"00000001",
  4698=>"11111101",
  4699=>"00000001",
  4700=>"11111101",
  4701=>"00000001",
  4702=>"11111110",
  4703=>"00000010",
  4704=>"11111111",
  4705=>"11111110",
  4706=>"11111111",
  4707=>"11111101",
  4708=>"11111111",
  4709=>"00000010",
  4710=>"00000000",
  4711=>"00000000",
  4712=>"11111100",
  4713=>"11111111",
  4714=>"00000001",
  4715=>"00000000",
  4716=>"11111101",
  4717=>"00000101",
  4718=>"11111110",
  4719=>"11111101",
  4720=>"00000000",
  4721=>"00000000",
  4722=>"11111101",
  4723=>"11111111",
  4724=>"11111110",
  4725=>"00000000",
  4726=>"00000000",
  4727=>"11111111",
  4728=>"11111101",
  4729=>"00000000",
  4730=>"11111111",
  4731=>"00000001",
  4732=>"11111101",
  4733=>"11111110",
  4734=>"11111100",
  4735=>"00000000",
  4736=>"00000001",
  4737=>"11111111",
  4738=>"00000010",
  4739=>"00000010",
  4740=>"11111110",
  4741=>"11111111",
  4742=>"00000011",
  4743=>"11111111",
  4744=>"11111101",
  4745=>"00000000",
  4746=>"00000000",
  4747=>"11111101",
  4748=>"00000000",
  4749=>"00000011",
  4750=>"11111110",
  4751=>"00000000",
  4752=>"11111111",
  4753=>"00000000",
  4754=>"00000011",
  4755=>"00000000",
  4756=>"11111110",
  4757=>"11111111",
  4758=>"00000011",
  4759=>"11111101",
  4760=>"11111101",
  4761=>"11111100",
  4762=>"11111110",
  4763=>"11111111",
  4764=>"11111101",
  4765=>"11111111",
  4766=>"00000011",
  4767=>"00000010",
  4768=>"00000010",
  4769=>"00000000",
  4770=>"00000100",
  4771=>"11111111",
  4772=>"00000010",
  4773=>"00000001",
  4774=>"00000001",
  4775=>"00000101",
  4776=>"11111110",
  4777=>"11111110",
  4778=>"11111101",
  4779=>"00000000",
  4780=>"11111111",
  4781=>"11111111",
  4782=>"00000010",
  4783=>"00000000",
  4784=>"11111100",
  4785=>"00000101",
  4786=>"11111110",
  4787=>"11111110",
  4788=>"11111110",
  4789=>"00000011",
  4790=>"11111111",
  4791=>"11111111",
  4792=>"00000010",
  4793=>"00000000",
  4794=>"00000000",
  4795=>"11111111",
  4796=>"11111101",
  4797=>"11111110",
  4798=>"11111101",
  4799=>"11111101",
  4800=>"11111101",
  4801=>"00000011",
  4802=>"11111110",
  4803=>"11111101",
  4804=>"00000000",
  4805=>"00000010",
  4806=>"00000100",
  4807=>"00000100",
  4808=>"11111101",
  4809=>"00000001",
  4810=>"11111111",
  4811=>"11111110",
  4812=>"11111111",
  4813=>"00000000",
  4814=>"00000010",
  4815=>"11111111",
  4816=>"11111110",
  4817=>"00000010",
  4818=>"00000000",
  4819=>"11111111",
  4820=>"00000001",
  4821=>"11111101",
  4822=>"00000001",
  4823=>"00000100",
  4824=>"00000011",
  4825=>"11111110",
  4826=>"11111110",
  4827=>"00000100",
  4828=>"00000010",
  4829=>"11111110",
  4830=>"00000011",
  4831=>"00000001",
  4832=>"11111111",
  4833=>"11111110",
  4834=>"00000100",
  4835=>"11111111",
  4836=>"11111101",
  4837=>"00000011",
  4838=>"00000000",
  4839=>"11111100",
  4840=>"00000100",
  4841=>"00000011",
  4842=>"11111110",
  4843=>"11111110",
  4844=>"00000000",
  4845=>"11111111",
  4846=>"00000000",
  4847=>"11111111",
  4848=>"11111110",
  4849=>"11111111",
  4850=>"11111101",
  4851=>"11111101",
  4852=>"11111110",
  4853=>"00000010",
  4854=>"00000011",
  4855=>"11111101",
  4856=>"11111101",
  4857=>"11111101",
  4858=>"00000010",
  4859=>"00000010",
  4860=>"11111111",
  4861=>"00000011",
  4862=>"00000010",
  4863=>"11111110",
  4864=>"11111100",
  4865=>"00000001",
  4866=>"11111101",
  4867=>"11111100",
  4868=>"00000000",
  4869=>"00000000",
  4870=>"11111101",
  4871=>"11111110",
  4872=>"11111111",
  4873=>"11111111",
  4874=>"11111111",
  4875=>"00000100",
  4876=>"00000001",
  4877=>"11111100",
  4878=>"00000000",
  4879=>"00000011",
  4880=>"11111110",
  4881=>"00000001",
  4882=>"11111100",
  4883=>"00000000",
  4884=>"00000001",
  4885=>"00000101",
  4886=>"00000000",
  4887=>"00000000",
  4888=>"00000100",
  4889=>"11111111",
  4890=>"11111110",
  4891=>"11111110",
  4892=>"11111110",
  4893=>"00000001",
  4894=>"00000000",
  4895=>"11111111",
  4896=>"00000001",
  4897=>"00000000",
  4898=>"11111111",
  4899=>"11111111",
  4900=>"11111101",
  4901=>"11111110",
  4902=>"00000000",
  4903=>"11111111",
  4904=>"00000010",
  4905=>"00000110",
  4906=>"00000000",
  4907=>"00000000",
  4908=>"00000010",
  4909=>"11111111",
  4910=>"11111111",
  4911=>"00000001",
  4912=>"00000101",
  4913=>"11111111",
  4914=>"00000101",
  4915=>"11111111",
  4916=>"00000000",
  4917=>"00000000",
  4918=>"11111111",
  4919=>"00000000",
  4920=>"00000100",
  4921=>"00000010",
  4922=>"00000001",
  4923=>"11111100",
  4924=>"11111110",
  4925=>"11111111",
  4926=>"11111111",
  4927=>"11111101",
  4928=>"00000100",
  4929=>"00000010",
  4930=>"00000001",
  4931=>"00000101",
  4932=>"00000010",
  4933=>"11111101",
  4934=>"11111110",
  4935=>"00000001",
  4936=>"11111010",
  4937=>"00000010",
  4938=>"11111111",
  4939=>"00000110",
  4940=>"11111110",
  4941=>"11111101",
  4942=>"11111110",
  4943=>"11111100",
  4944=>"00000001",
  4945=>"11111110",
  4946=>"00000001",
  4947=>"11111100",
  4948=>"00000001",
  4949=>"00000011",
  4950=>"00000001",
  4951=>"11111110",
  4952=>"00000011",
  4953=>"11111111",
  4954=>"00000000",
  4955=>"00000101",
  4956=>"00000000",
  4957=>"00000000",
  4958=>"00000010",
  4959=>"00000000",
  4960=>"11111111",
  4961=>"11111111",
  4962=>"11111110",
  4963=>"00000000",
  4964=>"11111111",
  4965=>"00000001",
  4966=>"11111111",
  4967=>"11111111",
  4968=>"00000001",
  4969=>"00000001",
  4970=>"00000000",
  4971=>"00000101",
  4972=>"00000010",
  4973=>"00000000",
  4974=>"00000111",
  4975=>"11111110",
  4976=>"00000101",
  4977=>"00000000",
  4978=>"11111111",
  4979=>"11111110",
  4980=>"00000001",
  4981=>"11111100",
  4982=>"00000010",
  4983=>"11111111",
  4984=>"11111110",
  4985=>"11111110",
  4986=>"11111101",
  4987=>"00000010",
  4988=>"00000011",
  4989=>"11111110",
  4990=>"11111110",
  4991=>"11111101",
  4992=>"00000000",
  4993=>"00000001",
  4994=>"00000010",
  4995=>"11111101",
  4996=>"11111110",
  4997=>"00000011",
  4998=>"00000011",
  4999=>"11111100",
  5000=>"00000000",
  5001=>"11111101",
  5002=>"00000010",
  5003=>"11111110",
  5004=>"00000010",
  5005=>"00000010",
  5006=>"00000100",
  5007=>"00000001",
  5008=>"00000000",
  5009=>"11111100",
  5010=>"11111111",
  5011=>"11111110",
  5012=>"11111101",
  5013=>"00000000",
  5014=>"11111111",
  5015=>"11111111",
  5016=>"00000011",
  5017=>"00000001",
  5018=>"11111110",
  5019=>"00000011",
  5020=>"00000011",
  5021=>"00000000",
  5022=>"11111100",
  5023=>"11111111",
  5024=>"11111101",
  5025=>"00000000",
  5026=>"00000000",
  5027=>"00000000",
  5028=>"00000000",
  5029=>"11111110",
  5030=>"00000001",
  5031=>"11111110",
  5032=>"00000001",
  5033=>"11111110",
  5034=>"00000000",
  5035=>"00000001",
  5036=>"11111101",
  5037=>"11111110",
  5038=>"11111110",
  5039=>"00000001",
  5040=>"11111111",
  5041=>"11111110",
  5042=>"00000100",
  5043=>"11111110",
  5044=>"11111111",
  5045=>"11111110",
  5046=>"00000001",
  5047=>"11111100",
  5048=>"00000011",
  5049=>"11111101",
  5050=>"00000001",
  5051=>"00000001",
  5052=>"00000001",
  5053=>"00000010",
  5054=>"11111110",
  5055=>"00000100",
  5056=>"00000001",
  5057=>"00000010",
  5058=>"11111110",
  5059=>"00000011",
  5060=>"11111110",
  5061=>"00000001",
  5062=>"11111110",
  5063=>"00000001",
  5064=>"11111101",
  5065=>"00000000",
  5066=>"11111110",
  5067=>"11111111",
  5068=>"00000010",
  5069=>"11111111",
  5070=>"11111100",
  5071=>"11111110",
  5072=>"00000001",
  5073=>"00000010",
  5074=>"00000000",
  5075=>"00000010",
  5076=>"11111110",
  5077=>"11111111",
  5078=>"00000011",
  5079=>"11111100",
  5080=>"00000001",
  5081=>"00000001",
  5082=>"00000001",
  5083=>"11111111",
  5084=>"11111111",
  5085=>"00000010",
  5086=>"11111110",
  5087=>"00000110",
  5088=>"00000001",
  5089=>"00000000",
  5090=>"00000001",
  5091=>"11111101",
  5092=>"11111110",
  5093=>"11111110",
  5094=>"00000010",
  5095=>"00000000",
  5096=>"00000010",
  5097=>"00000011",
  5098=>"00000001",
  5099=>"00000000",
  5100=>"11111111",
  5101=>"00000011",
  5102=>"11111101",
  5103=>"11111011",
  5104=>"00000001",
  5105=>"00000011",
  5106=>"11111101",
  5107=>"00000001",
  5108=>"00000000",
  5109=>"11111100",
  5110=>"00000000",
  5111=>"11111110",
  5112=>"00000010",
  5113=>"00000000",
  5114=>"00000000",
  5115=>"11111110",
  5116=>"11111111",
  5117=>"00000111",
  5118=>"11111101",
  5119=>"11111111",
  5120=>"11111111",
  5121=>"11111110",
  5122=>"11111110",
  5123=>"00000010",
  5124=>"11111101",
  5125=>"11111101",
  5126=>"11111111",
  5127=>"11111101",
  5128=>"00000011",
  5129=>"11111110",
  5130=>"00000010",
  5131=>"11111111",
  5132=>"00000001",
  5133=>"11111100",
  5134=>"00000000",
  5135=>"11111110",
  5136=>"00000011",
  5137=>"00000001",
  5138=>"00000101",
  5139=>"11111110",
  5140=>"11111111",
  5141=>"00000000",
  5142=>"11111111",
  5143=>"11111111",
  5144=>"11111101",
  5145=>"11111011",
  5146=>"11111111",
  5147=>"00000001",
  5148=>"11111101",
  5149=>"00000001",
  5150=>"00000101",
  5151=>"00000000",
  5152=>"11111111",
  5153=>"11111111",
  5154=>"11111110",
  5155=>"00000010",
  5156=>"11111110",
  5157=>"00000100",
  5158=>"00000010",
  5159=>"11111101",
  5160=>"00000001",
  5161=>"00000000",
  5162=>"00000001",
  5163=>"11111111",
  5164=>"00000000",
  5165=>"11111101",
  5166=>"00000010",
  5167=>"00000000",
  5168=>"00000001",
  5169=>"00000001",
  5170=>"00000011",
  5171=>"11111110",
  5172=>"00000000",
  5173=>"11111111",
  5174=>"00000000",
  5175=>"00000001",
  5176=>"11111111",
  5177=>"00000110",
  5178=>"11111110",
  5179=>"11111111",
  5180=>"00000000",
  5181=>"11111101",
  5182=>"11111101",
  5183=>"11111111",
  5184=>"11111110",
  5185=>"00000000",
  5186=>"11111101",
  5187=>"11111111",
  5188=>"11111111",
  5189=>"00000010",
  5190=>"00000001",
  5191=>"11111101",
  5192=>"11111111",
  5193=>"11111101",
  5194=>"00000001",
  5195=>"11111110",
  5196=>"11111101",
  5197=>"00000000",
  5198=>"00000001",
  5199=>"00000000",
  5200=>"11111111",
  5201=>"00000000",
  5202=>"00000001",
  5203=>"11111111",
  5204=>"11111110",
  5205=>"00000000",
  5206=>"00000001",
  5207=>"00000001",
  5208=>"11111110",
  5209=>"00000011",
  5210=>"11111111",
  5211=>"00000001",
  5212=>"00000101",
  5213=>"11111111",
  5214=>"00000011",
  5215=>"11111101",
  5216=>"11111101",
  5217=>"11111100",
  5218=>"11111111",
  5219=>"11111111",
  5220=>"00000010",
  5221=>"00000001",
  5222=>"00000000",
  5223=>"11111111",
  5224=>"00000010",
  5225=>"11111111",
  5226=>"00000001",
  5227=>"00000100",
  5228=>"00000101",
  5229=>"00000011",
  5230=>"11111111",
  5231=>"11111111",
  5232=>"11111110",
  5233=>"11111110",
  5234=>"11111111",
  5235=>"11111111",
  5236=>"00000000",
  5237=>"11111110",
  5238=>"11111111",
  5239=>"00000000",
  5240=>"11111100",
  5241=>"00000001",
  5242=>"11111111",
  5243=>"11111101",
  5244=>"11111101",
  5245=>"11111110",
  5246=>"11111110",
  5247=>"11111101",
  5248=>"11111110",
  5249=>"11111111",
  5250=>"00000010",
  5251=>"11111110",
  5252=>"11111101",
  5253=>"11111110",
  5254=>"00000001",
  5255=>"11111101",
  5256=>"00000010",
  5257=>"00000000",
  5258=>"11111110",
  5259=>"00000101",
  5260=>"11111100",
  5261=>"00000001",
  5262=>"11111101",
  5263=>"11111111",
  5264=>"00000100",
  5265=>"00000010",
  5266=>"00000010",
  5267=>"11111111",
  5268=>"00000100",
  5269=>"00000000",
  5270=>"11111101",
  5271=>"00000100",
  5272=>"00000111",
  5273=>"11111110",
  5274=>"00000010",
  5275=>"11111101",
  5276=>"00000001",
  5277=>"11111110",
  5278=>"11111111",
  5279=>"00000100",
  5280=>"00000000",
  5281=>"11111101",
  5282=>"11111101",
  5283=>"11111111",
  5284=>"00000000",
  5285=>"11111100",
  5286=>"00000001",
  5287=>"11111110",
  5288=>"11111111",
  5289=>"00000001",
  5290=>"00000010",
  5291=>"00000011",
  5292=>"11111111",
  5293=>"11111101",
  5294=>"11111110",
  5295=>"11111110",
  5296=>"00000011",
  5297=>"11111101",
  5298=>"11111111",
  5299=>"00000001",
  5300=>"00000010",
  5301=>"00000010",
  5302=>"00000011",
  5303=>"11111111",
  5304=>"11111101",
  5305=>"00000001",
  5306=>"00000000",
  5307=>"00000001",
  5308=>"00000001",
  5309=>"00000010",
  5310=>"00000000",
  5311=>"11111111",
  5312=>"11111101",
  5313=>"00000010",
  5314=>"11111111",
  5315=>"00000000",
  5316=>"00000010",
  5317=>"11111111",
  5318=>"00000010",
  5319=>"00000000",
  5320=>"11111110",
  5321=>"00000101",
  5322=>"00000000",
  5323=>"11111110",
  5324=>"00000101",
  5325=>"00000001",
  5326=>"00000000",
  5327=>"00000001",
  5328=>"00000101",
  5329=>"11111111",
  5330=>"11111111",
  5331=>"11111110",
  5332=>"00000010",
  5333=>"00000011",
  5334=>"00000011",
  5335=>"00000100",
  5336=>"11111111",
  5337=>"11111111",
  5338=>"00000000",
  5339=>"11111110",
  5340=>"00000000",
  5341=>"11111101",
  5342=>"00000000",
  5343=>"11111110",
  5344=>"11111101",
  5345=>"11111100",
  5346=>"00000001",
  5347=>"11111110",
  5348=>"00000001",
  5349=>"00000000",
  5350=>"00000001",
  5351=>"00000010",
  5352=>"11111111",
  5353=>"11111100",
  5354=>"11111110",
  5355=>"11111110",
  5356=>"00000001",
  5357=>"00000010",
  5358=>"00000011",
  5359=>"11111111",
  5360=>"11111101",
  5361=>"11111101",
  5362=>"00000010",
  5363=>"11111100",
  5364=>"11111110",
  5365=>"11111111",
  5366=>"00000011",
  5367=>"00000011",
  5368=>"00000100",
  5369=>"11111111",
  5370=>"11111101",
  5371=>"11111110",
  5372=>"00000001",
  5373=>"00000010",
  5374=>"00000000",
  5375=>"00000011",
  5376=>"00000001",
  5377=>"11111110",
  5378=>"00000011",
  5379=>"11111111",
  5380=>"11111101",
  5381=>"00000000",
  5382=>"11111111",
  5383=>"11111111",
  5384=>"00000001",
  5385=>"00000100",
  5386=>"00000001",
  5387=>"00000001",
  5388=>"00000000",
  5389=>"11111111",
  5390=>"00000010",
  5391=>"00000000",
  5392=>"00000001",
  5393=>"00000001",
  5394=>"00000000",
  5395=>"00000010",
  5396=>"11111101",
  5397=>"00000000",
  5398=>"00000000",
  5399=>"00000001",
  5400=>"11111100",
  5401=>"00000010",
  5402=>"00000010",
  5403=>"00000001",
  5404=>"00000000",
  5405=>"11111110",
  5406=>"00000000",
  5407=>"11111110",
  5408=>"00000001",
  5409=>"00000000",
  5410=>"00000010",
  5411=>"00000001",
  5412=>"11111110",
  5413=>"00000001",
  5414=>"11111101",
  5415=>"11111101",
  5416=>"00000011",
  5417=>"00000100",
  5418=>"11111111",
  5419=>"00000001",
  5420=>"11111111",
  5421=>"11111111",
  5422=>"11111101",
  5423=>"11111101",
  5424=>"11111101",
  5425=>"00000000",
  5426=>"11111101",
  5427=>"11111110",
  5428=>"11111110",
  5429=>"00000100",
  5430=>"11111110",
  5431=>"00000000",
  5432=>"00000001",
  5433=>"11111101",
  5434=>"11111101",
  5435=>"11111110",
  5436=>"00000000",
  5437=>"00000001",
  5438=>"00000000",
  5439=>"11111111",
  5440=>"11111111",
  5441=>"11111111",
  5442=>"11111111",
  5443=>"00000000",
  5444=>"00000001",
  5445=>"11111110",
  5446=>"00000010",
  5447=>"00000010",
  5448=>"11111101",
  5449=>"00000001",
  5450=>"11111101",
  5451=>"00000000",
  5452=>"00000010",
  5453=>"11111110",
  5454=>"00000001",
  5455=>"11111101",
  5456=>"00000010",
  5457=>"00000001",
  5458=>"11111111",
  5459=>"11111101",
  5460=>"00000001",
  5461=>"00000000",
  5462=>"11111111",
  5463=>"11111101",
  5464=>"00000001",
  5465=>"00000000",
  5466=>"00000000",
  5467=>"11111101",
  5468=>"11111111",
  5469=>"00000010",
  5470=>"00000000",
  5471=>"00000000",
  5472=>"11111110",
  5473=>"00000010",
  5474=>"11111110",
  5475=>"11111100",
  5476=>"00000010",
  5477=>"11111110",
  5478=>"00000001",
  5479=>"00000010",
  5480=>"00000000",
  5481=>"00000010",
  5482=>"00000001",
  5483=>"00000000",
  5484=>"11111110",
  5485=>"11111101",
  5486=>"11111111",
  5487=>"11111101",
  5488=>"00000001",
  5489=>"00000010",
  5490=>"11111111",
  5491=>"11111110",
  5492=>"11111111",
  5493=>"00000010",
  5494=>"11111111",
  5495=>"11111110",
  5496=>"00000000",
  5497=>"00000010",
  5498=>"11111110",
  5499=>"00000100",
  5500=>"00000000",
  5501=>"00000111",
  5502=>"11111111",
  5503=>"11111101",
  5504=>"00000001",
  5505=>"00000001",
  5506=>"11111101",
  5507=>"00000000",
  5508=>"00000000",
  5509=>"00000100",
  5510=>"11111111",
  5511=>"11111110",
  5512=>"00000010",
  5513=>"00000001",
  5514=>"00000001",
  5515=>"11111101",
  5516=>"00000010",
  5517=>"11111111",
  5518=>"11111101",
  5519=>"00000010",
  5520=>"11111111",
  5521=>"11111111",
  5522=>"11111101",
  5523=>"00000011",
  5524=>"11111101",
  5525=>"00000000",
  5526=>"11111101",
  5527=>"00000000",
  5528=>"11111110",
  5529=>"00000010",
  5530=>"11111100",
  5531=>"11111110",
  5532=>"00000000",
  5533=>"00000000",
  5534=>"11111101",
  5535=>"11111101",
  5536=>"00000100",
  5537=>"11111101",
  5538=>"11111111",
  5539=>"00000010",
  5540=>"11111110",
  5541=>"00000101",
  5542=>"00000001",
  5543=>"00000011",
  5544=>"00000101",
  5545=>"00000000",
  5546=>"00000011",
  5547=>"00000001",
  5548=>"00000011",
  5549=>"11111110",
  5550=>"00000010",
  5551=>"11111110",
  5552=>"00000001",
  5553=>"00000000",
  5554=>"11111101",
  5555=>"00000000",
  5556=>"11111101",
  5557=>"11111101",
  5558=>"11111100",
  5559=>"00000000",
  5560=>"00000000",
  5561=>"11111101",
  5562=>"00000001",
  5563=>"11111110",
  5564=>"00000001",
  5565=>"00000010",
  5566=>"11111111",
  5567=>"00000000",
  5568=>"00000001",
  5569=>"00000000",
  5570=>"11111110",
  5571=>"00000100",
  5572=>"00000000",
  5573=>"11111100",
  5574=>"00000011",
  5575=>"11111111",
  5576=>"00000001",
  5577=>"00000001",
  5578=>"11111110",
  5579=>"00000001",
  5580=>"00000011",
  5581=>"00000000",
  5582=>"00000010",
  5583=>"11111111",
  5584=>"11111111",
  5585=>"11111101",
  5586=>"00000100",
  5587=>"00000011",
  5588=>"11111101",
  5589=>"00000010",
  5590=>"11111111",
  5591=>"00000010",
  5592=>"11111110",
  5593=>"11111110",
  5594=>"00000011",
  5595=>"00000010",
  5596=>"00000010",
  5597=>"11111101",
  5598=>"11111110",
  5599=>"00000010",
  5600=>"00000001",
  5601=>"11111110",
  5602=>"00000001",
  5603=>"11111110",
  5604=>"11111111",
  5605=>"00000011",
  5606=>"00000010",
  5607=>"11111101",
  5608=>"00000000",
  5609=>"00000000",
  5610=>"00000010",
  5611=>"11111111",
  5612=>"11111111",
  5613=>"00000000",
  5614=>"00000010",
  5615=>"00000010",
  5616=>"00000001",
  5617=>"00000101",
  5618=>"11111111",
  5619=>"00000011",
  5620=>"00000001",
  5621=>"00000001",
  5622=>"00000001",
  5623=>"00000011",
  5624=>"00000001",
  5625=>"00000000",
  5626=>"11111111",
  5627=>"00000010",
  5628=>"11111111",
  5629=>"00000000",
  5630=>"11111111",
  5631=>"11111110",
  5632=>"11111101",
  5633=>"11111111",
  5634=>"00000010",
  5635=>"11111111",
  5636=>"11111101",
  5637=>"11111101",
  5638=>"00000001",
  5639=>"00000001",
  5640=>"00000001",
  5641=>"11111111",
  5642=>"11111110",
  5643=>"11111111",
  5644=>"00000101",
  5645=>"11111101",
  5646=>"00000100",
  5647=>"11111111",
  5648=>"00000011",
  5649=>"11111111",
  5650=>"11111111",
  5651=>"00000100",
  5652=>"11111110",
  5653=>"11111101",
  5654=>"11111111",
  5655=>"11111101",
  5656=>"00000010",
  5657=>"00000001",
  5658=>"00000010",
  5659=>"11111110",
  5660=>"11111111",
  5661=>"00000001",
  5662=>"11111111",
  5663=>"11111111",
  5664=>"00000001",
  5665=>"11111110",
  5666=>"00000010",
  5667=>"00000001",
  5668=>"11111110",
  5669=>"11111111",
  5670=>"00000000",
  5671=>"11111110",
  5672=>"00000001",
  5673=>"00000100",
  5674=>"11111111",
  5675=>"00000011",
  5676=>"00000001",
  5677=>"11111110",
  5678=>"11111110",
  5679=>"00000010",
  5680=>"00000001",
  5681=>"11111111",
  5682=>"11111110",
  5683=>"00000010",
  5684=>"00000000",
  5685=>"00000000",
  5686=>"00000010",
  5687=>"11111110",
  5688=>"11111111",
  5689=>"00000010",
  5690=>"11111111",
  5691=>"00000100",
  5692=>"11111111",
  5693=>"00000100",
  5694=>"11111111",
  5695=>"00000101",
  5696=>"00000011",
  5697=>"11111110",
  5698=>"00000001",
  5699=>"11111101",
  5700=>"00000000",
  5701=>"11111110",
  5702=>"11111110",
  5703=>"11111110",
  5704=>"11111110",
  5705=>"00000000",
  5706=>"11111110",
  5707=>"00001001",
  5708=>"00000001",
  5709=>"11111110",
  5710=>"00000001",
  5711=>"11111110",
  5712=>"00000010",
  5713=>"00000011",
  5714=>"11111110",
  5715=>"11111111",
  5716=>"00000000",
  5717=>"00000100",
  5718=>"00000010",
  5719=>"00000100",
  5720=>"11111111",
  5721=>"00000100",
  5722=>"00000001",
  5723=>"00000000",
  5724=>"00000001",
  5725=>"11111110",
  5726=>"00000001",
  5727=>"00000001",
  5728=>"11111110",
  5729=>"00000000",
  5730=>"00000001",
  5731=>"00000011",
  5732=>"11111101",
  5733=>"11111101",
  5734=>"11111110",
  5735=>"11111101",
  5736=>"00000000",
  5737=>"11111110",
  5738=>"11111110",
  5739=>"11111110",
  5740=>"00000010",
  5741=>"00000001",
  5742=>"00000001",
  5743=>"11111111",
  5744=>"00000000",
  5745=>"00000010",
  5746=>"00000010",
  5747=>"11111101",
  5748=>"00000001",
  5749=>"11111111",
  5750=>"00000100",
  5751=>"11111110",
  5752=>"11111111",
  5753=>"00000010",
  5754=>"11111110",
  5755=>"11111110",
  5756=>"00000001",
  5757=>"00000001",
  5758=>"00000101",
  5759=>"11111101",
  5760=>"11111111",
  5761=>"00000010",
  5762=>"11111100",
  5763=>"11111101",
  5764=>"00000011",
  5765=>"11111110",
  5766=>"11111111",
  5767=>"11111111",
  5768=>"00000000",
  5769=>"00000001",
  5770=>"00000000",
  5771=>"11111100",
  5772=>"11111111",
  5773=>"11111111",
  5774=>"11111111",
  5775=>"11111101",
  5776=>"11111111",
  5777=>"11111101",
  5778=>"11111110",
  5779=>"11111101",
  5780=>"00000010",
  5781=>"11111101",
  5782=>"11111111",
  5783=>"11111111",
  5784=>"00000101",
  5785=>"00000010",
  5786=>"11111101",
  5787=>"00000001",
  5788=>"11111100",
  5789=>"11111101",
  5790=>"00000010",
  5791=>"00000011",
  5792=>"00000001",
  5793=>"00000011",
  5794=>"00000110",
  5795=>"00000000",
  5796=>"11111110",
  5797=>"00000000",
  5798=>"00000100",
  5799=>"00000001",
  5800=>"11111100",
  5801=>"00000011",
  5802=>"00000010",
  5803=>"00000001",
  5804=>"11111111",
  5805=>"11111110",
  5806=>"00000000",
  5807=>"00000000",
  5808=>"11111111",
  5809=>"00000000",
  5810=>"00000001",
  5811=>"00000010",
  5812=>"00000010",
  5813=>"11111100",
  5814=>"00000010",
  5815=>"00000000",
  5816=>"11111111",
  5817=>"11111110",
  5818=>"11111111",
  5819=>"00000000",
  5820=>"11111111",
  5821=>"11111110",
  5822=>"11111100",
  5823=>"00000010",
  5824=>"11111110",
  5825=>"00000001",
  5826=>"11111111",
  5827=>"00000000",
  5828=>"11111110",
  5829=>"11111110",
  5830=>"11111101",
  5831=>"11111110",
  5832=>"00000001",
  5833=>"00000010",
  5834=>"00000000",
  5835=>"11111101",
  5836=>"00000101",
  5837=>"11111101",
  5838=>"00000001",
  5839=>"11111111",
  5840=>"11111101",
  5841=>"11111110",
  5842=>"11111110",
  5843=>"00000001",
  5844=>"11111110",
  5845=>"11111110",
  5846=>"00000000",
  5847=>"00000110",
  5848=>"11111111",
  5849=>"00000001",
  5850=>"11111110",
  5851=>"00000000",
  5852=>"00000000",
  5853=>"11111111",
  5854=>"00000001",
  5855=>"00000000",
  5856=>"11111101",
  5857=>"11111101",
  5858=>"00000000",
  5859=>"11111111",
  5860=>"00000000",
  5861=>"00000011",
  5862=>"00000000",
  5863=>"00000011",
  5864=>"00000010",
  5865=>"00000000",
  5866=>"00000001",
  5867=>"00000000",
  5868=>"00000010",
  5869=>"11111101",
  5870=>"00000011",
  5871=>"00000101",
  5872=>"00000000",
  5873=>"11111101",
  5874=>"00000001",
  5875=>"00000010",
  5876=>"11111110",
  5877=>"11111110",
  5878=>"00000000",
  5879=>"00000001",
  5880=>"11111100",
  5881=>"00000011",
  5882=>"11111110",
  5883=>"00000001",
  5884=>"11111110",
  5885=>"00000010",
  5886=>"00000010",
  5887=>"11111111",
  5888=>"00000011",
  5889=>"00000001",
  5890=>"00000010",
  5891=>"11111111",
  5892=>"00000000",
  5893=>"00000000",
  5894=>"00000000",
  5895=>"11111110",
  5896=>"11111100",
  5897=>"00000011",
  5898=>"00000010",
  5899=>"00000010",
  5900=>"11111110",
  5901=>"00000010",
  5902=>"00000100",
  5903=>"00000000",
  5904=>"00000001",
  5905=>"11111111",
  5906=>"11111110",
  5907=>"11111100",
  5908=>"00000010",
  5909=>"00000010",
  5910=>"00000010",
  5911=>"00000010",
  5912=>"00000001",
  5913=>"11111110",
  5914=>"00000000",
  5915=>"00000010",
  5916=>"00000001",
  5917=>"11111101",
  5918=>"11111101",
  5919=>"00000010",
  5920=>"11111100",
  5921=>"11111101",
  5922=>"11111110",
  5923=>"00000000",
  5924=>"00000000",
  5925=>"00000011",
  5926=>"00000011",
  5927=>"11111111",
  5928=>"00000001",
  5929=>"00000010",
  5930=>"00000001",
  5931=>"00000001",
  5932=>"11111111",
  5933=>"11111110",
  5934=>"00000000",
  5935=>"11111101",
  5936=>"00000010",
  5937=>"00000000",
  5938=>"11111101",
  5939=>"11111110",
  5940=>"00000000",
  5941=>"00000011",
  5942=>"11111111",
  5943=>"11111100",
  5944=>"11111100",
  5945=>"00000001",
  5946=>"11111101",
  5947=>"00000011",
  5948=>"11111110",
  5949=>"11111111",
  5950=>"00000001",
  5951=>"11111110",
  5952=>"00000000",
  5953=>"00000001",
  5954=>"00000001",
  5955=>"00000010",
  5956=>"00000000",
  5957=>"00000011",
  5958=>"11111111",
  5959=>"11111101",
  5960=>"11111110",
  5961=>"00000001",
  5962=>"00000011",
  5963=>"00000010",
  5964=>"11111110",
  5965=>"11111110",
  5966=>"11111110",
  5967=>"00000011",
  5968=>"00000011",
  5969=>"11111110",
  5970=>"00000000",
  5971=>"00000000",
  5972=>"11111111",
  5973=>"00000100",
  5974=>"00000001",
  5975=>"11111110",
  5976=>"00000010",
  5977=>"00000001",
  5978=>"11111111",
  5979=>"00000001",
  5980=>"11111110",
  5981=>"11111101",
  5982=>"00000010",
  5983=>"11111111",
  5984=>"00000010",
  5985=>"00000000",
  5986=>"11111111",
  5987=>"00000010",
  5988=>"11111111",
  5989=>"00000011",
  5990=>"00000000",
  5991=>"00000100",
  5992=>"00000011",
  5993=>"00000001",
  5994=>"00000001",
  5995=>"11111101",
  5996=>"00000001",
  5997=>"00000100",
  5998=>"11111100",
  5999=>"00000001",
  6000=>"11111101",
  6001=>"00000010",
  6002=>"11111101",
  6003=>"00000001",
  6004=>"00000000",
  6005=>"00000001",
  6006=>"00000001",
  6007=>"11111111",
  6008=>"00000000",
  6009=>"11111110",
  6010=>"00000100",
  6011=>"00000001",
  6012=>"11111101",
  6013=>"00000001",
  6014=>"11111101",
  6015=>"00000011",
  6016=>"11111111",
  6017=>"00000001",
  6018=>"00000000",
  6019=>"00000000",
  6020=>"00000010",
  6021=>"11111101",
  6022=>"11111111",
  6023=>"00000001",
  6024=>"00000000",
  6025=>"11111100",
  6026=>"00000001",
  6027=>"11111110",
  6028=>"00000010",
  6029=>"00000000",
  6030=>"11111101",
  6031=>"11111101",
  6032=>"11111111",
  6033=>"11111101",
  6034=>"11111111",
  6035=>"00000010",
  6036=>"00000001",
  6037=>"11111110",
  6038=>"11111101",
  6039=>"11111111",
  6040=>"00000001",
  6041=>"11111101",
  6042=>"11111101",
  6043=>"11111111",
  6044=>"00000010",
  6045=>"11111111",
  6046=>"00000000",
  6047=>"11111111",
  6048=>"11111101",
  6049=>"00000001",
  6050=>"11111101",
  6051=>"00000001",
  6052=>"00000001",
  6053=>"00000001",
  6054=>"11111101",
  6055=>"11111111",
  6056=>"00000001",
  6057=>"00000011",
  6058=>"00000001",
  6059=>"00000010",
  6060=>"00000000",
  6061=>"00000001",
  6062=>"00000001",
  6063=>"11111110",
  6064=>"00000001",
  6065=>"11111111",
  6066=>"11111110",
  6067=>"00000000",
  6068=>"00000000",
  6069=>"11111110",
  6070=>"11111101",
  6071=>"00000011",
  6072=>"11111111",
  6073=>"00000000",
  6074=>"11111111",
  6075=>"11111110",
  6076=>"00000000",
  6077=>"00000100",
  6078=>"00000000",
  6079=>"00000000",
  6080=>"11111110",
  6081=>"00000010",
  6082=>"11111110",
  6083=>"11111111",
  6084=>"11111111",
  6085=>"00000001",
  6086=>"00000100",
  6087=>"11111110",
  6088=>"11111111",
  6089=>"11111111",
  6090=>"11111101",
  6091=>"11111110",
  6092=>"11111110",
  6093=>"00000001",
  6094=>"11111111",
  6095=>"11111101",
  6096=>"11111110",
  6097=>"11111111",
  6098=>"00000000",
  6099=>"00000001",
  6100=>"00000000",
  6101=>"11111111",
  6102=>"00000000",
  6103=>"00000001",
  6104=>"11111111",
  6105=>"00000101",
  6106=>"11111101",
  6107=>"00000001",
  6108=>"00000001",
  6109=>"00000000",
  6110=>"11111110",
  6111=>"11111100",
  6112=>"11111111",
  6113=>"00000000",
  6114=>"11111111",
  6115=>"00000001",
  6116=>"11111110",
  6117=>"11111101",
  6118=>"11111100",
  6119=>"00000000",
  6120=>"00000000",
  6121=>"11111110",
  6122=>"00000100",
  6123=>"11111111",
  6124=>"00000100",
  6125=>"11111101",
  6126=>"00000000",
  6127=>"11111110",
  6128=>"00000100",
  6129=>"11111111",
  6130=>"00000100",
  6131=>"11111110",
  6132=>"00000001",
  6133=>"11111110",
  6134=>"00000101",
  6135=>"00000011",
  6136=>"11111111",
  6137=>"11111101",
  6138=>"00000000",
  6139=>"11111110",
  6140=>"00000010",
  6141=>"00000011",
  6142=>"11111111",
  6143=>"11111101",
  6144=>"00000010",
  6145=>"00000011",
  6146=>"00000001",
  6147=>"00000000",
  6148=>"00000111",
  6149=>"00000110",
  6150=>"11111110",
  6151=>"11111111",
  6152=>"11111111",
  6153=>"11111101",
  6154=>"00000011",
  6155=>"00000011",
  6156=>"11111110",
  6157=>"00000100",
  6158=>"11111011",
  6159=>"11111110",
  6160=>"11111110",
  6161=>"00000101",
  6162=>"00000011",
  6163=>"00000000",
  6164=>"00000000",
  6165=>"11111110",
  6166=>"11111110",
  6167=>"11111101",
  6168=>"11111111",
  6169=>"11111111",
  6170=>"00000000",
  6171=>"00001000",
  6172=>"00000001",
  6173=>"00000010",
  6174=>"11111101",
  6175=>"00000001",
  6176=>"11111111",
  6177=>"00000111",
  6178=>"11111111",
  6179=>"00000010",
  6180=>"00000011",
  6181=>"00000000",
  6182=>"00000100",
  6183=>"11111101",
  6184=>"11111101",
  6185=>"00000110",
  6186=>"11111011",
  6187=>"00000110",
  6188=>"00000001",
  6189=>"11111110",
  6190=>"11111101",
  6191=>"11111111",
  6192=>"11111101",
  6193=>"11111100",
  6194=>"11111110",
  6195=>"00000010",
  6196=>"11111111",
  6197=>"00000000",
  6198=>"00000001",
  6199=>"00000000",
  6200=>"00000000",
  6201=>"00000101",
  6202=>"00000010",
  6203=>"00000001",
  6204=>"00000000",
  6205=>"00000010",
  6206=>"00000000",
  6207=>"11111101",
  6208=>"00000100",
  6209=>"00000000",
  6210=>"00000101",
  6211=>"00000001",
  6212=>"11111111",
  6213=>"00000011",
  6214=>"00000100",
  6215=>"11111110",
  6216=>"11111111",
  6217=>"00000001",
  6218=>"11111101",
  6219=>"00000101",
  6220=>"00000011",
  6221=>"11111110",
  6222=>"00000000",
  6223=>"00000010",
  6224=>"11111111",
  6225=>"00000010",
  6226=>"00000001",
  6227=>"00000001",
  6228=>"11111101",
  6229=>"11111100",
  6230=>"00000001",
  6231=>"00000001",
  6232=>"00000010",
  6233=>"11111110",
  6234=>"11111111",
  6235=>"00000010",
  6236=>"00000001",
  6237=>"00000001",
  6238=>"00000001",
  6239=>"11111111",
  6240=>"00000000",
  6241=>"00000010",
  6242=>"00000100",
  6243=>"11111110",
  6244=>"11111111",
  6245=>"11111111",
  6246=>"00000001",
  6247=>"00000110",
  6248=>"11111101",
  6249=>"00000000",
  6250=>"00000110",
  6251=>"00000001",
  6252=>"00000001",
  6253=>"00000001",
  6254=>"00000011",
  6255=>"11111011",
  6256=>"11111011",
  6257=>"11111110",
  6258=>"00000011",
  6259=>"11111101",
  6260=>"11111101",
  6261=>"11111110",
  6262=>"11111110",
  6263=>"11111110",
  6264=>"11111101",
  6265=>"00000011",
  6266=>"00000001",
  6267=>"00000010",
  6268=>"11111101",
  6269=>"00000001",
  6270=>"11111110",
  6271=>"00000100",
  6272=>"00000010",
  6273=>"11111101",
  6274=>"11111111",
  6275=>"00000010",
  6276=>"00000000",
  6277=>"00000101",
  6278=>"00000010",
  6279=>"00000011",
  6280=>"00000001",
  6281=>"00000010",
  6282=>"00000000",
  6283=>"00000000",
  6284=>"11111111",
  6285=>"11111101",
  6286=>"11111110",
  6287=>"00000001",
  6288=>"00000001",
  6289=>"00000001",
  6290=>"00000001",
  6291=>"00000000",
  6292=>"00000001",
  6293=>"00000011",
  6294=>"00000001",
  6295=>"00000001",
  6296=>"00000001",
  6297=>"00000000",
  6298=>"00000000",
  6299=>"00000000",
  6300=>"11111110",
  6301=>"00000100",
  6302=>"11111111",
  6303=>"00000000",
  6304=>"00000001",
  6305=>"00000011",
  6306=>"00000001",
  6307=>"00000010",
  6308=>"00000000",
  6309=>"11111110",
  6310=>"11111101",
  6311=>"11111101",
  6312=>"11111101",
  6313=>"00000111",
  6314=>"11111110",
  6315=>"00000001",
  6316=>"11111101",
  6317=>"00000001",
  6318=>"00000011",
  6319=>"00000001",
  6320=>"00000001",
  6321=>"00000001",
  6322=>"11111011",
  6323=>"11111101",
  6324=>"00000101",
  6325=>"00000010",
  6326=>"00000000",
  6327=>"11111101",
  6328=>"00000010",
  6329=>"00000000",
  6330=>"00000000",
  6331=>"11111011",
  6332=>"00000111",
  6333=>"00000011",
  6334=>"00000001",
  6335=>"00000011",
  6336=>"00000010",
  6337=>"11111101",
  6338=>"11111110",
  6339=>"00000001",
  6340=>"00000000",
  6341=>"00000000",
  6342=>"00000001",
  6343=>"11111110",
  6344=>"11111111",
  6345=>"00000110",
  6346=>"00000001",
  6347=>"00000100",
  6348=>"00000001",
  6349=>"11111110",
  6350=>"11111110",
  6351=>"00000001",
  6352=>"00000011",
  6353=>"00000000",
  6354=>"00000000",
  6355=>"11111110",
  6356=>"00000010",
  6357=>"11111110",
  6358=>"00000001",
  6359=>"00000010",
  6360=>"11111111",
  6361=>"00000101",
  6362=>"00000010",
  6363=>"11111110",
  6364=>"00000000",
  6365=>"00000000",
  6366=>"11111100",
  6367=>"00000010",
  6368=>"11111111",
  6369=>"11111111",
  6370=>"11111101",
  6371=>"00000000",
  6372=>"00000011",
  6373=>"00000001",
  6374=>"11111101",
  6375=>"11111110",
  6376=>"00000001",
  6377=>"00000101",
  6378=>"00000001",
  6379=>"11111110",
  6380=>"11111101",
  6381=>"11111101",
  6382=>"00000001",
  6383=>"00000001",
  6384=>"00000000",
  6385=>"11111101",
  6386=>"00000100",
  6387=>"11111101",
  6388=>"11111110",
  6389=>"11111111",
  6390=>"00000010",
  6391=>"11111110",
  6392=>"11111111",
  6393=>"00000001",
  6394=>"11111111",
  6395=>"11111111",
  6396=>"00000011",
  6397=>"00000000",
  6398=>"00000100",
  6399=>"11111101",
  6400=>"00000010",
  6401=>"00000111",
  6402=>"11111011",
  6403=>"00000001",
  6404=>"00000001",
  6405=>"11111111",
  6406=>"11111101",
  6407=>"11111101",
  6408=>"00000011",
  6409=>"00000100",
  6410=>"00000000",
  6411=>"11111011",
  6412=>"11111101",
  6413=>"00000001",
  6414=>"00000000",
  6415=>"00000001",
  6416=>"00000100",
  6417=>"00000001",
  6418=>"11111111",
  6419=>"11111010",
  6420=>"11111111",
  6421=>"11111110",
  6422=>"00000000",
  6423=>"11111110",
  6424=>"11111101",
  6425=>"00000100",
  6426=>"00000001",
  6427=>"00000001",
  6428=>"11111111",
  6429=>"00000001",
  6430=>"00000100",
  6431=>"00000001",
  6432=>"11111111",
  6433=>"00000011",
  6434=>"11111101",
  6435=>"00000010",
  6436=>"11111111",
  6437=>"11111111",
  6438=>"00000011",
  6439=>"00000111",
  6440=>"11111110",
  6441=>"11111111",
  6442=>"11111101",
  6443=>"11111111",
  6444=>"00000000",
  6445=>"00000010",
  6446=>"00000001",
  6447=>"11111100",
  6448=>"00000000",
  6449=>"00000010",
  6450=>"11111100",
  6451=>"00000001",
  6452=>"00000011",
  6453=>"00000010",
  6454=>"00000010",
  6455=>"00000000",
  6456=>"11111110",
  6457=>"00000000",
  6458=>"11111110",
  6459=>"00000100",
  6460=>"11111110",
  6461=>"11111101",
  6462=>"11111101",
  6463=>"00000000",
  6464=>"11111110",
  6465=>"11111110",
  6466=>"11111110",
  6467=>"11111101",
  6468=>"11111111",
  6469=>"11111111",
  6470=>"11111100",
  6471=>"00000010",
  6472=>"00000001",
  6473=>"11111110",
  6474=>"11111111",
  6475=>"00000010",
  6476=>"00000101",
  6477=>"11111110",
  6478=>"00000100",
  6479=>"11111111",
  6480=>"00000011",
  6481=>"00000011",
  6482=>"00000001",
  6483=>"00000001",
  6484=>"11111110",
  6485=>"00000001",
  6486=>"11111100",
  6487=>"00000001",
  6488=>"11111011",
  6489=>"11111110",
  6490=>"00000001",
  6491=>"11111110",
  6492=>"11111111",
  6493=>"00000000",
  6494=>"11111111",
  6495=>"11111101",
  6496=>"00000011",
  6497=>"00000101",
  6498=>"00000000",
  6499=>"11111100",
  6500=>"11111110",
  6501=>"11111111",
  6502=>"00000010",
  6503=>"00000000",
  6504=>"00000010",
  6505=>"11111100",
  6506=>"11111111",
  6507=>"00000001",
  6508=>"00000001",
  6509=>"11111111",
  6510=>"00000001",
  6511=>"00000010",
  6512=>"11111110",
  6513=>"11111110",
  6514=>"00000000",
  6515=>"00000001",
  6516=>"00000010",
  6517=>"00000011",
  6518=>"11111110",
  6519=>"00000011",
  6520=>"00000011",
  6521=>"00000010",
  6522=>"00000111",
  6523=>"00000010",
  6524=>"11111111",
  6525=>"00000001",
  6526=>"00000000",
  6527=>"00000100",
  6528=>"11111100",
  6529=>"00000100",
  6530=>"00000010",
  6531=>"11111110",
  6532=>"11111111",
  6533=>"00000011",
  6534=>"00000010",
  6535=>"00000100",
  6536=>"00000000",
  6537=>"11111110",
  6538=>"00000000",
  6539=>"00000011",
  6540=>"00000000",
  6541=>"11111101",
  6542=>"00000001",
  6543=>"00000010",
  6544=>"11111111",
  6545=>"11111110",
  6546=>"11111001",
  6547=>"11111100",
  6548=>"00000101",
  6549=>"11111101",
  6550=>"11111101",
  6551=>"00000011",
  6552=>"00000101",
  6553=>"00000101",
  6554=>"00000001",
  6555=>"00000010",
  6556=>"00000000",
  6557=>"00000000",
  6558=>"00000110",
  6559=>"00000001",
  6560=>"00000011",
  6561=>"00000010",
  6562=>"00000011",
  6563=>"00000101",
  6564=>"11111111",
  6565=>"00000001",
  6566=>"00000011",
  6567=>"00000101",
  6568=>"00000010",
  6569=>"11111110",
  6570=>"00000000",
  6571=>"00000010",
  6572=>"11111110",
  6573=>"00000000",
  6574=>"00000101",
  6575=>"00000010",
  6576=>"00000110",
  6577=>"00000001",
  6578=>"00000010",
  6579=>"00000100",
  6580=>"11111110",
  6581=>"11111010",
  6582=>"00000000",
  6583=>"00000110",
  6584=>"11111010",
  6585=>"00000100",
  6586=>"00000010",
  6587=>"00000001",
  6588=>"00000000",
  6589=>"00000001",
  6590=>"00000010",
  6591=>"11111101",
  6592=>"11111111",
  6593=>"00000000",
  6594=>"00000110",
  6595=>"11111101",
  6596=>"11111100",
  6597=>"00000011",
  6598=>"11111011",
  6599=>"00000100",
  6600=>"11111110",
  6601=>"00000000",
  6602=>"00000000",
  6603=>"00000001",
  6604=>"00000111",
  6605=>"11111101",
  6606=>"11111111",
  6607=>"00000001",
  6608=>"11111101",
  6609=>"11111101",
  6610=>"00000010",
  6611=>"11111101",
  6612=>"00000001",
  6613=>"11111110",
  6614=>"11111101",
  6615=>"11111111",
  6616=>"11111111",
  6617=>"00000001",
  6618=>"00000000",
  6619=>"00000010",
  6620=>"11111100",
  6621=>"00000001",
  6622=>"00000010",
  6623=>"11111110",
  6624=>"11111010",
  6625=>"00000011",
  6626=>"00000011",
  6627=>"11111101",
  6628=>"00000001",
  6629=>"00000001",
  6630=>"00000011",
  6631=>"00000011",
  6632=>"00000000",
  6633=>"11111111",
  6634=>"11111110",
  6635=>"11111101",
  6636=>"11111011",
  6637=>"00000001",
  6638=>"00000010",
  6639=>"11111101",
  6640=>"00000001",
  6641=>"00000011",
  6642=>"00000000",
  6643=>"11111110",
  6644=>"00000010",
  6645=>"00000010",
  6646=>"00000010",
  6647=>"11111101",
  6648=>"00000000",
  6649=>"00000100",
  6650=>"00000100",
  6651=>"00000010",
  6652=>"00000011",
  6653=>"00000101",
  6654=>"11111100",
  6655=>"11111111",
  6656=>"00000000",
  6657=>"00000001",
  6658=>"00000001",
  6659=>"11111110",
  6660=>"00000010",
  6661=>"00000001",
  6662=>"00000110",
  6663=>"00000010",
  6664=>"00000001",
  6665=>"11111101",
  6666=>"00000001",
  6667=>"11111101",
  6668=>"00000011",
  6669=>"00000001",
  6670=>"11111111",
  6671=>"00000010",
  6672=>"11111110",
  6673=>"11111101",
  6674=>"00000010",
  6675=>"11111101",
  6676=>"00000101",
  6677=>"11111110",
  6678=>"00000001",
  6679=>"11111101",
  6680=>"00000001",
  6681=>"11111111",
  6682=>"00000101",
  6683=>"00000010",
  6684=>"00000010",
  6685=>"11111101",
  6686=>"11111111",
  6687=>"00000001",
  6688=>"00000100",
  6689=>"00000001",
  6690=>"11111111",
  6691=>"00000001",
  6692=>"11111111",
  6693=>"00000000",
  6694=>"11111111",
  6695=>"11111111",
  6696=>"00000001",
  6697=>"11111101",
  6698=>"00000000",
  6699=>"00000100",
  6700=>"00000101",
  6701=>"00000011",
  6702=>"00000000",
  6703=>"00000110",
  6704=>"00000000",
  6705=>"11111110",
  6706=>"11111101",
  6707=>"11111111",
  6708=>"00000000",
  6709=>"00000001",
  6710=>"00000000",
  6711=>"00000010",
  6712=>"00000100",
  6713=>"11111111",
  6714=>"00000000",
  6715=>"00000011",
  6716=>"00000001",
  6717=>"00000011",
  6718=>"11111110",
  6719=>"11111111",
  6720=>"00000100",
  6721=>"00000100",
  6722=>"00000100",
  6723=>"00000010",
  6724=>"11111101",
  6725=>"11111111",
  6726=>"11111111",
  6727=>"11111101",
  6728=>"11111111",
  6729=>"00000100",
  6730=>"00000101",
  6731=>"11111111",
  6732=>"00000000",
  6733=>"00000000",
  6734=>"11111101",
  6735=>"00000001",
  6736=>"00000011",
  6737=>"00000000",
  6738=>"00000001",
  6739=>"00000000",
  6740=>"00000010",
  6741=>"11111101",
  6742=>"11111110",
  6743=>"00000010",
  6744=>"00000000",
  6745=>"00000000",
  6746=>"00000001",
  6747=>"00000010",
  6748=>"11111110",
  6749=>"00000011",
  6750=>"11111100",
  6751=>"00000010",
  6752=>"00000000",
  6753=>"11111111",
  6754=>"00000100",
  6755=>"00000001",
  6756=>"00000000",
  6757=>"00000011",
  6758=>"11111101",
  6759=>"00000100",
  6760=>"00000001",
  6761=>"00000010",
  6762=>"11111110",
  6763=>"00000000",
  6764=>"00000000",
  6765=>"11111110",
  6766=>"00000011",
  6767=>"11111110",
  6768=>"00000000",
  6769=>"00000100",
  6770=>"00000010",
  6771=>"00000011",
  6772=>"11111101",
  6773=>"00000001",
  6774=>"11111111",
  6775=>"00000011",
  6776=>"11111110",
  6777=>"00000110",
  6778=>"00000000",
  6779=>"00000011",
  6780=>"00000001",
  6781=>"00000000",
  6782=>"00000010",
  6783=>"11111111",
  6784=>"00000010",
  6785=>"11111101",
  6786=>"11111101",
  6787=>"00000000",
  6788=>"11111101",
  6789=>"00000010",
  6790=>"00000000",
  6791=>"00000010",
  6792=>"11111100",
  6793=>"11111101",
  6794=>"00000010",
  6795=>"00000000",
  6796=>"00000001",
  6797=>"00000001",
  6798=>"00000100",
  6799=>"11111101",
  6800=>"00000010",
  6801=>"11111110",
  6802=>"00000101",
  6803=>"00000001",
  6804=>"11111100",
  6805=>"00000000",
  6806=>"11111110",
  6807=>"00000000",
  6808=>"11111110",
  6809=>"00000001",
  6810=>"00000000",
  6811=>"00000001",
  6812=>"00000001",
  6813=>"00000100",
  6814=>"11111101",
  6815=>"11111101",
  6816=>"00000011",
  6817=>"00000000",
  6818=>"11111111",
  6819=>"00000111",
  6820=>"00000011",
  6821=>"00000001",
  6822=>"00000010",
  6823=>"00000011",
  6824=>"11111111",
  6825=>"11111111",
  6826=>"11111110",
  6827=>"00000101",
  6828=>"11111110",
  6829=>"00000011",
  6830=>"11111110",
  6831=>"00000010",
  6832=>"11111111",
  6833=>"11111111",
  6834=>"00000001",
  6835=>"00000000",
  6836=>"11111110",
  6837=>"11111101",
  6838=>"00000001",
  6839=>"11111110",
  6840=>"00000101",
  6841=>"11111101",
  6842=>"11111111",
  6843=>"11111110",
  6844=>"00000100",
  6845=>"00000011",
  6846=>"11111101",
  6847=>"00000010",
  6848=>"00000011",
  6849=>"00000010",
  6850=>"00000000",
  6851=>"00000010",
  6852=>"00000001",
  6853=>"11111111",
  6854=>"11111111",
  6855=>"00000101",
  6856=>"00000000",
  6857=>"00000100",
  6858=>"00000100",
  6859=>"00000010",
  6860=>"00000011",
  6861=>"11111100",
  6862=>"00000000",
  6863=>"00000010",
  6864=>"11111111",
  6865=>"00000001",
  6866=>"00000000",
  6867=>"00000011",
  6868=>"11111101",
  6869=>"00000011",
  6870=>"11111110",
  6871=>"11111011",
  6872=>"11111101",
  6873=>"11111110",
  6874=>"11111111",
  6875=>"00000011",
  6876=>"00000101",
  6877=>"00000001",
  6878=>"11111111",
  6879=>"00000101",
  6880=>"00000011",
  6881=>"11111101",
  6882=>"11111101",
  6883=>"11111111",
  6884=>"11111110",
  6885=>"00000011",
  6886=>"11111110",
  6887=>"00000101",
  6888=>"00000010",
  6889=>"11111101",
  6890=>"00000011",
  6891=>"11111110",
  6892=>"11111111",
  6893=>"00000010",
  6894=>"11111011",
  6895=>"00000010",
  6896=>"00000001",
  6897=>"11111101",
  6898=>"11111110",
  6899=>"00000001",
  6900=>"11111110",
  6901=>"00000000",
  6902=>"00000011",
  6903=>"11111101",
  6904=>"00000110",
  6905=>"00000000",
  6906=>"00000010",
  6907=>"00000100",
  6908=>"00000001",
  6909=>"00000000",
  6910=>"11111111",
  6911=>"11111111",
  6912=>"00000000",
  6913=>"11111101",
  6914=>"00000001",
  6915=>"00000010",
  6916=>"00000010",
  6917=>"00000011",
  6918=>"00000010",
  6919=>"11111111",
  6920=>"00000010",
  6921=>"00000011",
  6922=>"00000000",
  6923=>"11111110",
  6924=>"00000000",
  6925=>"11111111",
  6926=>"00000100",
  6927=>"11111100",
  6928=>"00000101",
  6929=>"00000010",
  6930=>"00000100",
  6931=>"00000100",
  6932=>"11111111",
  6933=>"00000000",
  6934=>"00000011",
  6935=>"00000110",
  6936=>"11111101",
  6937=>"00000100",
  6938=>"00000100",
  6939=>"11111110",
  6940=>"00000001",
  6941=>"00000000",
  6942=>"00000010",
  6943=>"00000011",
  6944=>"00000000",
  6945=>"11111110",
  6946=>"00000010",
  6947=>"11111111",
  6948=>"11111101",
  6949=>"00000010",
  6950=>"11111110",
  6951=>"00000000",
  6952=>"00000011",
  6953=>"00000101",
  6954=>"11111110",
  6955=>"11111110",
  6956=>"00000000",
  6957=>"00000100",
  6958=>"11111101",
  6959=>"11111011",
  6960=>"00000011",
  6961=>"00000100",
  6962=>"11111111",
  6963=>"11111011",
  6964=>"11111111",
  6965=>"00000100",
  6966=>"11111101",
  6967=>"00000101",
  6968=>"00000100",
  6969=>"00000010",
  6970=>"11111111",
  6971=>"11111110",
  6972=>"11111110",
  6973=>"00000100",
  6974=>"11111110",
  6975=>"00000001",
  6976=>"11111111",
  6977=>"00000111",
  6978=>"00000011",
  6979=>"00000001",
  6980=>"11111101",
  6981=>"11111110",
  6982=>"00000011",
  6983=>"11111101",
  6984=>"11111011",
  6985=>"00000010",
  6986=>"11111111",
  6987=>"11111111",
  6988=>"00000001",
  6989=>"00000100",
  6990=>"00000011",
  6991=>"00000010",
  6992=>"11111111",
  6993=>"00000001",
  6994=>"00000010",
  6995=>"00000011",
  6996=>"00000011",
  6997=>"00000100",
  6998=>"00000001",
  6999=>"00000010",
  7000=>"00000001",
  7001=>"11111111",
  7002=>"00000101",
  7003=>"00000100",
  7004=>"11111110",
  7005=>"11111110",
  7006=>"11111111",
  7007=>"11111110",
  7008=>"00000100",
  7009=>"00000010",
  7010=>"11111101",
  7011=>"11111110",
  7012=>"11111110",
  7013=>"00000000",
  7014=>"00000000",
  7015=>"00000000",
  7016=>"00000000",
  7017=>"00000100",
  7018=>"00000001",
  7019=>"00000000",
  7020=>"00000100",
  7021=>"00000100",
  7022=>"11111110",
  7023=>"11111110",
  7024=>"00000010",
  7025=>"00000101",
  7026=>"11111110",
  7027=>"00000001",
  7028=>"00000010",
  7029=>"11111011",
  7030=>"11111100",
  7031=>"00000000",
  7032=>"00000001",
  7033=>"00000011",
  7034=>"11111101",
  7035=>"00000010",
  7036=>"11111100",
  7037=>"00000000",
  7038=>"11111110",
  7039=>"11111110",
  7040=>"11111111",
  7041=>"11111101",
  7042=>"00000000",
  7043=>"00000011",
  7044=>"00000001",
  7045=>"00000011",
  7046=>"00000010",
  7047=>"11111101",
  7048=>"00000101",
  7049=>"00000010",
  7050=>"00000000",
  7051=>"11111111",
  7052=>"11111011",
  7053=>"00000000",
  7054=>"11111100",
  7055=>"00000000",
  7056=>"00000000",
  7057=>"00000011",
  7058=>"00000011",
  7059=>"11111110",
  7060=>"00000000",
  7061=>"00000011",
  7062=>"11111111",
  7063=>"00000011",
  7064=>"00000100",
  7065=>"00000001",
  7066=>"00000001",
  7067=>"00000010",
  7068=>"11111110",
  7069=>"11111111",
  7070=>"00000101",
  7071=>"11111110",
  7072=>"00000001",
  7073=>"11111111",
  7074=>"00000100",
  7075=>"11111110",
  7076=>"00000000",
  7077=>"00000010",
  7078=>"11111111",
  7079=>"11111101",
  7080=>"00000100",
  7081=>"00000011",
  7082=>"11111111",
  7083=>"11111110",
  7084=>"00000000",
  7085=>"00000000",
  7086=>"00000001",
  7087=>"00000000",
  7088=>"00000110",
  7089=>"00000000",
  7090=>"00000001",
  7091=>"00000000",
  7092=>"11111100",
  7093=>"11111111",
  7094=>"11111111",
  7095=>"00000101",
  7096=>"00000010",
  7097=>"00000001",
  7098=>"00000010",
  7099=>"00000011",
  7100=>"11111111",
  7101=>"00000100",
  7102=>"00000000",
  7103=>"00000001",
  7104=>"11111100",
  7105=>"00000000",
  7106=>"00000110",
  7107=>"11111110",
  7108=>"00000010",
  7109=>"11111110",
  7110=>"00000001",
  7111=>"00000001",
  7112=>"11111100",
  7113=>"00000010",
  7114=>"00000011",
  7115=>"11111111",
  7116=>"11111110",
  7117=>"11111111",
  7118=>"11111110",
  7119=>"00000101",
  7120=>"00000001",
  7121=>"00000011",
  7122=>"00000000",
  7123=>"11111110",
  7124=>"11111111",
  7125=>"00000010",
  7126=>"11111110",
  7127=>"11111100",
  7128=>"11111110",
  7129=>"00000101",
  7130=>"11111110",
  7131=>"00000000",
  7132=>"00000000",
  7133=>"00000001",
  7134=>"11111110",
  7135=>"00000010",
  7136=>"00000100",
  7137=>"11111101",
  7138=>"00000011",
  7139=>"00000010",
  7140=>"00000000",
  7141=>"11111111",
  7142=>"11111111",
  7143=>"00000000",
  7144=>"11111110",
  7145=>"11111111",
  7146=>"00000001",
  7147=>"00000010",
  7148=>"11111101",
  7149=>"00000011",
  7150=>"11111111",
  7151=>"00000011",
  7152=>"00000100",
  7153=>"00000010",
  7154=>"00000010",
  7155=>"00000010",
  7156=>"11111110",
  7157=>"00000001",
  7158=>"00000011",
  7159=>"00000010",
  7160=>"00000101",
  7161=>"00000010",
  7162=>"00000011",
  7163=>"11111111",
  7164=>"00000011",
  7165=>"00000100",
  7166=>"11111110",
  7167=>"11111111",
  7168=>"11111101",
  7169=>"11111101",
  7170=>"00000100",
  7171=>"11111110",
  7172=>"00000001",
  7173=>"11111111",
  7174=>"00000001",
  7175=>"00000011",
  7176=>"11111110",
  7177=>"11111110",
  7178=>"11111111",
  7179=>"11111110",
  7180=>"00000000",
  7181=>"00000010",
  7182=>"11111100",
  7183=>"11111100",
  7184=>"11111111",
  7185=>"00000101",
  7186=>"00000100",
  7187=>"00000001",
  7188=>"00000101",
  7189=>"00000100",
  7190=>"00000001",
  7191=>"00000001",
  7192=>"00000010",
  7193=>"00000010",
  7194=>"11111110",
  7195=>"11111110",
  7196=>"00000010",
  7197=>"11111111",
  7198=>"11111111",
  7199=>"00000010",
  7200=>"11111110",
  7201=>"00000000",
  7202=>"11111101",
  7203=>"11111111",
  7204=>"00000100",
  7205=>"00000100",
  7206=>"11111111",
  7207=>"11111101",
  7208=>"11111110",
  7209=>"00000000",
  7210=>"11111110",
  7211=>"00000011",
  7212=>"11111110",
  7213=>"11111111",
  7214=>"00000000",
  7215=>"00000001",
  7216=>"00000000",
  7217=>"00000001",
  7218=>"11111110",
  7219=>"11111110",
  7220=>"11111111",
  7221=>"11111101",
  7222=>"11111110",
  7223=>"11111101",
  7224=>"00000010",
  7225=>"11111100",
  7226=>"11111101",
  7227=>"00000101",
  7228=>"11111111",
  7229=>"00000001",
  7230=>"00000000",
  7231=>"00000001",
  7232=>"11111110",
  7233=>"00000000",
  7234=>"11111101",
  7235=>"11111101",
  7236=>"00000000",
  7237=>"00000001",
  7238=>"11111101",
  7239=>"00000011",
  7240=>"00000000",
  7241=>"00000000",
  7242=>"00000000",
  7243=>"11111110",
  7244=>"00000010",
  7245=>"00000101",
  7246=>"00000010",
  7247=>"11111111",
  7248=>"00000010",
  7249=>"00000011",
  7250=>"11111110",
  7251=>"00000001",
  7252=>"11111110",
  7253=>"11111110",
  7254=>"00000010",
  7255=>"11111110",
  7256=>"11111111",
  7257=>"00000011",
  7258=>"00000010",
  7259=>"00000100",
  7260=>"00000001",
  7261=>"00000000",
  7262=>"00000010",
  7263=>"00000011",
  7264=>"00000011",
  7265=>"00000010",
  7266=>"00000010",
  7267=>"11111111",
  7268=>"00000001",
  7269=>"00000001",
  7270=>"11111101",
  7271=>"00000000",
  7272=>"11111110",
  7273=>"11111111",
  7274=>"11111110",
  7275=>"00000011",
  7276=>"11111111",
  7277=>"11111110",
  7278=>"11111101",
  7279=>"00000011",
  7280=>"11111110",
  7281=>"00000001",
  7282=>"00000011",
  7283=>"11111110",
  7284=>"00000011",
  7285=>"11111111",
  7286=>"11111101",
  7287=>"11111110",
  7288=>"11111110",
  7289=>"11111111",
  7290=>"11111111",
  7291=>"11111110",
  7292=>"11111110",
  7293=>"00000001",
  7294=>"00000001",
  7295=>"11111100",
  7296=>"00000001",
  7297=>"00000000",
  7298=>"11111111",
  7299=>"11111100",
  7300=>"11111101",
  7301=>"00000000",
  7302=>"00000000",
  7303=>"11111110",
  7304=>"00000010",
  7305=>"00000010",
  7306=>"11111110",
  7307=>"11111111",
  7308=>"00000100",
  7309=>"11111110",
  7310=>"11111111",
  7311=>"00000010",
  7312=>"00000000",
  7313=>"00000011",
  7314=>"00000100",
  7315=>"11111111",
  7316=>"00000000",
  7317=>"11111101",
  7318=>"00000000",
  7319=>"00000001",
  7320=>"11111101",
  7321=>"00000000",
  7322=>"00000010",
  7323=>"00000000",
  7324=>"11111110",
  7325=>"11111110",
  7326=>"00000001",
  7327=>"11111111",
  7328=>"00000010",
  7329=>"11111111",
  7330=>"00000011",
  7331=>"00000010",
  7332=>"00000010",
  7333=>"11111101",
  7334=>"11111110",
  7335=>"00000000",
  7336=>"00000100",
  7337=>"00000000",
  7338=>"00000000",
  7339=>"00000000",
  7340=>"00000010",
  7341=>"11111111",
  7342=>"11111111",
  7343=>"11111101",
  7344=>"00000100",
  7345=>"00000000",
  7346=>"00000011",
  7347=>"11111111",
  7348=>"00000000",
  7349=>"11111100",
  7350=>"11111101",
  7351=>"00000010",
  7352=>"11111111",
  7353=>"00000011",
  7354=>"11111111",
  7355=>"00000001",
  7356=>"11111111",
  7357=>"00000011",
  7358=>"11111110",
  7359=>"11111100",
  7360=>"11111100",
  7361=>"00000001",
  7362=>"00000110",
  7363=>"11111111",
  7364=>"00000001",
  7365=>"00000010",
  7366=>"11111101",
  7367=>"00000000",
  7368=>"11111111",
  7369=>"00000010",
  7370=>"00000101",
  7371=>"11111100",
  7372=>"00000011",
  7373=>"00000000",
  7374=>"11111111",
  7375=>"00000010",
  7376=>"00000010",
  7377=>"00000010",
  7378=>"11111111",
  7379=>"00000001",
  7380=>"00000011",
  7381=>"00000000",
  7382=>"11111110",
  7383=>"11111110",
  7384=>"00000000",
  7385=>"00000001",
  7386=>"00000011",
  7387=>"00000000",
  7388=>"00000010",
  7389=>"11111100",
  7390=>"00000000",
  7391=>"00000011",
  7392=>"00000001",
  7393=>"00000000",
  7394=>"00000000",
  7395=>"11111111",
  7396=>"11111111",
  7397=>"00000010",
  7398=>"00000010",
  7399=>"00000010",
  7400=>"00000000",
  7401=>"00000001",
  7402=>"00000001",
  7403=>"00000000",
  7404=>"11111110",
  7405=>"11111101",
  7406=>"00000000",
  7407=>"00000011",
  7408=>"00000011",
  7409=>"00000001",
  7410=>"00000000",
  7411=>"00000010",
  7412=>"11111110",
  7413=>"00000001",
  7414=>"11111110",
  7415=>"11111110",
  7416=>"00000001",
  7417=>"11111111",
  7418=>"00000001",
  7419=>"00000000",
  7420=>"11111110",
  7421=>"00000001",
  7422=>"11111101",
  7423=>"00000010",
  7424=>"11111110",
  7425=>"00000010",
  7426=>"11111100",
  7427=>"00000001",
  7428=>"11111110",
  7429=>"11111111",
  7430=>"11111111",
  7431=>"00000001",
  7432=>"11111110",
  7433=>"11111100",
  7434=>"00000010",
  7435=>"00000001",
  7436=>"11111110",
  7437=>"00000001",
  7438=>"11111111",
  7439=>"11111101",
  7440=>"11111101",
  7441=>"00000001",
  7442=>"00000100",
  7443=>"11111100",
  7444=>"00000001",
  7445=>"11111110",
  7446=>"00000001",
  7447=>"11111110",
  7448=>"11111111",
  7449=>"00000000",
  7450=>"00000010",
  7451=>"00000010",
  7452=>"11111101",
  7453=>"11111110",
  7454=>"00000001",
  7455=>"11111110",
  7456=>"00000011",
  7457=>"00000001",
  7458=>"00000010",
  7459=>"11111110",
  7460=>"11111110",
  7461=>"11111101",
  7462=>"00000001",
  7463=>"00000000",
  7464=>"11111101",
  7465=>"00000001",
  7466=>"00000001",
  7467=>"11111111",
  7468=>"11111110",
  7469=>"11111110",
  7470=>"00000000",
  7471=>"11111100",
  7472=>"00000001",
  7473=>"00000010",
  7474=>"11111101",
  7475=>"11111110",
  7476=>"00000010",
  7477=>"00000000",
  7478=>"00000010",
  7479=>"11111111",
  7480=>"11111101",
  7481=>"00000001",
  7482=>"11111101",
  7483=>"11111101",
  7484=>"00000000",
  7485=>"00000001",
  7486=>"00000000",
  7487=>"00000000",
  7488=>"11111111",
  7489=>"11111100",
  7490=>"00000000",
  7491=>"00000011",
  7492=>"11111111",
  7493=>"11111111",
  7494=>"11111101",
  7495=>"00000010",
  7496=>"00000101",
  7497=>"11111101",
  7498=>"00000001",
  7499=>"00000010",
  7500=>"11111101",
  7501=>"11111111",
  7502=>"00000011",
  7503=>"00000001",
  7504=>"00000001",
  7505=>"11111101",
  7506=>"11111101",
  7507=>"11111111",
  7508=>"00000001",
  7509=>"00000010",
  7510=>"00000100",
  7511=>"00000000",
  7512=>"11111101",
  7513=>"00000010",
  7514=>"00000010",
  7515=>"00000001",
  7516=>"11111110",
  7517=>"11111111",
  7518=>"11111111",
  7519=>"00000000",
  7520=>"11111101",
  7521=>"00000001",
  7522=>"11111111",
  7523=>"00000001",
  7524=>"11111111",
  7525=>"00000001",
  7526=>"00000000",
  7527=>"11111101",
  7528=>"11111111",
  7529=>"00000000",
  7530=>"11111110",
  7531=>"00000001",
  7532=>"00000010",
  7533=>"11111101",
  7534=>"11111101",
  7535=>"00000000",
  7536=>"11111110",
  7537=>"11111110",
  7538=>"00000010",
  7539=>"00000010",
  7540=>"11111101",
  7541=>"00000100",
  7542=>"00000000",
  7543=>"11111111",
  7544=>"11111111",
  7545=>"11111110",
  7546=>"00000111",
  7547=>"11111111",
  7548=>"00000001",
  7549=>"11111110",
  7550=>"11111110",
  7551=>"00000001",
  7552=>"11111101",
  7553=>"11111110",
  7554=>"00000011",
  7555=>"00000000",
  7556=>"00000011",
  7557=>"00000001",
  7558=>"00000000",
  7559=>"00000000",
  7560=>"11111111",
  7561=>"00000011",
  7562=>"00000011",
  7563=>"00000010",
  7564=>"00000000",
  7565=>"11111111",
  7566=>"11111111",
  7567=>"11111110",
  7568=>"00000001",
  7569=>"00000001",
  7570=>"11111110",
  7571=>"11111111",
  7572=>"00000001",
  7573=>"00000011",
  7574=>"00000010",
  7575=>"11111101",
  7576=>"11111011",
  7577=>"11111111",
  7578=>"00000010",
  7579=>"00000000",
  7580=>"00000010",
  7581=>"00000011",
  7582=>"11111110",
  7583=>"11111101",
  7584=>"11111101",
  7585=>"11111110",
  7586=>"11111111",
  7587=>"00000110",
  7588=>"00000010",
  7589=>"00000001",
  7590=>"11111111",
  7591=>"00000011",
  7592=>"11111110",
  7593=>"11111111",
  7594=>"00000101",
  7595=>"00000100",
  7596=>"00000000",
  7597=>"11111110",
  7598=>"11111110",
  7599=>"11111110",
  7600=>"11111111",
  7601=>"00000101",
  7602=>"00000010",
  7603=>"11111110",
  7604=>"00000001",
  7605=>"11111111",
  7606=>"11111110",
  7607=>"00000001",
  7608=>"11111111",
  7609=>"00000100",
  7610=>"11111110",
  7611=>"11111101",
  7612=>"00000001",
  7613=>"11111100",
  7614=>"11111100",
  7615=>"00000000",
  7616=>"11111110",
  7617=>"00000000",
  7618=>"11111111",
  7619=>"00000101",
  7620=>"11111111",
  7621=>"00000010",
  7622=>"00000011",
  7623=>"11111111",
  7624=>"11111101",
  7625=>"00000010",
  7626=>"11111111",
  7627=>"00000001",
  7628=>"11111101",
  7629=>"00000011",
  7630=>"00000001",
  7631=>"00000010",
  7632=>"00000010",
  7633=>"00000001",
  7634=>"00000010",
  7635=>"11111100",
  7636=>"00000010",
  7637=>"11111111",
  7638=>"00000001",
  7639=>"11111101",
  7640=>"00000011",
  7641=>"00000010",
  7642=>"11111111",
  7643=>"11111111",
  7644=>"00000010",
  7645=>"11111111",
  7646=>"00000010",
  7647=>"11111100",
  7648=>"00000011",
  7649=>"00000000",
  7650=>"11111110",
  7651=>"00000000",
  7652=>"11111110",
  7653=>"00000101",
  7654=>"00000010",
  7655=>"11111111",
  7656=>"00000000",
  7657=>"11111111",
  7658=>"00000010",
  7659=>"00000101",
  7660=>"00000011",
  7661=>"00000010",
  7662=>"11111111",
  7663=>"11111111",
  7664=>"11111110",
  7665=>"11111110",
  7666=>"00000000",
  7667=>"11111101",
  7668=>"11111111",
  7669=>"11111110",
  7670=>"11111101",
  7671=>"11111110",
  7672=>"11111110",
  7673=>"11111101",
  7674=>"00000000",
  7675=>"00000011",
  7676=>"11111111",
  7677=>"11111110",
  7678=>"11111110",
  7679=>"00000000",
  7680=>"00000001",
  7681=>"11111111",
  7682=>"11111101",
  7683=>"00000011",
  7684=>"00000100",
  7685=>"11111101",
  7686=>"11111110",
  7687=>"00000010",
  7688=>"00000000",
  7689=>"00000100",
  7690=>"00000001",
  7691=>"11111111",
  7692=>"00000000",
  7693=>"00000100",
  7694=>"00000001",
  7695=>"00000000",
  7696=>"11111101",
  7697=>"11111110",
  7698=>"11111111",
  7699=>"11111111",
  7700=>"11111111",
  7701=>"00000001",
  7702=>"00000000",
  7703=>"00000001",
  7704=>"00000010",
  7705=>"11111101",
  7706=>"00000001",
  7707=>"11111111",
  7708=>"11111111",
  7709=>"11111111",
  7710=>"00000100",
  7711=>"00000110",
  7712=>"00000001",
  7713=>"00000000",
  7714=>"00000100",
  7715=>"00000001",
  7716=>"00000000",
  7717=>"00000011",
  7718=>"11111111",
  7719=>"00000001",
  7720=>"00000010",
  7721=>"00000101",
  7722=>"11111111",
  7723=>"11111111",
  7724=>"00000101",
  7725=>"00000100",
  7726=>"11111110",
  7727=>"11111111",
  7728=>"11111101",
  7729=>"00000011",
  7730=>"00000001",
  7731=>"00000010",
  7732=>"00000000",
  7733=>"11111101",
  7734=>"11111111",
  7735=>"11111111",
  7736=>"11111110",
  7737=>"00000011",
  7738=>"00000000",
  7739=>"00000000",
  7740=>"00000000",
  7741=>"11111101",
  7742=>"00000001",
  7743=>"11111110",
  7744=>"11111111",
  7745=>"11111111",
  7746=>"00000010",
  7747=>"00000010",
  7748=>"11111101",
  7749=>"11111111",
  7750=>"00000001",
  7751=>"00000011",
  7752=>"11111101",
  7753=>"00000010",
  7754=>"00000000",
  7755=>"11111111",
  7756=>"00000011",
  7757=>"11111111",
  7758=>"00000000",
  7759=>"11111111",
  7760=>"00000100",
  7761=>"00000001",
  7762=>"00000010",
  7763=>"00000000",
  7764=>"00000011",
  7765=>"00000000",
  7766=>"00000010",
  7767=>"11111101",
  7768=>"11111101",
  7769=>"11111101",
  7770=>"00000000",
  7771=>"00000000",
  7772=>"11111111",
  7773=>"00000100",
  7774=>"00000011",
  7775=>"00000010",
  7776=>"11111111",
  7777=>"11111111",
  7778=>"00000000",
  7779=>"00000000",
  7780=>"00000010",
  7781=>"00000000",
  7782=>"11111111",
  7783=>"00000001",
  7784=>"00000000",
  7785=>"00000001",
  7786=>"00000011",
  7787=>"11111111",
  7788=>"00000011",
  7789=>"11111110",
  7790=>"00000000",
  7791=>"00000111",
  7792=>"00000011",
  7793=>"11111111",
  7794=>"11111111",
  7795=>"00000100",
  7796=>"00000010",
  7797=>"00000010",
  7798=>"00000101",
  7799=>"00000100",
  7800=>"11111101",
  7801=>"00000001",
  7802=>"00000000",
  7803=>"00000000",
  7804=>"00000000",
  7805=>"11111111",
  7806=>"11111110",
  7807=>"00000001",
  7808=>"00000010",
  7809=>"11111111",
  7810=>"00000010",
  7811=>"11111111",
  7812=>"00000100",
  7813=>"11111101",
  7814=>"11111111",
  7815=>"00000000",
  7816=>"00000101",
  7817=>"11111101",
  7818=>"00000011",
  7819=>"00000001",
  7820=>"00000000",
  7821=>"11111111",
  7822=>"00000000",
  7823=>"11111110",
  7824=>"00000010",
  7825=>"00000010",
  7826=>"11111110",
  7827=>"00000000",
  7828=>"00000100",
  7829=>"11111110",
  7830=>"11111111",
  7831=>"00000011",
  7832=>"11111111",
  7833=>"11111100",
  7834=>"00000000",
  7835=>"00000011",
  7836=>"00000000",
  7837=>"11111100",
  7838=>"00000000",
  7839=>"11111110",
  7840=>"00000010",
  7841=>"11111111",
  7842=>"00000001",
  7843=>"11111111",
  7844=>"00000000",
  7845=>"11111101",
  7846=>"00000010",
  7847=>"11111111",
  7848=>"11111110",
  7849=>"11111101",
  7850=>"11111100",
  7851=>"11111111",
  7852=>"00000011",
  7853=>"00000010",
  7854=>"00000010",
  7855=>"00000000",
  7856=>"00000000",
  7857=>"00000011",
  7858=>"00000011",
  7859=>"00000000",
  7860=>"11111101",
  7861=>"00000000",
  7862=>"11111111",
  7863=>"00000000",
  7864=>"00000000",
  7865=>"00000100",
  7866=>"00000001",
  7867=>"11111101",
  7868=>"11111101",
  7869=>"11111101",
  7870=>"11111111",
  7871=>"00000000",
  7872=>"00000001",
  7873=>"11111101",
  7874=>"00000001",
  7875=>"11111111",
  7876=>"11111101",
  7877=>"00000011",
  7878=>"00000000",
  7879=>"11111111",
  7880=>"00000010",
  7881=>"00000001",
  7882=>"00000000",
  7883=>"11111111",
  7884=>"11111111",
  7885=>"11111111",
  7886=>"00000100",
  7887=>"00000100",
  7888=>"11111111",
  7889=>"00000011",
  7890=>"11111111",
  7891=>"11111111",
  7892=>"11111110",
  7893=>"00000001",
  7894=>"00000100",
  7895=>"00000010",
  7896=>"11111111",
  7897=>"00000001",
  7898=>"00000011",
  7899=>"00000010",
  7900=>"00000011",
  7901=>"00000000",
  7902=>"11111110",
  7903=>"11111110",
  7904=>"11111101",
  7905=>"11111110",
  7906=>"11111110",
  7907=>"00000000",
  7908=>"00000010",
  7909=>"00000011",
  7910=>"00000000",
  7911=>"00000000",
  7912=>"00000000",
  7913=>"11111110",
  7914=>"00000100",
  7915=>"00000100",
  7916=>"00000000",
  7917=>"00000000",
  7918=>"00000010",
  7919=>"00000001",
  7920=>"00000000",
  7921=>"11111110",
  7922=>"11111111",
  7923=>"00000010",
  7924=>"00000001",
  7925=>"11111110",
  7926=>"00000000",
  7927=>"11111111",
  7928=>"00000010",
  7929=>"11111111",
  7930=>"11111110",
  7931=>"11111111",
  7932=>"00000010",
  7933=>"11111111",
  7934=>"00000000",
  7935=>"00000011",
  7936=>"11111111",
  7937=>"00000110",
  7938=>"11111111",
  7939=>"11111101",
  7940=>"00000011",
  7941=>"00000011",
  7942=>"00000000",
  7943=>"00000001",
  7944=>"00000100",
  7945=>"11111110",
  7946=>"11111111",
  7947=>"11111110",
  7948=>"00000010",
  7949=>"11111101",
  7950=>"11111110",
  7951=>"00000000",
  7952=>"11111110",
  7953=>"00000010",
  7954=>"11111101",
  7955=>"00000001",
  7956=>"00000011",
  7957=>"00000100",
  7958=>"11111110",
  7959=>"00000000",
  7960=>"11111110",
  7961=>"11111101",
  7962=>"11111101",
  7963=>"00000100",
  7964=>"00000001",
  7965=>"00000001",
  7966=>"00000111",
  7967=>"11111110",
  7968=>"00000000",
  7969=>"11111110",
  7970=>"11111110",
  7971=>"00000000",
  7972=>"00000010",
  7973=>"00000000",
  7974=>"00000110",
  7975=>"00000010",
  7976=>"00000010",
  7977=>"11111110",
  7978=>"00000100",
  7979=>"00000011",
  7980=>"00000000",
  7981=>"11111111",
  7982=>"11111111",
  7983=>"00000001",
  7984=>"00000010",
  7985=>"11111110",
  7986=>"11111111",
  7987=>"00000010",
  7988=>"00000011",
  7989=>"00000010",
  7990=>"00000001",
  7991=>"11111100",
  7992=>"11111100",
  7993=>"00000010",
  7994=>"11111110",
  7995=>"00000100",
  7996=>"00000000",
  7997=>"00000011",
  7998=>"00000101",
  7999=>"11111101",
  8000=>"11111110",
  8001=>"11111111",
  8002=>"00000000",
  8003=>"11111101",
  8004=>"00000110",
  8005=>"00000000",
  8006=>"00000001",
  8007=>"00000011",
  8008=>"00000010",
  8009=>"00000001",
  8010=>"00000010",
  8011=>"11111110",
  8012=>"00000100",
  8013=>"00000011",
  8014=>"11111101",
  8015=>"00000100",
  8016=>"00000010",
  8017=>"00000001",
  8018=>"00000010",
  8019=>"00000100",
  8020=>"11111111",
  8021=>"11111111",
  8022=>"00000010",
  8023=>"11111111",
  8024=>"11111101",
  8025=>"00000100",
  8026=>"11111100",
  8027=>"11111111",
  8028=>"00000100",
  8029=>"11111101",
  8030=>"00000000",
  8031=>"11111101",
  8032=>"11111110",
  8033=>"11111101",
  8034=>"11111110",
  8035=>"11111101",
  8036=>"00000010",
  8037=>"00000100",
  8038=>"00000010",
  8039=>"00000000",
  8040=>"00000001",
  8041=>"11111111",
  8042=>"00000101",
  8043=>"00000000",
  8044=>"11111111",
  8045=>"00000001",
  8046=>"11111111",
  8047=>"11111111",
  8048=>"00000001",
  8049=>"11111101",
  8050=>"11111110",
  8051=>"00000001",
  8052=>"00000000",
  8053=>"00000010",
  8054=>"11111110",
  8055=>"00000000",
  8056=>"00000010",
  8057=>"00000000",
  8058=>"11111110",
  8059=>"00000010",
  8060=>"11111111",
  8061=>"00000100",
  8062=>"00000010",
  8063=>"00000010",
  8064=>"00000010",
  8065=>"11111011",
  8066=>"00000001",
  8067=>"00000000",
  8068=>"00000010",
  8069=>"00000010",
  8070=>"00000010",
  8071=>"11111110",
  8072=>"11111110",
  8073=>"00000010",
  8074=>"00000010",
  8075=>"00000000",
  8076=>"00000011",
  8077=>"11111101",
  8078=>"00000101",
  8079=>"11111111",
  8080=>"11111111",
  8081=>"00000101",
  8082=>"11111111",
  8083=>"00000011",
  8084=>"00000100",
  8085=>"00000000",
  8086=>"11111111",
  8087=>"00000101",
  8088=>"00000001",
  8089=>"11111111",
  8090=>"00000001",
  8091=>"11111101",
  8092=>"00000001",
  8093=>"00000001",
  8094=>"00000010",
  8095=>"00000011",
  8096=>"00000000",
  8097=>"00000001",
  8098=>"11111100",
  8099=>"00000000",
  8100=>"11111111",
  8101=>"00000011",
  8102=>"00000010",
  8103=>"00000000",
  8104=>"00000010",
  8105=>"00000001",
  8106=>"11111110",
  8107=>"00000001",
  8108=>"11111111",
  8109=>"11111101",
  8110=>"00000011",
  8111=>"00000001",
  8112=>"11111101",
  8113=>"00000010",
  8114=>"11111111",
  8115=>"11111101",
  8116=>"00000000",
  8117=>"00000001",
  8118=>"00000101",
  8119=>"11111101",
  8120=>"11111110",
  8121=>"00000001",
  8122=>"11111110",
  8123=>"11111110",
  8124=>"11111110",
  8125=>"11111101",
  8126=>"00000010",
  8127=>"00000001",
  8128=>"00000001",
  8129=>"00000001",
  8130=>"11111101",
  8131=>"11111101",
  8132=>"00000010",
  8133=>"00000010",
  8134=>"00000011",
  8135=>"00000000",
  8136=>"11111101",
  8137=>"00000011",
  8138=>"00000011",
  8139=>"00000000",
  8140=>"00000011",
  8141=>"00000010",
  8142=>"00000000",
  8143=>"00000001",
  8144=>"00000010",
  8145=>"00000001",
  8146=>"00000010",
  8147=>"11111111",
  8148=>"00000001",
  8149=>"00000101",
  8150=>"11111110",
  8151=>"11111111",
  8152=>"11111111",
  8153=>"00000001",
  8154=>"00000010",
  8155=>"11111111",
  8156=>"00000011",
  8157=>"00000010",
  8158=>"11111110",
  8159=>"11111111",
  8160=>"11111111",
  8161=>"11111110",
  8162=>"11111111",
  8163=>"00000010",
  8164=>"00000010",
  8165=>"00000010",
  8166=>"11111110",
  8167=>"11111110",
  8168=>"00000001",
  8169=>"11111111",
  8170=>"00000001",
  8171=>"11111111",
  8172=>"11111110",
  8173=>"00000011",
  8174=>"11111110",
  8175=>"00000011",
  8176=>"00000001",
  8177=>"11111110",
  8178=>"11111101",
  8179=>"11111111",
  8180=>"11111101",
  8181=>"11111111",
  8182=>"00000010",
  8183=>"11111110",
  8184=>"00000100",
  8185=>"00000001",
  8186=>"00000100",
  8187=>"00000001",
  8188=>"11111101",
  8189=>"11111101",
  8190=>"00000101",
  8191=>"11111110",
  8192=>"00000000",
  8193=>"11111101",
  8194=>"11111111",
  8195=>"11111111",
  8196=>"11111100",
  8197=>"11111111",
  8198=>"11111110",
  8199=>"00000001",
  8200=>"00000001",
  8201=>"00000101",
  8202=>"11111111",
  8203=>"00000101",
  8204=>"00000010",
  8205=>"00000000",
  8206=>"00000011",
  8207=>"00000000",
  8208=>"00000100",
  8209=>"11111100",
  8210=>"00000000",
  8211=>"00000010",
  8212=>"11111111",
  8213=>"00000000",
  8214=>"00000010",
  8215=>"00000000",
  8216=>"11111101",
  8217=>"11111101",
  8218=>"00000001",
  8219=>"11111110",
  8220=>"11111110",
  8221=>"00000000",
  8222=>"11111111",
  8223=>"11111110",
  8224=>"00000011",
  8225=>"00000001",
  8226=>"00000000",
  8227=>"00000001",
  8228=>"11111110",
  8229=>"00000001",
  8230=>"00000010",
  8231=>"00000011",
  8232=>"00000001",
  8233=>"00000000",
  8234=>"00000001",
  8235=>"11111110",
  8236=>"11111111",
  8237=>"00000100",
  8238=>"00000001",
  8239=>"11111111",
  8240=>"00000010",
  8241=>"11111110",
  8242=>"11111101",
  8243=>"11111110",
  8244=>"00000010",
  8245=>"11111110",
  8246=>"00000001",
  8247=>"00000110",
  8248=>"00000001",
  8249=>"00000001",
  8250=>"11111110",
  8251=>"00000000",
  8252=>"11111111",
  8253=>"00000001",
  8254=>"11111110",
  8255=>"00000001",
  8256=>"11111110",
  8257=>"00000011",
  8258=>"00000011",
  8259=>"00000000",
  8260=>"00000010",
  8261=>"11111111",
  8262=>"11111110",
  8263=>"11111110",
  8264=>"00000110",
  8265=>"00000001",
  8266=>"11111111",
  8267=>"11111111",
  8268=>"00000011",
  8269=>"11111110",
  8270=>"00000000",
  8271=>"11111110",
  8272=>"11111110",
  8273=>"00000001",
  8274=>"00000011",
  8275=>"11111101",
  8276=>"11111110",
  8277=>"00000001",
  8278=>"11111110",
  8279=>"00000000",
  8280=>"00000010",
  8281=>"11111111",
  8282=>"11111111",
  8283=>"11111101",
  8284=>"11111101",
  8285=>"00000001",
  8286=>"11111101",
  8287=>"11111111",
  8288=>"11111111",
  8289=>"00000000",
  8290=>"11111100",
  8291=>"11111110",
  8292=>"00000010",
  8293=>"00000001",
  8294=>"00000000",
  8295=>"00000010",
  8296=>"11111100",
  8297=>"00000011",
  8298=>"11111110",
  8299=>"11111111",
  8300=>"11111100",
  8301=>"00000010",
  8302=>"00000011",
  8303=>"11111111",
  8304=>"00000001",
  8305=>"11111111",
  8306=>"00000010",
  8307=>"00000000",
  8308=>"00000001",
  8309=>"00000011",
  8310=>"00000011",
  8311=>"00000011",
  8312=>"11111111",
  8313=>"00000000",
  8314=>"00000001",
  8315=>"11111111",
  8316=>"11111111",
  8317=>"00000010",
  8318=>"00000010",
  8319=>"00000011",
  8320=>"00000010",
  8321=>"00000001",
  8322=>"00000001",
  8323=>"00000001",
  8324=>"11111111",
  8325=>"11111110",
  8326=>"00000001",
  8327=>"11111111",
  8328=>"11111110",
  8329=>"00000001",
  8330=>"00000100",
  8331=>"11111110",
  8332=>"00000000",
  8333=>"00000001",
  8334=>"00000000",
  8335=>"11111110",
  8336=>"00000010",
  8337=>"11111111",
  8338=>"00000010",
  8339=>"00000010",
  8340=>"11111111",
  8341=>"11111101",
  8342=>"11111111",
  8343=>"11111111",
  8344=>"00000010",
  8345=>"11111111",
  8346=>"00000011",
  8347=>"00000010",
  8348=>"11111110",
  8349=>"00000001",
  8350=>"00000001",
  8351=>"00000010",
  8352=>"00000000",
  8353=>"11111111",
  8354=>"00000001",
  8355=>"00000001",
  8356=>"00000001",
  8357=>"11111111",
  8358=>"11111110",
  8359=>"00000001",
  8360=>"00000011",
  8361=>"11111101",
  8362=>"00000110",
  8363=>"00000001",
  8364=>"00000011",
  8365=>"00000000",
  8366=>"00000010",
  8367=>"00000001",
  8368=>"00000011",
  8369=>"00000000",
  8370=>"11111111",
  8371=>"11111110",
  8372=>"00000000",
  8373=>"00000111",
  8374=>"00000000",
  8375=>"00000000",
  8376=>"11111111",
  8377=>"00000000",
  8378=>"00000000",
  8379=>"11111110",
  8380=>"11111111",
  8381=>"00000010",
  8382=>"11111111",
  8383=>"00000010",
  8384=>"11111110",
  8385=>"00000010",
  8386=>"00000011",
  8387=>"00000010",
  8388=>"11111101",
  8389=>"11111110",
  8390=>"00000000",
  8391=>"11111101",
  8392=>"00000001",
  8393=>"00000010",
  8394=>"00000001",
  8395=>"11111101",
  8396=>"11111101",
  8397=>"00000001",
  8398=>"00000011",
  8399=>"11111110",
  8400=>"11111110",
  8401=>"00000010",
  8402=>"00000000",
  8403=>"11111101",
  8404=>"11111111",
  8405=>"11111101",
  8406=>"00000000",
  8407=>"00000011",
  8408=>"00000001",
  8409=>"00000000",
  8410=>"11111101",
  8411=>"11111101",
  8412=>"00000001",
  8413=>"11111110",
  8414=>"00000111",
  8415=>"00000010",
  8416=>"11111111",
  8417=>"00000001",
  8418=>"00000001",
  8419=>"11111111",
  8420=>"11111110",
  8421=>"11111111",
  8422=>"11111110",
  8423=>"00000000",
  8424=>"11111110",
  8425=>"11111101",
  8426=>"00000010",
  8427=>"00000000",
  8428=>"00000001",
  8429=>"00000010",
  8430=>"00000000",
  8431=>"11111110",
  8432=>"11111111",
  8433=>"11111101",
  8434=>"11111101",
  8435=>"00000000",
  8436=>"11111101",
  8437=>"00000000",
  8438=>"11111110",
  8439=>"00000010",
  8440=>"11111110",
  8441=>"11111111",
  8442=>"00000110",
  8443=>"11111110",
  8444=>"00000001",
  8445=>"00000001",
  8446=>"00000011",
  8447=>"11111101",
  8448=>"00000001",
  8449=>"00000010",
  8450=>"00000001",
  8451=>"00000001",
  8452=>"11111111",
  8453=>"00000001",
  8454=>"00000000",
  8455=>"11111111",
  8456=>"00000010",
  8457=>"00000001",
  8458=>"00000010",
  8459=>"00000000",
  8460=>"00000001",
  8461=>"11111110",
  8462=>"00000010",
  8463=>"00000111",
  8464=>"00000000",
  8465=>"00000001",
  8466=>"00000000",
  8467=>"00000000",
  8468=>"11111111",
  8469=>"00000010",
  8470=>"11111111",
  8471=>"00000001",
  8472=>"11111110",
  8473=>"11111111",
  8474=>"00000010",
  8475=>"00000010",
  8476=>"11111101",
  8477=>"00000001",
  8478=>"11111101",
  8479=>"00000011",
  8480=>"00000010",
  8481=>"11111111",
  8482=>"00000010",
  8483=>"00000000",
  8484=>"11111101",
  8485=>"11111111",
  8486=>"11111111",
  8487=>"11111101",
  8488=>"00000010",
  8489=>"11111101",
  8490=>"00000001",
  8491=>"00000000",
  8492=>"11111110",
  8493=>"00000000",
  8494=>"11111111",
  8495=>"00000001",
  8496=>"00000000",
  8497=>"11111110",
  8498=>"11111110",
  8499=>"00000011",
  8500=>"00000001",
  8501=>"00000000",
  8502=>"00000000",
  8503=>"11111110",
  8504=>"00000010",
  8505=>"11111110",
  8506=>"11111110",
  8507=>"11111101",
  8508=>"11111110",
  8509=>"11111110",
  8510=>"00000010",
  8511=>"00000001",
  8512=>"00000000",
  8513=>"00000100",
  8514=>"00000001",
  8515=>"00000010",
  8516=>"11111110",
  8517=>"00000010",
  8518=>"00000011",
  8519=>"11111101",
  8520=>"00000110",
  8521=>"00000000",
  8522=>"00000000",
  8523=>"11111111",
  8524=>"11111110",
  8525=>"00000011",
  8526=>"11111101",
  8527=>"00000000",
  8528=>"00000100",
  8529=>"11111110",
  8530=>"11111111",
  8531=>"00000101",
  8532=>"00000010",
  8533=>"00000010",
  8534=>"11111101",
  8535=>"00000011",
  8536=>"11111111",
  8537=>"00000000",
  8538=>"00000010",
  8539=>"00000010",
  8540=>"00000000",
  8541=>"00000010",
  8542=>"00000000",
  8543=>"00000000",
  8544=>"00000000",
  8545=>"11111100",
  8546=>"11111110",
  8547=>"00000001",
  8548=>"11111101",
  8549=>"11111110",
  8550=>"00000010",
  8551=>"00000010",
  8552=>"00000001",
  8553=>"00000000",
  8554=>"11111111",
  8555=>"11111011",
  8556=>"00000000",
  8557=>"11111110",
  8558=>"00000101",
  8559=>"00000000",
  8560=>"00000001",
  8561=>"00000001",
  8562=>"11111111",
  8563=>"00000000",
  8564=>"00000100",
  8565=>"11111110",
  8566=>"11111111",
  8567=>"11111111",
  8568=>"00000010",
  8569=>"11111111",
  8570=>"11111101",
  8571=>"11111111",
  8572=>"11111101",
  8573=>"00000010",
  8574=>"00000010",
  8575=>"00000001",
  8576=>"00000000",
  8577=>"00000000",
  8578=>"00000001",
  8579=>"00000001",
  8580=>"00000010",
  8581=>"00000000",
  8582=>"00000000",
  8583=>"11111111",
  8584=>"11111111",
  8585=>"00000011",
  8586=>"00000011",
  8587=>"00000001",
  8588=>"11111111",
  8589=>"11111110",
  8590=>"11111111",
  8591=>"00000010",
  8592=>"11111111",
  8593=>"00000010",
  8594=>"00000011",
  8595=>"11111110",
  8596=>"11111110",
  8597=>"11111101",
  8598=>"00000000",
  8599=>"11111111",
  8600=>"11111110",
  8601=>"00000010",
  8602=>"00000001",
  8603=>"00000000",
  8604=>"11111110",
  8605=>"00000001",
  8606=>"00000000",
  8607=>"00000100",
  8608=>"11111101",
  8609=>"11111111",
  8610=>"00000011",
  8611=>"00000001",
  8612=>"00000010",
  8613=>"11111110",
  8614=>"00000011",
  8615=>"11111100",
  8616=>"11111110",
  8617=>"00000000",
  8618=>"00000011",
  8619=>"00000000",
  8620=>"11111111",
  8621=>"11111101",
  8622=>"11111111",
  8623=>"00000000",
  8624=>"00000011",
  8625=>"11111101",
  8626=>"00000001",
  8627=>"11111111",
  8628=>"11111111",
  8629=>"00000000",
  8630=>"00000010",
  8631=>"00000001",
  8632=>"11111111",
  8633=>"11111110",
  8634=>"11111110",
  8635=>"11111111",
  8636=>"00000010",
  8637=>"00000001",
  8638=>"11111111",
  8639=>"00000100",
  8640=>"11111110",
  8641=>"11111101",
  8642=>"00000001",
  8643=>"11111100",
  8644=>"11111110",
  8645=>"11111101",
  8646=>"11111101",
  8647=>"11111111",
  8648=>"11111110",
  8649=>"00000101",
  8650=>"11111110",
  8651=>"00000010",
  8652=>"00000011",
  8653=>"00000001",
  8654=>"11111111",
  8655=>"00000001",
  8656=>"00000010",
  8657=>"11111111",
  8658=>"00000010",
  8659=>"11111101",
  8660=>"00000000",
  8661=>"11111111",
  8662=>"00000010",
  8663=>"00000000",
  8664=>"00000010",
  8665=>"11111101",
  8666=>"11111110",
  8667=>"00000000",
  8668=>"11111101",
  8669=>"11111111",
  8670=>"11111111",
  8671=>"11111110",
  8672=>"11111111",
  8673=>"11111101",
  8674=>"11111111",
  8675=>"00000011",
  8676=>"11111111",
  8677=>"11111111",
  8678=>"00000000",
  8679=>"00000001",
  8680=>"11111101",
  8681=>"00000001",
  8682=>"11111111",
  8683=>"11111101",
  8684=>"00000001",
  8685=>"00000000",
  8686=>"00000001",
  8687=>"00000010",
  8688=>"00000010",
  8689=>"00000010",
  8690=>"00000001",
  8691=>"00000000",
  8692=>"11111111",
  8693=>"00000001",
  8694=>"11111101",
  8695=>"11111110",
  8696=>"00000011",
  8697=>"00000001",
  8698=>"00000001",
  8699=>"00000001",
  8700=>"00000010",
  8701=>"11111110",
  8702=>"11111101",
  8703=>"00000000",
  8704=>"11111110",
  8705=>"11111111",
  8706=>"11111110",
  8707=>"00000000",
  8708=>"00000000",
  8709=>"00000000",
  8710=>"11111110",
  8711=>"00000101",
  8712=>"00000000",
  8713=>"00000011",
  8714=>"00000011",
  8715=>"11111110",
  8716=>"11111111",
  8717=>"00000011",
  8718=>"00000000",
  8719=>"00000001",
  8720=>"00000010",
  8721=>"11111111",
  8722=>"00000001",
  8723=>"11111101",
  8724=>"11111101",
  8725=>"00000011",
  8726=>"11111111",
  8727=>"00000001",
  8728=>"11111110",
  8729=>"00000100",
  8730=>"00000001",
  8731=>"11111101",
  8732=>"11111101",
  8733=>"00000010",
  8734=>"11111111",
  8735=>"11111101",
  8736=>"11111111",
  8737=>"00000001",
  8738=>"00000000",
  8739=>"11111101",
  8740=>"11111111",
  8741=>"00000010",
  8742=>"00000010",
  8743=>"11111110",
  8744=>"00000001",
  8745=>"00000010",
  8746=>"11111101",
  8747=>"11111100",
  8748=>"00000001",
  8749=>"11111100",
  8750=>"11111111",
  8751=>"11111111",
  8752=>"00000000",
  8753=>"11111101",
  8754=>"00000001",
  8755=>"00000001",
  8756=>"11111100",
  8757=>"00000100",
  8758=>"00000011",
  8759=>"11111111",
  8760=>"00000001",
  8761=>"00000000",
  8762=>"11111111",
  8763=>"00000010",
  8764=>"11111111",
  8765=>"00000001",
  8766=>"11111110",
  8767=>"00000001",
  8768=>"11111111",
  8769=>"00000011",
  8770=>"00000001",
  8771=>"00000010",
  8772=>"00000101",
  8773=>"00000001",
  8774=>"11111101",
  8775=>"00000000",
  8776=>"00000001",
  8777=>"11111111",
  8778=>"11111111",
  8779=>"11111111",
  8780=>"00000000",
  8781=>"00000001",
  8782=>"11111100",
  8783=>"11111111",
  8784=>"00000001",
  8785=>"00000010",
  8786=>"00000100",
  8787=>"00000001",
  8788=>"00000001",
  8789=>"00000000",
  8790=>"11111101",
  8791=>"00000000",
  8792=>"11111110",
  8793=>"00000000",
  8794=>"00000000",
  8795=>"00000101",
  8796=>"00000001",
  8797=>"00000001",
  8798=>"00000100",
  8799=>"00000011",
  8800=>"00000000",
  8801=>"00000000",
  8802=>"00000010",
  8803=>"11111111",
  8804=>"11111111",
  8805=>"11111100",
  8806=>"00000011",
  8807=>"11111100",
  8808=>"00000001",
  8809=>"11111111",
  8810=>"00000001",
  8811=>"00000100",
  8812=>"11111110",
  8813=>"00000101",
  8814=>"11111101",
  8815=>"11111100",
  8816=>"00000000",
  8817=>"11111101",
  8818=>"00000010",
  8819=>"11111110",
  8820=>"00000010",
  8821=>"11111101",
  8822=>"00000010",
  8823=>"00000001",
  8824=>"00000001",
  8825=>"00000000",
  8826=>"00000000",
  8827=>"11111101",
  8828=>"11111110",
  8829=>"11111110",
  8830=>"11111100",
  8831=>"00000010",
  8832=>"00000001",
  8833=>"11111101",
  8834=>"00000000",
  8835=>"11111100",
  8836=>"11111101",
  8837=>"11111111",
  8838=>"11111101",
  8839=>"00000000",
  8840=>"00000001",
  8841=>"00000010",
  8842=>"00000000",
  8843=>"11111100",
  8844=>"00000010",
  8845=>"00000000",
  8846=>"11111101",
  8847=>"11111111",
  8848=>"00000001",
  8849=>"00000111",
  8850=>"11111111",
  8851=>"00000001",
  8852=>"11111100",
  8853=>"11111110",
  8854=>"00000010",
  8855=>"00000001",
  8856=>"00000001",
  8857=>"11111110",
  8858=>"00000111",
  8859=>"00000010",
  8860=>"11111110",
  8861=>"00000010",
  8862=>"00000110",
  8863=>"11111101",
  8864=>"00000010",
  8865=>"11111110",
  8866=>"11111101",
  8867=>"11111100",
  8868=>"00000010",
  8869=>"11111110",
  8870=>"11111110",
  8871=>"11111110",
  8872=>"11111110",
  8873=>"00000010",
  8874=>"00000000",
  8875=>"00000011",
  8876=>"00000000",
  8877=>"00000000",
  8878=>"11111101",
  8879=>"11111111",
  8880=>"11111111",
  8881=>"00000001",
  8882=>"00000001",
  8883=>"00000000",
  8884=>"00000001",
  8885=>"11111110",
  8886=>"11111111",
  8887=>"00000001",
  8888=>"11111111",
  8889=>"00000000",
  8890=>"00000001",
  8891=>"00000010",
  8892=>"00000001",
  8893=>"00000000",
  8894=>"00000010",
  8895=>"11111111",
  8896=>"00000001",
  8897=>"11111101",
  8898=>"11111110",
  8899=>"11111111",
  8900=>"11111111",
  8901=>"00000011",
  8902=>"00000010",
  8903=>"00000001",
  8904=>"00000001",
  8905=>"11111110",
  8906=>"11111111",
  8907=>"00000000",
  8908=>"00000000",
  8909=>"00000011",
  8910=>"00000001",
  8911=>"00000000",
  8912=>"11111110",
  8913=>"11111111",
  8914=>"11111101",
  8915=>"00000101",
  8916=>"00000001",
  8917=>"11111111",
  8918=>"00000000",
  8919=>"11111101",
  8920=>"00000110",
  8921=>"11111111",
  8922=>"00000100",
  8923=>"11111110",
  8924=>"00000000",
  8925=>"00000010",
  8926=>"00000000",
  8927=>"11111111",
  8928=>"00000010",
  8929=>"00000001",
  8930=>"00000101",
  8931=>"11111110",
  8932=>"00000010",
  8933=>"00000001",
  8934=>"11111101",
  8935=>"11111111",
  8936=>"11111101",
  8937=>"11111111",
  8938=>"00000001",
  8939=>"00000011",
  8940=>"11111110",
  8941=>"00000000",
  8942=>"11111110",
  8943=>"11111111",
  8944=>"11111110",
  8945=>"11111111",
  8946=>"11111110",
  8947=>"00000010",
  8948=>"00000001",
  8949=>"00000001",
  8950=>"11111101",
  8951=>"00000010",
  8952=>"11111100",
  8953=>"11111100",
  8954=>"00000010",
  8955=>"00000001",
  8956=>"00000010",
  8957=>"11111111",
  8958=>"11111111",
  8959=>"00000011",
  8960=>"11111110",
  8961=>"11111111",
  8962=>"11111110",
  8963=>"00000010",
  8964=>"11111110",
  8965=>"11111110",
  8966=>"00000000",
  8967=>"11111110",
  8968=>"00000010",
  8969=>"11111111",
  8970=>"11111101",
  8971=>"00000010",
  8972=>"11111111",
  8973=>"11111111",
  8974=>"11111101",
  8975=>"11111111",
  8976=>"00000010",
  8977=>"11111110",
  8978=>"11111110",
  8979=>"00000010",
  8980=>"11111100",
  8981=>"11111110",
  8982=>"11111111",
  8983=>"11111110",
  8984=>"11111111",
  8985=>"11111110",
  8986=>"11111110",
  8987=>"11111100",
  8988=>"00000010",
  8989=>"11111110",
  8990=>"00000000",
  8991=>"00000001",
  8992=>"11111100",
  8993=>"11111110",
  8994=>"00000100",
  8995=>"11111111",
  8996=>"11111111",
  8997=>"11111111",
  8998=>"11111110",
  8999=>"11111110",
  9000=>"00000010",
  9001=>"00000000",
  9002=>"11111011",
  9003=>"11111101",
  9004=>"11111110",
  9005=>"11111101",
  9006=>"11111111",
  9007=>"00000100",
  9008=>"11111110",
  9009=>"11111111",
  9010=>"00000001",
  9011=>"11111111",
  9012=>"00000001",
  9013=>"11111100",
  9014=>"00000000",
  9015=>"00000000",
  9016=>"11111110",
  9017=>"00000001",
  9018=>"00000010",
  9019=>"00000010",
  9020=>"11111111",
  9021=>"00000010",
  9022=>"00000010",
  9023=>"11111111",
  9024=>"11111100",
  9025=>"00000000",
  9026=>"00000000",
  9027=>"11111111",
  9028=>"11111101",
  9029=>"11111110",
  9030=>"11111111",
  9031=>"00000010",
  9032=>"00000100",
  9033=>"00000000",
  9034=>"11111110",
  9035=>"00000011",
  9036=>"00000001",
  9037=>"11111111",
  9038=>"00000001",
  9039=>"00000100",
  9040=>"00000010",
  9041=>"00000000",
  9042=>"11111111",
  9043=>"11111111",
  9044=>"11111111",
  9045=>"00000001",
  9046=>"11111111",
  9047=>"00000001",
  9048=>"00000000",
  9049=>"11111111",
  9050=>"11111111",
  9051=>"00000011",
  9052=>"11111101",
  9053=>"11111111",
  9054=>"11111110",
  9055=>"11111101",
  9056=>"00000010",
  9057=>"00000110",
  9058=>"00000000",
  9059=>"00000010",
  9060=>"00000011",
  9061=>"11111110",
  9062=>"00000011",
  9063=>"00000000",
  9064=>"00000010",
  9065=>"00000100",
  9066=>"11111111",
  9067=>"00000000",
  9068=>"11111111",
  9069=>"11111101",
  9070=>"00000000",
  9071=>"11111110",
  9072=>"00000000",
  9073=>"00000010",
  9074=>"00000001",
  9075=>"11111110",
  9076=>"00000011",
  9077=>"11111101",
  9078=>"11111101",
  9079=>"00000001",
  9080=>"00000000",
  9081=>"00000001",
  9082=>"00000000",
  9083=>"00000001",
  9084=>"00000110",
  9085=>"00000001",
  9086=>"00001000",
  9087=>"00000001",
  9088=>"00000001",
  9089=>"00000100",
  9090=>"00000010",
  9091=>"00000000",
  9092=>"00000001",
  9093=>"00000010",
  9094=>"11111111",
  9095=>"00000001",
  9096=>"00000001",
  9097=>"00000001",
  9098=>"11111110",
  9099=>"11111111",
  9100=>"11111101",
  9101=>"00000011",
  9102=>"00000000",
  9103=>"00000100",
  9104=>"00000001",
  9105=>"11111110",
  9106=>"11111101",
  9107=>"00000000",
  9108=>"11111111",
  9109=>"11111110",
  9110=>"00000010",
  9111=>"00000010",
  9112=>"11111100",
  9113=>"11111111",
  9114=>"00000000",
  9115=>"00000010",
  9116=>"11111110",
  9117=>"00000000",
  9118=>"00000001",
  9119=>"11111100",
  9120=>"11111110",
  9121=>"00000010",
  9122=>"00000000",
  9123=>"11111111",
  9124=>"00000001",
  9125=>"00000010",
  9126=>"00000011",
  9127=>"11111111",
  9128=>"00000000",
  9129=>"11111101",
  9130=>"00000000",
  9131=>"00000001",
  9132=>"00000011",
  9133=>"11111101",
  9134=>"00000001",
  9135=>"11111111",
  9136=>"11111110",
  9137=>"11111100",
  9138=>"00000101",
  9139=>"00000010",
  9140=>"11111111",
  9141=>"00000101",
  9142=>"00000000",
  9143=>"11111110",
  9144=>"11111111",
  9145=>"11111111",
  9146=>"11111111",
  9147=>"00000001",
  9148=>"11111101",
  9149=>"11111101",
  9150=>"00000001",
  9151=>"11111111",
  9152=>"11111110",
  9153=>"11111111",
  9154=>"11111110",
  9155=>"00000000",
  9156=>"11111110",
  9157=>"11111110",
  9158=>"11111101",
  9159=>"00000010",
  9160=>"11111110",
  9161=>"00000001",
  9162=>"00000000",
  9163=>"11111101",
  9164=>"00000001",
  9165=>"00000000",
  9166=>"00000000",
  9167=>"11111110",
  9168=>"11111111",
  9169=>"11111111",
  9170=>"11111100",
  9171=>"00000001",
  9172=>"11111111",
  9173=>"00000000",
  9174=>"11111101",
  9175=>"00000001",
  9176=>"11111110",
  9177=>"11111111",
  9178=>"00000000",
  9179=>"11111101",
  9180=>"00000000",
  9181=>"11111101",
  9182=>"11111111",
  9183=>"00000010",
  9184=>"11111111",
  9185=>"00000001",
  9186=>"11111111",
  9187=>"00000010",
  9188=>"00000011",
  9189=>"11111111",
  9190=>"00000000",
  9191=>"11111110",
  9192=>"11111110",
  9193=>"11111110",
  9194=>"11111101",
  9195=>"11111101",
  9196=>"00000000",
  9197=>"00000010",
  9198=>"11111110",
  9199=>"00000100",
  9200=>"00000010",
  9201=>"11111110",
  9202=>"00000001",
  9203=>"11111110",
  9204=>"11111101",
  9205=>"00000101",
  9206=>"00000010",
  9207=>"11111101",
  9208=>"11111101",
  9209=>"11111111",
  9210=>"11111101",
  9211=>"00000010",
  9212=>"11111111",
  9213=>"00000000",
  9214=>"00000000",
  9215=>"00000011",
  9216=>"11111101",
  9217=>"00000101",
  9218=>"00000000",
  9219=>"00000010",
  9220=>"11111111",
  9221=>"00000000",
  9222=>"11111101",
  9223=>"00000000",
  9224=>"11111111",
  9225=>"11111100",
  9226=>"00000000",
  9227=>"11111110",
  9228=>"00000010",
  9229=>"00000011",
  9230=>"11111100",
  9231=>"00000000",
  9232=>"11111101",
  9233=>"00000001",
  9234=>"00000001",
  9235=>"11111110",
  9236=>"11111111",
  9237=>"00000001",
  9238=>"11111111",
  9239=>"00000011",
  9240=>"11111101",
  9241=>"00000010",
  9242=>"00000101",
  9243=>"00000001",
  9244=>"11111110",
  9245=>"00000001",
  9246=>"00000000",
  9247=>"00000000",
  9248=>"11111111",
  9249=>"11111101",
  9250=>"11111101",
  9251=>"00000011",
  9252=>"00000000",
  9253=>"11111101",
  9254=>"11111111",
  9255=>"00000011",
  9256=>"11111101",
  9257=>"00000011",
  9258=>"00000010",
  9259=>"00000011",
  9260=>"00000011",
  9261=>"11111101",
  9262=>"11111111",
  9263=>"11111101",
  9264=>"00000010",
  9265=>"11111111",
  9266=>"11111110",
  9267=>"11111110",
  9268=>"00000011",
  9269=>"00000001",
  9270=>"11111111",
  9271=>"11111100",
  9272=>"11111100",
  9273=>"11111110",
  9274=>"00000001",
  9275=>"11111101",
  9276=>"00000100",
  9277=>"11111110",
  9278=>"11111110",
  9279=>"00000000",
  9280=>"11111111",
  9281=>"00000000",
  9282=>"11111101",
  9283=>"00000010",
  9284=>"00000000",
  9285=>"00000010",
  9286=>"00000001",
  9287=>"00000001",
  9288=>"00000001",
  9289=>"00000000",
  9290=>"00000001",
  9291=>"00000000",
  9292=>"00000000",
  9293=>"11111110",
  9294=>"00000001",
  9295=>"11111111",
  9296=>"11111111",
  9297=>"00000011",
  9298=>"00000111",
  9299=>"11111110",
  9300=>"00000010",
  9301=>"11111111",
  9302=>"11111110",
  9303=>"00000011",
  9304=>"00000010",
  9305=>"11111011",
  9306=>"00000000",
  9307=>"00000000",
  9308=>"11111101",
  9309=>"11111111",
  9310=>"11111111",
  9311=>"00000100",
  9312=>"11111100",
  9313=>"11111111",
  9314=>"00000010",
  9315=>"00000001",
  9316=>"11111101",
  9317=>"11111101",
  9318=>"00000010",
  9319=>"00000000",
  9320=>"00000001",
  9321=>"11111111",
  9322=>"11111111",
  9323=>"11111110",
  9324=>"00000010",
  9325=>"00000001",
  9326=>"00000010",
  9327=>"00000001",
  9328=>"00000010",
  9329=>"00000000",
  9330=>"11111100",
  9331=>"11111111",
  9332=>"11111110",
  9333=>"00000001",
  9334=>"11111101",
  9335=>"00000001",
  9336=>"00000010",
  9337=>"11111110",
  9338=>"00000000",
  9339=>"00000000",
  9340=>"00000001",
  9341=>"00000000",
  9342=>"11111110",
  9343=>"00000010",
  9344=>"11111100",
  9345=>"00000010",
  9346=>"11111111",
  9347=>"11111101",
  9348=>"00000010",
  9349=>"11111110",
  9350=>"00000010",
  9351=>"00000001",
  9352=>"11111110",
  9353=>"11111101",
  9354=>"00000010",
  9355=>"11111111",
  9356=>"11111110",
  9357=>"00000001",
  9358=>"00000010",
  9359=>"00000011",
  9360=>"11111111",
  9361=>"11111111",
  9362=>"11111110",
  9363=>"11111110",
  9364=>"11111100",
  9365=>"11111111",
  9366=>"00000001",
  9367=>"00000000",
  9368=>"00000010",
  9369=>"00000010",
  9370=>"11111110",
  9371=>"00000010",
  9372=>"00000000",
  9373=>"11111111",
  9374=>"11111111",
  9375=>"11111111",
  9376=>"00000001",
  9377=>"00000010",
  9378=>"00000001",
  9379=>"11111110",
  9380=>"00000010",
  9381=>"00000001",
  9382=>"00000111",
  9383=>"11111111",
  9384=>"11111110",
  9385=>"11111111",
  9386=>"11111101",
  9387=>"11111100",
  9388=>"11111111",
  9389=>"00000001",
  9390=>"00000010",
  9391=>"00000010",
  9392=>"11111111",
  9393=>"11111101",
  9394=>"11111101",
  9395=>"00000001",
  9396=>"00000000",
  9397=>"11111110",
  9398=>"00000100",
  9399=>"11111110",
  9400=>"11111111",
  9401=>"11111101",
  9402=>"11111110",
  9403=>"11111111",
  9404=>"00000001",
  9405=>"11111111",
  9406=>"11111110",
  9407=>"00000011",
  9408=>"11111101",
  9409=>"00000010",
  9410=>"11111110",
  9411=>"11111111",
  9412=>"00000000",
  9413=>"00000011",
  9414=>"00000001",
  9415=>"00000100",
  9416=>"00000000",
  9417=>"11111111",
  9418=>"00000010",
  9419=>"00000001",
  9420=>"00000001",
  9421=>"00000001",
  9422=>"00000000",
  9423=>"00000110",
  9424=>"00000100",
  9425=>"00000000",
  9426=>"11111111",
  9427=>"00000000",
  9428=>"11111110",
  9429=>"11111110",
  9430=>"00000011",
  9431=>"11111111",
  9432=>"00000001",
  9433=>"00000011",
  9434=>"00000001",
  9435=>"11111101",
  9436=>"11111110",
  9437=>"00000110",
  9438=>"11111101",
  9439=>"00000101",
  9440=>"00000010",
  9441=>"11111110",
  9442=>"11111101",
  9443=>"11111111",
  9444=>"11111110",
  9445=>"00000011",
  9446=>"11111101",
  9447=>"00000001",
  9448=>"00000000",
  9449=>"00000100",
  9450=>"11111110",
  9451=>"11111111",
  9452=>"00000001",
  9453=>"00000010",
  9454=>"11111110",
  9455=>"00000000",
  9456=>"00000000",
  9457=>"00000000",
  9458=>"11111101",
  9459=>"00000001",
  9460=>"00000010",
  9461=>"11111111",
  9462=>"00000001",
  9463=>"11111110",
  9464=>"11111100",
  9465=>"00000010",
  9466=>"11111111",
  9467=>"11111111",
  9468=>"11111111",
  9469=>"00000001",
  9470=>"11111111",
  9471=>"11111111",
  9472=>"00000010",
  9473=>"11111101",
  9474=>"00000001",
  9475=>"00000011",
  9476=>"00000010",
  9477=>"00000100",
  9478=>"00000000",
  9479=>"00000000",
  9480=>"00000010",
  9481=>"00000010",
  9482=>"00000000",
  9483=>"00000001",
  9484=>"00000010",
  9485=>"00000011",
  9486=>"00000000",
  9487=>"11111110",
  9488=>"00000000",
  9489=>"00000010",
  9490=>"00000000",
  9491=>"11111110",
  9492=>"00000010",
  9493=>"11111111",
  9494=>"11111111",
  9495=>"00000001",
  9496=>"00000001",
  9497=>"00000100",
  9498=>"00000010",
  9499=>"11111110",
  9500=>"11111111",
  9501=>"11111110",
  9502=>"00000001",
  9503=>"11111110",
  9504=>"11111110",
  9505=>"11111111",
  9506=>"11111110",
  9507=>"11111101",
  9508=>"11111110",
  9509=>"00000000",
  9510=>"00000001",
  9511=>"11111111",
  9512=>"11111111",
  9513=>"11111111",
  9514=>"00000011",
  9515=>"11111101",
  9516=>"11111111",
  9517=>"11111110",
  9518=>"00000001",
  9519=>"00000001",
  9520=>"00000000",
  9521=>"00000100",
  9522=>"00000001",
  9523=>"11111101",
  9524=>"00000000",
  9525=>"00000000",
  9526=>"11111111",
  9527=>"11111100",
  9528=>"11111110",
  9529=>"11111111",
  9530=>"11111110",
  9531=>"00000100",
  9532=>"00000010",
  9533=>"00000001",
  9534=>"00000010",
  9535=>"11111110",
  9536=>"11111101",
  9537=>"11111101",
  9538=>"11111110",
  9539=>"11111111",
  9540=>"00000010",
  9541=>"00000001",
  9542=>"00000001",
  9543=>"11111110",
  9544=>"11111111",
  9545=>"11111101",
  9546=>"00000011",
  9547=>"00000000",
  9548=>"11111101",
  9549=>"00000011",
  9550=>"11111111",
  9551=>"00000011",
  9552=>"00000001",
  9553=>"11111101",
  9554=>"00000001",
  9555=>"11111110",
  9556=>"11111111",
  9557=>"11111111",
  9558=>"11111101",
  9559=>"11111110",
  9560=>"11111101",
  9561=>"00000000",
  9562=>"11111111",
  9563=>"00000100",
  9564=>"11111101",
  9565=>"11111101",
  9566=>"00000011",
  9567=>"11111110",
  9568=>"11111101",
  9569=>"11111101",
  9570=>"00000000",
  9571=>"11111100",
  9572=>"11111101",
  9573=>"00000010",
  9574=>"00000000",
  9575=>"00000000",
  9576=>"00000000",
  9577=>"00000011",
  9578=>"11111110",
  9579=>"00000001",
  9580=>"00000000",
  9581=>"11111111",
  9582=>"00000001",
  9583=>"00000001",
  9584=>"00000000",
  9585=>"11111110",
  9586=>"00000001",
  9587=>"00000100",
  9588=>"00000010",
  9589=>"00000010",
  9590=>"11111111",
  9591=>"00000010",
  9592=>"11111110",
  9593=>"11111111",
  9594=>"11111111",
  9595=>"11111111",
  9596=>"11111111",
  9597=>"00000000",
  9598=>"00000001",
  9599=>"00000011",
  9600=>"11111111",
  9601=>"00000000",
  9602=>"00000001",
  9603=>"00000000",
  9604=>"11111101",
  9605=>"11111110",
  9606=>"00000011",
  9607=>"00000000",
  9608=>"11111101",
  9609=>"11111101",
  9610=>"00000001",
  9611=>"00000001",
  9612=>"11111111",
  9613=>"11111110",
  9614=>"11111110",
  9615=>"00000101",
  9616=>"11111111",
  9617=>"11111101",
  9618=>"00000001",
  9619=>"11111110",
  9620=>"00000101",
  9621=>"00000000",
  9622=>"00000010",
  9623=>"11111111",
  9624=>"00000001",
  9625=>"00000001",
  9626=>"00000010",
  9627=>"11111111",
  9628=>"00000010",
  9629=>"11111110",
  9630=>"11111101",
  9631=>"11111110",
  9632=>"00000010",
  9633=>"11111101",
  9634=>"00000010",
  9635=>"00000010",
  9636=>"11111110",
  9637=>"00000010",
  9638=>"11111101",
  9639=>"00000000",
  9640=>"00000010",
  9641=>"00000001",
  9642=>"11111110",
  9643=>"11111111",
  9644=>"00000010",
  9645=>"00000000",
  9646=>"11111101",
  9647=>"11111111",
  9648=>"00000010",
  9649=>"00000011",
  9650=>"11111111",
  9651=>"11111111",
  9652=>"00000000",
  9653=>"11111101",
  9654=>"00000001",
  9655=>"00000010",
  9656=>"00000010",
  9657=>"00000001",
  9658=>"00000010",
  9659=>"00000001",
  9660=>"11111111",
  9661=>"11111110",
  9662=>"11111100",
  9663=>"11111110",
  9664=>"11111100",
  9665=>"00000110",
  9666=>"00000100",
  9667=>"11111111",
  9668=>"00000000",
  9669=>"11111110",
  9670=>"00000011",
  9671=>"11111110",
  9672=>"00000001",
  9673=>"11111101",
  9674=>"00000010",
  9675=>"00000010",
  9676=>"00000011",
  9677=>"00000010",
  9678=>"00000010",
  9679=>"00000000",
  9680=>"00000010",
  9681=>"11111110",
  9682=>"00000010",
  9683=>"00000001",
  9684=>"00000000",
  9685=>"00000010",
  9686=>"00000000",
  9687=>"11111111",
  9688=>"00000000",
  9689=>"00000000",
  9690=>"00000001",
  9691=>"00000000",
  9692=>"00000100",
  9693=>"00000011",
  9694=>"00000010",
  9695=>"00000001",
  9696=>"00000011",
  9697=>"00000001",
  9698=>"11111111",
  9699=>"00000000",
  9700=>"00000001",
  9701=>"11111101",
  9702=>"00000010",
  9703=>"00000001",
  9704=>"11111111",
  9705=>"00000001",
  9706=>"11111110",
  9707=>"11111101",
  9708=>"00000000",
  9709=>"11111101",
  9710=>"00000000",
  9711=>"11111111",
  9712=>"00000001",
  9713=>"00000001",
  9714=>"11111110",
  9715=>"11111110",
  9716=>"00000000",
  9717=>"00000010",
  9718=>"00000000",
  9719=>"00000011",
  9720=>"11111111",
  9721=>"11111111",
  9722=>"00000000",
  9723=>"00000001",
  9724=>"11111111",
  9725=>"00000001",
  9726=>"00000000",
  9727=>"11111110",
  9728=>"11111110",
  9729=>"00000110",
  9730=>"00000000",
  9731=>"00000001",
  9732=>"11111101",
  9733=>"11111111",
  9734=>"00000010",
  9735=>"00000000",
  9736=>"00000010",
  9737=>"00000100",
  9738=>"00000001",
  9739=>"11111110",
  9740=>"11111110",
  9741=>"00000000",
  9742=>"00000000",
  9743=>"00000100",
  9744=>"11111101",
  9745=>"00000000",
  9746=>"00000011",
  9747=>"11111111",
  9748=>"00000000",
  9749=>"11111110",
  9750=>"11111110",
  9751=>"00000001",
  9752=>"00000000",
  9753=>"00000010",
  9754=>"00000000",
  9755=>"00000001",
  9756=>"00000000",
  9757=>"11111110",
  9758=>"00000010",
  9759=>"00000010",
  9760=>"11111110",
  9761=>"11111111",
  9762=>"11111110",
  9763=>"11111110",
  9764=>"00000001",
  9765=>"11111101",
  9766=>"00000010",
  9767=>"11111111",
  9768=>"00000100",
  9769=>"00000000",
  9770=>"00000010",
  9771=>"11111101",
  9772=>"11111101",
  9773=>"11111110",
  9774=>"11111101",
  9775=>"11111101",
  9776=>"00000100",
  9777=>"00000001",
  9778=>"00000001",
  9779=>"11111101",
  9780=>"11111110",
  9781=>"00000111",
  9782=>"11111101",
  9783=>"00000010",
  9784=>"00000010",
  9785=>"00000000",
  9786=>"00000010",
  9787=>"11111110",
  9788=>"00000001",
  9789=>"00000001",
  9790=>"00000011",
  9791=>"11111100",
  9792=>"11111100",
  9793=>"11111110",
  9794=>"11111101",
  9795=>"00000010",
  9796=>"11111111",
  9797=>"11111101",
  9798=>"11111110",
  9799=>"11111110",
  9800=>"00000001",
  9801=>"00000001",
  9802=>"00000010",
  9803=>"00000011",
  9804=>"11111110",
  9805=>"00000001",
  9806=>"11111100",
  9807=>"00000011",
  9808=>"11111111",
  9809=>"00000001",
  9810=>"11111110",
  9811=>"00000001",
  9812=>"00000000",
  9813=>"11111110",
  9814=>"00000001",
  9815=>"11111111",
  9816=>"00000011",
  9817=>"11111110",
  9818=>"00000011",
  9819=>"00000001",
  9820=>"00000111",
  9821=>"00000001",
  9822=>"00000011",
  9823=>"11111110",
  9824=>"11111101",
  9825=>"11111110",
  9826=>"00000011",
  9827=>"11111110",
  9828=>"11111110",
  9829=>"00000001",
  9830=>"00000001",
  9831=>"11111110",
  9832=>"00000010",
  9833=>"11111110",
  9834=>"00000010",
  9835=>"00000011",
  9836=>"00000000",
  9837=>"00000010",
  9838=>"00000000",
  9839=>"11111111",
  9840=>"11111111",
  9841=>"00000000",
  9842=>"00000011",
  9843=>"00000000",
  9844=>"00000010",
  9845=>"00000000",
  9846=>"00000001",
  9847=>"00000011",
  9848=>"00000101",
  9849=>"00000000",
  9850=>"11111111",
  9851=>"00000010",
  9852=>"11111111",
  9853=>"11111111",
  9854=>"00000110",
  9855=>"00000000",
  9856=>"11111111",
  9857=>"00000001",
  9858=>"00000110",
  9859=>"00000101",
  9860=>"11111110",
  9861=>"00000001",
  9862=>"00000001",
  9863=>"11111110",
  9864=>"00000011",
  9865=>"00000110",
  9866=>"00000100",
  9867=>"00000000",
  9868=>"00000000",
  9869=>"00000000",
  9870=>"00000001",
  9871=>"11111101",
  9872=>"00000000",
  9873=>"00000001",
  9874=>"11111101",
  9875=>"11111111",
  9876=>"11111111",
  9877=>"00000100",
  9878=>"11111110",
  9879=>"11111101",
  9880=>"11111111",
  9881=>"00000010",
  9882=>"11111110",
  9883=>"00000011",
  9884=>"11111101",
  9885=>"11111111",
  9886=>"11111111",
  9887=>"00000001",
  9888=>"00000010",
  9889=>"11111110",
  9890=>"11111110",
  9891=>"00000000",
  9892=>"11111101",
  9893=>"11111110",
  9894=>"00000000",
  9895=>"11111101",
  9896=>"00000000",
  9897=>"11111111",
  9898=>"00000011",
  9899=>"00000000",
  9900=>"11111110",
  9901=>"00000000",
  9902=>"00000000",
  9903=>"00000000",
  9904=>"00000100",
  9905=>"00000010",
  9906=>"00000001",
  9907=>"00000000",
  9908=>"00000001",
  9909=>"00000100",
  9910=>"00000010",
  9911=>"00000001",
  9912=>"11111111",
  9913=>"11111110",
  9914=>"11111111",
  9915=>"00000000",
  9916=>"00000000",
  9917=>"00000011",
  9918=>"11111101",
  9919=>"11111111",
  9920=>"11111111",
  9921=>"00000010",
  9922=>"00000010",
  9923=>"11111111",
  9924=>"00000001",
  9925=>"11111111",
  9926=>"00000001",
  9927=>"00000000",
  9928=>"11111110",
  9929=>"11111111",
  9930=>"00000011",
  9931=>"11111110",
  9932=>"00000010",
  9933=>"11111110",
  9934=>"00000000",
  9935=>"11111100",
  9936=>"11111111",
  9937=>"11111110",
  9938=>"00000100",
  9939=>"00000111",
  9940=>"11111110",
  9941=>"00000000",
  9942=>"11111111",
  9943=>"11111111",
  9944=>"11111101",
  9945=>"00000001",
  9946=>"11111110",
  9947=>"00000000",
  9948=>"00000001",
  9949=>"00000000",
  9950=>"00000011",
  9951=>"00000101",
  9952=>"11111110",
  9953=>"00000000",
  9954=>"11111110",
  9955=>"11111110",
  9956=>"11111111",
  9957=>"00000001",
  9958=>"00000001",
  9959=>"11111110",
  9960=>"00000000",
  9961=>"00000010",
  9962=>"00000001",
  9963=>"11111110",
  9964=>"11111110",
  9965=>"11111110",
  9966=>"11111110",
  9967=>"11111111",
  9968=>"00000000",
  9969=>"11111110",
  9970=>"11111111",
  9971=>"00000001",
  9972=>"00000110",
  9973=>"00000100",
  9974=>"11111110",
  9975=>"00000011",
  9976=>"00000010",
  9977=>"11111110",
  9978=>"00000000",
  9979=>"00000101",
  9980=>"00000010",
  9981=>"11111110",
  9982=>"00000100",
  9983=>"11111110",
  9984=>"11111100",
  9985=>"11111110",
  9986=>"11111110",
  9987=>"11111101",
  9988=>"11111110",
  9989=>"11111101",
  9990=>"11111110",
  9991=>"00000001",
  9992=>"00000111",
  9993=>"00000100",
  9994=>"00000010",
  9995=>"00000011",
  9996=>"00000010",
  9997=>"00000010",
  9998=>"11111110",
  9999=>"00000000",
  10000=>"00000010",
  10001=>"00000000",
  10002=>"11111101",
  10003=>"00000011",
  10004=>"11111111",
  10005=>"11111110",
  10006=>"00000011",
  10007=>"00000001",
  10008=>"00000001",
  10009=>"00000000",
  10010=>"00000101",
  10011=>"00000001",
  10012=>"00000000",
  10013=>"00000001",
  10014=>"00001000",
  10015=>"00000001",
  10016=>"11111100",
  10017=>"11111110",
  10018=>"00000010",
  10019=>"11111111",
  10020=>"11111111",
  10021=>"11111101",
  10022=>"00000001",
  10023=>"11111111",
  10024=>"11111100",
  10025=>"11111111",
  10026=>"11111100",
  10027=>"00000010",
  10028=>"11111111",
  10029=>"11111111",
  10030=>"00000000",
  10031=>"11111111",
  10032=>"11111110",
  10033=>"00000000",
  10034=>"11111110",
  10035=>"00000001",
  10036=>"00000001",
  10037=>"11111101",
  10038=>"00000000",
  10039=>"00000000",
  10040=>"11111111",
  10041=>"11111111",
  10042=>"11111110",
  10043=>"11111101",
  10044=>"11111101",
  10045=>"00000010",
  10046=>"00000010",
  10047=>"11111110",
  10048=>"11111101",
  10049=>"00000010",
  10050=>"11111111",
  10051=>"11111111",
  10052=>"11111110",
  10053=>"11111101",
  10054=>"00000011",
  10055=>"11111101",
  10056=>"00000100",
  10057=>"00000001",
  10058=>"11111101",
  10059=>"11111101",
  10060=>"11111110",
  10061=>"00000001",
  10062=>"11111111",
  10063=>"11111110",
  10064=>"11111110",
  10065=>"00000001",
  10066=>"00000000",
  10067=>"00000000",
  10068=>"00000100",
  10069=>"11111110",
  10070=>"00000000",
  10071=>"00000001",
  10072=>"11111111",
  10073=>"11111110",
  10074=>"00000000",
  10075=>"11111111",
  10076=>"11111110",
  10077=>"00000100",
  10078=>"00000001",
  10079=>"11111110",
  10080=>"00000010",
  10081=>"11111111",
  10082=>"00000011",
  10083=>"00000000",
  10084=>"00000001",
  10085=>"00000001",
  10086=>"00000010",
  10087=>"11111110",
  10088=>"11111111",
  10089=>"00000000",
  10090=>"11111111",
  10091=>"11111111",
  10092=>"11111111",
  10093=>"00000011",
  10094=>"11111111",
  10095=>"11111110",
  10096=>"00000011",
  10097=>"11111111",
  10098=>"11111110",
  10099=>"00000001",
  10100=>"00000000",
  10101=>"11111110",
  10102=>"11111100",
  10103=>"11111101",
  10104=>"00000010",
  10105=>"00000000",
  10106=>"00000001",
  10107=>"00000010",
  10108=>"11111110",
  10109=>"00000001",
  10110=>"11111101",
  10111=>"00000001",
  10112=>"11111101",
  10113=>"00000001",
  10114=>"00000001",
  10115=>"11111111",
  10116=>"00000001",
  10117=>"11111110",
  10118=>"00000001",
  10119=>"11111100",
  10120=>"00000110",
  10121=>"11111110",
  10122=>"11111111",
  10123=>"11111110",
  10124=>"11111101",
  10125=>"00000010",
  10126=>"00000000",
  10127=>"00000010",
  10128=>"00000010",
  10129=>"00000011",
  10130=>"00000001",
  10131=>"11111111",
  10132=>"00000100",
  10133=>"00000100",
  10134=>"00000000",
  10135=>"00000000",
  10136=>"11111101",
  10137=>"11111110",
  10138=>"00000000",
  10139=>"00000000",
  10140=>"11111101",
  10141=>"00000010",
  10142=>"11111110",
  10143=>"11111101",
  10144=>"00000011",
  10145=>"00000010",
  10146=>"00000101",
  10147=>"00000001",
  10148=>"00000010",
  10149=>"11111111",
  10150=>"00000010",
  10151=>"00000011",
  10152=>"00000001",
  10153=>"00000011",
  10154=>"00000100",
  10155=>"00000011",
  10156=>"00000010",
  10157=>"11111111",
  10158=>"00000001",
  10159=>"00000011",
  10160=>"11111101",
  10161=>"11111111",
  10162=>"11111110",
  10163=>"11111110",
  10164=>"00000001",
  10165=>"00000100",
  10166=>"00000000",
  10167=>"11111100",
  10168=>"00000011",
  10169=>"11111101",
  10170=>"11111111",
  10171=>"11111101",
  10172=>"00000001",
  10173=>"00000010",
  10174=>"11111110",
  10175=>"11111111",
  10176=>"00000011",
  10177=>"00000001",
  10178=>"11111101",
  10179=>"00000000",
  10180=>"11111110",
  10181=>"00000001",
  10182=>"00000000",
  10183=>"11111101",
  10184=>"00000010",
  10185=>"11111111",
  10186=>"00000100",
  10187=>"00000000",
  10188=>"00000001",
  10189=>"00000001",
  10190=>"11111110",
  10191=>"00000011",
  10192=>"11111110",
  10193=>"11111111",
  10194=>"00000100",
  10195=>"00000011",
  10196=>"00000010",
  10197=>"00000010",
  10198=>"00000001",
  10199=>"00000010",
  10200=>"00000001",
  10201=>"11111110",
  10202=>"11111101",
  10203=>"00000000",
  10204=>"00000000",
  10205=>"11111111",
  10206=>"00000011",
  10207=>"00000010",
  10208=>"00000001",
  10209=>"00000010",
  10210=>"11111111",
  10211=>"11111110",
  10212=>"00000001",
  10213=>"00000010",
  10214=>"11111101",
  10215=>"11111111",
  10216=>"00000010",
  10217=>"11111111",
  10218=>"00000100",
  10219=>"00000010",
  10220=>"00000010",
  10221=>"11111101",
  10222=>"00000001",
  10223=>"00000001",
  10224=>"00000000",
  10225=>"11111111",
  10226=>"00000001",
  10227=>"11111111",
  10228=>"11111100",
  10229=>"00000100",
  10230=>"11111111",
  10231=>"00000010",
  10232=>"11111111",
  10233=>"00000001",
  10234=>"11111101",
  10235=>"11111111",
  10236=>"00000001",
  10237=>"11111100",
  10238=>"11111111",
  10239=>"00000001",
  10240=>"11111101",
  10241=>"00000010",
  10242=>"00000000",
  10243=>"00000011",
  10244=>"00000000",
  10245=>"00000011",
  10246=>"11111110",
  10247=>"00000001",
  10248=>"00000010",
  10249=>"11111101",
  10250=>"11111110",
  10251=>"00000011",
  10252=>"11111101",
  10253=>"11111111",
  10254=>"00000101",
  10255=>"11111111",
  10256=>"00000001",
  10257=>"00000000",
  10258=>"11111101",
  10259=>"00000101",
  10260=>"11111111",
  10261=>"00000000",
  10262=>"00000000",
  10263=>"00000000",
  10264=>"00000110",
  10265=>"00000010",
  10266=>"11111110",
  10267=>"11111111",
  10268=>"11111101",
  10269=>"00000000",
  10270=>"00000010",
  10271=>"11111101",
  10272=>"00000100",
  10273=>"00000001",
  10274=>"00000010",
  10275=>"11111110",
  10276=>"00000000",
  10277=>"11111101",
  10278=>"00000001",
  10279=>"00000000",
  10280=>"11111101",
  10281=>"00000000",
  10282=>"00000000",
  10283=>"11111110",
  10284=>"11111110",
  10285=>"11111110",
  10286=>"00000001",
  10287=>"11111110",
  10288=>"00000001",
  10289=>"00000001",
  10290=>"00000111",
  10291=>"11111101",
  10292=>"11111111",
  10293=>"00000000",
  10294=>"00000001",
  10295=>"11111110",
  10296=>"00000001",
  10297=>"00000000",
  10298=>"00000000",
  10299=>"00000000",
  10300=>"11111111",
  10301=>"00000000",
  10302=>"00000001",
  10303=>"11111101",
  10304=>"11111110",
  10305=>"00000000",
  10306=>"11111110",
  10307=>"00000000",
  10308=>"00000001",
  10309=>"00000010",
  10310=>"00000010",
  10311=>"00000100",
  10312=>"00000100",
  10313=>"11111110",
  10314=>"00000011",
  10315=>"11111101",
  10316=>"11111111",
  10317=>"00000010",
  10318=>"11111110",
  10319=>"11111110",
  10320=>"00000000",
  10321=>"11111101",
  10322=>"11111110",
  10323=>"00000010",
  10324=>"00000010",
  10325=>"00000011",
  10326=>"11111111",
  10327=>"11111110",
  10328=>"00000001",
  10329=>"11111110",
  10330=>"00000100",
  10331=>"11111101",
  10332=>"11111111",
  10333=>"00000000",
  10334=>"11111101",
  10335=>"00000000",
  10336=>"11111110",
  10337=>"11111101",
  10338=>"11111101",
  10339=>"00000100",
  10340=>"11111110",
  10341=>"11111101",
  10342=>"00000010",
  10343=>"11111101",
  10344=>"00000000",
  10345=>"00000001",
  10346=>"11111101",
  10347=>"00000001",
  10348=>"11111111",
  10349=>"11111111",
  10350=>"00000010",
  10351=>"00000000",
  10352=>"11111110",
  10353=>"11111101",
  10354=>"11111110",
  10355=>"00000101",
  10356=>"11111110",
  10357=>"00000001",
  10358=>"11111111",
  10359=>"00000001",
  10360=>"00000001",
  10361=>"11111101",
  10362=>"00000101",
  10363=>"11111111",
  10364=>"00000001",
  10365=>"00000010",
  10366=>"11111101",
  10367=>"00000011",
  10368=>"11111101",
  10369=>"11111111",
  10370=>"00000110",
  10371=>"00000000",
  10372=>"00000010",
  10373=>"11111111",
  10374=>"00000001",
  10375=>"00000011",
  10376=>"11111111",
  10377=>"00000001",
  10378=>"00000011",
  10379=>"11111111",
  10380=>"00000110",
  10381=>"00000001",
  10382=>"00000011",
  10383=>"00000000",
  10384=>"11111101",
  10385=>"11111101",
  10386=>"11111110",
  10387=>"11111110",
  10388=>"00000010",
  10389=>"00000001",
  10390=>"00000001",
  10391=>"00000000",
  10392=>"00000001",
  10393=>"00000000",
  10394=>"11111110",
  10395=>"00000000",
  10396=>"00000000",
  10397=>"11111110",
  10398=>"11111110",
  10399=>"00000011",
  10400=>"00000000",
  10401=>"11111100",
  10402=>"11111101",
  10403=>"11111101",
  10404=>"00000001",
  10405=>"00000001",
  10406=>"11111101",
  10407=>"00000001",
  10408=>"00000000",
  10409=>"00000001",
  10410=>"11111110",
  10411=>"00000011",
  10412=>"00000010",
  10413=>"00000100",
  10414=>"00000100",
  10415=>"00000001",
  10416=>"11111101",
  10417=>"11111100",
  10418=>"00000010",
  10419=>"00000010",
  10420=>"00000011",
  10421=>"00000001",
  10422=>"00000010",
  10423=>"00001000",
  10424=>"11111101",
  10425=>"00000001",
  10426=>"11111101",
  10427=>"00000010",
  10428=>"11111101",
  10429=>"11111111",
  10430=>"00000000",
  10431=>"00000011",
  10432=>"11111110",
  10433=>"00000001",
  10434=>"00000001",
  10435=>"00000100",
  10436=>"11111111",
  10437=>"00000011",
  10438=>"00000010",
  10439=>"11111110",
  10440=>"00000010",
  10441=>"11111110",
  10442=>"00000001",
  10443=>"00000000",
  10444=>"11111110",
  10445=>"00000001",
  10446=>"11111111",
  10447=>"00000000",
  10448=>"00000010",
  10449=>"11111110",
  10450=>"00000000",
  10451=>"11111110",
  10452=>"00000001",
  10453=>"11111110",
  10454=>"11111101",
  10455=>"00000100",
  10456=>"00000001",
  10457=>"11111111",
  10458=>"00000001",
  10459=>"00000110",
  10460=>"00000000",
  10461=>"11111110",
  10462=>"00000001",
  10463=>"00000000",
  10464=>"00000110",
  10465=>"00000001",
  10466=>"00000010",
  10467=>"00000000",
  10468=>"00000010",
  10469=>"11111101",
  10470=>"00000100",
  10471=>"00000000",
  10472=>"00000000",
  10473=>"00000000",
  10474=>"00000011",
  10475=>"11111111",
  10476=>"11111111",
  10477=>"11111111",
  10478=>"00000010",
  10479=>"11111110",
  10480=>"11111110",
  10481=>"11111111",
  10482=>"11111110",
  10483=>"11111101",
  10484=>"11111111",
  10485=>"00000000",
  10486=>"11111101",
  10487=>"11111110",
  10488=>"00000010",
  10489=>"00000001",
  10490=>"11111111",
  10491=>"00000000",
  10492=>"00000110",
  10493=>"00000001",
  10494=>"11111111",
  10495=>"00000011",
  10496=>"11111111",
  10497=>"11111101",
  10498=>"00000010",
  10499=>"00000011",
  10500=>"11111110",
  10501=>"00000000",
  10502=>"11111111",
  10503=>"00000010",
  10504=>"00000010",
  10505=>"11111101",
  10506=>"11111111",
  10507=>"11111110",
  10508=>"11111110",
  10509=>"11111110",
  10510=>"11111111",
  10511=>"00000010",
  10512=>"00000000",
  10513=>"00000001",
  10514=>"00000001",
  10515=>"00000100",
  10516=>"11111101",
  10517=>"00000000",
  10518=>"11111101",
  10519=>"11111110",
  10520=>"11111111",
  10521=>"11111101",
  10522=>"00000001",
  10523=>"11111111",
  10524=>"00000110",
  10525=>"11111101",
  10526=>"11111110",
  10527=>"11111110",
  10528=>"11111110",
  10529=>"00000000",
  10530=>"11111110",
  10531=>"11111111",
  10532=>"00000010",
  10533=>"11111111",
  10534=>"11111110",
  10535=>"00000010",
  10536=>"00000011",
  10537=>"00000000",
  10538=>"00000001",
  10539=>"00000001",
  10540=>"00000000",
  10541=>"11111110",
  10542=>"11111101",
  10543=>"11111111",
  10544=>"00000000",
  10545=>"00000000",
  10546=>"11111100",
  10547=>"00000001",
  10548=>"11111110",
  10549=>"11111110",
  10550=>"00000010",
  10551=>"11111111",
  10552=>"00000000",
  10553=>"11111111",
  10554=>"00000001",
  10555=>"11111111",
  10556=>"00000000",
  10557=>"00000011",
  10558=>"00000001",
  10559=>"00000001",
  10560=>"00000000",
  10561=>"00000000",
  10562=>"11111101",
  10563=>"00000000",
  10564=>"11111101",
  10565=>"11111111",
  10566=>"11111100",
  10567=>"11111110",
  10568=>"00000011",
  10569=>"11111101",
  10570=>"00000101",
  10571=>"00000000",
  10572=>"11111101",
  10573=>"11111110",
  10574=>"00000001",
  10575=>"00000001",
  10576=>"00000010",
  10577=>"00000010",
  10578=>"00000000",
  10579=>"00000001",
  10580=>"11111100",
  10581=>"00000000",
  10582=>"11111111",
  10583=>"11111101",
  10584=>"11111110",
  10585=>"11111110",
  10586=>"00000000",
  10587=>"00000001",
  10588=>"11111101",
  10589=>"11111110",
  10590=>"11111111",
  10591=>"00000001",
  10592=>"00000000",
  10593=>"11111111",
  10594=>"00000110",
  10595=>"00000011",
  10596=>"00000010",
  10597=>"11111110",
  10598=>"11111101",
  10599=>"00000001",
  10600=>"11111101",
  10601=>"11111101",
  10602=>"11111111",
  10603=>"11111101",
  10604=>"11111101",
  10605=>"11111111",
  10606=>"00000010",
  10607=>"00000011",
  10608=>"11111111",
  10609=>"00000000",
  10610=>"00000010",
  10611=>"11111101",
  10612=>"11111101",
  10613=>"11111101",
  10614=>"11111111",
  10615=>"11111111",
  10616=>"00000010",
  10617=>"00000011",
  10618=>"11111100",
  10619=>"00000000",
  10620=>"00000010",
  10621=>"00000000",
  10622=>"00000010",
  10623=>"00000000",
  10624=>"11111110",
  10625=>"00000101",
  10626=>"11111111",
  10627=>"11111101",
  10628=>"00000100",
  10629=>"00000000",
  10630=>"00000010",
  10631=>"00000010",
  10632=>"00000000",
  10633=>"11111101",
  10634=>"11111101",
  10635=>"00000010",
  10636=>"00000000",
  10637=>"00000011",
  10638=>"00000000",
  10639=>"00000000",
  10640=>"00000000",
  10641=>"00000000",
  10642=>"00000010",
  10643=>"00000011",
  10644=>"00000010",
  10645=>"11111110",
  10646=>"00000010",
  10647=>"11111110",
  10648=>"11111110",
  10649=>"00000100",
  10650=>"11111111",
  10651=>"11111110",
  10652=>"00000001",
  10653=>"11111111",
  10654=>"00000001",
  10655=>"00000010",
  10656=>"11111110",
  10657=>"00000000",
  10658=>"00000001",
  10659=>"11111100",
  10660=>"00000010",
  10661=>"00000000",
  10662=>"00000010",
  10663=>"00000000",
  10664=>"00000011",
  10665=>"00000010",
  10666=>"11111101",
  10667=>"11111101",
  10668=>"00000011",
  10669=>"00000100",
  10670=>"00000100",
  10671=>"11111111",
  10672=>"11111111",
  10673=>"00000011",
  10674=>"11111110",
  10675=>"11111111",
  10676=>"00000001",
  10677=>"00000010",
  10678=>"11111111",
  10679=>"11111101",
  10680=>"00000011",
  10681=>"11111101",
  10682=>"11111111",
  10683=>"00000000",
  10684=>"00000000",
  10685=>"11111101",
  10686=>"00000000",
  10687=>"00000001",
  10688=>"11111111",
  10689=>"11111100",
  10690=>"00000001",
  10691=>"11111100",
  10692=>"11111111",
  10693=>"00000001",
  10694=>"11111111",
  10695=>"11111110",
  10696=>"00000001",
  10697=>"00000000",
  10698=>"11111111",
  10699=>"00000001",
  10700=>"00000000",
  10701=>"11111110",
  10702=>"11111101",
  10703=>"00000001",
  10704=>"00000010",
  10705=>"11111110",
  10706=>"11111111",
  10707=>"00000001",
  10708=>"11111101",
  10709=>"00000011",
  10710=>"00000010",
  10711=>"00000011",
  10712=>"00000010",
  10713=>"11111101",
  10714=>"00000000",
  10715=>"00000001",
  10716=>"11111110",
  10717=>"00000001",
  10718=>"11111101",
  10719=>"00000000",
  10720=>"00000001",
  10721=>"00000010",
  10722=>"00000001",
  10723=>"11111111",
  10724=>"00000010",
  10725=>"11111110",
  10726=>"00000011",
  10727=>"00000000",
  10728=>"11111101",
  10729=>"00000010",
  10730=>"11111111",
  10731=>"00000000",
  10732=>"11111110",
  10733=>"11111100",
  10734=>"00000000",
  10735=>"00000010",
  10736=>"11111111",
  10737=>"00000000",
  10738=>"00000000",
  10739=>"00000010",
  10740=>"11111101",
  10741=>"00000001",
  10742=>"11111110",
  10743=>"11111110",
  10744=>"00000000",
  10745=>"00000100",
  10746=>"00000000",
  10747=>"00000010",
  10748=>"11111111",
  10749=>"00000010",
  10750=>"00000011",
  10751=>"11111111",
  10752=>"00000001",
  10753=>"11111111",
  10754=>"00000000",
  10755=>"00000000",
  10756=>"00000000",
  10757=>"11111110",
  10758=>"00000110",
  10759=>"11111111",
  10760=>"11111111",
  10761=>"11111101",
  10762=>"11111110",
  10763=>"11111110",
  10764=>"11111101",
  10765=>"11111101",
  10766=>"00000001",
  10767=>"11111111",
  10768=>"11111111",
  10769=>"00000100",
  10770=>"00000011",
  10771=>"11111111",
  10772=>"11111111",
  10773=>"11111111",
  10774=>"00000000",
  10775=>"11111110",
  10776=>"11111111",
  10777=>"11111110",
  10778=>"11111110",
  10779=>"00000000",
  10780=>"00000011",
  10781=>"00000001",
  10782=>"11111110",
  10783=>"11111111",
  10784=>"00000111",
  10785=>"00000001",
  10786=>"00000010",
  10787=>"00000001",
  10788=>"00000011",
  10789=>"00000101",
  10790=>"11111110",
  10791=>"00000000",
  10792=>"00000101",
  10793=>"00000000",
  10794=>"00000000",
  10795=>"11111100",
  10796=>"11111111",
  10797=>"11111111",
  10798=>"00000001",
  10799=>"00000000",
  10800=>"11111111",
  10801=>"11111111",
  10802=>"11111110",
  10803=>"11111100",
  10804=>"00000100",
  10805=>"00000010",
  10806=>"11111110",
  10807=>"00000001",
  10808=>"11111101",
  10809=>"11111111",
  10810=>"11111111",
  10811=>"00000010",
  10812=>"11111110",
  10813=>"11111110",
  10814=>"00000000",
  10815=>"11111110",
  10816=>"11111110",
  10817=>"11111111",
  10818=>"11111111",
  10819=>"11111110",
  10820=>"11111110",
  10821=>"00000001",
  10822=>"00000000",
  10823=>"11111111",
  10824=>"00000100",
  10825=>"00000010",
  10826=>"11111101",
  10827=>"00000000",
  10828=>"11111110",
  10829=>"00000001",
  10830=>"11111101",
  10831=>"00000010",
  10832=>"11111101",
  10833=>"00000000",
  10834=>"00000010",
  10835=>"00000000",
  10836=>"11111110",
  10837=>"11111111",
  10838=>"11111110",
  10839=>"11111110",
  10840=>"11111111",
  10841=>"00000100",
  10842=>"11111111",
  10843=>"00000001",
  10844=>"11111101",
  10845=>"00000000",
  10846=>"00000001",
  10847=>"11111111",
  10848=>"00000011",
  10849=>"11111111",
  10850=>"00000000",
  10851=>"11111101",
  10852=>"11111110",
  10853=>"00000001",
  10854=>"11111110",
  10855=>"11111101",
  10856=>"00000001",
  10857=>"11111111",
  10858=>"00000000",
  10859=>"11111101",
  10860=>"00000001",
  10861=>"11111111",
  10862=>"00000001",
  10863=>"00000011",
  10864=>"00000010",
  10865=>"00000001",
  10866=>"00000000",
  10867=>"11111100",
  10868=>"00000001",
  10869=>"00000110",
  10870=>"11111111",
  10871=>"11111111",
  10872=>"00000000",
  10873=>"11111111",
  10874=>"11111101",
  10875=>"00000011",
  10876=>"11111110",
  10877=>"00000000",
  10878=>"11111100",
  10879=>"11111110",
  10880=>"11111110",
  10881=>"00000001",
  10882=>"11111110",
  10883=>"00000001",
  10884=>"00000100",
  10885=>"11111111",
  10886=>"00000000",
  10887=>"00000000",
  10888=>"00000010",
  10889=>"00000010",
  10890=>"00000000",
  10891=>"00000001",
  10892=>"11111111",
  10893=>"11111111",
  10894=>"00000010",
  10895=>"11111110",
  10896=>"11111110",
  10897=>"11111110",
  10898=>"11111101",
  10899=>"00000010",
  10900=>"11111101",
  10901=>"00000001",
  10902=>"11111110",
  10903=>"00000011",
  10904=>"11111101",
  10905=>"00000001",
  10906=>"00000000",
  10907=>"11111110",
  10908=>"11111101",
  10909=>"00000001",
  10910=>"11111101",
  10911=>"11111111",
  10912=>"11111111",
  10913=>"11111111",
  10914=>"00000010",
  10915=>"11111100",
  10916=>"00000010",
  10917=>"11111101",
  10918=>"00000000",
  10919=>"00000010",
  10920=>"00000010",
  10921=>"00000011",
  10922=>"11111110",
  10923=>"11111110",
  10924=>"11111110",
  10925=>"11111101",
  10926=>"00000000",
  10927=>"11111110",
  10928=>"11111110",
  10929=>"00000010",
  10930=>"11111110",
  10931=>"00000001",
  10932=>"00000000",
  10933=>"00000000",
  10934=>"11111110",
  10935=>"11111101",
  10936=>"00000010",
  10937=>"00000000",
  10938=>"11111111",
  10939=>"00000100",
  10940=>"11111110",
  10941=>"11111111",
  10942=>"11111101",
  10943=>"00000000",
  10944=>"00000011",
  10945=>"00000010",
  10946=>"00000001",
  10947=>"00000101",
  10948=>"00000010",
  10949=>"11111101",
  10950=>"00000000",
  10951=>"11111111",
  10952=>"00000010",
  10953=>"00000011",
  10954=>"00000010",
  10955=>"00000011",
  10956=>"11111101",
  10957=>"11111111",
  10958=>"11111110",
  10959=>"00000001",
  10960=>"00000010",
  10961=>"00000000",
  10962=>"00000001",
  10963=>"11111101",
  10964=>"00000010",
  10965=>"11111101",
  10966=>"11111110",
  10967=>"00000010",
  10968=>"00000001",
  10969=>"00000000",
  10970=>"11111111",
  10971=>"11111110",
  10972=>"11111110",
  10973=>"00000001",
  10974=>"00000001",
  10975=>"11111100",
  10976=>"11111111",
  10977=>"11111111",
  10978=>"00000100",
  10979=>"11111101",
  10980=>"11111110",
  10981=>"00000010",
  10982=>"00000000",
  10983=>"11111101",
  10984=>"11111111",
  10985=>"00000001",
  10986=>"11111101",
  10987=>"00000001",
  10988=>"00000010",
  10989=>"00000000",
  10990=>"00000011",
  10991=>"00000010",
  10992=>"00000000",
  10993=>"00000001",
  10994=>"00000100",
  10995=>"00000000",
  10996=>"00000010",
  10997=>"11111101",
  10998=>"11111101",
  10999=>"00000001",
  11000=>"00000001",
  11001=>"00000011",
  11002=>"00000000",
  11003=>"00000001",
  11004=>"11111110",
  11005=>"00000000",
  11006=>"00000010",
  11007=>"00000000",
  11008=>"11111111",
  11009=>"00000010",
  11010=>"00000100",
  11011=>"00000100",
  11012=>"00000011",
  11013=>"00000000",
  11014=>"11111110",
  11015=>"11111101",
  11016=>"11111110",
  11017=>"11111101",
  11018=>"00000001",
  11019=>"11111101",
  11020=>"11111111",
  11021=>"00000011",
  11022=>"00000101",
  11023=>"11111101",
  11024=>"11111111",
  11025=>"00000001",
  11026=>"00000000",
  11027=>"11111110",
  11028=>"00000100",
  11029=>"11111111",
  11030=>"00000001",
  11031=>"00000001",
  11032=>"00000000",
  11033=>"00000000",
  11034=>"00000010",
  11035=>"11111110",
  11036=>"00000000",
  11037=>"00000001",
  11038=>"00000001",
  11039=>"00000000",
  11040=>"11111111",
  11041=>"00000011",
  11042=>"11111110",
  11043=>"11111101",
  11044=>"00000010",
  11045=>"11111110",
  11046=>"11111101",
  11047=>"11111101",
  11048=>"11111111",
  11049=>"00000011",
  11050=>"11111100",
  11051=>"00000010",
  11052=>"11111111",
  11053=>"11111111",
  11054=>"00000010",
  11055=>"00000001",
  11056=>"00000010",
  11057=>"11111111",
  11058=>"11111101",
  11059=>"00000010",
  11060=>"11111110",
  11061=>"00000111",
  11062=>"00000001",
  11063=>"11111101",
  11064=>"11111101",
  11065=>"11111111",
  11066=>"11111111",
  11067=>"11111101",
  11068=>"00000010",
  11069=>"11111101",
  11070=>"11111111",
  11071=>"11111111",
  11072=>"11111111",
  11073=>"11111111",
  11074=>"11111111",
  11075=>"00000000",
  11076=>"00000010",
  11077=>"00000001",
  11078=>"11111111",
  11079=>"11111110",
  11080=>"11111110",
  11081=>"00000001",
  11082=>"11111101",
  11083=>"00000001",
  11084=>"00000010",
  11085=>"00000010",
  11086=>"11111111",
  11087=>"00000001",
  11088=>"11111111",
  11089=>"00000001",
  11090=>"00000000",
  11091=>"11111111",
  11092=>"11111111",
  11093=>"11111110",
  11094=>"00000000",
  11095=>"00000001",
  11096=>"00000000",
  11097=>"00000011",
  11098=>"00000010",
  11099=>"00000000",
  11100=>"00000011",
  11101=>"11111111",
  11102=>"00000011",
  11103=>"11111110",
  11104=>"00000011",
  11105=>"11111111",
  11106=>"00000110",
  11107=>"00000000",
  11108=>"00000011",
  11109=>"11111110",
  11110=>"00000101",
  11111=>"11111110",
  11112=>"00000100",
  11113=>"00000011",
  11114=>"00000001",
  11115=>"00000000",
  11116=>"00000010",
  11117=>"11111110",
  11118=>"11111110",
  11119=>"11111111",
  11120=>"00000010",
  11121=>"00000001",
  11122=>"00000010",
  11123=>"11111111",
  11124=>"11111101",
  11125=>"00000000",
  11126=>"00000011",
  11127=>"00000000",
  11128=>"11111110",
  11129=>"00000010",
  11130=>"11111101",
  11131=>"11111111",
  11132=>"11111101",
  11133=>"00000100",
  11134=>"00000000",
  11135=>"00000100",
  11136=>"11111111",
  11137=>"11111111",
  11138=>"00000000",
  11139=>"11111101",
  11140=>"00000001",
  11141=>"00000000",
  11142=>"00000000",
  11143=>"11111111",
  11144=>"00000000",
  11145=>"11111100",
  11146=>"11111101",
  11147=>"11111111",
  11148=>"00000000",
  11149=>"11111111",
  11150=>"00000001",
  11151=>"11111101",
  11152=>"11111110",
  11153=>"00000001",
  11154=>"11111101",
  11155=>"11111111",
  11156=>"11111111",
  11157=>"11111101",
  11158=>"00000101",
  11159=>"00000000",
  11160=>"00000101",
  11161=>"00000011",
  11162=>"00000010",
  11163=>"00000010",
  11164=>"00000100",
  11165=>"00000000",
  11166=>"00000100",
  11167=>"11111110",
  11168=>"11111101",
  11169=>"00000001",
  11170=>"11111111",
  11171=>"00000000",
  11172=>"11111111",
  11173=>"00000100",
  11174=>"11111101",
  11175=>"00000010",
  11176=>"00000100",
  11177=>"11111110",
  11178=>"00000001",
  11179=>"11111111",
  11180=>"11111111",
  11181=>"11111111",
  11182=>"11111111",
  11183=>"00000000",
  11184=>"00000001",
  11185=>"00000010",
  11186=>"00000000",
  11187=>"11111101",
  11188=>"00000001",
  11189=>"00000000",
  11190=>"00000000",
  11191=>"11111111",
  11192=>"00000000",
  11193=>"00000000",
  11194=>"00000000",
  11195=>"00000000",
  11196=>"11111110",
  11197=>"11111110",
  11198=>"00000000",
  11199=>"11111110",
  11200=>"11111101",
  11201=>"11111111",
  11202=>"00000001",
  11203=>"11111111",
  11204=>"00000011",
  11205=>"00000010",
  11206=>"11111110",
  11207=>"00000010",
  11208=>"00000110",
  11209=>"00000100",
  11210=>"11111110",
  11211=>"00000010",
  11212=>"00000010",
  11213=>"00000100",
  11214=>"00000010",
  11215=>"00000001",
  11216=>"11111111",
  11217=>"00000000",
  11218=>"11111011",
  11219=>"11111110",
  11220=>"11111110",
  11221=>"00000000",
  11222=>"00000110",
  11223=>"00000001",
  11224=>"11111110",
  11225=>"00000000",
  11226=>"11111101",
  11227=>"00000001",
  11228=>"00000100",
  11229=>"11111111",
  11230=>"11111111",
  11231=>"11111101",
  11232=>"00000001",
  11233=>"11111111",
  11234=>"00000000",
  11235=>"00000001",
  11236=>"00000101",
  11237=>"00000010",
  11238=>"00000011",
  11239=>"00000001",
  11240=>"00000000",
  11241=>"11111110",
  11242=>"11111110",
  11243=>"11111110",
  11244=>"00000010",
  11245=>"11111110",
  11246=>"11111110",
  11247=>"11111111",
  11248=>"00000100",
  11249=>"11111101",
  11250=>"00000000",
  11251=>"11111101",
  11252=>"00000011",
  11253=>"11111111",
  11254=>"00000001",
  11255=>"11111100",
  11256=>"00000010",
  11257=>"00000010",
  11258=>"11111110",
  11259=>"00000001",
  11260=>"11111110",
  11261=>"00000000",
  11262=>"00000010",
  11263=>"11111111",
  11264=>"00000001",
  11265=>"11111110",
  11266=>"00000010",
  11267=>"00000010",
  11268=>"11111100",
  11269=>"00000100",
  11270=>"00000001",
  11271=>"00000001",
  11272=>"00000110",
  11273=>"00000011",
  11274=>"00000011",
  11275=>"00000010",
  11276=>"11111110",
  11277=>"11111101",
  11278=>"11111101",
  11279=>"11111111",
  11280=>"11111110",
  11281=>"00000010",
  11282=>"11111110",
  11283=>"11111110",
  11284=>"00000011",
  11285=>"00000010",
  11286=>"11111110",
  11287=>"00000000",
  11288=>"00000011",
  11289=>"00000000",
  11290=>"11111110",
  11291=>"11111101",
  11292=>"11111110",
  11293=>"00000010",
  11294=>"00000000",
  11295=>"00000010",
  11296=>"11111111",
  11297=>"11111110",
  11298=>"00000000",
  11299=>"00000000",
  11300=>"11111110",
  11301=>"11111110",
  11302=>"11111100",
  11303=>"00000011",
  11304=>"11111101",
  11305=>"00000100",
  11306=>"00000101",
  11307=>"11111110",
  11308=>"11111100",
  11309=>"00000010",
  11310=>"00000000",
  11311=>"11111110",
  11312=>"11111111",
  11313=>"00000001",
  11314=>"00000010",
  11315=>"11111100",
  11316=>"00000001",
  11317=>"00000000",
  11318=>"00000001",
  11319=>"00000000",
  11320=>"00000100",
  11321=>"00000000",
  11322=>"00000001",
  11323=>"11111101",
  11324=>"00000001",
  11325=>"00000011",
  11326=>"00000101",
  11327=>"11111101",
  11328=>"11111101",
  11329=>"11111111",
  11330=>"00000001",
  11331=>"11111110",
  11332=>"00000001",
  11333=>"00000001",
  11334=>"11111110",
  11335=>"00000010",
  11336=>"00000000",
  11337=>"00000010",
  11338=>"11111110",
  11339=>"00000000",
  11340=>"00000000",
  11341=>"00000010",
  11342=>"00000010",
  11343=>"00000011",
  11344=>"00000010",
  11345=>"11111110",
  11346=>"11111101",
  11347=>"11111111",
  11348=>"00000001",
  11349=>"00000001",
  11350=>"00000001",
  11351=>"00000010",
  11352=>"00000000",
  11353=>"11111110",
  11354=>"00000011",
  11355=>"11111100",
  11356=>"11111101",
  11357=>"00000010",
  11358=>"11111110",
  11359=>"11111111",
  11360=>"11111111",
  11361=>"00000100",
  11362=>"00000001",
  11363=>"00000101",
  11364=>"11111111",
  11365=>"00000010",
  11366=>"00000101",
  11367=>"00000100",
  11368=>"00000001",
  11369=>"11111101",
  11370=>"00000001",
  11371=>"11111110",
  11372=>"00000000",
  11373=>"11111111",
  11374=>"11111110",
  11375=>"11111111",
  11376=>"00000000",
  11377=>"11111101",
  11378=>"00000000",
  11379=>"00000000",
  11380=>"00000001",
  11381=>"11111111",
  11382=>"11111101",
  11383=>"11111110",
  11384=>"00000001",
  11385=>"00000011",
  11386=>"11111101",
  11387=>"00000011",
  11388=>"00000001",
  11389=>"00000000",
  11390=>"11111111",
  11391=>"00000010",
  11392=>"11111110",
  11393=>"00000011",
  11394=>"00000100",
  11395=>"00000100",
  11396=>"00000100",
  11397=>"00000001",
  11398=>"00000001",
  11399=>"11111111",
  11400=>"00000110",
  11401=>"11111110",
  11402=>"00000100",
  11403=>"11111111",
  11404=>"00000000",
  11405=>"00000011",
  11406=>"00000010",
  11407=>"11111110",
  11408=>"11111110",
  11409=>"00000000",
  11410=>"00000000",
  11411=>"00000010",
  11412=>"00000001",
  11413=>"00000000",
  11414=>"11111100",
  11415=>"00000000",
  11416=>"11111111",
  11417=>"11111111",
  11418=>"11111111",
  11419=>"11111110",
  11420=>"00000010",
  11421=>"00000001",
  11422=>"11111110",
  11423=>"11111110",
  11424=>"00000010",
  11425=>"11111110",
  11426=>"00000001",
  11427=>"00000010",
  11428=>"00000011",
  11429=>"00000001",
  11430=>"00000100",
  11431=>"00000010",
  11432=>"00000001",
  11433=>"00000000",
  11434=>"11111111",
  11435=>"11111111",
  11436=>"11111111",
  11437=>"11111111",
  11438=>"00000000",
  11439=>"00000001",
  11440=>"00000001",
  11441=>"11111110",
  11442=>"00000000",
  11443=>"00000010",
  11444=>"00000000",
  11445=>"00000011",
  11446=>"11111110",
  11447=>"11111110",
  11448=>"11111100",
  11449=>"11111111",
  11450=>"11111111",
  11451=>"00000110",
  11452=>"11111110",
  11453=>"00000000",
  11454=>"00000100",
  11455=>"00000010",
  11456=>"00000000",
  11457=>"00000010",
  11458=>"11111110",
  11459=>"11111111",
  11460=>"00000000",
  11461=>"11111101",
  11462=>"11111111",
  11463=>"11111101",
  11464=>"00000001",
  11465=>"00000010",
  11466=>"11111110",
  11467=>"00000001",
  11468=>"11111101",
  11469=>"00000011",
  11470=>"11111110",
  11471=>"00000010",
  11472=>"11111100",
  11473=>"00000001",
  11474=>"00000000",
  11475=>"00000001",
  11476=>"11111111",
  11477=>"11111111",
  11478=>"00000001",
  11479=>"11111111",
  11480=>"00000110",
  11481=>"11111111",
  11482=>"11111110",
  11483=>"11111110",
  11484=>"00000100",
  11485=>"11111111",
  11486=>"00000010",
  11487=>"00000000",
  11488=>"11111101",
  11489=>"11111110",
  11490=>"11111101",
  11491=>"11111111",
  11492=>"00000000",
  11493=>"00000001",
  11494=>"11111110",
  11495=>"00000000",
  11496=>"11111111",
  11497=>"00000001",
  11498=>"00000011",
  11499=>"00000000",
  11500=>"00000001",
  11501=>"00000011",
  11502=>"00000000",
  11503=>"00000010",
  11504=>"11111111",
  11505=>"00000011",
  11506=>"00000001",
  11507=>"00000010",
  11508=>"00000000",
  11509=>"11111110",
  11510=>"11111110",
  11511=>"11111111",
  11512=>"11111111",
  11513=>"00000000",
  11514=>"11111111",
  11515=>"11111111",
  11516=>"00000000",
  11517=>"11111111",
  11518=>"11111111",
  11519=>"00000011",
  11520=>"00000001",
  11521=>"00000010",
  11522=>"11111101",
  11523=>"11111111",
  11524=>"11111111",
  11525=>"00000001",
  11526=>"00000010",
  11527=>"00000001",
  11528=>"11111111",
  11529=>"00000010",
  11530=>"11111101",
  11531=>"00000010",
  11532=>"11111110",
  11533=>"00000001",
  11534=>"00000000",
  11535=>"00000000",
  11536=>"11111101",
  11537=>"00000010",
  11538=>"11111111",
  11539=>"00000000",
  11540=>"11111110",
  11541=>"11111111",
  11542=>"00000001",
  11543=>"00000001",
  11544=>"00000001",
  11545=>"11111111",
  11546=>"00000011",
  11547=>"00000000",
  11548=>"11111111",
  11549=>"00000001",
  11550=>"11111111",
  11551=>"11111111",
  11552=>"11111111",
  11553=>"11111111",
  11554=>"00000001",
  11555=>"00000001",
  11556=>"00000011",
  11557=>"11111111",
  11558=>"11111110",
  11559=>"11111101",
  11560=>"00000001",
  11561=>"11111110",
  11562=>"00000011",
  11563=>"11111101",
  11564=>"00000001",
  11565=>"00000001",
  11566=>"00000001",
  11567=>"00000011",
  11568=>"00000001",
  11569=>"00000011",
  11570=>"11111111",
  11571=>"00000001",
  11572=>"00000000",
  11573=>"11111110",
  11574=>"00000000",
  11575=>"11111110",
  11576=>"00000001",
  11577=>"00000001",
  11578=>"00000010",
  11579=>"11111101",
  11580=>"11111110",
  11581=>"00000101",
  11582=>"00000010",
  11583=>"00000010",
  11584=>"11111111",
  11585=>"11111111",
  11586=>"11111111",
  11587=>"11111110",
  11588=>"00000010",
  11589=>"00000011",
  11590=>"11111100",
  11591=>"00000000",
  11592=>"11111101",
  11593=>"11111110",
  11594=>"00000011",
  11595=>"00000010",
  11596=>"00000001",
  11597=>"11111111",
  11598=>"00000010",
  11599=>"11111111",
  11600=>"11111111",
  11601=>"11111111",
  11602=>"00000011",
  11603=>"00000000",
  11604=>"00000011",
  11605=>"00000001",
  11606=>"00000011",
  11607=>"11111110",
  11608=>"00000011",
  11609=>"00000001",
  11610=>"00000000",
  11611=>"11111110",
  11612=>"00000010",
  11613=>"11111111",
  11614=>"00000001",
  11615=>"00000011",
  11616=>"00000001",
  11617=>"11111101",
  11618=>"00000010",
  11619=>"11111111",
  11620=>"11111101",
  11621=>"00000011",
  11622=>"11111100",
  11623=>"11111110",
  11624=>"00000011",
  11625=>"00000001",
  11626=>"11111110",
  11627=>"00000000",
  11628=>"11111101",
  11629=>"00000100",
  11630=>"00000000",
  11631=>"11111111",
  11632=>"11111111",
  11633=>"00000010",
  11634=>"11111110",
  11635=>"00000011",
  11636=>"11111110",
  11637=>"00000010",
  11638=>"11111101",
  11639=>"11111101",
  11640=>"00000000",
  11641=>"11111111",
  11642=>"11111111",
  11643=>"11111110",
  11644=>"00000001",
  11645=>"11111101",
  11646=>"11111101",
  11647=>"00000000",
  11648=>"00000001",
  11649=>"00000011",
  11650=>"00000001",
  11651=>"00000000",
  11652=>"00000010",
  11653=>"00000000",
  11654=>"00000000",
  11655=>"00000011",
  11656=>"11111111",
  11657=>"00000001",
  11658=>"11111111",
  11659=>"00000000",
  11660=>"00000001",
  11661=>"11111110",
  11662=>"00000101",
  11663=>"00000011",
  11664=>"00000010",
  11665=>"00000001",
  11666=>"00000001",
  11667=>"00000010",
  11668=>"00000001",
  11669=>"00000010",
  11670=>"00000100",
  11671=>"00000010",
  11672=>"11111111",
  11673=>"11111100",
  11674=>"00000001",
  11675=>"11111101",
  11676=>"11111111",
  11677=>"00000010",
  11678=>"11111111",
  11679=>"00000000",
  11680=>"00000000",
  11681=>"11111110",
  11682=>"11111100",
  11683=>"11111111",
  11684=>"00000001",
  11685=>"00000010",
  11686=>"11111110",
  11687=>"11111101",
  11688=>"11111101",
  11689=>"00000000",
  11690=>"00000001",
  11691=>"00000011",
  11692=>"00000010",
  11693=>"11111111",
  11694=>"00000011",
  11695=>"00000001",
  11696=>"11111111",
  11697=>"00000000",
  11698=>"11111111",
  11699=>"11111110",
  11700=>"11111110",
  11701=>"11111110",
  11702=>"00000000",
  11703=>"11111111",
  11704=>"11111110",
  11705=>"00000011",
  11706=>"00000001",
  11707=>"00000001",
  11708=>"11111110",
  11709=>"00000001",
  11710=>"11111101",
  11711=>"00000010",
  11712=>"00000110",
  11713=>"11111101",
  11714=>"11111110",
  11715=>"11111110",
  11716=>"00000001",
  11717=>"11111111",
  11718=>"00000000",
  11719=>"11111100",
  11720=>"00000011",
  11721=>"11111111",
  11722=>"00000010",
  11723=>"00000000",
  11724=>"00000010",
  11725=>"00000001",
  11726=>"11111110",
  11727=>"11111100",
  11728=>"00000011",
  11729=>"00000000",
  11730=>"11111110",
  11731=>"11111111",
  11732=>"00000010",
  11733=>"11111101",
  11734=>"00000000",
  11735=>"11111100",
  11736=>"00000000",
  11737=>"11111110",
  11738=>"00000010",
  11739=>"00000000",
  11740=>"00000101",
  11741=>"00000010",
  11742=>"11111111",
  11743=>"00000011",
  11744=>"00000010",
  11745=>"00000000",
  11746=>"00000000",
  11747=>"00000000",
  11748=>"00000011",
  11749=>"11111110",
  11750=>"00000000",
  11751=>"00000011",
  11752=>"00000001",
  11753=>"00000000",
  11754=>"00000100",
  11755=>"11111110",
  11756=>"11111110",
  11757=>"00000011",
  11758=>"00000000",
  11759=>"11111101",
  11760=>"00000000",
  11761=>"00000001",
  11762=>"11111110",
  11763=>"11111101",
  11764=>"00000011",
  11765=>"00000001",
  11766=>"11111110",
  11767=>"11111101",
  11768=>"00000010",
  11769=>"00000010",
  11770=>"00000011",
  11771=>"00000010",
  11772=>"11111111",
  11773=>"11111111",
  11774=>"00000011",
  11775=>"00000000",
  11776=>"00000011",
  11777=>"11111111",
  11778=>"11111101",
  11779=>"00000010",
  11780=>"11111111",
  11781=>"00000010",
  11782=>"00000010",
  11783=>"11111100",
  11784=>"00000000",
  11785=>"11111111",
  11786=>"00000000",
  11787=>"00000001",
  11788=>"11111110",
  11789=>"00000011",
  11790=>"00000001",
  11791=>"00000010",
  11792=>"00000001",
  11793=>"00000010",
  11794=>"00000001",
  11795=>"11111101",
  11796=>"00000010",
  11797=>"00000100",
  11798=>"11111111",
  11799=>"00000001",
  11800=>"00000001",
  11801=>"11111110",
  11802=>"00000000",
  11803=>"11111110",
  11804=>"00000001",
  11805=>"00000010",
  11806=>"00000011",
  11807=>"00000010",
  11808=>"00000011",
  11809=>"00000010",
  11810=>"11111110",
  11811=>"11111101",
  11812=>"00000010",
  11813=>"11111100",
  11814=>"11111111",
  11815=>"00000011",
  11816=>"00000010",
  11817=>"00000000",
  11818=>"11111111",
  11819=>"00000010",
  11820=>"11111111",
  11821=>"11111101",
  11822=>"11111111",
  11823=>"00000011",
  11824=>"00000100",
  11825=>"11111110",
  11826=>"11111110",
  11827=>"00000000",
  11828=>"11111101",
  11829=>"11111111",
  11830=>"11111110",
  11831=>"00000011",
  11832=>"00000011",
  11833=>"00000011",
  11834=>"11111111",
  11835=>"11111111",
  11836=>"11111111",
  11837=>"00000011",
  11838=>"11111101",
  11839=>"11111111",
  11840=>"00000000",
  11841=>"11111110",
  11842=>"00000000",
  11843=>"11111111",
  11844=>"00000000",
  11845=>"00000110",
  11846=>"00000001",
  11847=>"00000010",
  11848=>"00000011",
  11849=>"00000001",
  11850=>"00000000",
  11851=>"11111100",
  11852=>"00000000",
  11853=>"00000110",
  11854=>"00000101",
  11855=>"00000001",
  11856=>"11111110",
  11857=>"11111100",
  11858=>"11111110",
  11859=>"11111111",
  11860=>"00000001",
  11861=>"11111111",
  11862=>"00000000",
  11863=>"11111111",
  11864=>"11111111",
  11865=>"00000000",
  11866=>"11111111",
  11867=>"00000011",
  11868=>"11111111",
  11869=>"11111110",
  11870=>"11111101",
  11871=>"11111110",
  11872=>"00000000",
  11873=>"00000000",
  11874=>"00000010",
  11875=>"00000110",
  11876=>"00000001",
  11877=>"11111100",
  11878=>"00000011",
  11879=>"11111101",
  11880=>"00000001",
  11881=>"11111110",
  11882=>"11111110",
  11883=>"11111111",
  11884=>"11111110",
  11885=>"11111110",
  11886=>"11111110",
  11887=>"11111111",
  11888=>"11111110",
  11889=>"11111110",
  11890=>"00000010",
  11891=>"00000011",
  11892=>"00000001",
  11893=>"00000100",
  11894=>"11111111",
  11895=>"11111100",
  11896=>"00000000",
  11897=>"00000000",
  11898=>"00000000",
  11899=>"11111101",
  11900=>"00000010",
  11901=>"00000011",
  11902=>"11111110",
  11903=>"11111111",
  11904=>"00000000",
  11905=>"11111101",
  11906=>"11111101",
  11907=>"00000100",
  11908=>"11111110",
  11909=>"11111101",
  11910=>"11111101",
  11911=>"00000010",
  11912=>"11111111",
  11913=>"11111111",
  11914=>"00000001",
  11915=>"11111111",
  11916=>"11111111",
  11917=>"00000000",
  11918=>"00000011",
  11919=>"11111111",
  11920=>"00000000",
  11921=>"00000000",
  11922=>"11111110",
  11923=>"11111111",
  11924=>"00000000",
  11925=>"00000011",
  11926=>"11111111",
  11927=>"11111100",
  11928=>"11111110",
  11929=>"11111101",
  11930=>"11111101",
  11931=>"00000010",
  11932=>"11111101",
  11933=>"00000001",
  11934=>"11111101",
  11935=>"00000000",
  11936=>"00000001",
  11937=>"11111111",
  11938=>"11111111",
  11939=>"00000100",
  11940=>"00000000",
  11941=>"00000000",
  11942=>"00000001",
  11943=>"00000010",
  11944=>"00000011",
  11945=>"11111101",
  11946=>"11111110",
  11947=>"11111101",
  11948=>"00000001",
  11949=>"11111110",
  11950=>"00000010",
  11951=>"11111110",
  11952=>"00000010",
  11953=>"00000010",
  11954=>"00000000",
  11955=>"11111111",
  11956=>"00000000",
  11957=>"00000011",
  11958=>"00000000",
  11959=>"00000010",
  11960=>"11111111",
  11961=>"00000001",
  11962=>"00000000",
  11963=>"11111101",
  11964=>"11111110",
  11965=>"00000001",
  11966=>"00000001",
  11967=>"00000011",
  11968=>"11111110",
  11969=>"11111101",
  11970=>"00000001",
  11971=>"00000000",
  11972=>"00000001",
  11973=>"00000000",
  11974=>"11111111",
  11975=>"11111111",
  11976=>"00000010",
  11977=>"00000001",
  11978=>"00000011",
  11979=>"11111110",
  11980=>"00000001",
  11981=>"11111111",
  11982=>"11111111",
  11983=>"11111111",
  11984=>"00000000",
  11985=>"00000010",
  11986=>"00000010",
  11987=>"11111101",
  11988=>"00000101",
  11989=>"11111111",
  11990=>"00000010",
  11991=>"00000011",
  11992=>"00000010",
  11993=>"11111111",
  11994=>"11111110",
  11995=>"11111101",
  11996=>"11111100",
  11997=>"00000010",
  11998=>"11111110",
  11999=>"11111110",
  12000=>"00000011",
  12001=>"00000011",
  12002=>"00000001",
  12003=>"00000001",
  12004=>"00000000",
  12005=>"11111101",
  12006=>"00000011",
  12007=>"11111101",
  12008=>"00000000",
  12009=>"00000010",
  12010=>"11111101",
  12011=>"11111110",
  12012=>"11111101",
  12013=>"11111111",
  12014=>"00000000",
  12015=>"11111110",
  12016=>"00000000",
  12017=>"11111111",
  12018=>"11111111",
  12019=>"11111111",
  12020=>"00000010",
  12021=>"11111101",
  12022=>"11111111",
  12023=>"00000001",
  12024=>"11111111",
  12025=>"11111111",
  12026=>"00000010",
  12027=>"00000000",
  12028=>"11111111",
  12029=>"11111101",
  12030=>"00000011",
  12031=>"11111110",
  12032=>"00000011",
  12033=>"00000001",
  12034=>"00000001",
  12035=>"11111111",
  12036=>"00000001",
  12037=>"00000000",
  12038=>"11111111",
  12039=>"11111111",
  12040=>"11111110",
  12041=>"00000001",
  12042=>"00000000",
  12043=>"11111110",
  12044=>"11111110",
  12045=>"00000100",
  12046=>"00000000",
  12047=>"00000001",
  12048=>"11111111",
  12049=>"00000011",
  12050=>"00000011",
  12051=>"00000011",
  12052=>"00000000",
  12053=>"11111110",
  12054=>"11111111",
  12055=>"00000001",
  12056=>"00000000",
  12057=>"11111111",
  12058=>"11111101",
  12059=>"00000011",
  12060=>"00000000",
  12061=>"11111110",
  12062=>"00000100",
  12063=>"00000000",
  12064=>"00000100",
  12065=>"00000001",
  12066=>"00000010",
  12067=>"00000001",
  12068=>"00000011",
  12069=>"11111100",
  12070=>"00000010",
  12071=>"11111110",
  12072=>"00000000",
  12073=>"11111110",
  12074=>"11111110",
  12075=>"00000010",
  12076=>"11111110",
  12077=>"00000010",
  12078=>"00000001",
  12079=>"00000011",
  12080=>"00000001",
  12081=>"00000000",
  12082=>"00000000",
  12083=>"00000110",
  12084=>"00000011",
  12085=>"11111101",
  12086=>"00000010",
  12087=>"00000000",
  12088=>"00000001",
  12089=>"00000010",
  12090=>"00000001",
  12091=>"00000011",
  12092=>"11111110",
  12093=>"11111111",
  12094=>"11111110",
  12095=>"11111101",
  12096=>"00000100",
  12097=>"11111101",
  12098=>"00000000",
  12099=>"00000101",
  12100=>"11111110",
  12101=>"00000000",
  12102=>"11111101",
  12103=>"00000100",
  12104=>"00000101",
  12105=>"11111111",
  12106=>"00000001",
  12107=>"11111110",
  12108=>"11111110",
  12109=>"11111111",
  12110=>"00000011",
  12111=>"00000001",
  12112=>"00000011",
  12113=>"00000000",
  12114=>"00000011",
  12115=>"00000001",
  12116=>"00000001",
  12117=>"11111111",
  12118=>"11111111",
  12119=>"00000000",
  12120=>"00000000",
  12121=>"00000100",
  12122=>"11111101",
  12123=>"00000000",
  12124=>"00000000",
  12125=>"11111111",
  12126=>"00000001",
  12127=>"00000000",
  12128=>"00000000",
  12129=>"11111111",
  12130=>"11111111",
  12131=>"00000000",
  12132=>"11111110",
  12133=>"11111111",
  12134=>"00000000",
  12135=>"11111101",
  12136=>"00000010",
  12137=>"11111110",
  12138=>"11111111",
  12139=>"11111101",
  12140=>"00000001",
  12141=>"11111101",
  12142=>"11111101",
  12143=>"00000010",
  12144=>"00000001",
  12145=>"00000010",
  12146=>"00000001",
  12147=>"00000001",
  12148=>"00000000",
  12149=>"00000011",
  12150=>"00000011",
  12151=>"11111110",
  12152=>"00000011",
  12153=>"00000010",
  12154=>"00000001",
  12155=>"11111111",
  12156=>"11111111",
  12157=>"00000000",
  12158=>"00000001",
  12159=>"00000010",
  12160=>"00000011",
  12161=>"11111110",
  12162=>"00000000",
  12163=>"00000010",
  12164=>"00000010",
  12165=>"11111101",
  12166=>"11111101",
  12167=>"00000010",
  12168=>"11111110",
  12169=>"11111111",
  12170=>"00000010",
  12171=>"11111100",
  12172=>"00000001",
  12173=>"00000001",
  12174=>"00000000",
  12175=>"00000000",
  12176=>"00000001",
  12177=>"11111101",
  12178=>"11111101",
  12179=>"11111111",
  12180=>"11111110",
  12181=>"00000011",
  12182=>"11111111",
  12183=>"00000010",
  12184=>"00000010",
  12185=>"00000011",
  12186=>"11111111",
  12187=>"11111111",
  12188=>"11111111",
  12189=>"11111101",
  12190=>"11111101",
  12191=>"00000000",
  12192=>"00000000",
  12193=>"00000010",
  12194=>"11111111",
  12195=>"11111111",
  12196=>"00000011",
  12197=>"11111111",
  12198=>"00000001",
  12199=>"11111110",
  12200=>"00000001",
  12201=>"00000000",
  12202=>"11111110",
  12203=>"00000000",
  12204=>"11111110",
  12205=>"00000011",
  12206=>"11111110",
  12207=>"00000011",
  12208=>"00000110",
  12209=>"11111111",
  12210=>"11111101",
  12211=>"11111101",
  12212=>"11111110",
  12213=>"11111111",
  12214=>"11111101",
  12215=>"11111101",
  12216=>"11111111",
  12217=>"11111111",
  12218=>"00000000",
  12219=>"00000010",
  12220=>"00000000",
  12221=>"00000010",
  12222=>"11111111",
  12223=>"00000100",
  12224=>"00000001",
  12225=>"00000000",
  12226=>"11111110",
  12227=>"11111111",
  12228=>"11111110",
  12229=>"11111110",
  12230=>"00000001",
  12231=>"00000010",
  12232=>"00000001",
  12233=>"00000011",
  12234=>"11111110",
  12235=>"00000011",
  12236=>"00000000",
  12237=>"00000000",
  12238=>"00000010",
  12239=>"00000000",
  12240=>"00000001",
  12241=>"00000010",
  12242=>"00000010",
  12243=>"00000100",
  12244=>"11111111",
  12245=>"00000000",
  12246=>"11111111",
  12247=>"00000010",
  12248=>"11111110",
  12249=>"00000001",
  12250=>"00000000",
  12251=>"00000000",
  12252=>"11111111",
  12253=>"00000000",
  12254=>"00000010",
  12255=>"11111110",
  12256=>"11111110",
  12257=>"00000001",
  12258=>"00000000",
  12259=>"11111110",
  12260=>"00000000",
  12261=>"11111101",
  12262=>"11111100",
  12263=>"11111110",
  12264=>"00000011",
  12265=>"11111111",
  12266=>"11111101",
  12267=>"00000001",
  12268=>"00000001",
  12269=>"00000001",
  12270=>"11111111",
  12271=>"00000000",
  12272=>"00000000",
  12273=>"00000011",
  12274=>"00000000",
  12275=>"00000011",
  12276=>"00000001",
  12277=>"00000100",
  12278=>"00000000",
  12279=>"00000001",
  12280=>"00000001",
  12281=>"00000011",
  12282=>"11111101",
  12283=>"00000010",
  12284=>"00000000",
  12285=>"00000000",
  12286=>"00000011",
  12287=>"00000011",
  12288=>"11111110",
  12289=>"00000000",
  12290=>"11111110",
  12291=>"00000001",
  12292=>"00000001",
  12293=>"11111111",
  12294=>"00000010",
  12295=>"00000001",
  12296=>"11111111",
  12297=>"11111111",
  12298=>"11111111",
  12299=>"11111111",
  12300=>"00000001",
  12301=>"00000001",
  12302=>"00000001",
  12303=>"00000001",
  12304=>"11111111",
  12305=>"00000000",
  12306=>"00000001",
  12307=>"00000001",
  12308=>"11111111",
  12309=>"11111111",
  12310=>"00000000",
  12311=>"00000001",
  12312=>"11111111",
  12313=>"00000001",
  12314=>"00000001",
  12315=>"00000001",
  12316=>"11111111",
  12317=>"00000000",
  12318=>"00000000",
  12319=>"00000000",
  12320=>"11111111",
  12321=>"00000000",
  12322=>"11111111",
  12323=>"00000001",
  12324=>"00000001",
  12325=>"11111111",
  12326=>"00000000",
  12327=>"00000001",
  12328=>"11111110",
  12329=>"00000001",
  12330=>"11111111",
  12331=>"00000010",
  12332=>"11111111",
  12333=>"11111100",
  12334=>"00000000",
  12335=>"00000001",
  12336=>"00000000",
  12337=>"11111110",
  12338=>"00000000",
  12339=>"00000001",
  12340=>"11111101",
  12341=>"11111111",
  12342=>"00000000",
  12343=>"00000000",
  12344=>"00000001",
  12345=>"00000001",
  12346=>"11111110",
  12347=>"11111111",
  12348=>"11111111",
  12349=>"00000000",
  12350=>"11111111",
  12351=>"00000000",
  12352=>"11111110",
  12353=>"00000000",
  12354=>"11111111",
  12355=>"00000001",
  12356=>"00000000",
  12357=>"00000010",
  12358=>"00000000",
  12359=>"00000000",
  12360=>"00000001",
  12361=>"00000010",
  12362=>"00000000",
  12363=>"00000010",
  12364=>"00000010",
  12365=>"00000001",
  12366=>"00000000",
  12367=>"00000000",
  12368=>"00000001",
  12369=>"11111111",
  12370=>"11111111",
  12371=>"11111110",
  12372=>"00000000",
  12373=>"00000000",
  12374=>"00000000",
  12375=>"11111111",
  12376=>"00000000",
  12377=>"00000000",
  12378=>"11111111",
  12379=>"11111111",
  12380=>"00000010",
  12381=>"00000001",
  12382=>"00000000",
  12383=>"11111110",
  12384=>"11111110",
  12385=>"00000001",
  12386=>"00000001",
  12387=>"11111111",
  12388=>"00000001",
  12389=>"11111111",
  12390=>"00000001",
  12391=>"00000000",
  12392=>"00000000",
  12393=>"11111111",
  12394=>"11111110",
  12395=>"11111111",
  12396=>"00000001",
  12397=>"00000001",
  12398=>"00000001",
  12399=>"00000001",
  12400=>"11111111",
  12401=>"11111111",
  12402=>"00000001",
  12403=>"00000000",
  12404=>"00000000",
  12405=>"00000001",
  12406=>"00000010",
  12407=>"00000000",
  12408=>"00000000",
  12409=>"11111111",
  12410=>"00000000",
  12411=>"11111111",
  12412=>"00000001",
  12413=>"00000010",
  12414=>"11111111",
  12415=>"00000010",
  12416=>"00000001",
  12417=>"11111110",
  12418=>"11111110",
  12419=>"00000001",
  12420=>"00000000",
  12421=>"00000010",
  12422=>"00000010",
  12423=>"00000001",
  12424=>"11111111",
  12425=>"11111111",
  12426=>"11111111",
  12427=>"00000010",
  12428=>"11111111",
  12429=>"00000001",
  12430=>"00000001",
  12431=>"11111111",
  12432=>"00000011",
  12433=>"11111111",
  12434=>"00000001",
  12435=>"00000000",
  12436=>"00000000",
  12437=>"00000001",
  12438=>"11111111",
  12439=>"00000001",
  12440=>"00000001",
  12441=>"00000000",
  12442=>"00000001",
  12443=>"00000001",
  12444=>"11111111",
  12445=>"00000000",
  12446=>"00000000",
  12447=>"11111110",
  12448=>"11111111",
  12449=>"00000000",
  12450=>"00000000",
  12451=>"00000001",
  12452=>"00000001",
  12453=>"00000001",
  12454=>"00000000",
  12455=>"00000000",
  12456=>"00000001",
  12457=>"00000000",
  12458=>"00000000",
  12459=>"00000010",
  12460=>"00000000",
  12461=>"11111111",
  12462=>"11111111",
  12463=>"00000000",
  12464=>"11111111",
  12465=>"00000001",
  12466=>"11111111",
  12467=>"00000001",
  12468=>"00000000",
  12469=>"11111111",
  12470=>"11111111",
  12471=>"11111111",
  12472=>"00000000",
  12473=>"11111111",
  12474=>"11111110",
  12475=>"00000001",
  12476=>"11111111",
  12477=>"11111111",
  12478=>"00000001",
  12479=>"00000001",
  12480=>"00000010",
  12481=>"00000000",
  12482=>"00000000",
  12483=>"00000001",
  12484=>"11111111",
  12485=>"11111111",
  12486=>"11111111",
  12487=>"00000001",
  12488=>"00000001",
  12489=>"00000001",
  12490=>"00000001",
  12491=>"11111110",
  12492=>"11111111",
  12493=>"00000001",
  12494=>"00000000",
  12495=>"00000000",
  12496=>"00000001",
  12497=>"00000001",
  12498=>"11111111",
  12499=>"11111111",
  12500=>"00000000",
  12501=>"00000000",
  12502=>"00000001",
  12503=>"11111111",
  12504=>"00000001",
  12505=>"00000001",
  12506=>"00000001",
  12507=>"11111111",
  12508=>"11111110",
  12509=>"00000001",
  12510=>"11111110",
  12511=>"11111111",
  12512=>"11111111",
  12513=>"00000000",
  12514=>"00000001",
  12515=>"11111111",
  12516=>"00000001",
  12517=>"00000001",
  12518=>"00000000",
  12519=>"11111111",
  12520=>"00000000",
  12521=>"00000010",
  12522=>"00000000",
  12523=>"00000001",
  12524=>"00000001",
  12525=>"00000001",
  12526=>"11111111",
  12527=>"11111111",
  12528=>"11111111",
  12529=>"00000000",
  12530=>"00000000",
  12531=>"00000010",
  12532=>"11111110",
  12533=>"11111111",
  12534=>"00000010",
  12535=>"00000001",
  12536=>"00000010",
  12537=>"00000001",
  12538=>"11111111",
  12539=>"00000010",
  12540=>"11111111",
  12541=>"11111111",
  12542=>"00000010",
  12543=>"00000000",
  12544=>"00000001",
  12545=>"00000000",
  12546=>"00000010",
  12547=>"11111111",
  12548=>"11111111",
  12549=>"11111110",
  12550=>"00000001",
  12551=>"00000010",
  12552=>"11111110",
  12553=>"00000001",
  12554=>"00000001",
  12555=>"00000001",
  12556=>"00000001",
  12557=>"00000001",
  12558=>"11111110",
  12559=>"11111111",
  12560=>"11111111",
  12561=>"00000000",
  12562=>"00000010",
  12563=>"00000000",
  12564=>"00000001",
  12565=>"00000001",
  12566=>"11111111",
  12567=>"00000010",
  12568=>"00000000",
  12569=>"11111110",
  12570=>"00000011",
  12571=>"11111111",
  12572=>"00000000",
  12573=>"00000010",
  12574=>"00000001",
  12575=>"11111111",
  12576=>"00000000",
  12577=>"00000000",
  12578=>"00000000",
  12579=>"00000001",
  12580=>"00000010",
  12581=>"00000010",
  12582=>"00000001",
  12583=>"00000010",
  12584=>"00000010",
  12585=>"00000001",
  12586=>"00000010",
  12587=>"00000001",
  12588=>"11111111",
  12589=>"00000001",
  12590=>"00000000",
  12591=>"00000000",
  12592=>"00000000",
  12593=>"00000000",
  12594=>"00000001",
  12595=>"11111111",
  12596=>"00000001",
  12597=>"11111110",
  12598=>"00000000",
  12599=>"00000000",
  12600=>"00000000",
  12601=>"11111111",
  12602=>"00000010",
  12603=>"00000001",
  12604=>"11111111",
  12605=>"00000000",
  12606=>"11111110",
  12607=>"00000000",
  12608=>"11111111",
  12609=>"00000000",
  12610=>"00000000",
  12611=>"11111111",
  12612=>"11111111",
  12613=>"11111111",
  12614=>"00000000",
  12615=>"11111111",
  12616=>"00000000",
  12617=>"00000010",
  12618=>"00000001",
  12619=>"00000000",
  12620=>"00000000",
  12621=>"00000000",
  12622=>"11111110",
  12623=>"11111111",
  12624=>"11111110",
  12625=>"00000001",
  12626=>"00000001",
  12627=>"00000001",
  12628=>"00000001",
  12629=>"11111111",
  12630=>"11111110",
  12631=>"11111110",
  12632=>"00000000",
  12633=>"00000001",
  12634=>"11111110",
  12635=>"00000000",
  12636=>"11111110",
  12637=>"11111110",
  12638=>"00000010",
  12639=>"11111111",
  12640=>"00000000",
  12641=>"11111111",
  12642=>"00000000",
  12643=>"00000001",
  12644=>"11111111",
  12645=>"00000001",
  12646=>"11111111",
  12647=>"00000000",
  12648=>"00000001",
  12649=>"11111111",
  12650=>"11111111",
  12651=>"00000001",
  12652=>"00000000",
  12653=>"11111111",
  12654=>"00000001",
  12655=>"00000001",
  12656=>"11111110",
  12657=>"00000000",
  12658=>"11111111",
  12659=>"00000010",
  12660=>"00000000",
  12661=>"00000000",
  12662=>"11111111",
  12663=>"00000010",
  12664=>"00000001",
  12665=>"11111110",
  12666=>"00000000",
  12667=>"11111110",
  12668=>"11111111",
  12669=>"00000000",
  12670=>"00000000",
  12671=>"00000001",
  12672=>"00000001",
  12673=>"00000010",
  12674=>"00000000",
  12675=>"11111110",
  12676=>"00000001",
  12677=>"00000001",
  12678=>"00000001",
  12679=>"00000000",
  12680=>"11111111",
  12681=>"00000010",
  12682=>"00000010",
  12683=>"00000001",
  12684=>"11111111",
  12685=>"00000001",
  12686=>"00000000",
  12687=>"11111111",
  12688=>"11111110",
  12689=>"00000001",
  12690=>"11111111",
  12691=>"00000001",
  12692=>"11111111",
  12693=>"11111111",
  12694=>"00000001",
  12695=>"11111111",
  12696=>"00000000",
  12697=>"11111111",
  12698=>"11111111",
  12699=>"00000001",
  12700=>"00000001",
  12701=>"00000001",
  12702=>"11111111",
  12703=>"11111111",
  12704=>"00000001",
  12705=>"00000010",
  12706=>"00000000",
  12707=>"11111111",
  12708=>"00000010",
  12709=>"11111110",
  12710=>"00000001",
  12711=>"00000001",
  12712=>"11111111",
  12713=>"00000000",
  12714=>"00000000",
  12715=>"11111110",
  12716=>"11111111",
  12717=>"00000001",
  12718=>"11111111",
  12719=>"11111111",
  12720=>"00000000",
  12721=>"00000000",
  12722=>"11111110",
  12723=>"00000001",
  12724=>"00000000",
  12725=>"00000001",
  12726=>"00000001",
  12727=>"11111111",
  12728=>"00000001",
  12729=>"11111110",
  12730=>"00000001",
  12731=>"00000000",
  12732=>"00000001",
  12733=>"11111110",
  12734=>"00000010",
  12735=>"11111111",
  12736=>"00000010",
  12737=>"00000000",
  12738=>"00000000",
  12739=>"00000001",
  12740=>"00000000",
  12741=>"11111111",
  12742=>"00000001",
  12743=>"00000000",
  12744=>"00000001",
  12745=>"11111110",
  12746=>"00000001",
  12747=>"11111111",
  12748=>"00000011",
  12749=>"11111111",
  12750=>"11111111",
  12751=>"00000000",
  12752=>"00000001",
  12753=>"00000000",
  12754=>"00000000",
  12755=>"11111111",
  12756=>"11111110",
  12757=>"00000000",
  12758=>"00000000",
  12759=>"11111110",
  12760=>"11111111",
  12761=>"11111111",
  12762=>"00000001",
  12763=>"00000000",
  12764=>"11111111",
  12765=>"00000000",
  12766=>"00000000",
  12767=>"11111111",
  12768=>"11111110",
  12769=>"11111111",
  12770=>"00000010",
  12771=>"11111111",
  12772=>"00000000",
  12773=>"00000000",
  12774=>"11111111",
  12775=>"11111110",
  12776=>"00000001",
  12777=>"00000001",
  12778=>"00000000",
  12779=>"00000000",
  12780=>"00000001",
  12781=>"00000010",
  12782=>"11111111",
  12783=>"00000000",
  12784=>"11111111",
  12785=>"00000000",
  12786=>"00000001",
  12787=>"11111111",
  12788=>"00000001",
  12789=>"00000000",
  12790=>"00000000",
  12791=>"11111111",
  12792=>"00000000",
  12793=>"11111111",
  12794=>"00000000",
  12795=>"00000001",
  12796=>"00000001",
  12797=>"00000001",
  12798=>"11111110",
  12799=>"00000001",
  12800=>"00000010",
  12801=>"00000010",
  12802=>"11111111",
  12803=>"11111111",
  12804=>"00000000",
  12805=>"00000000",
  12806=>"00000000",
  12807=>"11111110",
  12808=>"11111111",
  12809=>"00000010",
  12810=>"00000000",
  12811=>"11111110",
  12812=>"00000000",
  12813=>"00000000",
  12814=>"00000000",
  12815=>"00000001",
  12816=>"00000010",
  12817=>"00000000",
  12818=>"11111111",
  12819=>"00000000",
  12820=>"00000001",
  12821=>"00000000",
  12822=>"00000010",
  12823=>"11111111",
  12824=>"00000001",
  12825=>"11111111",
  12826=>"11111101",
  12827=>"11111111",
  12828=>"11111110",
  12829=>"11111111",
  12830=>"00000001",
  12831=>"11111110",
  12832=>"11111110",
  12833=>"11111110",
  12834=>"00000000",
  12835=>"00000000",
  12836=>"00000000",
  12837=>"00000001",
  12838=>"00000001",
  12839=>"00000001",
  12840=>"00000001",
  12841=>"00000010",
  12842=>"00000001",
  12843=>"11111111",
  12844=>"00000000",
  12845=>"00000000",
  12846=>"00000001",
  12847=>"00000000",
  12848=>"00000001",
  12849=>"00000001",
  12850=>"11111110",
  12851=>"00000000",
  12852=>"00000000",
  12853=>"11111111",
  12854=>"00000001",
  12855=>"11111111",
  12856=>"11111111",
  12857=>"00000000",
  12858=>"00000010",
  12859=>"00000000",
  12860=>"00000010",
  12861=>"00000000",
  12862=>"00000001",
  12863=>"00000000",
  12864=>"00000000",
  12865=>"11111111",
  12866=>"11111111",
  12867=>"11111111",
  12868=>"00000010",
  12869=>"00000001",
  12870=>"00000001",
  12871=>"00000000",
  12872=>"00000010",
  12873=>"00000001",
  12874=>"00000000",
  12875=>"00000000",
  12876=>"00000000",
  12877=>"00000000",
  12878=>"00000001",
  12879=>"00000001",
  12880=>"11111111",
  12881=>"00000001",
  12882=>"00000000",
  12883=>"00000001",
  12884=>"11111110",
  12885=>"00000010",
  12886=>"00000010",
  12887=>"11111110",
  12888=>"00000001",
  12889=>"00000001",
  12890=>"00000010",
  12891=>"00000000",
  12892=>"00000000",
  12893=>"00000000",
  12894=>"00000000",
  12895=>"11111111",
  12896=>"00000000",
  12897=>"00000001",
  12898=>"11111111",
  12899=>"00000000",
  12900=>"00000000",
  12901=>"00000001",
  12902=>"11111111",
  12903=>"00000000",
  12904=>"00000001",
  12905=>"00000010",
  12906=>"00000010",
  12907=>"00000000",
  12908=>"00000000",
  12909=>"00000001",
  12910=>"00000000",
  12911=>"00000001",
  12912=>"00000001",
  12913=>"00000001",
  12914=>"11111111",
  12915=>"00000001",
  12916=>"00000001",
  12917=>"11111111",
  12918=>"11111111",
  12919=>"00000000",
  12920=>"11111111",
  12921=>"00000010",
  12922=>"00000001",
  12923=>"00000000",
  12924=>"11111111",
  12925=>"00000000",
  12926=>"00000000",
  12927=>"11111110",
  12928=>"11111111",
  12929=>"00000001",
  12930=>"00000000",
  12931=>"00000000",
  12932=>"00000001",
  12933=>"00000001",
  12934=>"11111111",
  12935=>"11111111",
  12936=>"00000010",
  12937=>"00000001",
  12938=>"00000001",
  12939=>"11111111",
  12940=>"00000000",
  12941=>"11111110",
  12942=>"00000001",
  12943=>"11111111",
  12944=>"00000001",
  12945=>"11111111",
  12946=>"00000010",
  12947=>"00000000",
  12948=>"00000000",
  12949=>"00000010",
  12950=>"00000001",
  12951=>"00000001",
  12952=>"00000010",
  12953=>"00000001",
  12954=>"11111111",
  12955=>"11111111",
  12956=>"11111111",
  12957=>"00000001",
  12958=>"11111111",
  12959=>"00000000",
  12960=>"00000000",
  12961=>"00000001",
  12962=>"11111110",
  12963=>"11111111",
  12964=>"00000010",
  12965=>"11111111",
  12966=>"11111111",
  12967=>"00000001",
  12968=>"11111111",
  12969=>"00000001",
  12970=>"11111110",
  12971=>"00000011",
  12972=>"11111110",
  12973=>"00000010",
  12974=>"00000001",
  12975=>"00000001",
  12976=>"11111111",
  12977=>"00000010",
  12978=>"11111111",
  12979=>"00000001",
  12980=>"00000010",
  12981=>"11111111",
  12982=>"11111111",
  12983=>"00000001",
  12984=>"11111110",
  12985=>"11111111",
  12986=>"11111111",
  12987=>"00000000",
  12988=>"00000001",
  12989=>"11111111",
  12990=>"00000001",
  12991=>"11111111",
  12992=>"11111111",
  12993=>"00000001",
  12994=>"00000000",
  12995=>"11111110",
  12996=>"00000010",
  12997=>"00000001",
  12998=>"00000010",
  12999=>"00000010",
  13000=>"00000000",
  13001=>"00000001",
  13002=>"00000000",
  13003=>"00000001",
  13004=>"00000001",
  13005=>"00000001",
  13006=>"00000000",
  13007=>"11111110",
  13008=>"00000001",
  13009=>"00000010",
  13010=>"00000001",
  13011=>"00000000",
  13012=>"00000010",
  13013=>"00000001",
  13014=>"11111111",
  13015=>"11111110",
  13016=>"11111110",
  13017=>"11111111",
  13018=>"00000000",
  13019=>"11111110",
  13020=>"00000001",
  13021=>"11111110",
  13022=>"00000000",
  13023=>"00000010",
  13024=>"00000001",
  13025=>"11111111",
  13026=>"00000010",
  13027=>"00000001",
  13028=>"00000010",
  13029=>"00000010",
  13030=>"11111111",
  13031=>"00000000",
  13032=>"00000000",
  13033=>"11111111",
  13034=>"00000000",
  13035=>"00000001",
  13036=>"00000001",
  13037=>"00000001",
  13038=>"00000001",
  13039=>"00000000",
  13040=>"00000001",
  13041=>"11111111",
  13042=>"00000010",
  13043=>"00000000",
  13044=>"11111111",
  13045=>"11111111",
  13046=>"00000000",
  13047=>"11111110",
  13048=>"00000000",
  13049=>"11111110",
  13050=>"11111110",
  13051=>"11111111",
  13052=>"11111111",
  13053=>"00000000",
  13054=>"11111110",
  13055=>"00000001",
  13056=>"00000001",
  13057=>"11111111",
  13058=>"00000001",
  13059=>"00000000",
  13060=>"00000010",
  13061=>"11111110",
  13062=>"11111111",
  13063=>"00000001",
  13064=>"00000000",
  13065=>"00000000",
  13066=>"11111111",
  13067=>"11111110",
  13068=>"11111110",
  13069=>"00000001",
  13070=>"11111111",
  13071=>"00000001",
  13072=>"11111110",
  13073=>"11111111",
  13074=>"00000000",
  13075=>"11111111",
  13076=>"00000000",
  13077=>"11111110",
  13078=>"11111111",
  13079=>"11111111",
  13080=>"11111111",
  13081=>"00000000",
  13082=>"00000000",
  13083=>"11111111",
  13084=>"00000010",
  13085=>"00000000",
  13086=>"00000000",
  13087=>"00000000",
  13088=>"11111111",
  13089=>"00000010",
  13090=>"11111111",
  13091=>"11111111",
  13092=>"00000001",
  13093=>"11111111",
  13094=>"00000001",
  13095=>"11111111",
  13096=>"00000001",
  13097=>"11111111",
  13098=>"11111111",
  13099=>"00000010",
  13100=>"11111110",
  13101=>"00000000",
  13102=>"00000001",
  13103=>"11111111",
  13104=>"00000001",
  13105=>"11111110",
  13106=>"11111111",
  13107=>"11111111",
  13108=>"11111110",
  13109=>"00000001",
  13110=>"11111110",
  13111=>"11111111",
  13112=>"00000010",
  13113=>"00000000",
  13114=>"00000000",
  13115=>"00000010",
  13116=>"00000001",
  13117=>"00000011",
  13118=>"00000000",
  13119=>"11111110",
  13120=>"00000001",
  13121=>"00000001",
  13122=>"00000000",
  13123=>"00000000",
  13124=>"00000001",
  13125=>"00000000",
  13126=>"00000000",
  13127=>"00000001",
  13128=>"00000000",
  13129=>"00000010",
  13130=>"00000000",
  13131=>"00000000",
  13132=>"11111111",
  13133=>"11111110",
  13134=>"00000001",
  13135=>"11111111",
  13136=>"11111110",
  13137=>"11111111",
  13138=>"11111111",
  13139=>"11111111",
  13140=>"00000000",
  13141=>"00000001",
  13142=>"00000001",
  13143=>"00000001",
  13144=>"11111111",
  13145=>"11111111",
  13146=>"00000000",
  13147=>"11111110",
  13148=>"11111111",
  13149=>"00000000",
  13150=>"11111111",
  13151=>"00000010",
  13152=>"00000001",
  13153=>"00000001",
  13154=>"00000000",
  13155=>"00000010",
  13156=>"11111111",
  13157=>"11111111",
  13158=>"00000000",
  13159=>"00000000",
  13160=>"11111111",
  13161=>"11111111",
  13162=>"11111111",
  13163=>"00000001",
  13164=>"11111111",
  13165=>"00000001",
  13166=>"00000001",
  13167=>"11111111",
  13168=>"11111110",
  13169=>"11111111",
  13170=>"00000000",
  13171=>"00000001",
  13172=>"00000010",
  13173=>"11111110",
  13174=>"00000000",
  13175=>"11111110",
  13176=>"11111111",
  13177=>"11111111",
  13178=>"11111111",
  13179=>"11111111",
  13180=>"00000000",
  13181=>"00000000",
  13182=>"11111111",
  13183=>"00000000",
  13184=>"11111111",
  13185=>"00000000",
  13186=>"11111111",
  13187=>"00000000",
  13188=>"11111111",
  13189=>"11111110",
  13190=>"00000010",
  13191=>"11111111",
  13192=>"11111111",
  13193=>"11111111",
  13194=>"00000010",
  13195=>"00000000",
  13196=>"11111110",
  13197=>"11111111",
  13198=>"00000001",
  13199=>"11111110",
  13200=>"00000010",
  13201=>"11111111",
  13202=>"00000001",
  13203=>"00000001",
  13204=>"11111111",
  13205=>"00000000",
  13206=>"00000001",
  13207=>"00000000",
  13208=>"00000000",
  13209=>"11111110",
  13210=>"00000001",
  13211=>"00000001",
  13212=>"00000000",
  13213=>"00000001",
  13214=>"00000000",
  13215=>"00000001",
  13216=>"00000000",
  13217=>"00000001",
  13218=>"11111111",
  13219=>"00000001",
  13220=>"00000010",
  13221=>"11111111",
  13222=>"11111110",
  13223=>"11111111",
  13224=>"11111111",
  13225=>"00000010",
  13226=>"00000000",
  13227=>"11111111",
  13228=>"00000000",
  13229=>"11111110",
  13230=>"11111111",
  13231=>"11111111",
  13232=>"11111111",
  13233=>"11111110",
  13234=>"11111111",
  13235=>"00000000",
  13236=>"00000000",
  13237=>"11111111",
  13238=>"11111111",
  13239=>"11111111",
  13240=>"00000000",
  13241=>"00000010",
  13242=>"11111101",
  13243=>"00000011",
  13244=>"00000010",
  13245=>"00000000",
  13246=>"00000001",
  13247=>"00000000",
  13248=>"00000000",
  13249=>"00000010",
  13250=>"11111111",
  13251=>"11111111",
  13252=>"11111110",
  13253=>"11111111",
  13254=>"11111111",
  13255=>"11111111",
  13256=>"11111111",
  13257=>"00000000",
  13258=>"00000001",
  13259=>"00000010",
  13260=>"00000000",
  13261=>"00000010",
  13262=>"00000000",
  13263=>"00000010",
  13264=>"00000001",
  13265=>"00000000",
  13266=>"00000000",
  13267=>"00000000",
  13268=>"00000010",
  13269=>"00000001",
  13270=>"00000000",
  13271=>"11111111",
  13272=>"11111111",
  13273=>"00000000",
  13274=>"11111110",
  13275=>"11111110",
  13276=>"11111110",
  13277=>"00000010",
  13278=>"00000001",
  13279=>"00000000",
  13280=>"00000010",
  13281=>"00000001",
  13282=>"11111111",
  13283=>"11111110",
  13284=>"11111111",
  13285=>"00000000",
  13286=>"11111111",
  13287=>"00000000",
  13288=>"00000001",
  13289=>"00000001",
  13290=>"11111111",
  13291=>"11111111",
  13292=>"00000000",
  13293=>"00000001",
  13294=>"11111111",
  13295=>"00000000",
  13296=>"11111111",
  13297=>"00000000",
  13298=>"11111110",
  13299=>"11111111",
  13300=>"00000010",
  13301=>"00000000",
  13302=>"00000000",
  13303=>"11111110",
  13304=>"11111111",
  13305=>"00000000",
  13306=>"00000000",
  13307=>"00000000",
  13308=>"00000000",
  13309=>"00000001",
  13310=>"00000001",
  13311=>"00000000",
  13312=>"00000010",
  13313=>"00000011",
  13314=>"00000000",
  13315=>"00000010",
  13316=>"00000000",
  13317=>"00000001",
  13318=>"00000001",
  13319=>"11111110",
  13320=>"00000000",
  13321=>"00000001",
  13322=>"00000001",
  13323=>"11111110",
  13324=>"11111111",
  13325=>"00000001",
  13326=>"00000001",
  13327=>"00000001",
  13328=>"00000000",
  13329=>"00000001",
  13330=>"00000001",
  13331=>"11111111",
  13332=>"11111111",
  13333=>"11111111",
  13334=>"00000000",
  13335=>"00000000",
  13336=>"00000010",
  13337=>"00000001",
  13338=>"00000001",
  13339=>"11111111",
  13340=>"00000010",
  13341=>"00000001",
  13342=>"00000001",
  13343=>"00000000",
  13344=>"00000000",
  13345=>"00000000",
  13346=>"00000000",
  13347=>"00000001",
  13348=>"00000000",
  13349=>"00000001",
  13350=>"11111110",
  13351=>"00000001",
  13352=>"00000001",
  13353=>"00000000",
  13354=>"00000010",
  13355=>"11111110",
  13356=>"00000000",
  13357=>"00000000",
  13358=>"00000001",
  13359=>"00000010",
  13360=>"11111111",
  13361=>"00000010",
  13362=>"11111110",
  13363=>"00000000",
  13364=>"11111101",
  13365=>"00000001",
  13366=>"11111110",
  13367=>"00000001",
  13368=>"11111111",
  13369=>"00000010",
  13370=>"11111111",
  13371=>"11111111",
  13372=>"00000000",
  13373=>"11111111",
  13374=>"00000001",
  13375=>"00000010",
  13376=>"00000010",
  13377=>"11111110",
  13378=>"00000001",
  13379=>"00000000",
  13380=>"00000000",
  13381=>"00000010",
  13382=>"11111110",
  13383=>"00000011",
  13384=>"00000000",
  13385=>"11111110",
  13386=>"00000001",
  13387=>"11111111",
  13388=>"00000000",
  13389=>"00000000",
  13390=>"11111110",
  13391=>"00000010",
  13392=>"00000000",
  13393=>"11111111",
  13394=>"00000000",
  13395=>"11111111",
  13396=>"00000001",
  13397=>"00000000",
  13398=>"00000000",
  13399=>"11111110",
  13400=>"00000000",
  13401=>"00000010",
  13402=>"11111110",
  13403=>"00000001",
  13404=>"00000000",
  13405=>"00000010",
  13406=>"00000010",
  13407=>"11111111",
  13408=>"11111111",
  13409=>"00000001",
  13410=>"00000000",
  13411=>"11111111",
  13412=>"00000001",
  13413=>"00000001",
  13414=>"11111111",
  13415=>"11111111",
  13416=>"00000001",
  13417=>"11111111",
  13418=>"11111111",
  13419=>"11111111",
  13420=>"11111110",
  13421=>"00000001",
  13422=>"11111110",
  13423=>"11111111",
  13424=>"00000000",
  13425=>"00000001",
  13426=>"00000010",
  13427=>"11111111",
  13428=>"00000010",
  13429=>"11111111",
  13430=>"11111111",
  13431=>"00000000",
  13432=>"11111111",
  13433=>"00000000",
  13434=>"11111111",
  13435=>"00000001",
  13436=>"00000000",
  13437=>"00000000",
  13438=>"00000010",
  13439=>"00000001",
  13440=>"11111110",
  13441=>"11111111",
  13442=>"11111110",
  13443=>"00000001",
  13444=>"00000011",
  13445=>"00000000",
  13446=>"11111110",
  13447=>"00000001",
  13448=>"00000001",
  13449=>"00000001",
  13450=>"00000010",
  13451=>"00000001",
  13452=>"11111111",
  13453=>"00000010",
  13454=>"11111111",
  13455=>"00000010",
  13456=>"11111111",
  13457=>"11111111",
  13458=>"11111111",
  13459=>"00000000",
  13460=>"00000000",
  13461=>"00000000",
  13462=>"00000010",
  13463=>"00000001",
  13464=>"11111101",
  13465=>"11111111",
  13466=>"00000000",
  13467=>"11111111",
  13468=>"00000001",
  13469=>"11111111",
  13470=>"11111110",
  13471=>"00000010",
  13472=>"00000001",
  13473=>"11111111",
  13474=>"00000010",
  13475=>"00000001",
  13476=>"00000001",
  13477=>"00000001",
  13478=>"11111111",
  13479=>"11111111",
  13480=>"00000000",
  13481=>"00000000",
  13482=>"11111110",
  13483=>"00000001",
  13484=>"11111111",
  13485=>"00000000",
  13486=>"11111111",
  13487=>"00000001",
  13488=>"00000000",
  13489=>"00000001",
  13490=>"11111111",
  13491=>"00000010",
  13492=>"11111111",
  13493=>"11111110",
  13494=>"00000001",
  13495=>"11111111",
  13496=>"00000000",
  13497=>"11111111",
  13498=>"00000010",
  13499=>"11111110",
  13500=>"00000001",
  13501=>"11111110",
  13502=>"11111110",
  13503=>"00000001",
  13504=>"11111111",
  13505=>"00000001",
  13506=>"00000000",
  13507=>"00000010",
  13508=>"00000000",
  13509=>"11111110",
  13510=>"11111111",
  13511=>"11111110",
  13512=>"11111111",
  13513=>"00000000",
  13514=>"00000001",
  13515=>"00000001",
  13516=>"00000010",
  13517=>"11111111",
  13518=>"00000000",
  13519=>"11111111",
  13520=>"11111111",
  13521=>"00000001",
  13522=>"11111111",
  13523=>"00000001",
  13524=>"00000001",
  13525=>"11111111",
  13526=>"11111110",
  13527=>"11111111",
  13528=>"00000000",
  13529=>"11111110",
  13530=>"11111111",
  13531=>"00000000",
  13532=>"11111110",
  13533=>"00000000",
  13534=>"11111111",
  13535=>"11111111",
  13536=>"00000100",
  13537=>"00000001",
  13538=>"00000000",
  13539=>"00000000",
  13540=>"00000010",
  13541=>"00000001",
  13542=>"00000000",
  13543=>"11111110",
  13544=>"00000000",
  13545=>"00000000",
  13546=>"00000010",
  13547=>"11111110",
  13548=>"00000000",
  13549=>"11111111",
  13550=>"11111111",
  13551=>"00000010",
  13552=>"11111110",
  13553=>"00000001",
  13554=>"11111111",
  13555=>"00000001",
  13556=>"00000001",
  13557=>"00000001",
  13558=>"00000010",
  13559=>"11111111",
  13560=>"00000000",
  13561=>"11111110",
  13562=>"00000000",
  13563=>"00000010",
  13564=>"00000000",
  13565=>"00000000",
  13566=>"11111111",
  13567=>"00000000",
  13568=>"11111111",
  13569=>"00000001",
  13570=>"00000011",
  13571=>"11111111",
  13572=>"11111111",
  13573=>"00000000",
  13574=>"11111110",
  13575=>"00000001",
  13576=>"00000000",
  13577=>"11111111",
  13578=>"00000001",
  13579=>"11111111",
  13580=>"00000010",
  13581=>"00000010",
  13582=>"11111110",
  13583=>"00000001",
  13584=>"00000000",
  13585=>"00000000",
  13586=>"00000001",
  13587=>"11111110",
  13588=>"11111111",
  13589=>"00000000",
  13590=>"00000000",
  13591=>"00000001",
  13592=>"00000001",
  13593=>"00000001",
  13594=>"00000001",
  13595=>"00000000",
  13596=>"00000000",
  13597=>"00000010",
  13598=>"00000001",
  13599=>"00000001",
  13600=>"00000000",
  13601=>"00000001",
  13602=>"00000010",
  13603=>"00000001",
  13604=>"11111111",
  13605=>"11111111",
  13606=>"00000000",
  13607=>"00000010",
  13608=>"00000001",
  13609=>"00000000",
  13610=>"11111111",
  13611=>"11111111",
  13612=>"11111110",
  13613=>"00000000",
  13614=>"11111101",
  13615=>"00000000",
  13616=>"11111110",
  13617=>"00000010",
  13618=>"00000001",
  13619=>"11111111",
  13620=>"00000000",
  13621=>"11111110",
  13622=>"11111111",
  13623=>"11111111",
  13624=>"00000001",
  13625=>"00000001",
  13626=>"00000000",
  13627=>"11111111",
  13628=>"00000000",
  13629=>"11111111",
  13630=>"11111110",
  13631=>"11111110",
  13632=>"00000000",
  13633=>"00000010",
  13634=>"00000010",
  13635=>"00000000",
  13636=>"11111111",
  13637=>"00000000",
  13638=>"00000000",
  13639=>"00000010",
  13640=>"00000000",
  13641=>"00000000",
  13642=>"11111111",
  13643=>"00000000",
  13644=>"11111111",
  13645=>"00000001",
  13646=>"11111111",
  13647=>"00000000",
  13648=>"00000001",
  13649=>"00000001",
  13650=>"00000001",
  13651=>"11111110",
  13652=>"11111101",
  13653=>"00000001",
  13654=>"11111110",
  13655=>"00000001",
  13656=>"00000001",
  13657=>"11111101",
  13658=>"11111110",
  13659=>"11111111",
  13660=>"00000000",
  13661=>"11111111",
  13662=>"00000000",
  13663=>"00000011",
  13664=>"11111111",
  13665=>"00000000",
  13666=>"00000001",
  13667=>"00000001",
  13668=>"00000001",
  13669=>"11111110",
  13670=>"00000000",
  13671=>"11111111",
  13672=>"11111111",
  13673=>"00000011",
  13674=>"00000010",
  13675=>"00000000",
  13676=>"00000000",
  13677=>"11111110",
  13678=>"00000000",
  13679=>"11111110",
  13680=>"11111111",
  13681=>"11111111",
  13682=>"11111110",
  13683=>"11111111",
  13684=>"00000000",
  13685=>"11111111",
  13686=>"11111110",
  13687=>"11111110",
  13688=>"00000000",
  13689=>"11111101",
  13690=>"11111111",
  13691=>"00000010",
  13692=>"11111111",
  13693=>"11111110",
  13694=>"00000001",
  13695=>"00000010",
  13696=>"00000000",
  13697=>"00000000",
  13698=>"11111110",
  13699=>"11111111",
  13700=>"00000001",
  13701=>"00000000",
  13702=>"00000010",
  13703=>"00000001",
  13704=>"11111111",
  13705=>"00000010",
  13706=>"00000010",
  13707=>"00000011",
  13708=>"11111110",
  13709=>"00000001",
  13710=>"00000010",
  13711=>"11111110",
  13712=>"11111110",
  13713=>"00000010",
  13714=>"00000000",
  13715=>"00000000",
  13716=>"00000000",
  13717=>"00000000",
  13718=>"00000001",
  13719=>"00000001",
  13720=>"00000000",
  13721=>"11111111",
  13722=>"00000001",
  13723=>"11111101",
  13724=>"11111111",
  13725=>"00000000",
  13726=>"00000000",
  13727=>"00000010",
  13728=>"00000001",
  13729=>"00000001",
  13730=>"11111111",
  13731=>"11111111",
  13732=>"11111111",
  13733=>"11111111",
  13734=>"00000010",
  13735=>"00000001",
  13736=>"00000010",
  13737=>"00000001",
  13738=>"00000000",
  13739=>"11111110",
  13740=>"00000001",
  13741=>"11111111",
  13742=>"00000000",
  13743=>"00000000",
  13744=>"11111111",
  13745=>"00000000",
  13746=>"11111110",
  13747=>"00000001",
  13748=>"11111111",
  13749=>"00000001",
  13750=>"11111111",
  13751=>"00000000",
  13752=>"11111110",
  13753=>"00000010",
  13754=>"00000001",
  13755=>"00000000",
  13756=>"11111111",
  13757=>"00000000",
  13758=>"11111111",
  13759=>"11111111",
  13760=>"11111110",
  13761=>"00000000",
  13762=>"00000001",
  13763=>"11111111",
  13764=>"00000001",
  13765=>"00000001",
  13766=>"00000000",
  13767=>"00000000",
  13768=>"11111111",
  13769=>"11111110",
  13770=>"00000000",
  13771=>"11111111",
  13772=>"00000000",
  13773=>"00000010",
  13774=>"00000001",
  13775=>"00000001",
  13776=>"00000000",
  13777=>"11111110",
  13778=>"11111111",
  13779=>"00000000",
  13780=>"00000001",
  13781=>"00000000",
  13782=>"11111110",
  13783=>"11111110",
  13784=>"00000000",
  13785=>"00000001",
  13786=>"11111110",
  13787=>"00000001",
  13788=>"11111111",
  13789=>"00000000",
  13790=>"11111110",
  13791=>"11111110",
  13792=>"00000010",
  13793=>"00000001",
  13794=>"00000000",
  13795=>"11111111",
  13796=>"11111110",
  13797=>"11111110",
  13798=>"11111110",
  13799=>"00000001",
  13800=>"00000000",
  13801=>"00000001",
  13802=>"00000000",
  13803=>"00000001",
  13804=>"00000001",
  13805=>"00000001",
  13806=>"00000001",
  13807=>"00000010",
  13808=>"00000010",
  13809=>"00000010",
  13810=>"00000000",
  13811=>"00000001",
  13812=>"00000000",
  13813=>"00000001",
  13814=>"00000001",
  13815=>"11111111",
  13816=>"11111111",
  13817=>"11111111",
  13818=>"00000001",
  13819=>"00000001",
  13820=>"00000001",
  13821=>"11111110",
  13822=>"00000010",
  13823=>"00000001",
  13824=>"00000010",
  13825=>"00000000",
  13826=>"11111111",
  13827=>"11111110",
  13828=>"00000000",
  13829=>"00000000",
  13830=>"00000001",
  13831=>"00000001",
  13832=>"11111111",
  13833=>"00000001",
  13834=>"00000001",
  13835=>"00000001",
  13836=>"00000000",
  13837=>"11111111",
  13838=>"00000000",
  13839=>"11111110",
  13840=>"11111111",
  13841=>"11111110",
  13842=>"00000010",
  13843=>"00000010",
  13844=>"00000001",
  13845=>"00000001",
  13846=>"00000010",
  13847=>"11111110",
  13848=>"11111110",
  13849=>"00000010",
  13850=>"00000010",
  13851=>"00000001",
  13852=>"00000010",
  13853=>"00000000",
  13854=>"00000000",
  13855=>"00000010",
  13856=>"00000010",
  13857=>"00000001",
  13858=>"00000001",
  13859=>"11111111",
  13860=>"00000000",
  13861=>"00000000",
  13862=>"11111111",
  13863=>"00000000",
  13864=>"11111111",
  13865=>"00000010",
  13866=>"00000000",
  13867=>"11111111",
  13868=>"11111111",
  13869=>"00000010",
  13870=>"00000000",
  13871=>"00000000",
  13872=>"00000001",
  13873=>"00000000",
  13874=>"11111111",
  13875=>"00000001",
  13876=>"11111111",
  13877=>"11111111",
  13878=>"00000001",
  13879=>"00000000",
  13880=>"00000000",
  13881=>"00000001",
  13882=>"11111111",
  13883=>"11111110",
  13884=>"11111110",
  13885=>"00000001",
  13886=>"00000001",
  13887=>"11111111",
  13888=>"00000001",
  13889=>"11111111",
  13890=>"00000001",
  13891=>"11111111",
  13892=>"00000001",
  13893=>"00000010",
  13894=>"00000001",
  13895=>"00000001",
  13896=>"00000001",
  13897=>"00000010",
  13898=>"00000000",
  13899=>"00000010",
  13900=>"00000001",
  13901=>"11111111",
  13902=>"00000000",
  13903=>"00000010",
  13904=>"00000010",
  13905=>"00000001",
  13906=>"00000000",
  13907=>"00000000",
  13908=>"11111110",
  13909=>"11111111",
  13910=>"00000010",
  13911=>"00000000",
  13912=>"00000001",
  13913=>"11111111",
  13914=>"00000000",
  13915=>"11111110",
  13916=>"11111110",
  13917=>"11111011",
  13918=>"11111111",
  13919=>"00000010",
  13920=>"00000000",
  13921=>"00000001",
  13922=>"11111111",
  13923=>"11111110",
  13924=>"00000001",
  13925=>"00000001",
  13926=>"11111111",
  13927=>"00000000",
  13928=>"00000000",
  13929=>"00000010",
  13930=>"11111111",
  13931=>"00000001",
  13932=>"11111110",
  13933=>"00000000",
  13934=>"00000000",
  13935=>"11111111",
  13936=>"00000000",
  13937=>"00000010",
  13938=>"00000001",
  13939=>"00000001",
  13940=>"11111111",
  13941=>"11111111",
  13942=>"11111110",
  13943=>"11111111",
  13944=>"11111111",
  13945=>"11111111",
  13946=>"11111101",
  13947=>"00000000",
  13948=>"00000000",
  13949=>"00000000",
  13950=>"11111111",
  13951=>"11111111",
  13952=>"11111110",
  13953=>"00000000",
  13954=>"11111111",
  13955=>"00000001",
  13956=>"11111111",
  13957=>"00000000",
  13958=>"11111110",
  13959=>"00000010",
  13960=>"11111111",
  13961=>"00000000",
  13962=>"00000001",
  13963=>"00000000",
  13964=>"11111111",
  13965=>"00000011",
  13966=>"11111111",
  13967=>"00000010",
  13968=>"00000001",
  13969=>"00000010",
  13970=>"00000000",
  13971=>"11111110",
  13972=>"11111111",
  13973=>"00000001",
  13974=>"11111111",
  13975=>"00000001",
  13976=>"00000000",
  13977=>"11111111",
  13978=>"00000000",
  13979=>"00000011",
  13980=>"00000001",
  13981=>"00000001",
  13982=>"00000010",
  13983=>"00000000",
  13984=>"00000000",
  13985=>"11111110",
  13986=>"11111111",
  13987=>"00000000",
  13988=>"00000001",
  13989=>"11111111",
  13990=>"00000000",
  13991=>"11111110",
  13992=>"00000001",
  13993=>"11111110",
  13994=>"00000000",
  13995=>"00000001",
  13996=>"00000010",
  13997=>"00000001",
  13998=>"00000010",
  13999=>"00000001",
  14000=>"00000001",
  14001=>"00000001",
  14002=>"00000010",
  14003=>"11111111",
  14004=>"11111111",
  14005=>"11111110",
  14006=>"00000010",
  14007=>"00000000",
  14008=>"11111111",
  14009=>"11111111",
  14010=>"00000000",
  14011=>"00000010",
  14012=>"11111110",
  14013=>"11111111",
  14014=>"00000000",
  14015=>"00000000",
  14016=>"00000010",
  14017=>"00000001",
  14018=>"11111101",
  14019=>"00000001",
  14020=>"11111111",
  14021=>"00000000",
  14022=>"00000001",
  14023=>"11111110",
  14024=>"00000001",
  14025=>"11111111",
  14026=>"11111110",
  14027=>"00000000",
  14028=>"11111110",
  14029=>"00000001",
  14030=>"00000000",
  14031=>"00000001",
  14032=>"00000000",
  14033=>"00000000",
  14034=>"00000010",
  14035=>"00000001",
  14036=>"00000000",
  14037=>"00000001",
  14038=>"00000000",
  14039=>"00000010",
  14040=>"11111111",
  14041=>"11111110",
  14042=>"00000001",
  14043=>"00000000",
  14044=>"00000001",
  14045=>"11111111",
  14046=>"00000001",
  14047=>"00000000",
  14048=>"11111110",
  14049=>"00000011",
  14050=>"11111111",
  14051=>"00000000",
  14052=>"00000001",
  14053=>"11111110",
  14054=>"11111111",
  14055=>"11111111",
  14056=>"11111111",
  14057=>"00000000",
  14058=>"00000001",
  14059=>"11111111",
  14060=>"00000000",
  14061=>"11111110",
  14062=>"11111111",
  14063=>"00000010",
  14064=>"00000000",
  14065=>"11111111",
  14066=>"00000001",
  14067=>"11111110",
  14068=>"00000011",
  14069=>"11111111",
  14070=>"00000011",
  14071=>"11111110",
  14072=>"11111111",
  14073=>"00000001",
  14074=>"00000001",
  14075=>"00000010",
  14076=>"00000000",
  14077=>"00000000",
  14078=>"00000000",
  14079=>"00000001",
  14080=>"00000000",
  14081=>"00000001",
  14082=>"11111101",
  14083=>"11111110",
  14084=>"11111110",
  14085=>"00000000",
  14086=>"11111111",
  14087=>"11111111",
  14088=>"11111110",
  14089=>"00000010",
  14090=>"00000000",
  14091=>"00000000",
  14092=>"11111111",
  14093=>"00000000",
  14094=>"11111111",
  14095=>"00000010",
  14096=>"00000001",
  14097=>"11111101",
  14098=>"00000001",
  14099=>"00000001",
  14100=>"11111111",
  14101=>"00000001",
  14102=>"00000001",
  14103=>"00000000",
  14104=>"00000000",
  14105=>"11111111",
  14106=>"00000000",
  14107=>"11111111",
  14108=>"00000010",
  14109=>"11111111",
  14110=>"00000010",
  14111=>"11111111",
  14112=>"11111101",
  14113=>"11111101",
  14114=>"11111111",
  14115=>"00000000",
  14116=>"00000000",
  14117=>"00000001",
  14118=>"11111111",
  14119=>"00000001",
  14120=>"00000000",
  14121=>"00000001",
  14122=>"11111110",
  14123=>"00000010",
  14124=>"00000000",
  14125=>"00000000",
  14126=>"11111111",
  14127=>"11111111",
  14128=>"00000001",
  14129=>"00000000",
  14130=>"00000010",
  14131=>"00000000",
  14132=>"11111111",
  14133=>"00000000",
  14134=>"11111111",
  14135=>"00000010",
  14136=>"11111110",
  14137=>"00000001",
  14138=>"00000010",
  14139=>"00000001",
  14140=>"00000000",
  14141=>"00000011",
  14142=>"11111110",
  14143=>"00000000",
  14144=>"00000001",
  14145=>"00000000",
  14146=>"11111111",
  14147=>"00000000",
  14148=>"11111111",
  14149=>"00000010",
  14150=>"11111111",
  14151=>"00000001",
  14152=>"00000001",
  14153=>"11111111",
  14154=>"00000000",
  14155=>"11111110",
  14156=>"00000010",
  14157=>"11111110",
  14158=>"11111110",
  14159=>"11111111",
  14160=>"00000001",
  14161=>"11111110",
  14162=>"11111110",
  14163=>"00000001",
  14164=>"00000001",
  14165=>"00000001",
  14166=>"00000000",
  14167=>"00000001",
  14168=>"00000010",
  14169=>"11111111",
  14170=>"00000000",
  14171=>"00000000",
  14172=>"11111111",
  14173=>"00000000",
  14174=>"11111111",
  14175=>"11111111",
  14176=>"11111111",
  14177=>"00000001",
  14178=>"00000001",
  14179=>"00000001",
  14180=>"00000000",
  14181=>"11111111",
  14182=>"11111111",
  14183=>"11111110",
  14184=>"00000000",
  14185=>"00000001",
  14186=>"11111111",
  14187=>"00000000",
  14188=>"11111110",
  14189=>"00000000",
  14190=>"00000010",
  14191=>"00000000",
  14192=>"00000000",
  14193=>"11111101",
  14194=>"00000000",
  14195=>"11111110",
  14196=>"11111111",
  14197=>"00000010",
  14198=>"00000001",
  14199=>"00000000",
  14200=>"11111111",
  14201=>"00000001",
  14202=>"00000000",
  14203=>"00000000",
  14204=>"11111111",
  14205=>"00000001",
  14206=>"00000000",
  14207=>"00000001",
  14208=>"11111111",
  14209=>"00000000",
  14210=>"11111111",
  14211=>"00000010",
  14212=>"00000000",
  14213=>"00000001",
  14214=>"11111110",
  14215=>"11111111",
  14216=>"00000000",
  14217=>"11111111",
  14218=>"00000001",
  14219=>"00000000",
  14220=>"00000000",
  14221=>"11111111",
  14222=>"11111111",
  14223=>"00000000",
  14224=>"00000000",
  14225=>"00000001",
  14226=>"00000000",
  14227=>"00000010",
  14228=>"00000000",
  14229=>"11111111",
  14230=>"11111110",
  14231=>"00000001",
  14232=>"00000010",
  14233=>"00000010",
  14234=>"00000000",
  14235=>"11111111",
  14236=>"00000001",
  14237=>"11111110",
  14238=>"00000010",
  14239=>"00000011",
  14240=>"00000000",
  14241=>"11111111",
  14242=>"00000010",
  14243=>"11111111",
  14244=>"00000011",
  14245=>"00000001",
  14246=>"11111111",
  14247=>"00000001",
  14248=>"11111110",
  14249=>"00000010",
  14250=>"11111110",
  14251=>"00000001",
  14252=>"11111111",
  14253=>"11111111",
  14254=>"00000010",
  14255=>"00000010",
  14256=>"00000001",
  14257=>"11111111",
  14258=>"00000001",
  14259=>"11111111",
  14260=>"00000001",
  14261=>"11111110",
  14262=>"11111101",
  14263=>"00000010",
  14264=>"00000010",
  14265=>"00000000",
  14266=>"00000010",
  14267=>"11111111",
  14268=>"00000000",
  14269=>"00000010",
  14270=>"00000000",
  14271=>"11111110",
  14272=>"11111111",
  14273=>"11111110",
  14274=>"11111111",
  14275=>"11111110",
  14276=>"11111110",
  14277=>"00000000",
  14278=>"00000001",
  14279=>"11111110",
  14280=>"11111111",
  14281=>"00000010",
  14282=>"00000001",
  14283=>"00000000",
  14284=>"00000001",
  14285=>"00000010",
  14286=>"00000000",
  14287=>"00000001",
  14288=>"11111110",
  14289=>"00000000",
  14290=>"11111110",
  14291=>"00000010",
  14292=>"00000000",
  14293=>"11111110",
  14294=>"00000001",
  14295=>"11111111",
  14296=>"00000000",
  14297=>"00000000",
  14298=>"00000001",
  14299=>"00000001",
  14300=>"11111111",
  14301=>"11111111",
  14302=>"00000001",
  14303=>"00000001",
  14304=>"00000000",
  14305=>"11111110",
  14306=>"00000001",
  14307=>"00000000",
  14308=>"00000010",
  14309=>"00000001",
  14310=>"00000000",
  14311=>"00000000",
  14312=>"00000000",
  14313=>"11111111",
  14314=>"00000001",
  14315=>"11111111",
  14316=>"11111111",
  14317=>"11111111",
  14318=>"00000010",
  14319=>"00000000",
  14320=>"00000001",
  14321=>"11111110",
  14322=>"11111111",
  14323=>"11111111",
  14324=>"11111110",
  14325=>"00000001",
  14326=>"00000001",
  14327=>"11111111",
  14328=>"00000000",
  14329=>"00000000",
  14330=>"11111111",
  14331=>"00000010",
  14332=>"00000000",
  14333=>"11111111",
  14334=>"00000001",
  14335=>"00000000",
  14336=>"11111111",
  14337=>"00000000",
  14338=>"00000000",
  14339=>"00000000",
  14340=>"00000000",
  14341=>"00000000",
  14342=>"00000000",
  14343=>"00000000",
  14344=>"00000000",
  14345=>"00000000",
  14346=>"00000000",
  14347=>"00000000",
  14348=>"00000000",
  14349=>"00000000",
  14350=>"00000000",
  14351=>"00000000",
  14352=>"00000000",
  14353=>"00000000",
  14354=>"00000000",
  14355=>"00000000",
  14356=>"00000000",
  14357=>"00000000",
  14358=>"00000000",
  14359=>"00000000",
  14360=>"00000000",
  14361=>"00000000",
  14362=>"00000000",
  14363=>"00000000",
  14364=>"00000000",
  14365=>"00000000",
  14366=>"00000000",
  14367=>"00000000",
  14368=>"00000000",
  14369=>"00000000",
  14370=>"00000000",
  14371=>"00000000",
  14372=>"00000000",
  14373=>"00000000",
  14374=>"00000000",
  14375=>"00000000",
  14376=>"00000000",
  14377=>"00000000",
  14378=>"00000000",
  14379=>"00000000",
  14380=>"00000000",
  14381=>"11111111",
  14382=>"11111111",
  14383=>"00000000",
  14384=>"00000000",
  14385=>"00000000",
  14386=>"00000000",
  14387=>"00000000",
  14388=>"00000000",
  14389=>"00000000",
  14390=>"00000000",
  14391=>"00000000",
  14392=>"00000000",
  14393=>"00000000",
  14394=>"00000000",
  14395=>"00000000",
  14396=>"00000000",
  14397=>"00000000",
  14398=>"00000000",
  14399=>"00000000",
  14400=>"00000000",
  14401=>"00000000",
  14402=>"00000000",
  14403=>"00000000",
  14404=>"00000000",
  14405=>"00000000",
  14406=>"00000000",
  14407=>"00000000",
  14408=>"00000000",
  14409=>"00000000",
  14410=>"00000000",
  14411=>"00000000",
  14412=>"00000000",
  14413=>"00000000",
  14414=>"00000000",
  14415=>"00000000",
  14416=>"11111111",
  14417=>"00000000",
  14418=>"00000000",
  14419=>"00000000",
  14420=>"00000000",
  14421=>"00000000",
  14422=>"00000000",
  14423=>"00000000",
  14424=>"00000000",
  14425=>"00000000",
  14426=>"00000000",
  14427=>"00000000",
  14428=>"00000000",
  14429=>"00000000",
  14430=>"00000000",
  14431=>"00000000",
  14432=>"00000000",
  14433=>"00000000",
  14434=>"00000000",
  14435=>"00000000",
  14436=>"00000000",
  14437=>"00000001",
  14438=>"00000000",
  14439=>"11111111",
  14440=>"00000000",
  14441=>"00000000",
  14442=>"00000000",
  14443=>"00000000",
  14444=>"00000000",
  14445=>"00000000",
  14446=>"00000000",
  14447=>"00000000",
  14448=>"00000000",
  14449=>"00000000",
  14450=>"00000000",
  14451=>"00000000",
  14452=>"00000000",
  14453=>"00000000",
  14454=>"00000000",
  14455=>"00000000",
  14456=>"00000000",
  14457=>"00000000",
  14458=>"00000000",
  14459=>"00000000",
  14460=>"00000000",
  14461=>"00000000",
  14462=>"00000000",
  14463=>"00000000",
  14464=>"00000000",
  14465=>"00000000",
  14466=>"11111111",
  14467=>"11111111",
  14468=>"00000000",
  14469=>"00000000",
  14470=>"00000000",
  14471=>"00000000",
  14472=>"00000000",
  14473=>"00000000",
  14474=>"00000000",
  14475=>"00000000",
  14476=>"00000000",
  14477=>"00000001",
  14478=>"00000000",
  14479=>"00000000",
  14480=>"00000000",
  14481=>"00000000",
  14482=>"00000000",
  14483=>"00000000",
  14484=>"00000000",
  14485=>"00000000",
  14486=>"00000000",
  14487=>"00000000",
  14488=>"00000000",
  14489=>"00000000",
  14490=>"00000000",
  14491=>"00000000",
  14492=>"00000000",
  14493=>"00000000",
  14494=>"00000000",
  14495=>"00000000",
  14496=>"11111111",
  14497=>"00000000",
  14498=>"00000000",
  14499=>"00000000",
  14500=>"11111111",
  14501=>"00000000",
  14502=>"00000000",
  14503=>"00000000",
  14504=>"00000000",
  14505=>"00000000",
  14506=>"00000000",
  14507=>"00000000",
  14508=>"00000000",
  14509=>"00000000",
  14510=>"00000000",
  14511=>"00000000",
  14512=>"00000000",
  14513=>"00000000",
  14514=>"00000000",
  14515=>"00000000",
  14516=>"00000000",
  14517=>"00000000",
  14518=>"00000000",
  14519=>"00000000",
  14520=>"00000000",
  14521=>"00000000",
  14522=>"00000000",
  14523=>"00000000",
  14524=>"00000000",
  14525=>"00000000",
  14526=>"00000000",
  14527=>"00000000",
  14528=>"00000000",
  14529=>"00000001",
  14530=>"00000000",
  14531=>"00000000",
  14532=>"00000000",
  14533=>"00000000",
  14534=>"00000000",
  14535=>"00000000",
  14536=>"00000000",
  14537=>"00000000",
  14538=>"11111111",
  14539=>"00000000",
  14540=>"00000000",
  14541=>"00000000",
  14542=>"00000001",
  14543=>"00000000",
  14544=>"00000000",
  14545=>"00000000",
  14546=>"00000000",
  14547=>"00000000",
  14548=>"00000000",
  14549=>"00000000",
  14550=>"00000000",
  14551=>"00000000",
  14552=>"00000001",
  14553=>"00000000",
  14554=>"00000001",
  14555=>"00000000",
  14556=>"00000000",
  14557=>"00000000",
  14558=>"00000000",
  14559=>"00000000",
  14560=>"00000000",
  14561=>"00000000",
  14562=>"00000000",
  14563=>"00000001",
  14564=>"00000000",
  14565=>"00000000",
  14566=>"00000000",
  14567=>"00000000",
  14568=>"00000000",
  14569=>"00000000",
  14570=>"00000001",
  14571=>"00000001",
  14572=>"00000000",
  14573=>"00000000",
  14574=>"00000000",
  14575=>"11111111",
  14576=>"00000000",
  14577=>"00000000",
  14578=>"00000000",
  14579=>"00000000",
  14580=>"00000000",
  14581=>"00000000",
  14582=>"00000001",
  14583=>"00000000",
  14584=>"00000000",
  14585=>"00000000",
  14586=>"00000000",
  14587=>"00000000",
  14588=>"00000001",
  14589=>"00000000",
  14590=>"00000000",
  14591=>"00000000",
  14592=>"00000001",
  14593=>"00000000",
  14594=>"00000000",
  14595=>"00000000",
  14596=>"00000001",
  14597=>"00000000",
  14598=>"00000000",
  14599=>"00000000",
  14600=>"00000001",
  14601=>"00000000",
  14602=>"00000000",
  14603=>"00000000",
  14604=>"00000000",
  14605=>"00000000",
  14606=>"00000000",
  14607=>"00000000",
  14608=>"00000000",
  14609=>"00000000",
  14610=>"00000001",
  14611=>"00000000",
  14612=>"00000000",
  14613=>"00000000",
  14614=>"00000000",
  14615=>"00000000",
  14616=>"00000000",
  14617=>"00000000",
  14618=>"00000000",
  14619=>"11111111",
  14620=>"00000001",
  14621=>"00000000",
  14622=>"00000000",
  14623=>"00000000",
  14624=>"00000000",
  14625=>"11111111",
  14626=>"00000001",
  14627=>"00000000",
  14628=>"00000000",
  14629=>"00000000",
  14630=>"00000000",
  14631=>"00000000",
  14632=>"00000000",
  14633=>"00000000",
  14634=>"00000000",
  14635=>"00000000",
  14636=>"00000000",
  14637=>"00000001",
  14638=>"00000000",
  14639=>"00000000",
  14640=>"00000000",
  14641=>"00000000",
  14642=>"00000000",
  14643=>"00000000",
  14644=>"00000000",
  14645=>"00000000",
  14646=>"00000000",
  14647=>"00000000",
  14648=>"00000000",
  14649=>"00000000",
  14650=>"00000000",
  14651=>"00000000",
  14652=>"00000001",
  14653=>"00000000",
  14654=>"00000000",
  14655=>"00000000",
  14656=>"00000000",
  14657=>"00000000",
  14658=>"00000000",
  14659=>"00000000",
  14660=>"11111111",
  14661=>"00000000",
  14662=>"00000000",
  14663=>"00000000",
  14664=>"00000000",
  14665=>"00000000",
  14666=>"00000000",
  14667=>"00000000",
  14668=>"00000000",
  14669=>"00000000",
  14670=>"00000000",
  14671=>"00000000",
  14672=>"00000000",
  14673=>"00000000",
  14674=>"00000000",
  14675=>"00000000",
  14676=>"00000000",
  14677=>"00000000",
  14678=>"00000000",
  14679=>"00000000",
  14680=>"00000000",
  14681=>"00000000",
  14682=>"00000000",
  14683=>"00000000",
  14684=>"00000000",
  14685=>"00000001",
  14686=>"00000000",
  14687=>"00000000",
  14688=>"00000000",
  14689=>"00000000",
  14690=>"00000000",
  14691=>"00000000",
  14692=>"00000001",
  14693=>"11111111",
  14694=>"00000000",
  14695=>"00000000",
  14696=>"00000000",
  14697=>"00000000",
  14698=>"00000000",
  14699=>"00000000",
  14700=>"00000000",
  14701=>"00000000",
  14702=>"00000000",
  14703=>"00000001",
  14704=>"00000001",
  14705=>"00000000",
  14706=>"11111111",
  14707=>"00000000",
  14708=>"00000000",
  14709=>"00000000",
  14710=>"00000000",
  14711=>"11111111",
  14712=>"00000000",
  14713=>"00000000",
  14714=>"00000000",
  14715=>"00000000",
  14716=>"11111111",
  14717=>"00000000",
  14718=>"00000000",
  14719=>"00000000",
  14720=>"00000000",
  14721=>"11111111",
  14722=>"00000000",
  14723=>"00000000",
  14724=>"00000001",
  14725=>"00000000",
  14726=>"00000000",
  14727=>"00000000",
  14728=>"00000000",
  14729=>"00000000",
  14730=>"00000000",
  14731=>"00000000",
  14732=>"00000000",
  14733=>"00000000",
  14734=>"00000000",
  14735=>"00000000",
  14736=>"00000000",
  14737=>"00000000",
  14738=>"00000000",
  14739=>"00000000",
  14740=>"00000000",
  14741=>"00000000",
  14742=>"00000000",
  14743=>"00000000",
  14744=>"00000000",
  14745=>"00000000",
  14746=>"00000000",
  14747=>"00000000",
  14748=>"00000000",
  14749=>"00000000",
  14750=>"11111111",
  14751=>"00000000",
  14752=>"00000000",
  14753=>"00000000",
  14754=>"11111111",
  14755=>"00000000",
  14756=>"00000000",
  14757=>"00000000",
  14758=>"00000000",
  14759=>"00000000",
  14760=>"00000000",
  14761=>"00000000",
  14762=>"00000000",
  14763=>"00000000",
  14764=>"11111111",
  14765=>"00000000",
  14766=>"11111111",
  14767=>"00000000",
  14768=>"00000000",
  14769=>"00000000",
  14770=>"00000000",
  14771=>"11111111",
  14772=>"00000000",
  14773=>"00000000",
  14774=>"00000000",
  14775=>"00000000",
  14776=>"00000000",
  14777=>"00000000",
  14778=>"00000000",
  14779=>"00000000",
  14780=>"00000000",
  14781=>"00000000",
  14782=>"00000000",
  14783=>"00000000",
  14784=>"00000000",
  14785=>"00000000",
  14786=>"00000000",
  14787=>"00000000",
  14788=>"00000000",
  14789=>"00000000",
  14790=>"00000000",
  14791=>"00000000",
  14792=>"00000000",
  14793=>"00000000",
  14794=>"00000000",
  14795=>"00000000",
  14796=>"00000000",
  14797=>"00000000",
  14798=>"00000000",
  14799=>"00000000",
  14800=>"00000000",
  14801=>"00000000",
  14802=>"00000000",
  14803=>"00000000",
  14804=>"00000000",
  14805=>"00000000",
  14806=>"00000000",
  14807=>"00000000",
  14808=>"00000000",
  14809=>"00000000",
  14810=>"00000000",
  14811=>"00000000",
  14812=>"00000000",
  14813=>"00000000",
  14814=>"00000000",
  14815=>"00000000",
  14816=>"00000000",
  14817=>"00000000",
  14818=>"00000000",
  14819=>"00000000",
  14820=>"00000000",
  14821=>"00000000",
  14822=>"11111111",
  14823=>"00000000",
  14824=>"00000000",
  14825=>"00000000",
  14826=>"00000000",
  14827=>"00000000",
  14828=>"11111111",
  14829=>"00000000",
  14830=>"00000000",
  14831=>"00000000",
  14832=>"00000001",
  14833=>"00000000",
  14834=>"00000001",
  14835=>"00000000",
  14836=>"00000000",
  14837=>"00000000",
  14838=>"00000000",
  14839=>"00000000",
  14840=>"00000000",
  14841=>"00000000",
  14842=>"00000000",
  14843=>"00000000",
  14844=>"00000000",
  14845=>"00000000",
  14846=>"00000000",
  14847=>"00000000",
  14848=>"00000001",
  14849=>"00000000",
  14850=>"00000000",
  14851=>"00000000",
  14852=>"00000000",
  14853=>"00000000",
  14854=>"00000000",
  14855=>"00000000",
  14856=>"00000000",
  14857=>"00000000",
  14858=>"00000000",
  14859=>"00000000",
  14860=>"00000000",
  14861=>"11111111",
  14862=>"00000000",
  14863=>"00000000",
  14864=>"00000000",
  14865=>"00000000",
  14866=>"00000000",
  14867=>"00000000",
  14868=>"00000000",
  14869=>"00000000",
  14870=>"00000000",
  14871=>"00000000",
  14872=>"00000000",
  14873=>"00000000",
  14874=>"00000000",
  14875=>"00000000",
  14876=>"00000000",
  14877=>"00000000",
  14878=>"00000000",
  14879=>"00000000",
  14880=>"00000000",
  14881=>"00000000",
  14882=>"11111111",
  14883=>"00000000",
  14884=>"00000000",
  14885=>"00000000",
  14886=>"00000000",
  14887=>"00000000",
  14888=>"00000000",
  14889=>"00000001",
  14890=>"00000000",
  14891=>"00000000",
  14892=>"00000000",
  14893=>"00000000",
  14894=>"00000000",
  14895=>"11111111",
  14896=>"00000000",
  14897=>"00000000",
  14898=>"00000000",
  14899=>"11111111",
  14900=>"00000000",
  14901=>"00000000",
  14902=>"00000001",
  14903=>"00000000",
  14904=>"00000000",
  14905=>"00000000",
  14906=>"00000000",
  14907=>"00000000",
  14908=>"00000000",
  14909=>"00000000",
  14910=>"00000000",
  14911=>"00000000",
  14912=>"00000000",
  14913=>"00000000",
  14914=>"00000000",
  14915=>"00000000",
  14916=>"00000000",
  14917=>"00000000",
  14918=>"00000000",
  14919=>"00000000",
  14920=>"00000000",
  14921=>"00000000",
  14922=>"00000000",
  14923=>"00000000",
  14924=>"00000000",
  14925=>"00000000",
  14926=>"00000000",
  14927=>"00000000",
  14928=>"00000000",
  14929=>"00000000",
  14930=>"00000000",
  14931=>"00000000",
  14932=>"00000000",
  14933=>"00000000",
  14934=>"00000000",
  14935=>"00000000",
  14936=>"00000000",
  14937=>"00000000",
  14938=>"00000000",
  14939=>"00000000",
  14940=>"00000000",
  14941=>"00000000",
  14942=>"00000000",
  14943=>"00000000",
  14944=>"00000000",
  14945=>"00000000",
  14946=>"00000001",
  14947=>"00000000",
  14948=>"00000000",
  14949=>"00000000",
  14950=>"00000001",
  14951=>"00000000",
  14952=>"00000000",
  14953=>"00000000",
  14954=>"00000000",
  14955=>"00000000",
  14956=>"00000000",
  14957=>"00000000",
  14958=>"00000000",
  14959=>"00000000",
  14960=>"00000000",
  14961=>"00000000",
  14962=>"00000000",
  14963=>"00000000",
  14964=>"00000000",
  14965=>"00000000",
  14966=>"00000000",
  14967=>"00000000",
  14968=>"00000000",
  14969=>"00000000",
  14970=>"00000000",
  14971=>"00000000",
  14972=>"00000001",
  14973=>"00000000",
  14974=>"00000000",
  14975=>"00000000",
  14976=>"00000000",
  14977=>"11111111",
  14978=>"00000000",
  14979=>"00000000",
  14980=>"00000000",
  14981=>"00000000",
  14982=>"00000000",
  14983=>"00000000",
  14984=>"00000000",
  14985=>"00000000",
  14986=>"00000000",
  14987=>"00000000",
  14988=>"00000000",
  14989=>"00000000",
  14990=>"00000000",
  14991=>"00000000",
  14992=>"00000000",
  14993=>"00000000",
  14994=>"00000000",
  14995=>"00000000",
  14996=>"00000000",
  14997=>"00000000",
  14998=>"00000001",
  14999=>"00000000",
  15000=>"00000000",
  15001=>"00000000",
  15002=>"11111111",
  15003=>"00000001",
  15004=>"00000000",
  15005=>"00000000",
  15006=>"00000000",
  15007=>"00000000",
  15008=>"00000000",
  15009=>"00000000",
  15010=>"00000000",
  15011=>"00000000",
  15012=>"00000000",
  15013=>"00000000",
  15014=>"00000000",
  15015=>"00000000",
  15016=>"00000000",
  15017=>"00000000",
  15018=>"00000000",
  15019=>"00000000",
  15020=>"00000000",
  15021=>"00000000",
  15022=>"00000000",
  15023=>"00000000",
  15024=>"00000000",
  15025=>"00000000",
  15026=>"00000000",
  15027=>"00000000",
  15028=>"00000000",
  15029=>"00000000",
  15030=>"00000001",
  15031=>"00000000",
  15032=>"00000000",
  15033=>"00000000",
  15034=>"00000001",
  15035=>"00000000",
  15036=>"00000000",
  15037=>"00000000",
  15038=>"00000000",
  15039=>"00000000",
  15040=>"00000000",
  15041=>"00000000",
  15042=>"00000000",
  15043=>"00000000",
  15044=>"00000000",
  15045=>"00000000",
  15046=>"00000000",
  15047=>"00000001",
  15048=>"00000000",
  15049=>"00000000",
  15050=>"00000000",
  15051=>"00000000",
  15052=>"00000000",
  15053=>"00000000",
  15054=>"00000000",
  15055=>"00000000",
  15056=>"00000000",
  15057=>"00000000",
  15058=>"00000000",
  15059=>"00000000",
  15060=>"00000000",
  15061=>"00000000",
  15062=>"00000000",
  15063=>"00000000",
  15064=>"00000000",
  15065=>"00000000",
  15066=>"00000001",
  15067=>"00000000",
  15068=>"00000000",
  15069=>"00000000",
  15070=>"00000000",
  15071=>"00000000",
  15072=>"00000000",
  15073=>"00000000",
  15074=>"00000000",
  15075=>"00000000",
  15076=>"00000000",
  15077=>"11111111",
  15078=>"00000000",
  15079=>"00000000",
  15080=>"00000000",
  15081=>"00000000",
  15082=>"00000000",
  15083=>"00000000",
  15084=>"00000000",
  15085=>"00000000",
  15086=>"00000000",
  15087=>"00000000",
  15088=>"00000000",
  15089=>"00000000",
  15090=>"00000000",
  15091=>"00000000",
  15092=>"00000000",
  15093=>"00000000",
  15094=>"00000000",
  15095=>"00000000",
  15096=>"00000000",
  15097=>"00000000",
  15098=>"00000000",
  15099=>"00000000",
  15100=>"00000000",
  15101=>"00000000",
  15102=>"00000000",
  15103=>"00000001",
  15104=>"00000000",
  15105=>"00000000",
  15106=>"00000000",
  15107=>"00000000",
  15108=>"00000000",
  15109=>"00000000",
  15110=>"00000001",
  15111=>"00000000",
  15112=>"00000000",
  15113=>"00000000",
  15114=>"00000000",
  15115=>"00000000",
  15116=>"00000000",
  15117=>"00000000",
  15118=>"00000000",
  15119=>"00000000",
  15120=>"00000000",
  15121=>"00000000",
  15122=>"00000000",
  15123=>"00000000",
  15124=>"00000001",
  15125=>"11111111",
  15126=>"00000000",
  15127=>"00000000",
  15128=>"00000000",
  15129=>"00000000",
  15130=>"00000000",
  15131=>"00000000",
  15132=>"00000000",
  15133=>"00000000",
  15134=>"00000000",
  15135=>"00000000",
  15136=>"00000000",
  15137=>"00000000",
  15138=>"00000000",
  15139=>"00000000",
  15140=>"00000000",
  15141=>"00000000",
  15142=>"00000000",
  15143=>"00000000",
  15144=>"00000000",
  15145=>"00000000",
  15146=>"00000000",
  15147=>"00000000",
  15148=>"00000000",
  15149=>"00000000",
  15150=>"00000000",
  15151=>"11111111",
  15152=>"00000000",
  15153=>"00000000",
  15154=>"00000000",
  15155=>"00000000",
  15156=>"00000000",
  15157=>"00000000",
  15158=>"00000000",
  15159=>"00000000",
  15160=>"00000000",
  15161=>"00000001",
  15162=>"11111111",
  15163=>"00000000",
  15164=>"00000000",
  15165=>"00000000",
  15166=>"00000000",
  15167=>"00000000",
  15168=>"00000000",
  15169=>"00000000",
  15170=>"00000000",
  15171=>"00000000",
  15172=>"00000000",
  15173=>"00000000",
  15174=>"00000000",
  15175=>"00000000",
  15176=>"00000000",
  15177=>"00000000",
  15178=>"00000000",
  15179=>"00000000",
  15180=>"00000001",
  15181=>"00000000",
  15182=>"00000000",
  15183=>"00000001",
  15184=>"00000000",
  15185=>"00000000",
  15186=>"00000000",
  15187=>"00000000",
  15188=>"00000000",
  15189=>"00000000",
  15190=>"00000000",
  15191=>"00000000",
  15192=>"00000000",
  15193=>"00000000",
  15194=>"00000000",
  15195=>"00000000",
  15196=>"00000000",
  15197=>"00000000",
  15198=>"00000000",
  15199=>"00000000",
  15200=>"00000000",
  15201=>"00000000",
  15202=>"00000000",
  15203=>"00000000",
  15204=>"00000001",
  15205=>"00000000",
  15206=>"00000000",
  15207=>"00000000",
  15208=>"00000000",
  15209=>"00000000",
  15210=>"00000000",
  15211=>"00000000",
  15212=>"00000000",
  15213=>"00000000",
  15214=>"00000000",
  15215=>"00000000",
  15216=>"00000000",
  15217=>"00000000",
  15218=>"00000000",
  15219=>"00000000",
  15220=>"00000000",
  15221=>"00000000",
  15222=>"00000000",
  15223=>"00000000",
  15224=>"00000000",
  15225=>"00000000",
  15226=>"00000000",
  15227=>"00000000",
  15228=>"00000000",
  15229=>"00000000",
  15230=>"00000000",
  15231=>"00000000",
  15232=>"11111111",
  15233=>"00000000",
  15234=>"00000000",
  15235=>"00000000",
  15236=>"00000000",
  15237=>"00000000",
  15238=>"00000000",
  15239=>"00000000",
  15240=>"00000000",
  15241=>"00000000",
  15242=>"00000001",
  15243=>"00000000",
  15244=>"00000000",
  15245=>"00000000",
  15246=>"00000000",
  15247=>"00000000",
  15248=>"00000000",
  15249=>"00000001",
  15250=>"00000000",
  15251=>"00000000",
  15252=>"00000000",
  15253=>"00000000",
  15254=>"00000000",
  15255=>"00000000",
  15256=>"00000000",
  15257=>"00000000",
  15258=>"00000000",
  15259=>"00000000",
  15260=>"00000000",
  15261=>"00000000",
  15262=>"00000000",
  15263=>"11111111",
  15264=>"00000000",
  15265=>"00000000",
  15266=>"00000000",
  15267=>"00000000",
  15268=>"00000000",
  15269=>"00000000",
  15270=>"00000000",
  15271=>"00000000",
  15272=>"00000000",
  15273=>"00000000",
  15274=>"00000000",
  15275=>"00000000",
  15276=>"00000000",
  15277=>"00000000",
  15278=>"00000000",
  15279=>"00000000",
  15280=>"00000000",
  15281=>"00000000",
  15282=>"00000000",
  15283=>"00000000",
  15284=>"00000001",
  15285=>"00000000",
  15286=>"00000000",
  15287=>"00000000",
  15288=>"00000000",
  15289=>"00000000",
  15290=>"00000000",
  15291=>"11111111",
  15292=>"00000000",
  15293=>"00000000",
  15294=>"00000000",
  15295=>"00000000",
  15296=>"00000000",
  15297=>"00000000",
  15298=>"00000000",
  15299=>"00000000",
  15300=>"00000000",
  15301=>"00000000",
  15302=>"00000000",
  15303=>"00000000",
  15304=>"00000000",
  15305=>"00000000",
  15306=>"00000000",
  15307=>"00000000",
  15308=>"00000000",
  15309=>"00000000",
  15310=>"00000000",
  15311=>"00000000",
  15312=>"00000000",
  15313=>"00000000",
  15314=>"00000000",
  15315=>"00000000",
  15316=>"00000000",
  15317=>"00000000",
  15318=>"00000000",
  15319=>"00000000",
  15320=>"00000000",
  15321=>"00000000",
  15322=>"00000000",
  15323=>"00000000",
  15324=>"00000000",
  15325=>"00000000",
  15326=>"00000000",
  15327=>"00000000",
  15328=>"00000000",
  15329=>"00000000",
  15330=>"00000000",
  15331=>"00000000",
  15332=>"00000000",
  15333=>"00000000",
  15334=>"00000000",
  15335=>"00000000",
  15336=>"00000000",
  15337=>"00000000",
  15338=>"00000000",
  15339=>"00000000",
  15340=>"00000000",
  15341=>"11111111",
  15342=>"00000000",
  15343=>"00000000",
  15344=>"00000000",
  15345=>"00000000",
  15346=>"00000000",
  15347=>"00000000",
  15348=>"00000000",
  15349=>"00000000",
  15350=>"00000000",
  15351=>"00000000",
  15352=>"00000000",
  15353=>"00000000",
  15354=>"00000000",
  15355=>"00000000",
  15356=>"00000000",
  15357=>"00000000",
  15358=>"00000000",
  15359=>"00000000",
  15360=>"00000000",
  15361=>"00000000",
  15362=>"00000001",
  15363=>"00000000",
  15364=>"00000000",
  15365=>"00000000",
  15366=>"00000000",
  15367=>"00000000",
  15368=>"00000000",
  15369=>"00000000",
  15370=>"11111111",
  15371=>"11111111",
  15372=>"00000001",
  15373=>"00000000",
  15374=>"00000000",
  15375=>"00000000",
  15376=>"00000000",
  15377=>"00000000",
  15378=>"00000000",
  15379=>"00000000",
  15380=>"00000000",
  15381=>"00000001",
  15382=>"00000000",
  15383=>"00000000",
  15384=>"00000000",
  15385=>"00000000",
  15386=>"00000000",
  15387=>"00000000",
  15388=>"00000000",
  15389=>"11111111",
  15390=>"00000000",
  15391=>"00000000",
  15392=>"00000000",
  15393=>"00000000",
  15394=>"00000000",
  15395=>"00000000",
  15396=>"00000000",
  15397=>"00000000",
  15398=>"00000000",
  15399=>"00000000",
  15400=>"00000000",
  15401=>"00000000",
  15402=>"00000000",
  15403=>"00000000",
  15404=>"00000000",
  15405=>"00000000",
  15406=>"00000000",
  15407=>"00000000",
  15408=>"00000000",
  15409=>"00000000",
  15410=>"00000000",
  15411=>"00000000",
  15412=>"00000000",
  15413=>"00000000",
  15414=>"11111110",
  15415=>"00000001",
  15416=>"00000000",
  15417=>"00000000",
  15418=>"00000000",
  15419=>"00000000",
  15420=>"00000001",
  15421=>"00000000",
  15422=>"00000000",
  15423=>"00000001",
  15424=>"00000000",
  15425=>"00000000",
  15426=>"00000000",
  15427=>"00000000",
  15428=>"00000000",
  15429=>"00000001",
  15430=>"00000000",
  15431=>"00000000",
  15432=>"00000001",
  15433=>"00000000",
  15434=>"00000000",
  15435=>"00000000",
  15436=>"00000000",
  15437=>"00000000",
  15438=>"00000000",
  15439=>"00000001",
  15440=>"00000000",
  15441=>"00000000",
  15442=>"00000000",
  15443=>"00000000",
  15444=>"00000000",
  15445=>"00000000",
  15446=>"00000000",
  15447=>"00000000",
  15448=>"00000000",
  15449=>"00000000",
  15450=>"00000000",
  15451=>"00000000",
  15452=>"00000000",
  15453=>"00000000",
  15454=>"00000000",
  15455=>"00000000",
  15456=>"00000000",
  15457=>"00000001",
  15458=>"00000000",
  15459=>"00000000",
  15460=>"00000000",
  15461=>"00000000",
  15462=>"00000000",
  15463=>"00000000",
  15464=>"00000000",
  15465=>"00000000",
  15466=>"00000000",
  15467=>"00000000",
  15468=>"00000000",
  15469=>"00000000",
  15470=>"00000000",
  15471=>"00000000",
  15472=>"00000000",
  15473=>"00000001",
  15474=>"00000000",
  15475=>"00000000",
  15476=>"00000000",
  15477=>"00000000",
  15478=>"00000000",
  15479=>"00000000",
  15480=>"00000000",
  15481=>"00000000",
  15482=>"00000000",
  15483=>"00000000",
  15484=>"00000000",
  15485=>"11111111",
  15486=>"00000000",
  15487=>"00000000",
  15488=>"00000000",
  15489=>"00000000",
  15490=>"00000000",
  15491=>"00000000",
  15492=>"00000000",
  15493=>"00000000",
  15494=>"00000000",
  15495=>"00000000",
  15496=>"00000000",
  15497=>"00000000",
  15498=>"00000000",
  15499=>"00000001",
  15500=>"00000000",
  15501=>"00000000",
  15502=>"00000000",
  15503=>"00000000",
  15504=>"00000000",
  15505=>"00000000",
  15506=>"11111111",
  15507=>"00000000",
  15508=>"00000000",
  15509=>"00000000",
  15510=>"00000000",
  15511=>"00000000",
  15512=>"00000000",
  15513=>"00000000",
  15514=>"00000000",
  15515=>"00000000",
  15516=>"11111111",
  15517=>"00000000",
  15518=>"00000000",
  15519=>"00000000",
  15520=>"11111111",
  15521=>"11111111",
  15522=>"00000000",
  15523=>"00000000",
  15524=>"11111111",
  15525=>"00000000",
  15526=>"00000000",
  15527=>"00000000",
  15528=>"00000000",
  15529=>"00000000",
  15530=>"00000000",
  15531=>"00000000",
  15532=>"00000000",
  15533=>"00000000",
  15534=>"11111111",
  15535=>"00000000",
  15536=>"00000000",
  15537=>"00000000",
  15538=>"00000001",
  15539=>"00000001",
  15540=>"00000000",
  15541=>"00000000",
  15542=>"00000000",
  15543=>"00000000",
  15544=>"00000000",
  15545=>"00000000",
  15546=>"00000000",
  15547=>"00000000",
  15548=>"00000000",
  15549=>"11111011",
  15550=>"00000000",
  15551=>"00000000",
  15552=>"00000000",
  15553=>"11111110",
  15554=>"00000001",
  15555=>"00000000",
  15556=>"00000000",
  15557=>"00000000",
  15558=>"00000000",
  15559=>"00000001",
  15560=>"00000000",
  15561=>"00000000",
  15562=>"00000000",
  15563=>"00000000",
  15564=>"00000000",
  15565=>"00000000",
  15566=>"11111110",
  15567=>"00000000",
  15568=>"00000000",
  15569=>"00000000",
  15570=>"11111110",
  15571=>"00000000",
  15572=>"00000001",
  15573=>"00000000",
  15574=>"00000001",
  15575=>"00000000",
  15576=>"00000001",
  15577=>"11111111",
  15578=>"00000001",
  15579=>"11111111",
  15580=>"00000000",
  15581=>"00000000",
  15582=>"00000000",
  15583=>"00000000",
  15584=>"00000001",
  15585=>"00000000",
  15586=>"00000000",
  15587=>"00000000",
  15588=>"00000000",
  15589=>"11111111",
  15590=>"00000000",
  15591=>"00000000",
  15592=>"00000000",
  15593=>"00000000",
  15594=>"00000001",
  15595=>"11111110",
  15596=>"11111111",
  15597=>"00000001",
  15598=>"00000000",
  15599=>"00000000",
  15600=>"00000000",
  15601=>"00000000",
  15602=>"00000000",
  15603=>"00000000",
  15604=>"00000000",
  15605=>"00000000",
  15606=>"00000000",
  15607=>"00000000",
  15608=>"00000000",
  15609=>"00000000",
  15610=>"00000000",
  15611=>"00000000",
  15612=>"00000000",
  15613=>"00000000",
  15614=>"00000000",
  15615=>"00000000",
  15616=>"00000000",
  15617=>"00000000",
  15618=>"00000000",
  15619=>"00000000",
  15620=>"11111100",
  15621=>"00000000",
  15622=>"00000000",
  15623=>"00000000",
  15624=>"11111110",
  15625=>"00000001",
  15626=>"00000000",
  15627=>"00000000",
  15628=>"00000001",
  15629=>"00000000",
  15630=>"11111111",
  15631=>"00000000",
  15632=>"00000000",
  15633=>"00000000",
  15634=>"00000000",
  15635=>"00000000",
  15636=>"00000000",
  15637=>"11111111",
  15638=>"11111110",
  15639=>"00000000",
  15640=>"00000000",
  15641=>"00000000",
  15642=>"00000000",
  15643=>"00000000",
  15644=>"00000000",
  15645=>"00000000",
  15646=>"00000000",
  15647=>"00000000",
  15648=>"00000000",
  15649=>"00000000",
  15650=>"11111101",
  15651=>"00000000",
  15652=>"00000000",
  15653=>"00000000",
  15654=>"00000000",
  15655=>"00000000",
  15656=>"00000000",
  15657=>"00000000",
  15658=>"00000000",
  15659=>"00000000",
  15660=>"00000000",
  15661=>"00000000",
  15662=>"00000000",
  15663=>"00000000",
  15664=>"11111111",
  15665=>"11111111",
  15666=>"00000000",
  15667=>"00000000",
  15668=>"00000000",
  15669=>"00000000",
  15670=>"00000000",
  15671=>"11111111",
  15672=>"00000000",
  15673=>"11111111",
  15674=>"00000000",
  15675=>"00000001",
  15676=>"00000000",
  15677=>"11111111",
  15678=>"00000000",
  15679=>"11111110",
  15680=>"11111111",
  15681=>"00000000",
  15682=>"00000000",
  15683=>"00000001",
  15684=>"00000000",
  15685=>"00000000",
  15686=>"00000000",
  15687=>"00000000",
  15688=>"00000000",
  15689=>"00000000",
  15690=>"00000000",
  15691=>"11111111",
  15692=>"00000000",
  15693=>"11111111",
  15694=>"00000000",
  15695=>"00000000",
  15696=>"00000000",
  15697=>"00000000",
  15698=>"00000000",
  15699=>"00000000",
  15700=>"11111110",
  15701=>"00000000",
  15702=>"00000000",
  15703=>"00000000",
  15704=>"00000000",
  15705=>"00000000",
  15706=>"00000000",
  15707=>"00000000",
  15708=>"00000000",
  15709=>"11111111",
  15710=>"00000000",
  15711=>"11111111",
  15712=>"00000000",
  15713=>"00000000",
  15714=>"00000000",
  15715=>"00000000",
  15716=>"00000000",
  15717=>"00000000",
  15718=>"00000000",
  15719=>"00000000",
  15720=>"11111111",
  15721=>"00000000",
  15722=>"00000000",
  15723=>"00000000",
  15724=>"00000000",
  15725=>"00000000",
  15726=>"00000000",
  15727=>"11111111",
  15728=>"00000001",
  15729=>"00000000",
  15730=>"00000000",
  15731=>"00000000",
  15732=>"00000000",
  15733=>"00000000",
  15734=>"00000000",
  15735=>"11111111",
  15736=>"00000000",
  15737=>"00000000",
  15738=>"00000000",
  15739=>"00000000",
  15740=>"00000000",
  15741=>"00000000",
  15742=>"00000000",
  15743=>"00000000",
  15744=>"00000000",
  15745=>"00000000",
  15746=>"00000000",
  15747=>"00000000",
  15748=>"00000000",
  15749=>"00000000",
  15750=>"00000000",
  15751=>"00000001",
  15752=>"00000000",
  15753=>"00000000",
  15754=>"00000000",
  15755=>"00000001",
  15756=>"00000000",
  15757=>"11111111",
  15758=>"00000000",
  15759=>"00000000",
  15760=>"00000000",
  15761=>"00000000",
  15762=>"00000000",
  15763=>"00000000",
  15764=>"00000000",
  15765=>"00000000",
  15766=>"00000000",
  15767=>"00000000",
  15768=>"00000001",
  15769=>"00000000",
  15770=>"00000000",
  15771=>"00000000",
  15772=>"00000000",
  15773=>"00000000",
  15774=>"00000000",
  15775=>"00000000",
  15776=>"00000000",
  15777=>"00000001",
  15778=>"00000000",
  15779=>"00000000",
  15780=>"11111111",
  15781=>"00000000",
  15782=>"00000000",
  15783=>"00000000",
  15784=>"00000001",
  15785=>"00000000",
  15786=>"00000000",
  15787=>"00000000",
  15788=>"00000000",
  15789=>"00000000",
  15790=>"00000000",
  15791=>"00000000",
  15792=>"00000000",
  15793=>"00000000",
  15794=>"00000000",
  15795=>"00000000",
  15796=>"00000000",
  15797=>"00000000",
  15798=>"00000000",
  15799=>"00000000",
  15800=>"00000000",
  15801=>"00000000",
  15802=>"00000000",
  15803=>"00000000",
  15804=>"00000000",
  15805=>"00000000",
  15806=>"00000000",
  15807=>"00000000",
  15808=>"00000000",
  15809=>"00000000",
  15810=>"00000000",
  15811=>"00000000",
  15812=>"00000000",
  15813=>"00000000",
  15814=>"00000000",
  15815=>"00000000",
  15816=>"00000000",
  15817=>"00000000",
  15818=>"00000000",
  15819=>"00000000",
  15820=>"00000000",
  15821=>"00000000",
  15822=>"00000000",
  15823=>"00000000",
  15824=>"00000000",
  15825=>"00000000",
  15826=>"00000000",
  15827=>"00000000",
  15828=>"00000000",
  15829=>"00000000",
  15830=>"00000000",
  15831=>"00000000",
  15832=>"00000000",
  15833=>"00000000",
  15834=>"00000000",
  15835=>"00000000",
  15836=>"00000000",
  15837=>"00000001",
  15838=>"00000001",
  15839=>"00000000",
  15840=>"00000000",
  15841=>"00000000",
  15842=>"00000000",
  15843=>"00000000",
  15844=>"00000000",
  15845=>"00000000",
  15846=>"00000001",
  15847=>"00000001",
  15848=>"00000000",
  15849=>"00000000",
  15850=>"00000000",
  15851=>"00000000",
  15852=>"00000000",
  15853=>"00000000",
  15854=>"00000000",
  15855=>"00000000",
  15856=>"11111111",
  15857=>"00000000",
  15858=>"11111111",
  15859=>"00000000",
  15860=>"00000001",
  15861=>"00000000",
  15862=>"00000000",
  15863=>"00000000",
  15864=>"11111111",
  15865=>"00000000",
  15866=>"00000000",
  15867=>"00000000",
  15868=>"00000000",
  15869=>"00000000",
  15870=>"00000000",
  15871=>"11111111",
  15872=>"11111111",
  15873=>"00000000",
  15874=>"00000000",
  15875=>"00000000",
  15876=>"00000000",
  15877=>"00000000",
  15878=>"00000000",
  15879=>"00000000",
  15880=>"00000000",
  15881=>"00000000",
  15882=>"00000001",
  15883=>"11111111",
  15884=>"00000000",
  15885=>"00000001",
  15886=>"00000000",
  15887=>"00000000",
  15888=>"00000000",
  15889=>"00000000",
  15890=>"00000000",
  15891=>"00000000",
  15892=>"00000000",
  15893=>"00000000",
  15894=>"00000000",
  15895=>"00000000",
  15896=>"11111111",
  15897=>"11111111",
  15898=>"00000000",
  15899=>"00000000",
  15900=>"00000000",
  15901=>"00000000",
  15902=>"00000000",
  15903=>"00000000",
  15904=>"00000000",
  15905=>"11111111",
  15906=>"00000000",
  15907=>"00000000",
  15908=>"00000000",
  15909=>"00000000",
  15910=>"00000000",
  15911=>"00000000",
  15912=>"11111111",
  15913=>"00000001",
  15914=>"00000000",
  15915=>"00000000",
  15916=>"00000000",
  15917=>"00000000",
  15918=>"00000000",
  15919=>"00000000",
  15920=>"00000000",
  15921=>"00000000",
  15922=>"00000000",
  15923=>"00000001",
  15924=>"00000000",
  15925=>"00000000",
  15926=>"00000000",
  15927=>"00000000",
  15928=>"11111111",
  15929=>"00000000",
  15930=>"00000000",
  15931=>"00000000",
  15932=>"11111111",
  15933=>"00000000",
  15934=>"00000000",
  15935=>"00000000",
  15936=>"00000000",
  15937=>"00000000",
  15938=>"11111111",
  15939=>"00000000",
  15940=>"00000000",
  15941=>"00000001",
  15942=>"00000000",
  15943=>"00000000",
  15944=>"00000000",
  15945=>"11111111",
  15946=>"00000000",
  15947=>"00000000",
  15948=>"00000000",
  15949=>"00000000",
  15950=>"00000000",
  15951=>"00000000",
  15952=>"00000000",
  15953=>"00000000",
  15954=>"00000000",
  15955=>"00000001",
  15956=>"11111111",
  15957=>"00000000",
  15958=>"00000000",
  15959=>"00000000",
  15960=>"00000000",
  15961=>"00000000",
  15962=>"00000001",
  15963=>"00000000",
  15964=>"00000000",
  15965=>"00000000",
  15966=>"00000000",
  15967=>"00000000",
  15968=>"00000000",
  15969=>"00000000",
  15970=>"00000000",
  15971=>"00000001",
  15972=>"00000000",
  15973=>"00000001",
  15974=>"00000000",
  15975=>"00000000",
  15976=>"00000000",
  15977=>"00000000",
  15978=>"00000000",
  15979=>"00000000",
  15980=>"00000000",
  15981=>"00000000",
  15982=>"00000000",
  15983=>"00000000",
  15984=>"00000000",
  15985=>"00000000",
  15986=>"00000000",
  15987=>"00000000",
  15988=>"00000000",
  15989=>"00000000",
  15990=>"00000000",
  15991=>"00000000",
  15992=>"00000000",
  15993=>"11111111",
  15994=>"00000000",
  15995=>"00000000",
  15996=>"00000000",
  15997=>"00000001",
  15998=>"00000000",
  15999=>"00000000",
  16000=>"11111111",
  16001=>"00000000",
  16002=>"00000000",
  16003=>"00000000",
  16004=>"00000000",
  16005=>"00000000",
  16006=>"00000000",
  16007=>"11111111",
  16008=>"00000000",
  16009=>"00000000",
  16010=>"11111111",
  16011=>"00000000",
  16012=>"00000001",
  16013=>"11111111",
  16014=>"00000001",
  16015=>"00000000",
  16016=>"00000000",
  16017=>"00000000",
  16018=>"00000000",
  16019=>"11111111",
  16020=>"00000000",
  16021=>"00000000",
  16022=>"00000000",
  16023=>"00000000",
  16024=>"00000000",
  16025=>"00000000",
  16026=>"00000000",
  16027=>"00000000",
  16028=>"00000000",
  16029=>"00000000",
  16030=>"00000000",
  16031=>"00000000",
  16032=>"11111111",
  16033=>"00000000",
  16034=>"00000000",
  16035=>"00000000",
  16036=>"00000000",
  16037=>"00000000",
  16038=>"00000000",
  16039=>"00000000",
  16040=>"00000000",
  16041=>"00000000",
  16042=>"00000000",
  16043=>"00000000",
  16044=>"00000000",
  16045=>"00000000",
  16046=>"00000000",
  16047=>"00000000",
  16048=>"00000000",
  16049=>"00000000",
  16050=>"00000000",
  16051=>"00000000",
  16052=>"11111111",
  16053=>"00000000",
  16054=>"00000000",
  16055=>"00000000",
  16056=>"00000000",
  16057=>"00000000",
  16058=>"11111111",
  16059=>"00000000",
  16060=>"00000000",
  16061=>"00000000",
  16062=>"00000000",
  16063=>"11111111",
  16064=>"00000000",
  16065=>"00000000",
  16066=>"00000000",
  16067=>"11111111",
  16068=>"00000000",
  16069=>"00000000",
  16070=>"00000000",
  16071=>"00000000",
  16072=>"00000000",
  16073=>"00000000",
  16074=>"00000000",
  16075=>"00000000",
  16076=>"00000001",
  16077=>"00000000",
  16078=>"00000000",
  16079=>"00000000",
  16080=>"11111110",
  16081=>"00000000",
  16082=>"00000000",
  16083=>"00000000",
  16084=>"00000000",
  16085=>"00000000",
  16086=>"00000000",
  16087=>"00000000",
  16088=>"00000000",
  16089=>"00000000",
  16090=>"00000001",
  16091=>"00000000",
  16092=>"00000000",
  16093=>"11111110",
  16094=>"11111111",
  16095=>"00000000",
  16096=>"00000001",
  16097=>"00000000",
  16098=>"00000000",
  16099=>"00000001",
  16100=>"00000000",
  16101=>"00000000",
  16102=>"00000000",
  16103=>"00000000",
  16104=>"00000000",
  16105=>"00000000",
  16106=>"00000000",
  16107=>"11111111",
  16108=>"11111111",
  16109=>"00000000",
  16110=>"00000000",
  16111=>"00000000",
  16112=>"00000000",
  16113=>"00000000",
  16114=>"11111111",
  16115=>"11111111",
  16116=>"00000000",
  16117=>"00000000",
  16118=>"00000000",
  16119=>"00000000",
  16120=>"00000000",
  16121=>"00000000",
  16122=>"00000000",
  16123=>"00000000",
  16124=>"00000000",
  16125=>"00000000",
  16126=>"00000000",
  16127=>"00000000",
  16128=>"00000000",
  16129=>"00000000",
  16130=>"00000000",
  16131=>"00000000",
  16132=>"00000000",
  16133=>"00000000",
  16134=>"00000000",
  16135=>"00000000",
  16136=>"00000000",
  16137=>"00000000",
  16138=>"00000001",
  16139=>"00000000",
  16140=>"00000000",
  16141=>"00000000",
  16142=>"00000000",
  16143=>"00000000",
  16144=>"00000000",
  16145=>"11111111",
  16146=>"00000000",
  16147=>"00000000",
  16148=>"00000000",
  16149=>"00000000",
  16150=>"00000000",
  16151=>"00000000",
  16152=>"00000000",
  16153=>"00000000",
  16154=>"00000000",
  16155=>"00000000",
  16156=>"00000000",
  16157=>"00000000",
  16158=>"00000000",
  16159=>"00000000",
  16160=>"00000000",
  16161=>"00000000",
  16162=>"11111111",
  16163=>"00000000",
  16164=>"00000000",
  16165=>"00000000",
  16166=>"00000000",
  16167=>"11111111",
  16168=>"00000000",
  16169=>"00000000",
  16170=>"00000000",
  16171=>"11111111",
  16172=>"00000000",
  16173=>"00000001",
  16174=>"00000000",
  16175=>"00000000",
  16176=>"00000000",
  16177=>"00000000",
  16178=>"00000000",
  16179=>"00000000",
  16180=>"00000010",
  16181=>"00000000",
  16182=>"00000001",
  16183=>"00000000",
  16184=>"00000000",
  16185=>"11111111",
  16186=>"11111111",
  16187=>"00000000",
  16188=>"00000000",
  16189=>"00000000",
  16190=>"00000000",
  16191=>"00000000",
  16192=>"00000000",
  16193=>"00000000",
  16194=>"00000000",
  16195=>"00000000",
  16196=>"00000000",
  16197=>"00000000",
  16198=>"00000000",
  16199=>"00000000",
  16200=>"00000000",
  16201=>"00000000",
  16202=>"00000000",
  16203=>"00000000",
  16204=>"00000000",
  16205=>"00000000",
  16206=>"00000000",
  16207=>"00000000",
  16208=>"00000000",
  16209=>"00000000",
  16210=>"00000000",
  16211=>"00000000",
  16212=>"00000000",
  16213=>"00000000",
  16214=>"00000000",
  16215=>"00000000",
  16216=>"00000000",
  16217=>"00000000",
  16218=>"00000001",
  16219=>"00000000",
  16220=>"00000000",
  16221=>"00000000",
  16222=>"00000000",
  16223=>"00000000",
  16224=>"00000000",
  16225=>"00000000",
  16226=>"00000000",
  16227=>"00000000",
  16228=>"00000001",
  16229=>"00000000",
  16230=>"00000000",
  16231=>"00000000",
  16232=>"00000000",
  16233=>"00000000",
  16234=>"11111111",
  16235=>"00000000",
  16236=>"00000000",
  16237=>"00000000",
  16238=>"00000001",
  16239=>"00000000",
  16240=>"00000000",
  16241=>"00000000",
  16242=>"00000000",
  16243=>"00000000",
  16244=>"00000000",
  16245=>"00000000",
  16246=>"00000000",
  16247=>"00000000",
  16248=>"00000000",
  16249=>"00000000",
  16250=>"00000000",
  16251=>"11111111",
  16252=>"00000000",
  16253=>"11111111",
  16254=>"00000000",
  16255=>"00000001",
  16256=>"11111111",
  16257=>"00000000",
  16258=>"00000001",
  16259=>"00000000",
  16260=>"11111111",
  16261=>"00000000",
  16262=>"00000000",
  16263=>"00000000",
  16264=>"00000000",
  16265=>"00000000",
  16266=>"11111111",
  16267=>"00000000",
  16268=>"00000000",
  16269=>"00000001",
  16270=>"00000000",
  16271=>"00000000",
  16272=>"00000000",
  16273=>"00000000",
  16274=>"00000000",
  16275=>"11111111",
  16276=>"11111111",
  16277=>"00000000",
  16278=>"00000000",
  16279=>"00000000",
  16280=>"11111111",
  16281=>"00000000",
  16282=>"00000000",
  16283=>"00000000",
  16284=>"00000000",
  16285=>"00000000",
  16286=>"00000000",
  16287=>"00000000",
  16288=>"00000000",
  16289=>"11111111",
  16290=>"00000000",
  16291=>"00000000",
  16292=>"11111111",
  16293=>"00000000",
  16294=>"00000000",
  16295=>"00000000",
  16296=>"00000001",
  16297=>"00000000",
  16298=>"00000000",
  16299=>"00000001",
  16300=>"00000000",
  16301=>"00000000",
  16302=>"00000000",
  16303=>"00000000",
  16304=>"00000000",
  16305=>"00000000",
  16306=>"00000000",
  16307=>"00000000",
  16308=>"00000001",
  16309=>"00000000",
  16310=>"00000001",
  16311=>"00000000",
  16312=>"00000000",
  16313=>"00000000",
  16314=>"00000000",
  16315=>"00000001",
  16316=>"00000000",
  16317=>"00000000",
  16318=>"00000000",
  16319=>"00000000",
  16320=>"00000000",
  16321=>"00000000",
  16322=>"00000000",
  16323=>"00000000",
  16324=>"00000000",
  16325=>"00000000",
  16326=>"00000000",
  16327=>"11111111",
  16328=>"00000000",
  16329=>"00000001",
  16330=>"00000000",
  16331=>"00000000",
  16332=>"00000000",
  16333=>"11111111",
  16334=>"00000000",
  16335=>"00000000",
  16336=>"00000000",
  16337=>"00000000",
  16338=>"00000000",
  16339=>"00000000",
  16340=>"00000000",
  16341=>"00000000",
  16342=>"00000000",
  16343=>"00000000",
  16344=>"00000000",
  16345=>"00000000",
  16346=>"00000000",
  16347=>"00000000",
  16348=>"00000000",
  16349=>"00000000",
  16350=>"00000000",
  16351=>"00000000",
  16352=>"00000000",
  16353=>"00000000",
  16354=>"00000000",
  16355=>"00000000",
  16356=>"00000000",
  16357=>"00000000",
  16358=>"00000000",
  16359=>"00000000",
  16360=>"00000000",
  16361=>"00000000",
  16362=>"00000000",
  16363=>"00000000",
  16364=>"00000000",
  16365=>"00000000",
  16366=>"00000000",
  16367=>"00000000",
  16368=>"00000001",
  16369=>"00000000",
  16370=>"00000000",
  16371=>"00000000",
  16372=>"00000000",
  16373=>"00000000",
  16374=>"00000000",
  16375=>"11111111",
  16376=>"00000000",
  16377=>"00000000",
  16378=>"00000000",
  16379=>"00000000",
  16380=>"00000000",
  16381=>"00000000",
  16382=>"00000000",
  16383=>"00000000",
  16384=>"11111110",
  16385=>"11111110",
  16386=>"11111010",
  16387=>"11111011",
  16388=>"00000100",
  16389=>"00000011",
  16390=>"11111011",
  16391=>"00000011",
  16392=>"11111110",
  16393=>"00000010",
  16394=>"11111101",
  16395=>"11111110",
  16396=>"00000100",
  16397=>"00000011",
  16398=>"00000101",
  16399=>"00000000",
  16400=>"00000000",
  16401=>"00000100",
  16402=>"00000001",
  16403=>"00000100",
  16404=>"00000011",
  16405=>"00000000",
  16406=>"00000010",
  16407=>"11111001",
  16408=>"11111100",
  16409=>"11111111",
  16410=>"00000011",
  16411=>"00000000",
  16412=>"11111001",
  16413=>"00000010",
  16414=>"11111110",
  16415=>"11111110",
  16416=>"11111111",
  16417=>"11111110",
  16418=>"11111111",
  16419=>"11111011",
  16420=>"11111111",
  16421=>"11111111",
  16422=>"11111011",
  16423=>"00000000",
  16424=>"00000011",
  16425=>"00000000",
  16426=>"11111101",
  16427=>"11111111",
  16428=>"11111110",
  16429=>"11110110",
  16430=>"11111101",
  16431=>"00000010",
  16432=>"11111011",
  16433=>"11111100",
  16434=>"00000000",
  16435=>"11111010",
  16436=>"11110100",
  16437=>"11111111",
  16438=>"11111100",
  16439=>"11111010",
  16440=>"00000001",
  16441=>"11111110",
  16442=>"11111100",
  16443=>"00000101",
  16444=>"00000010",
  16445=>"11111100",
  16446=>"11111110",
  16447=>"11111100",
  16448=>"00000010",
  16449=>"00000100",
  16450=>"11111011",
  16451=>"11110011",
  16452=>"11111111",
  16453=>"11111100",
  16454=>"00000001",
  16455=>"11111110",
  16456=>"11111111",
  16457=>"11111011",
  16458=>"00000001",
  16459=>"00000001",
  16460=>"11111111",
  16461=>"11111111",
  16462=>"11111111",
  16463=>"11111011",
  16464=>"11111111",
  16465=>"11111010",
  16466=>"00000010",
  16467=>"00000011",
  16468=>"11111111",
  16469=>"00000011",
  16470=>"11111111",
  16471=>"11111010",
  16472=>"00000011",
  16473=>"00000011",
  16474=>"00000001",
  16475=>"00000010",
  16476=>"00000000",
  16477=>"11111011",
  16478=>"00000010",
  16479=>"00000101",
  16480=>"00000000",
  16481=>"11111100",
  16482=>"00000011",
  16483=>"00000000",
  16484=>"00000000",
  16485=>"00000010",
  16486=>"00000001",
  16487=>"11111001",
  16488=>"00000110",
  16489=>"00000000",
  16490=>"00000010",
  16491=>"11111100",
  16492=>"00000010",
  16493=>"00000000",
  16494=>"00000001",
  16495=>"11111101",
  16496=>"00000011",
  16497=>"11111110",
  16498=>"00000001",
  16499=>"00000011",
  16500=>"11111110",
  16501=>"11111111",
  16502=>"11111111",
  16503=>"11111100",
  16504=>"11111110",
  16505=>"00000110",
  16506=>"00000010",
  16507=>"11111111",
  16508=>"11111111",
  16509=>"11111110",
  16510=>"11111110",
  16511=>"11111010",
  16512=>"00000101",
  16513=>"11111101",
  16514=>"11111111",
  16515=>"11111110",
  16516=>"00000011",
  16517=>"11111101",
  16518=>"11111100",
  16519=>"00000010",
  16520=>"00000010",
  16521=>"11111110",
  16522=>"00000111",
  16523=>"00000010",
  16524=>"00000010",
  16525=>"11111110",
  16526=>"00000100",
  16527=>"11111111",
  16528=>"11111100",
  16529=>"00000001",
  16530=>"11111001",
  16531=>"11111100",
  16532=>"00000010",
  16533=>"00000000",
  16534=>"11111111",
  16535=>"11111101",
  16536=>"00000001",
  16537=>"11111111",
  16538=>"00000000",
  16539=>"00000001",
  16540=>"11111111",
  16541=>"11111110",
  16542=>"11111011",
  16543=>"00000001",
  16544=>"11111111",
  16545=>"00000010",
  16546=>"00000001",
  16547=>"00000001",
  16548=>"11111010",
  16549=>"11111111",
  16550=>"00000000",
  16551=>"00000101",
  16552=>"00000010",
  16553=>"11111001",
  16554=>"00000000",
  16555=>"00000000",
  16556=>"11111101",
  16557=>"11111011",
  16558=>"00000010",
  16559=>"00000000",
  16560=>"00000011",
  16561=>"11111100",
  16562=>"11111111",
  16563=>"00000000",
  16564=>"00000010",
  16565=>"00000001",
  16566=>"00000001",
  16567=>"11111111",
  16568=>"00000010",
  16569=>"11111101",
  16570=>"00000000",
  16571=>"00000001",
  16572=>"00000000",
  16573=>"11111010",
  16574=>"11111100",
  16575=>"11111110",
  16576=>"11111011",
  16577=>"11111011",
  16578=>"11111111",
  16579=>"00000001",
  16580=>"11111111",
  16581=>"00000011",
  16582=>"11111100",
  16583=>"00000001",
  16584=>"00000011",
  16585=>"00000100",
  16586=>"11111011",
  16587=>"00000000",
  16588=>"00000011",
  16589=>"11111010",
  16590=>"11111101",
  16591=>"11111110",
  16592=>"00000001",
  16593=>"11111111",
  16594=>"11111100",
  16595=>"11111110",
  16596=>"11111010",
  16597=>"00000001",
  16598=>"11111110",
  16599=>"00000001",
  16600=>"00000011",
  16601=>"11111001",
  16602=>"11111101",
  16603=>"00000000",
  16604=>"11111110",
  16605=>"00000010",
  16606=>"00000001",
  16607=>"00000011",
  16608=>"11111011",
  16609=>"00000001",
  16610=>"11111100",
  16611=>"11111111",
  16612=>"11111111",
  16613=>"11111101",
  16614=>"11111111",
  16615=>"11111011",
  16616=>"11110111",
  16617=>"00000000",
  16618=>"00000001",
  16619=>"11111010",
  16620=>"11111011",
  16621=>"11111110",
  16622=>"00000001",
  16623=>"11111011",
  16624=>"00000011",
  16625=>"00000000",
  16626=>"11111100",
  16627=>"11111001",
  16628=>"11111011",
  16629=>"00000011",
  16630=>"00000000",
  16631=>"11111010",
  16632=>"00000010",
  16633=>"11111100",
  16634=>"00000011",
  16635=>"11111100",
  16636=>"00000111",
  16637=>"00000011",
  16638=>"11111110",
  16639=>"00000100",
  16640=>"11111011",
  16641=>"11111111",
  16642=>"00000100",
  16643=>"00000001",
  16644=>"11111110",
  16645=>"11111111",
  16646=>"00000011",
  16647=>"00000001",
  16648=>"11111110",
  16649=>"00000001",
  16650=>"00000011",
  16651=>"11111111",
  16652=>"11111110",
  16653=>"00000001",
  16654=>"11111110",
  16655=>"00000000",
  16656=>"00000000",
  16657=>"00000010",
  16658=>"11111111",
  16659=>"11111110",
  16660=>"00000011",
  16661=>"11111111",
  16662=>"11111110",
  16663=>"00000001",
  16664=>"00000100",
  16665=>"11111000",
  16666=>"11111101",
  16667=>"11111110",
  16668=>"00000110",
  16669=>"11111010",
  16670=>"00000000",
  16671=>"11111111",
  16672=>"11111101",
  16673=>"00000001",
  16674=>"11111111",
  16675=>"11111011",
  16676=>"00000010",
  16677=>"00000011",
  16678=>"00000000",
  16679=>"00000000",
  16680=>"11111100",
  16681=>"11111111",
  16682=>"11111110",
  16683=>"00000100",
  16684=>"11111011",
  16685=>"11111110",
  16686=>"00000000",
  16687=>"00000010",
  16688=>"11111101",
  16689=>"11111010",
  16690=>"00000111",
  16691=>"11111100",
  16692=>"00000001",
  16693=>"11111100",
  16694=>"00000000",
  16695=>"11111100",
  16696=>"11111110",
  16697=>"00000000",
  16698=>"11110111",
  16699=>"11111111",
  16700=>"00000001",
  16701=>"11111110",
  16702=>"11111111",
  16703=>"00000000",
  16704=>"11111011",
  16705=>"11111111",
  16706=>"11111011",
  16707=>"11111000",
  16708=>"11111011",
  16709=>"00000001",
  16710=>"00000011",
  16711=>"00000000",
  16712=>"11111111",
  16713=>"00000011",
  16714=>"00000000",
  16715=>"11111101",
  16716=>"00000000",
  16717=>"11111100",
  16718=>"00000000",
  16719=>"11111110",
  16720=>"11111101",
  16721=>"11111111",
  16722=>"11111101",
  16723=>"00000100",
  16724=>"00000000",
  16725=>"00000110",
  16726=>"11111111",
  16727=>"11111101",
  16728=>"00000000",
  16729=>"00000000",
  16730=>"11111100",
  16731=>"00000000",
  16732=>"11111010",
  16733=>"11111010",
  16734=>"11111110",
  16735=>"11111101",
  16736=>"11111101",
  16737=>"11111111",
  16738=>"11111101",
  16739=>"11111111",
  16740=>"00000001",
  16741=>"11111011",
  16742=>"00001001",
  16743=>"11111001",
  16744=>"11111011",
  16745=>"11111110",
  16746=>"11110110",
  16747=>"00000000",
  16748=>"00000001",
  16749=>"00000001",
  16750=>"00000010",
  16751=>"00000001",
  16752=>"11111100",
  16753=>"11111101",
  16754=>"00000001",
  16755=>"00000010",
  16756=>"11111110",
  16757=>"00000100",
  16758=>"11111110",
  16759=>"11111100",
  16760=>"00000000",
  16761=>"00000000",
  16762=>"00000100",
  16763=>"11111100",
  16764=>"00000001",
  16765=>"11111111",
  16766=>"11111101",
  16767=>"11111110",
  16768=>"11111110",
  16769=>"00000011",
  16770=>"11111100",
  16771=>"11111010",
  16772=>"00000001",
  16773=>"11111110",
  16774=>"11111110",
  16775=>"00000000",
  16776=>"11111110",
  16777=>"00000010",
  16778=>"00000000",
  16779=>"11110100",
  16780=>"11111011",
  16781=>"00000010",
  16782=>"00000010",
  16783=>"00000001",
  16784=>"11111001",
  16785=>"11111110",
  16786=>"11111111",
  16787=>"11111100",
  16788=>"11111111",
  16789=>"00000001",
  16790=>"11111000",
  16791=>"11111110",
  16792=>"11111101",
  16793=>"00000010",
  16794=>"11111110",
  16795=>"11111101",
  16796=>"11110111",
  16797=>"00000110",
  16798=>"11111011",
  16799=>"11111110",
  16800=>"00000010",
  16801=>"11111100",
  16802=>"00000001",
  16803=>"11111111",
  16804=>"11110101",
  16805=>"11111100",
  16806=>"00000000",
  16807=>"11111010",
  16808=>"00000000",
  16809=>"11111110",
  16810=>"11111011",
  16811=>"11111011",
  16812=>"11111101",
  16813=>"00000001",
  16814=>"00000011",
  16815=>"11111101",
  16816=>"11111110",
  16817=>"11111111",
  16818=>"11111011",
  16819=>"00000001",
  16820=>"11111111",
  16821=>"11111110",
  16822=>"00000001",
  16823=>"11111101",
  16824=>"00000000",
  16825=>"11111111",
  16826=>"11111011",
  16827=>"11111011",
  16828=>"11111100",
  16829=>"00000000",
  16830=>"00000001",
  16831=>"11111010",
  16832=>"00000110",
  16833=>"00000010",
  16834=>"00000001",
  16835=>"00000001",
  16836=>"00000011",
  16837=>"11111101",
  16838=>"00000000",
  16839=>"00000001",
  16840=>"00000000",
  16841=>"00000001",
  16842=>"00000001",
  16843=>"00000001",
  16844=>"00000000",
  16845=>"11111010",
  16846=>"00000001",
  16847=>"00000001",
  16848=>"11111100",
  16849=>"00000010",
  16850=>"11111110",
  16851=>"00000000",
  16852=>"11111101",
  16853=>"00000000",
  16854=>"11111110",
  16855=>"11111111",
  16856=>"11111100",
  16857=>"11111110",
  16858=>"11111110",
  16859=>"11111111",
  16860=>"00000001",
  16861=>"11111100",
  16862=>"11111101",
  16863=>"00000000",
  16864=>"11111111",
  16865=>"11111010",
  16866=>"11111101",
  16867=>"00000000",
  16868=>"11111000",
  16869=>"11111001",
  16870=>"11111111",
  16871=>"11111010",
  16872=>"00000100",
  16873=>"11111001",
  16874=>"00000011",
  16875=>"00000001",
  16876=>"00000100",
  16877=>"00000000",
  16878=>"11111111",
  16879=>"11111110",
  16880=>"11111100",
  16881=>"00000010",
  16882=>"11111011",
  16883=>"11111110",
  16884=>"11111010",
  16885=>"00000000",
  16886=>"11111000",
  16887=>"00000100",
  16888=>"00000100",
  16889=>"00000011",
  16890=>"11111011",
  16891=>"00000000",
  16892=>"11111000",
  16893=>"00000011",
  16894=>"00000000",
  16895=>"11111001",
  16896=>"11111110",
  16897=>"00000001",
  16898=>"11111101",
  16899=>"11111100",
  16900=>"00000000",
  16901=>"11111101",
  16902=>"11111111",
  16903=>"00000010",
  16904=>"00000001",
  16905=>"00000010",
  16906=>"11111010",
  16907=>"11111101",
  16908=>"11111110",
  16909=>"11111110",
  16910=>"00000010",
  16911=>"00000000",
  16912=>"00000000",
  16913=>"00000001",
  16914=>"11111110",
  16915=>"00000001",
  16916=>"11111101",
  16917=>"11111010",
  16918=>"11111110",
  16919=>"11111100",
  16920=>"11111101",
  16921=>"00000011",
  16922=>"11111110",
  16923=>"11110111",
  16924=>"11111101",
  16925=>"11111110",
  16926=>"11111110",
  16927=>"00000001",
  16928=>"00000101",
  16929=>"00000010",
  16930=>"11111111",
  16931=>"00000010",
  16932=>"11111101",
  16933=>"00000010",
  16934=>"11111011",
  16935=>"00000001",
  16936=>"00000001",
  16937=>"00000000",
  16938=>"11111110",
  16939=>"00000010",
  16940=>"00000011",
  16941=>"00000001",
  16942=>"00000000",
  16943=>"11111111",
  16944=>"00000011",
  16945=>"00000101",
  16946=>"11111010",
  16947=>"11111100",
  16948=>"11111111",
  16949=>"00000000",
  16950=>"11111100",
  16951=>"00000001",
  16952=>"11111101",
  16953=>"11111000",
  16954=>"11111010",
  16955=>"11111111",
  16956=>"11111110",
  16957=>"00000010",
  16958=>"11111110",
  16959=>"11111010",
  16960=>"00000000",
  16961=>"11111101",
  16962=>"11111110",
  16963=>"11111100",
  16964=>"11111111",
  16965=>"11111111",
  16966=>"00000001",
  16967=>"00000100",
  16968=>"11111111",
  16969=>"11111011",
  16970=>"00000011",
  16971=>"00000011",
  16972=>"11111100",
  16973=>"00000000",
  16974=>"11111111",
  16975=>"11111100",
  16976=>"11111010",
  16977=>"11111111",
  16978=>"11111011",
  16979=>"11111101",
  16980=>"00000000",
  16981=>"11111101",
  16982=>"11111011",
  16983=>"11111010",
  16984=>"00000001",
  16985=>"11111110",
  16986=>"11111101",
  16987=>"00000001",
  16988=>"11111111",
  16989=>"11111110",
  16990=>"11111110",
  16991=>"11111111",
  16992=>"11111101",
  16993=>"11111011",
  16994=>"00000001",
  16995=>"11111111",
  16996=>"00000001",
  16997=>"11111001",
  16998=>"11111001",
  16999=>"11111110",
  17000=>"00000001",
  17001=>"00000010",
  17002=>"11111010",
  17003=>"11111101",
  17004=>"11111110",
  17005=>"11111110",
  17006=>"00000001",
  17007=>"00000010",
  17008=>"00000100",
  17009=>"11111111",
  17010=>"11111110",
  17011=>"11111111",
  17012=>"11111010",
  17013=>"11111101",
  17014=>"00000000",
  17015=>"00000010",
  17016=>"00000010",
  17017=>"11111010",
  17018=>"00000000",
  17019=>"00000011",
  17020=>"11111010",
  17021=>"11111010",
  17022=>"11111111",
  17023=>"11111100",
  17024=>"11111100",
  17025=>"11111010",
  17026=>"11111111",
  17027=>"00000100",
  17028=>"11111101",
  17029=>"00000010",
  17030=>"11111111",
  17031=>"00000010",
  17032=>"11111101",
  17033=>"00000011",
  17034=>"11111101",
  17035=>"00000001",
  17036=>"11111000",
  17037=>"11111100",
  17038=>"11111100",
  17039=>"00000011",
  17040=>"11111110",
  17041=>"00000001",
  17042=>"11111101",
  17043=>"11111100",
  17044=>"00000001",
  17045=>"00000000",
  17046=>"11111111",
  17047=>"00000000",
  17048=>"00000010",
  17049=>"00000001",
  17050=>"11111100",
  17051=>"11111011",
  17052=>"11111110",
  17053=>"00000000",
  17054=>"11111111",
  17055=>"11111110",
  17056=>"11111100",
  17057=>"00000011",
  17058=>"11111101",
  17059=>"00000001",
  17060=>"11111101",
  17061=>"00000000",
  17062=>"00000001",
  17063=>"00000010",
  17064=>"00000001",
  17065=>"00000010",
  17066=>"11111110",
  17067=>"11111101",
  17068=>"11111011",
  17069=>"11111001",
  17070=>"11110111",
  17071=>"00000100",
  17072=>"00000000",
  17073=>"00000000",
  17074=>"11111101",
  17075=>"11110111",
  17076=>"11111011",
  17077=>"00000010",
  17078=>"11111101",
  17079=>"00000111",
  17080=>"00000000",
  17081=>"11111010",
  17082=>"11110111",
  17083=>"11111110",
  17084=>"00000010",
  17085=>"11111111",
  17086=>"00000011",
  17087=>"11111001",
  17088=>"11111010",
  17089=>"00000001",
  17090=>"11111110",
  17091=>"11111100",
  17092=>"11111110",
  17093=>"00000011",
  17094=>"11111011",
  17095=>"00000100",
  17096=>"11111111",
  17097=>"00000000",
  17098=>"00000001",
  17099=>"00000000",
  17100=>"00000000",
  17101=>"00000011",
  17102=>"11111011",
  17103=>"11111100",
  17104=>"11111011",
  17105=>"11111110",
  17106=>"00000001",
  17107=>"00000001",
  17108=>"11111110",
  17109=>"00000001",
  17110=>"11111011",
  17111=>"11111110",
  17112=>"00000010",
  17113=>"11111111",
  17114=>"11111100",
  17115=>"11111110",
  17116=>"00000010",
  17117=>"11111001",
  17118=>"00000001",
  17119=>"00000011",
  17120=>"11111111",
  17121=>"11111111",
  17122=>"00000000",
  17123=>"00000010",
  17124=>"11111100",
  17125=>"11111101",
  17126=>"00000010",
  17127=>"11111100",
  17128=>"11111000",
  17129=>"11111100",
  17130=>"00000010",
  17131=>"11111111",
  17132=>"11111110",
  17133=>"00000001",
  17134=>"11111101",
  17135=>"00000001",
  17136=>"11111101",
  17137=>"11111110",
  17138=>"11111011",
  17139=>"11111101",
  17140=>"11111111",
  17141=>"00000000",
  17142=>"11111110",
  17143=>"11111101",
  17144=>"11111110",
  17145=>"00000010",
  17146=>"00000000",
  17147=>"00000010",
  17148=>"11111001",
  17149=>"00000001",
  17150=>"00000011",
  17151=>"11111110",
  17152=>"11111011",
  17153=>"11111100",
  17154=>"11111100",
  17155=>"11111101",
  17156=>"11111111",
  17157=>"11111010",
  17158=>"11111101",
  17159=>"11111111",
  17160=>"00000000",
  17161=>"00000011",
  17162=>"11111011",
  17163=>"11111111",
  17164=>"00000001",
  17165=>"00000000",
  17166=>"11111111",
  17167=>"11111010",
  17168=>"11111110",
  17169=>"11111111",
  17170=>"11111111",
  17171=>"11111110",
  17172=>"11111010",
  17173=>"00000000",
  17174=>"00000000",
  17175=>"11111110",
  17176=>"00000011",
  17177=>"11111101",
  17178=>"11111111",
  17179=>"11111111",
  17180=>"00000000",
  17181=>"11111111",
  17182=>"11111110",
  17183=>"11111101",
  17184=>"11111110",
  17185=>"00000000",
  17186=>"11111101",
  17187=>"11111101",
  17188=>"00000001",
  17189=>"00000011",
  17190=>"11111111",
  17191=>"00000100",
  17192=>"00000011",
  17193=>"00000011",
  17194=>"00000000",
  17195=>"11111111",
  17196=>"00000000",
  17197=>"11111000",
  17198=>"00000010",
  17199=>"00000100",
  17200=>"00000000",
  17201=>"00000001",
  17202=>"11111110",
  17203=>"00000100",
  17204=>"11111010",
  17205=>"00000010",
  17206=>"11111111",
  17207=>"00000000",
  17208=>"11111111",
  17209=>"11111100",
  17210=>"11111111",
  17211=>"00000011",
  17212=>"11111101",
  17213=>"11111101",
  17214=>"11111101",
  17215=>"00000000",
  17216=>"00000010",
  17217=>"00000000",
  17218=>"11111101",
  17219=>"11111110",
  17220=>"00000000",
  17221=>"11111101",
  17222=>"11111111",
  17223=>"00000001",
  17224=>"00000001",
  17225=>"11111001",
  17226=>"11111111",
  17227=>"00000011",
  17228=>"11111010",
  17229=>"11111010",
  17230=>"00000001",
  17231=>"00000011",
  17232=>"00000000",
  17233=>"11111011",
  17234=>"11111110",
  17235=>"00000011",
  17236=>"11111010",
  17237=>"11111110",
  17238=>"11111111",
  17239=>"00000001",
  17240=>"00000001",
  17241=>"11111001",
  17242=>"11111101",
  17243=>"11111111",
  17244=>"11111100",
  17245=>"00000010",
  17246=>"11111110",
  17247=>"00000001",
  17248=>"00000000",
  17249=>"11111100",
  17250=>"00000001",
  17251=>"11111110",
  17252=>"00000010",
  17253=>"11111001",
  17254=>"11111111",
  17255=>"11111110",
  17256=>"11111011",
  17257=>"00000010",
  17258=>"11111011",
  17259=>"11111101",
  17260=>"11111010",
  17261=>"00000001",
  17262=>"00000101",
  17263=>"11111111",
  17264=>"00000100",
  17265=>"00000000",
  17266=>"11111101",
  17267=>"00000001",
  17268=>"11111001",
  17269=>"11111111",
  17270=>"11111111",
  17271=>"00000000",
  17272=>"00000001",
  17273=>"00000001",
  17274=>"11111110",
  17275=>"11111100",
  17276=>"00000000",
  17277=>"00000000",
  17278=>"11111110",
  17279=>"00000010",
  17280=>"11111010",
  17281=>"11111111",
  17282=>"11111000",
  17283=>"00000001",
  17284=>"11111101",
  17285=>"11111101",
  17286=>"11111010",
  17287=>"11111111",
  17288=>"00000000",
  17289=>"11111111",
  17290=>"11111101",
  17291=>"00000010",
  17292=>"11111110",
  17293=>"11111101",
  17294=>"00000011",
  17295=>"11111001",
  17296=>"11110110",
  17297=>"00000000",
  17298=>"00000010",
  17299=>"11111010",
  17300=>"11111100",
  17301=>"11111110",
  17302=>"00000010",
  17303=>"11111110",
  17304=>"11111100",
  17305=>"11111101",
  17306=>"11111111",
  17307=>"00000001",
  17308=>"11111101",
  17309=>"11111001",
  17310=>"00000000",
  17311=>"11111010",
  17312=>"00000000",
  17313=>"11111101",
  17314=>"00000100",
  17315=>"11111011",
  17316=>"11111101",
  17317=>"00000001",
  17318=>"00000011",
  17319=>"00000000",
  17320=>"11111000",
  17321=>"11111100",
  17322=>"11111110",
  17323=>"11111011",
  17324=>"11111101",
  17325=>"11111100",
  17326=>"11111101",
  17327=>"11111011",
  17328=>"00000011",
  17329=>"11111101",
  17330=>"11111111",
  17331=>"00000000",
  17332=>"11111101",
  17333=>"00000010",
  17334=>"11111101",
  17335=>"00000001",
  17336=>"11111111",
  17337=>"11111001",
  17338=>"11111110",
  17339=>"11111010",
  17340=>"11111101",
  17341=>"00000001",
  17342=>"11111101",
  17343=>"11111110",
  17344=>"00000001",
  17345=>"11111101",
  17346=>"11111001",
  17347=>"11111011",
  17348=>"11111001",
  17349=>"11111010",
  17350=>"11111111",
  17351=>"11111001",
  17352=>"00000011",
  17353=>"11111100",
  17354=>"11111110",
  17355=>"11111111",
  17356=>"11111101",
  17357=>"00000001",
  17358=>"00000001",
  17359=>"11111110",
  17360=>"11111110",
  17361=>"00000010",
  17362=>"00000001",
  17363=>"11111001",
  17364=>"11111101",
  17365=>"11111101",
  17366=>"11111100",
  17367=>"00000100",
  17368=>"11111010",
  17369=>"11111110",
  17370=>"11111101",
  17371=>"11111111",
  17372=>"11111001",
  17373=>"00000011",
  17374=>"00000001",
  17375=>"00000001",
  17376=>"00000000",
  17377=>"11111111",
  17378=>"11111101",
  17379=>"11111110",
  17380=>"11111011",
  17381=>"11111110",
  17382=>"00000010",
  17383=>"00000010",
  17384=>"11111110",
  17385=>"11111010",
  17386=>"00000011",
  17387=>"00000001",
  17388=>"00000001",
  17389=>"11111011",
  17390=>"00000110",
  17391=>"11111110",
  17392=>"11111110",
  17393=>"11111101",
  17394=>"00000011",
  17395=>"11111010",
  17396=>"11111101",
  17397=>"00000101",
  17398=>"00000100",
  17399=>"11111110",
  17400=>"11111011",
  17401=>"11110111",
  17402=>"00000001",
  17403=>"11111111",
  17404=>"00000100",
  17405=>"00000000",
  17406=>"11111110",
  17407=>"11111110",
  17408=>"11111111",
  17409=>"00000010",
  17410=>"00000010",
  17411=>"00000000",
  17412=>"11111100",
  17413=>"11111111",
  17414=>"11111110",
  17415=>"00000001",
  17416=>"00000001",
  17417=>"00000001",
  17418=>"00000001",
  17419=>"00000000",
  17420=>"11111101",
  17421=>"00000000",
  17422=>"00000010",
  17423=>"11111110",
  17424=>"11111111",
  17425=>"00000010",
  17426=>"11111111",
  17427=>"00000010",
  17428=>"11111111",
  17429=>"11111111",
  17430=>"11111111",
  17431=>"00000001",
  17432=>"00000000",
  17433=>"00000001",
  17434=>"11111110",
  17435=>"11111100",
  17436=>"11111110",
  17437=>"11111110",
  17438=>"11111110",
  17439=>"00000100",
  17440=>"11111100",
  17441=>"11111110",
  17442=>"11111111",
  17443=>"11111110",
  17444=>"00000010",
  17445=>"00000011",
  17446=>"11111101",
  17447=>"11111111",
  17448=>"00000000",
  17449=>"00000000",
  17450=>"00000010",
  17451=>"00000000",
  17452=>"11111110",
  17453=>"00000010",
  17454=>"00000001",
  17455=>"00000010",
  17456=>"00000001",
  17457=>"11111110",
  17458=>"11111110",
  17459=>"11111101",
  17460=>"00000000",
  17461=>"00000010",
  17462=>"00000010",
  17463=>"00000010",
  17464=>"11111111",
  17465=>"00000001",
  17466=>"11111101",
  17467=>"00000011",
  17468=>"11111101",
  17469=>"11111111",
  17470=>"00000000",
  17471=>"11111101",
  17472=>"11111110",
  17473=>"11111100",
  17474=>"11111111",
  17475=>"11111110",
  17476=>"00000001",
  17477=>"11111111",
  17478=>"11111111",
  17479=>"11111101",
  17480=>"11111101",
  17481=>"00000000",
  17482=>"00000001",
  17483=>"11111111",
  17484=>"11111111",
  17485=>"00000000",
  17486=>"00000011",
  17487=>"00000010",
  17488=>"00000000",
  17489=>"11111110",
  17490=>"11111101",
  17491=>"11111101",
  17492=>"11111101",
  17493=>"00000010",
  17494=>"11111110",
  17495=>"00000001",
  17496=>"00000100",
  17497=>"11111101",
  17498=>"11111110",
  17499=>"11111101",
  17500=>"11111111",
  17501=>"00000011",
  17502=>"11111110",
  17503=>"00000100",
  17504=>"00000100",
  17505=>"00000000",
  17506=>"11111101",
  17507=>"00000010",
  17508=>"00000100",
  17509=>"00000010",
  17510=>"00000010",
  17511=>"11111110",
  17512=>"11111111",
  17513=>"00000100",
  17514=>"00000000",
  17515=>"00000010",
  17516=>"11111111",
  17517=>"00000000",
  17518=>"00000001",
  17519=>"00000011",
  17520=>"00000000",
  17521=>"00000010",
  17522=>"11111101",
  17523=>"00000010",
  17524=>"00000001",
  17525=>"11111101",
  17526=>"11111111",
  17527=>"00000100",
  17528=>"11111110",
  17529=>"00000000",
  17530=>"00000011",
  17531=>"00000011",
  17532=>"00000000",
  17533=>"00000011",
  17534=>"00000001",
  17535=>"00000000",
  17536=>"11111110",
  17537=>"00000010",
  17538=>"11111111",
  17539=>"11111111",
  17540=>"00000001",
  17541=>"11111110",
  17542=>"00000000",
  17543=>"00000101",
  17544=>"00000010",
  17545=>"11111101",
  17546=>"00000010",
  17547=>"11111100",
  17548=>"11111111",
  17549=>"00000000",
  17550=>"11111100",
  17551=>"11111101",
  17552=>"00000001",
  17553=>"11111110",
  17554=>"00000001",
  17555=>"11111111",
  17556=>"11111110",
  17557=>"00000011",
  17558=>"11111101",
  17559=>"11111111",
  17560=>"11111111",
  17561=>"00000010",
  17562=>"11111111",
  17563=>"11111110",
  17564=>"00000010",
  17565=>"11111110",
  17566=>"00000001",
  17567=>"11111111",
  17568=>"00000011",
  17569=>"00000100",
  17570=>"00000001",
  17571=>"11111111",
  17572=>"11111101",
  17573=>"11111111",
  17574=>"11111111",
  17575=>"11111110",
  17576=>"11111111",
  17577=>"11111111",
  17578=>"11111101",
  17579=>"00000010",
  17580=>"00000010",
  17581=>"11111111",
  17582=>"00000011",
  17583=>"00000000",
  17584=>"11111110",
  17585=>"00000000",
  17586=>"00000010",
  17587=>"00000000",
  17588=>"00000000",
  17589=>"11111101",
  17590=>"11111110",
  17591=>"11111110",
  17592=>"00000011",
  17593=>"00000000",
  17594=>"11111110",
  17595=>"00000001",
  17596=>"00000001",
  17597=>"00000010",
  17598=>"11111110",
  17599=>"00000001",
  17600=>"00000001",
  17601=>"00000001",
  17602=>"11111110",
  17603=>"00000010",
  17604=>"11111110",
  17605=>"00000010",
  17606=>"00000110",
  17607=>"11111111",
  17608=>"11111101",
  17609=>"11111100",
  17610=>"11111111",
  17611=>"11111110",
  17612=>"11111101",
  17613=>"11111110",
  17614=>"00000001",
  17615=>"00000010",
  17616=>"00000001",
  17617=>"11111111",
  17618=>"00000010",
  17619=>"11111111",
  17620=>"00000000",
  17621=>"11111101",
  17622=>"11111111",
  17623=>"00000000",
  17624=>"00000000",
  17625=>"00000001",
  17626=>"11111111",
  17627=>"00000000",
  17628=>"00000001",
  17629=>"00000000",
  17630=>"00000011",
  17631=>"11111110",
  17632=>"11111111",
  17633=>"11111110",
  17634=>"11111111",
  17635=>"00000000",
  17636=>"11111101",
  17637=>"11111110",
  17638=>"11111110",
  17639=>"11111110",
  17640=>"11111110",
  17641=>"11111110",
  17642=>"00000010",
  17643=>"11111111",
  17644=>"00000000",
  17645=>"11111101",
  17646=>"00000001",
  17647=>"11111111",
  17648=>"11111111",
  17649=>"00000010",
  17650=>"11111111",
  17651=>"11111110",
  17652=>"00000010",
  17653=>"00000010",
  17654=>"00000000",
  17655=>"00000000",
  17656=>"00000011",
  17657=>"00000010",
  17658=>"00000001",
  17659=>"11111110",
  17660=>"11111111",
  17661=>"00000100",
  17662=>"11111111",
  17663=>"00000100",
  17664=>"00000100",
  17665=>"00000000",
  17666=>"11111101",
  17667=>"00000010",
  17668=>"00000001",
  17669=>"00000000",
  17670=>"11111101",
  17671=>"00000101",
  17672=>"00000001",
  17673=>"11111111",
  17674=>"00000000",
  17675=>"11111111",
  17676=>"00000000",
  17677=>"11111101",
  17678=>"00000001",
  17679=>"11111101",
  17680=>"00000010",
  17681=>"11111111",
  17682=>"11111110",
  17683=>"00000001",
  17684=>"11111110",
  17685=>"00000011",
  17686=>"11111111",
  17687=>"00000001",
  17688=>"00000011",
  17689=>"11111110",
  17690=>"00000010",
  17691=>"11111110",
  17692=>"00000110",
  17693=>"00000001",
  17694=>"00000010",
  17695=>"00000100",
  17696=>"11111101",
  17697=>"11111101",
  17698=>"00000010",
  17699=>"00000010",
  17700=>"00000000",
  17701=>"11111101",
  17702=>"00000001",
  17703=>"11111111",
  17704=>"00000001",
  17705=>"11111101",
  17706=>"00000110",
  17707=>"11111101",
  17708=>"11111101",
  17709=>"00000001",
  17710=>"11111110",
  17711=>"11111101",
  17712=>"00000100",
  17713=>"11111111",
  17714=>"00000101",
  17715=>"11111101",
  17716=>"11111110",
  17717=>"11111110",
  17718=>"00000100",
  17719=>"00000010",
  17720=>"11111111",
  17721=>"00000010",
  17722=>"11111110",
  17723=>"11111111",
  17724=>"11111100",
  17725=>"11111110",
  17726=>"11111111",
  17727=>"11111101",
  17728=>"00000000",
  17729=>"11111110",
  17730=>"00000011",
  17731=>"11111110",
  17732=>"11111111",
  17733=>"00000010",
  17734=>"00000011",
  17735=>"00000010",
  17736=>"00000000",
  17737=>"00000011",
  17738=>"11111110",
  17739=>"00000010",
  17740=>"11111101",
  17741=>"00000000",
  17742=>"00000011",
  17743=>"11111101",
  17744=>"00000010",
  17745=>"00000010",
  17746=>"11111110",
  17747=>"11111110",
  17748=>"11111101",
  17749=>"11111101",
  17750=>"11111101",
  17751=>"11111111",
  17752=>"00000100",
  17753=>"11111101",
  17754=>"00000001",
  17755=>"00000010",
  17756=>"11111110",
  17757=>"11111101",
  17758=>"00000010",
  17759=>"00000001",
  17760=>"00000000",
  17761=>"00000010",
  17762=>"00000011",
  17763=>"00000001",
  17764=>"00000000",
  17765=>"00000000",
  17766=>"00000001",
  17767=>"11111111",
  17768=>"11111101",
  17769=>"00000011",
  17770=>"11111111",
  17771=>"11111110",
  17772=>"11111111",
  17773=>"00000000",
  17774=>"11111110",
  17775=>"11111110",
  17776=>"11111110",
  17777=>"00000001",
  17778=>"11111110",
  17779=>"11111101",
  17780=>"00000001",
  17781=>"11111111",
  17782=>"00000000",
  17783=>"00000000",
  17784=>"00000001",
  17785=>"11111111",
  17786=>"11111111",
  17787=>"11111101",
  17788=>"00000000",
  17789=>"11111110",
  17790=>"00000011",
  17791=>"11111101",
  17792=>"11111110",
  17793=>"00000000",
  17794=>"00000001",
  17795=>"00000011",
  17796=>"11111110",
  17797=>"11111111",
  17798=>"11111101",
  17799=>"11111101",
  17800=>"11111111",
  17801=>"11111111",
  17802=>"00000000",
  17803=>"00000010",
  17804=>"00000010",
  17805=>"00000000",
  17806=>"11111101",
  17807=>"00000010",
  17808=>"11111110",
  17809=>"00000000",
  17810=>"11111100",
  17811=>"00000010",
  17812=>"11111100",
  17813=>"00000000",
  17814=>"11111111",
  17815=>"00000000",
  17816=>"11111110",
  17817=>"00000010",
  17818=>"00000001",
  17819=>"00000011",
  17820=>"00000010",
  17821=>"00000001",
  17822=>"00000010",
  17823=>"11111111",
  17824=>"11111101",
  17825=>"00000001",
  17826=>"11111101",
  17827=>"11111110",
  17828=>"11111111",
  17829=>"11111110",
  17830=>"11111110",
  17831=>"00000001",
  17832=>"00000100",
  17833=>"00000000",
  17834=>"00000000",
  17835=>"00000000",
  17836=>"11111101",
  17837=>"00000000",
  17838=>"11111111",
  17839=>"11111110",
  17840=>"11111110",
  17841=>"11111101",
  17842=>"00000100",
  17843=>"11111101",
  17844=>"11111110",
  17845=>"00000000",
  17846=>"00000001",
  17847=>"11111111",
  17848=>"00000100",
  17849=>"00000001",
  17850=>"11111101",
  17851=>"00000001",
  17852=>"11111111",
  17853=>"00000010",
  17854=>"00000001",
  17855=>"00000001",
  17856=>"00000000",
  17857=>"00000100",
  17858=>"00000001",
  17859=>"00000011",
  17860=>"11111111",
  17861=>"11111101",
  17862=>"11111111",
  17863=>"11111101",
  17864=>"00000000",
  17865=>"00000100",
  17866=>"00000000",
  17867=>"00000000",
  17868=>"00000000",
  17869=>"00000010",
  17870=>"00000101",
  17871=>"00000010",
  17872=>"11111111",
  17873=>"00000010",
  17874=>"00000010",
  17875=>"11111111",
  17876=>"11111101",
  17877=>"00000000",
  17878=>"00000110",
  17879=>"00000000",
  17880=>"00000000",
  17881=>"00000101",
  17882=>"11111111",
  17883=>"00000110",
  17884=>"00000011",
  17885=>"11111111",
  17886=>"00000000",
  17887=>"11111111",
  17888=>"11111111",
  17889=>"11111111",
  17890=>"11111110",
  17891=>"00000000",
  17892=>"00000001",
  17893=>"00000010",
  17894=>"00000011",
  17895=>"11111110",
  17896=>"00000000",
  17897=>"11111111",
  17898=>"00000101",
  17899=>"11111111",
  17900=>"11111111",
  17901=>"00000011",
  17902=>"00000100",
  17903=>"00000001",
  17904=>"00000001",
  17905=>"00000000",
  17906=>"11111110",
  17907=>"00000001",
  17908=>"00000000",
  17909=>"11111110",
  17910=>"11111111",
  17911=>"00000101",
  17912=>"11111101",
  17913=>"00000010",
  17914=>"00000001",
  17915=>"00000101",
  17916=>"11111110",
  17917=>"11111111",
  17918=>"00000000",
  17919=>"00000000",
  17920=>"00000001",
  17921=>"00000000",
  17922=>"11111110",
  17923=>"11111111",
  17924=>"00000010",
  17925=>"00000100",
  17926=>"00000000",
  17927=>"11111110",
  17928=>"11111110",
  17929=>"00000000",
  17930=>"11111111",
  17931=>"00000001",
  17932=>"11111111",
  17933=>"11111110",
  17934=>"11111111",
  17935=>"11111101",
  17936=>"00000011",
  17937=>"00000110",
  17938=>"00000001",
  17939=>"11111110",
  17940=>"00000010",
  17941=>"11111110",
  17942=>"11111110",
  17943=>"00000110",
  17944=>"11111101",
  17945=>"11111110",
  17946=>"00000100",
  17947=>"11111111",
  17948=>"00000000",
  17949=>"11111110",
  17950=>"00000010",
  17951=>"11111110",
  17952=>"11111100",
  17953=>"11111110",
  17954=>"11111111",
  17955=>"00000010",
  17956=>"11111101",
  17957=>"00000010",
  17958=>"00000000",
  17959=>"11111101",
  17960=>"11111111",
  17961=>"00000001",
  17962=>"00000011",
  17963=>"00000001",
  17964=>"00000011",
  17965=>"11111111",
  17966=>"00000111",
  17967=>"00000001",
  17968=>"11111101",
  17969=>"00000001",
  17970=>"11111110",
  17971=>"00000011",
  17972=>"00000010",
  17973=>"11111111",
  17974=>"00000011",
  17975=>"00000001",
  17976=>"00000000",
  17977=>"00000001",
  17978=>"11111111",
  17979=>"00000011",
  17980=>"11111101",
  17981=>"11111101",
  17982=>"11111101",
  17983=>"11111101",
  17984=>"11111110",
  17985=>"11111111",
  17986=>"00000000",
  17987=>"11111110",
  17988=>"11111111",
  17989=>"00000010",
  17990=>"00000000",
  17991=>"00000100",
  17992=>"00000011",
  17993=>"00000001",
  17994=>"11111111",
  17995=>"00000001",
  17996=>"00000011",
  17997=>"11111111",
  17998=>"11111110",
  17999=>"00000010",
  18000=>"00000010",
  18001=>"00000000",
  18002=>"00000011",
  18003=>"00000010",
  18004=>"11111101",
  18005=>"00000010",
  18006=>"00000000",
  18007=>"00000011",
  18008=>"00000001",
  18009=>"00000011",
  18010=>"00000000",
  18011=>"00000000",
  18012=>"00000001",
  18013=>"00000000",
  18014=>"00000000",
  18015=>"11111101",
  18016=>"00000100",
  18017=>"11111101",
  18018=>"11111111",
  18019=>"00000010",
  18020=>"00000010",
  18021=>"00000010",
  18022=>"11111110",
  18023=>"00000011",
  18024=>"11111110",
  18025=>"00000010",
  18026=>"11111110",
  18027=>"11111110",
  18028=>"11111100",
  18029=>"00000000",
  18030=>"11111110",
  18031=>"11111101",
  18032=>"11111101",
  18033=>"11111110",
  18034=>"00000001",
  18035=>"11111111",
  18036=>"00000011",
  18037=>"00000000",
  18038=>"00000010",
  18039=>"00000000",
  18040=>"11111111",
  18041=>"11111111",
  18042=>"00000101",
  18043=>"00000101",
  18044=>"00000010",
  18045=>"11111111",
  18046=>"11111101",
  18047=>"00000100",
  18048=>"00000000",
  18049=>"11111111",
  18050=>"11111111",
  18051=>"11111110",
  18052=>"11111111",
  18053=>"00000001",
  18054=>"11111110",
  18055=>"00000001",
  18056=>"11111111",
  18057=>"11111110",
  18058=>"00000011",
  18059=>"11111111",
  18060=>"00000001",
  18061=>"11111111",
  18062=>"11111110",
  18063=>"11111101",
  18064=>"00000000",
  18065=>"11111101",
  18066=>"11111110",
  18067=>"11111111",
  18068=>"11111111",
  18069=>"11111110",
  18070=>"00000010",
  18071=>"00000011",
  18072=>"00000011",
  18073=>"00000001",
  18074=>"00000000",
  18075=>"00000010",
  18076=>"11111110",
  18077=>"11111111",
  18078=>"00000000",
  18079=>"00000000",
  18080=>"11111101",
  18081=>"00000100",
  18082=>"11111100",
  18083=>"00000001",
  18084=>"00000000",
  18085=>"11111110",
  18086=>"11111101",
  18087=>"00000100",
  18088=>"11111101",
  18089=>"11111101",
  18090=>"11111101",
  18091=>"11111101",
  18092=>"11111110",
  18093=>"00000000",
  18094=>"11111101",
  18095=>"00000010",
  18096=>"00000010",
  18097=>"11111111",
  18098=>"11111101",
  18099=>"11111101",
  18100=>"00000001",
  18101=>"00000101",
  18102=>"00000011",
  18103=>"11111101",
  18104=>"00000000",
  18105=>"11111110",
  18106=>"00000010",
  18107=>"00000001",
  18108=>"00000001",
  18109=>"00000000",
  18110=>"11111110",
  18111=>"00000001",
  18112=>"11111111",
  18113=>"11111110",
  18114=>"11111110",
  18115=>"00000100",
  18116=>"11111111",
  18117=>"11111101",
  18118=>"00000000",
  18119=>"11111111",
  18120=>"11111101",
  18121=>"00000001",
  18122=>"00000000",
  18123=>"11111111",
  18124=>"11111111",
  18125=>"11111111",
  18126=>"11111101",
  18127=>"11111110",
  18128=>"00000010",
  18129=>"11111110",
  18130=>"11111101",
  18131=>"11111111",
  18132=>"00000010",
  18133=>"00000001",
  18134=>"00000010",
  18135=>"11111111",
  18136=>"00000000",
  18137=>"00000000",
  18138=>"11111110",
  18139=>"00000001",
  18140=>"00000011",
  18141=>"11111111",
  18142=>"11111111",
  18143=>"11111111",
  18144=>"00000001",
  18145=>"11111111",
  18146=>"11111110",
  18147=>"00000101",
  18148=>"11111111",
  18149=>"00000001",
  18150=>"00000000",
  18151=>"11111111",
  18152=>"00000001",
  18153=>"11111101",
  18154=>"00000011",
  18155=>"11111100",
  18156=>"00000000",
  18157=>"00000101",
  18158=>"11111110",
  18159=>"00000010",
  18160=>"00000100",
  18161=>"11111110",
  18162=>"11111110",
  18163=>"00000001",
  18164=>"00000001",
  18165=>"00000001",
  18166=>"11111101",
  18167=>"00000001",
  18168=>"11111110",
  18169=>"11111110",
  18170=>"00000000",
  18171=>"11111110",
  18172=>"00000000",
  18173=>"00000011",
  18174=>"11111111",
  18175=>"11111110",
  18176=>"00000111",
  18177=>"00000001",
  18178=>"11111110",
  18179=>"11111110",
  18180=>"00000001",
  18181=>"00000001",
  18182=>"00000010",
  18183=>"11111111",
  18184=>"00000001",
  18185=>"00000000",
  18186=>"11111111",
  18187=>"11111111",
  18188=>"11111111",
  18189=>"00000000",
  18190=>"11111101",
  18191=>"11111111",
  18192=>"00000001",
  18193=>"11111101",
  18194=>"11111101",
  18195=>"00000000",
  18196=>"00000010",
  18197=>"11111110",
  18198=>"11111111",
  18199=>"11111110",
  18200=>"11111111",
  18201=>"00000010",
  18202=>"00000011",
  18203=>"11111101",
  18204=>"11111111",
  18205=>"11111110",
  18206=>"11111110",
  18207=>"00000000",
  18208=>"00000010",
  18209=>"00000001",
  18210=>"00000001",
  18211=>"00000000",
  18212=>"11111111",
  18213=>"00000001",
  18214=>"00000101",
  18215=>"11111100",
  18216=>"11111110",
  18217=>"11111101",
  18218=>"00000000",
  18219=>"00000011",
  18220=>"00000000",
  18221=>"00000001",
  18222=>"00000000",
  18223=>"11111110",
  18224=>"00000100",
  18225=>"11111110",
  18226=>"00000011",
  18227=>"00000000",
  18228=>"00000000",
  18229=>"00000000",
  18230=>"00000010",
  18231=>"11111101",
  18232=>"11111111",
  18233=>"00000000",
  18234=>"11111101",
  18235=>"00000011",
  18236=>"11111111",
  18237=>"11111110",
  18238=>"11111110",
  18239=>"11111110",
  18240=>"00000101",
  18241=>"11111100",
  18242=>"00000001",
  18243=>"00000011",
  18244=>"00000000",
  18245=>"00000000",
  18246=>"11111101",
  18247=>"00000100",
  18248=>"00000010",
  18249=>"00000000",
  18250=>"00000010",
  18251=>"11111110",
  18252=>"11111101",
  18253=>"11111101",
  18254=>"00000001",
  18255=>"00000010",
  18256=>"11111111",
  18257=>"00000000",
  18258=>"00000000",
  18259=>"00000001",
  18260=>"11111101",
  18261=>"00000001",
  18262=>"11111101",
  18263=>"11111111",
  18264=>"00000010",
  18265=>"11111110",
  18266=>"11111110",
  18267=>"11111110",
  18268=>"00000000",
  18269=>"11111111",
  18270=>"11111111",
  18271=>"11111110",
  18272=>"00000001",
  18273=>"11111110",
  18274=>"11111110",
  18275=>"11111101",
  18276=>"00000011",
  18277=>"11111110",
  18278=>"11111110",
  18279=>"00000000",
  18280=>"00000011",
  18281=>"00000110",
  18282=>"00000010",
  18283=>"00000010",
  18284=>"11111110",
  18285=>"00000000",
  18286=>"00000010",
  18287=>"00000000",
  18288=>"11111110",
  18289=>"11111111",
  18290=>"00000000",
  18291=>"11111111",
  18292=>"00000001",
  18293=>"00000000",
  18294=>"00000011",
  18295=>"00000001",
  18296=>"00000000",
  18297=>"11111101",
  18298=>"00000000",
  18299=>"11111101",
  18300=>"11111111",
  18301=>"11111110",
  18302=>"11111110",
  18303=>"11111100",
  18304=>"00000000",
  18305=>"11111111",
  18306=>"11111110",
  18307=>"11111110",
  18308=>"00000001",
  18309=>"11111111",
  18310=>"00000010",
  18311=>"11111111",
  18312=>"11111111",
  18313=>"00000011",
  18314=>"11111111",
  18315=>"11111110",
  18316=>"00000011",
  18317=>"11111101",
  18318=>"00000010",
  18319=>"00000001",
  18320=>"00000000",
  18321=>"11111110",
  18322=>"11111111",
  18323=>"11111111",
  18324=>"00000001",
  18325=>"00000010",
  18326=>"00000011",
  18327=>"11111111",
  18328=>"11111110",
  18329=>"00000001",
  18330=>"11111110",
  18331=>"11111111",
  18332=>"00000000",
  18333=>"00000001",
  18334=>"00000001",
  18335=>"11111101",
  18336=>"11111101",
  18337=>"00000001",
  18338=>"00000000",
  18339=>"00000000",
  18340=>"11111101",
  18341=>"00000001",
  18342=>"11111101",
  18343=>"00000001",
  18344=>"00000000",
  18345=>"00000000",
  18346=>"00000001",
  18347=>"00000010",
  18348=>"00000000",
  18349=>"00000000",
  18350=>"00000000",
  18351=>"11111101",
  18352=>"00000010",
  18353=>"00000000",
  18354=>"11111111",
  18355=>"11111111",
  18356=>"00000000",
  18357=>"11111101",
  18358=>"00000001",
  18359=>"00000100",
  18360=>"00000000",
  18361=>"11111111",
  18362=>"11111110",
  18363=>"11111110",
  18364=>"00000100",
  18365=>"00000101",
  18366=>"00000000",
  18367=>"00000010",
  18368=>"00000010",
  18369=>"00000010",
  18370=>"00000000",
  18371=>"00000001",
  18372=>"11111110",
  18373=>"00000001",
  18374=>"11111101",
  18375=>"11111111",
  18376=>"11111101",
  18377=>"00000010",
  18378=>"00000011",
  18379=>"00000011",
  18380=>"00000000",
  18381=>"00000010",
  18382=>"00000011",
  18383=>"11111111",
  18384=>"11111101",
  18385=>"00000000",
  18386=>"00000101",
  18387=>"00000010",
  18388=>"11111111",
  18389=>"00000001",
  18390=>"00000000",
  18391=>"11111100",
  18392=>"11111110",
  18393=>"00000001",
  18394=>"11111110",
  18395=>"00000011",
  18396=>"00000000",
  18397=>"00000001",
  18398=>"00000001",
  18399=>"11111110",
  18400=>"11111111",
  18401=>"00000000",
  18402=>"00000010",
  18403=>"00000000",
  18404=>"11111110",
  18405=>"11111101",
  18406=>"00000011",
  18407=>"11111110",
  18408=>"00000011",
  18409=>"00000010",
  18410=>"11111100",
  18411=>"00000000",
  18412=>"11111111",
  18413=>"00000010",
  18414=>"00000110",
  18415=>"00000000",
  18416=>"00000000",
  18417=>"00000010",
  18418=>"00000001",
  18419=>"00000001",
  18420=>"00000011",
  18421=>"00000010",
  18422=>"00000000",
  18423=>"00000001",
  18424=>"00000001",
  18425=>"00000010",
  18426=>"00000001",
  18427=>"00000000",
  18428=>"00000010",
  18429=>"00000001",
  18430=>"00000011",
  18431=>"11111101",
  18432=>"00000010",
  18433=>"00000000",
  18434=>"00000001",
  18435=>"11111110",
  18436=>"00000011",
  18437=>"00000000",
  18438=>"11111111",
  18439=>"11111111",
  18440=>"00000000",
  18441=>"11111111",
  18442=>"11111101",
  18443=>"00000011",
  18444=>"11111110",
  18445=>"11111100",
  18446=>"00000001",
  18447=>"11111111",
  18448=>"11111100",
  18449=>"00000101",
  18450=>"11111110",
  18451=>"00000010",
  18452=>"00000101",
  18453=>"00000010",
  18454=>"00000001",
  18455=>"00000000",
  18456=>"00000010",
  18457=>"00000010",
  18458=>"11111100",
  18459=>"00000000",
  18460=>"11111101",
  18461=>"00000000",
  18462=>"00000001",
  18463=>"11111100",
  18464=>"11111101",
  18465=>"00000010",
  18466=>"11111101",
  18467=>"00000001",
  18468=>"11111110",
  18469=>"11111111",
  18470=>"11111111",
  18471=>"00000001",
  18472=>"00000001",
  18473=>"11111111",
  18474=>"00000001",
  18475=>"11111110",
  18476=>"11111111",
  18477=>"11111111",
  18478=>"00000001",
  18479=>"00000010",
  18480=>"11111110",
  18481=>"00000010",
  18482=>"11111111",
  18483=>"11111110",
  18484=>"00000010",
  18485=>"11111110",
  18486=>"00000001",
  18487=>"00000010",
  18488=>"00000011",
  18489=>"00000010",
  18490=>"00000000",
  18491=>"00000101",
  18492=>"11111111",
  18493=>"11111101",
  18494=>"00000001",
  18495=>"00000000",
  18496=>"00000001",
  18497=>"00000001",
  18498=>"11111110",
  18499=>"00000000",
  18500=>"11111110",
  18501=>"00000000",
  18502=>"11111111",
  18503=>"00000010",
  18504=>"00000010",
  18505=>"11111111",
  18506=>"11111110",
  18507=>"00000000",
  18508=>"11111111",
  18509=>"00000000",
  18510=>"11111101",
  18511=>"00000001",
  18512=>"00000001",
  18513=>"00000000",
  18514=>"00000001",
  18515=>"00000011",
  18516=>"00000001",
  18517=>"00000001",
  18518=>"11111110",
  18519=>"00000001",
  18520=>"11111110",
  18521=>"00000000",
  18522=>"00000000",
  18523=>"00000010",
  18524=>"00000101",
  18525=>"11111111",
  18526=>"11111100",
  18527=>"11111101",
  18528=>"11111110",
  18529=>"00000000",
  18530=>"00000000",
  18531=>"00000000",
  18532=>"11111110",
  18533=>"11111101",
  18534=>"11111111",
  18535=>"11111101",
  18536=>"11111110",
  18537=>"00000000",
  18538=>"11111111",
  18539=>"00000010",
  18540=>"11111111",
  18541=>"00000100",
  18542=>"11111111",
  18543=>"11111101",
  18544=>"11111110",
  18545=>"11111110",
  18546=>"00000001",
  18547=>"11111110",
  18548=>"00000001",
  18549=>"11111101",
  18550=>"11111101",
  18551=>"11111101",
  18552=>"00000001",
  18553=>"00000010",
  18554=>"00000010",
  18555=>"00000000",
  18556=>"00000010",
  18557=>"00000010",
  18558=>"00000001",
  18559=>"11111110",
  18560=>"11111111",
  18561=>"11111111",
  18562=>"00000001",
  18563=>"00000000",
  18564=>"11111111",
  18565=>"11111110",
  18566=>"00000000",
  18567=>"00000000",
  18568=>"00000001",
  18569=>"11111101",
  18570=>"00000000",
  18571=>"00000011",
  18572=>"00000000",
  18573=>"00000011",
  18574=>"11111100",
  18575=>"11111101",
  18576=>"11111101",
  18577=>"00000000",
  18578=>"00000000",
  18579=>"00000001",
  18580=>"00000010",
  18581=>"11111111",
  18582=>"00000001",
  18583=>"11111110",
  18584=>"00000000",
  18585=>"00000000",
  18586=>"00000010",
  18587=>"11111101",
  18588=>"00000001",
  18589=>"00000001",
  18590=>"11111111",
  18591=>"11111101",
  18592=>"00000010",
  18593=>"00000110",
  18594=>"00000001",
  18595=>"11111111",
  18596=>"11111110",
  18597=>"11111111",
  18598=>"11111101",
  18599=>"00000011",
  18600=>"11111110",
  18601=>"00000001",
  18602=>"00000010",
  18603=>"11111101",
  18604=>"00000001",
  18605=>"00000001",
  18606=>"11111110",
  18607=>"00000010",
  18608=>"11111110",
  18609=>"00000001",
  18610=>"11111111",
  18611=>"11111101",
  18612=>"00000000",
  18613=>"00000000",
  18614=>"11111111",
  18615=>"00000000",
  18616=>"11111110",
  18617=>"11111110",
  18618=>"11111111",
  18619=>"00000010",
  18620=>"00000001",
  18621=>"00000010",
  18622=>"00000011",
  18623=>"00000001",
  18624=>"00000001",
  18625=>"00000001",
  18626=>"00000100",
  18627=>"00000000",
  18628=>"00000001",
  18629=>"11111101",
  18630=>"00000001",
  18631=>"00000001",
  18632=>"00000100",
  18633=>"11111111",
  18634=>"11111110",
  18635=>"00000000",
  18636=>"11111101",
  18637=>"11111110",
  18638=>"00000000",
  18639=>"11111111",
  18640=>"00000011",
  18641=>"11111101",
  18642=>"00000000",
  18643=>"11111110",
  18644=>"00000001",
  18645=>"00000100",
  18646=>"00000001",
  18647=>"00000001",
  18648=>"11111110",
  18649=>"11111101",
  18650=>"00000001",
  18651=>"11111101",
  18652=>"00000001",
  18653=>"00000000",
  18654=>"00000000",
  18655=>"11111111",
  18656=>"11111110",
  18657=>"00000000",
  18658=>"11111111",
  18659=>"00000010",
  18660=>"00000000",
  18661=>"00000010",
  18662=>"00000001",
  18663=>"00000001",
  18664=>"11111110",
  18665=>"00000001",
  18666=>"11111111",
  18667=>"11111110",
  18668=>"11111101",
  18669=>"00000001",
  18670=>"00000001",
  18671=>"00000010",
  18672=>"11111100",
  18673=>"11111101",
  18674=>"11111111",
  18675=>"00000010",
  18676=>"11111110",
  18677=>"00000001",
  18678=>"00000011",
  18679=>"00000000",
  18680=>"00000100",
  18681=>"11111111",
  18682=>"11111110",
  18683=>"00000001",
  18684=>"00000100",
  18685=>"00000010",
  18686=>"11111101",
  18687=>"11111100",
  18688=>"00000000",
  18689=>"11111111",
  18690=>"00000011",
  18691=>"11111101",
  18692=>"00000000",
  18693=>"00000000",
  18694=>"00000001",
  18695=>"00000000",
  18696=>"00000000",
  18697=>"11111110",
  18698=>"00000000",
  18699=>"00000000",
  18700=>"11111110",
  18701=>"11111111",
  18702=>"11111111",
  18703=>"11111110",
  18704=>"11111110",
  18705=>"00000000",
  18706=>"00000100",
  18707=>"11111110",
  18708=>"11111111",
  18709=>"00000001",
  18710=>"00000010",
  18711=>"11111111",
  18712=>"11111110",
  18713=>"11111101",
  18714=>"11111101",
  18715=>"00000011",
  18716=>"11111101",
  18717=>"11111111",
  18718=>"11111101",
  18719=>"00000000",
  18720=>"00000010",
  18721=>"00000100",
  18722=>"00000001",
  18723=>"11111110",
  18724=>"00000000",
  18725=>"00000000",
  18726=>"00000011",
  18727=>"11111100",
  18728=>"00000001",
  18729=>"00000010",
  18730=>"11111111",
  18731=>"00000011",
  18732=>"00000001",
  18733=>"00000010",
  18734=>"11111101",
  18735=>"11111101",
  18736=>"00000000",
  18737=>"11111110",
  18738=>"00000010",
  18739=>"00000010",
  18740=>"00000000",
  18741=>"11111110",
  18742=>"11111110",
  18743=>"00000010",
  18744=>"00000000",
  18745=>"11111111",
  18746=>"00000010",
  18747=>"11111111",
  18748=>"00000001",
  18749=>"00000001",
  18750=>"00000010",
  18751=>"00000001",
  18752=>"00000010",
  18753=>"00000000",
  18754=>"00000011",
  18755=>"11111111",
  18756=>"11111111",
  18757=>"00000001",
  18758=>"11111110",
  18759=>"11111111",
  18760=>"11111101",
  18761=>"11111100",
  18762=>"11111100",
  18763=>"00000010",
  18764=>"00000101",
  18765=>"11111111",
  18766=>"00000100",
  18767=>"11111111",
  18768=>"11111111",
  18769=>"00000001",
  18770=>"11111111",
  18771=>"11111101",
  18772=>"00000001",
  18773=>"00000000",
  18774=>"00000011",
  18775=>"11111110",
  18776=>"00000100",
  18777=>"00000000",
  18778=>"00000010",
  18779=>"11111111",
  18780=>"00000001",
  18781=>"00000001",
  18782=>"11111101",
  18783=>"11111111",
  18784=>"11111110",
  18785=>"11111110",
  18786=>"00000001",
  18787=>"00000000",
  18788=>"00000000",
  18789=>"11111111",
  18790=>"00000010",
  18791=>"00000010",
  18792=>"00000000",
  18793=>"00000011",
  18794=>"00000001",
  18795=>"00000000",
  18796=>"11111110",
  18797=>"00000000",
  18798=>"00000010",
  18799=>"11111111",
  18800=>"11111110",
  18801=>"11111110",
  18802=>"00000011",
  18803=>"00000101",
  18804=>"00000010",
  18805=>"11111111",
  18806=>"11111110",
  18807=>"00000010",
  18808=>"11111111",
  18809=>"00000101",
  18810=>"11111110",
  18811=>"00000101",
  18812=>"11111111",
  18813=>"11111111",
  18814=>"11111111",
  18815=>"00000100",
  18816=>"00000001",
  18817=>"11111101",
  18818=>"00000000",
  18819=>"11111110",
  18820=>"00000000",
  18821=>"00000100",
  18822=>"11111100",
  18823=>"00000011",
  18824=>"00000001",
  18825=>"00000001",
  18826=>"11111110",
  18827=>"00000001",
  18828=>"11111111",
  18829=>"11111101",
  18830=>"11111101",
  18831=>"00000001",
  18832=>"11111111",
  18833=>"00000010",
  18834=>"00000000",
  18835=>"11111110",
  18836=>"11111111",
  18837=>"00000010",
  18838=>"00000011",
  18839=>"00000011",
  18840=>"00000000",
  18841=>"11111101",
  18842=>"00000001",
  18843=>"11111110",
  18844=>"00000010",
  18845=>"00000000",
  18846=>"11111101",
  18847=>"11111111",
  18848=>"00000011",
  18849=>"00000001",
  18850=>"11111111",
  18851=>"11111110",
  18852=>"11111111",
  18853=>"11111111",
  18854=>"11111110",
  18855=>"00000001",
  18856=>"00000000",
  18857=>"11111111",
  18858=>"11111111",
  18859=>"00000010",
  18860=>"11111111",
  18861=>"00000000",
  18862=>"11111111",
  18863=>"00000001",
  18864=>"11111111",
  18865=>"11111110",
  18866=>"11111110",
  18867=>"00000011",
  18868=>"00000101",
  18869=>"00000100",
  18870=>"00000001",
  18871=>"11111111",
  18872=>"11111110",
  18873=>"00000001",
  18874=>"00000010",
  18875=>"11111101",
  18876=>"11111110",
  18877=>"00000011",
  18878=>"11111110",
  18879=>"00000000",
  18880=>"00000000",
  18881=>"00000011",
  18882=>"00000001",
  18883=>"00000010",
  18884=>"00000000",
  18885=>"00000010",
  18886=>"11111111",
  18887=>"00000100",
  18888=>"11111111",
  18889=>"00000010",
  18890=>"00000010",
  18891=>"00000010",
  18892=>"11111111",
  18893=>"11111111",
  18894=>"00000001",
  18895=>"00000001",
  18896=>"11111111",
  18897=>"00000001",
  18898=>"00000010",
  18899=>"00000001",
  18900=>"00000001",
  18901=>"00000001",
  18902=>"00000011",
  18903=>"11111101",
  18904=>"11111111",
  18905=>"00000101",
  18906=>"11111101",
  18907=>"00000000",
  18908=>"00000000",
  18909=>"11111111",
  18910=>"11111110",
  18911=>"00000000",
  18912=>"11111111",
  18913=>"00000010",
  18914=>"11111110",
  18915=>"00000010",
  18916=>"00000010",
  18917=>"00000011",
  18918=>"00000000",
  18919=>"11111110",
  18920=>"00000101",
  18921=>"11111111",
  18922=>"11111100",
  18923=>"11111101",
  18924=>"00000001",
  18925=>"00000001",
  18926=>"11111101",
  18927=>"11111110",
  18928=>"00000001",
  18929=>"00000010",
  18930=>"00000010",
  18931=>"00000000",
  18932=>"00000000",
  18933=>"11111111",
  18934=>"00000000",
  18935=>"11111101",
  18936=>"11111110",
  18937=>"00000000",
  18938=>"00000010",
  18939=>"00000010",
  18940=>"00000010",
  18941=>"00000010",
  18942=>"11111110",
  18943=>"11111110",
  18944=>"00000001",
  18945=>"11111111",
  18946=>"00000110",
  18947=>"00000001",
  18948=>"11111110",
  18949=>"00000000",
  18950=>"00000110",
  18951=>"00000001",
  18952=>"11111101",
  18953=>"00000001",
  18954=>"11111110",
  18955=>"00000010",
  18956=>"11111111",
  18957=>"11111110",
  18958=>"11111100",
  18959=>"11111110",
  18960=>"00000010",
  18961=>"00000010",
  18962=>"00000010",
  18963=>"00000011",
  18964=>"11111111",
  18965=>"11111110",
  18966=>"00000001",
  18967=>"00000001",
  18968=>"11111111",
  18969=>"11111110",
  18970=>"00000001",
  18971=>"00000001",
  18972=>"11111110",
  18973=>"00000100",
  18974=>"00000001",
  18975=>"11111101",
  18976=>"00000000",
  18977=>"00000000",
  18978=>"00000001",
  18979=>"00000001",
  18980=>"11111101",
  18981=>"11111111",
  18982=>"00000001",
  18983=>"11111111",
  18984=>"11111110",
  18985=>"00000010",
  18986=>"11111100",
  18987=>"00000001",
  18988=>"00000010",
  18989=>"11111110",
  18990=>"00000001",
  18991=>"00000101",
  18992=>"00000010",
  18993=>"11111111",
  18994=>"00000000",
  18995=>"00000001",
  18996=>"00000000",
  18997=>"11111101",
  18998=>"00000011",
  18999=>"11111111",
  19000=>"11111111",
  19001=>"00000001",
  19002=>"00000010",
  19003=>"00000011",
  19004=>"00000010",
  19005=>"11111111",
  19006=>"00000001",
  19007=>"11111101",
  19008=>"11111101",
  19009=>"11111110",
  19010=>"00000010",
  19011=>"11111110",
  19012=>"00000010",
  19013=>"00000000",
  19014=>"11111111",
  19015=>"11111101",
  19016=>"11111111",
  19017=>"00000000",
  19018=>"00000011",
  19019=>"11111101",
  19020=>"00000000",
  19021=>"00000010",
  19022=>"11111110",
  19023=>"00000000",
  19024=>"11111111",
  19025=>"11111111",
  19026=>"00000010",
  19027=>"11111101",
  19028=>"00000000",
  19029=>"00000100",
  19030=>"11111110",
  19031=>"11111110",
  19032=>"00000001",
  19033=>"11111101",
  19034=>"00000001",
  19035=>"11111110",
  19036=>"11111111",
  19037=>"00000000",
  19038=>"11111111",
  19039=>"00000000",
  19040=>"00000101",
  19041=>"11111111",
  19042=>"00000001",
  19043=>"00000001",
  19044=>"00000011",
  19045=>"11111110",
  19046=>"00000011",
  19047=>"11111110",
  19048=>"00000000",
  19049=>"00000011",
  19050=>"00000000",
  19051=>"11111111",
  19052=>"00000011",
  19053=>"00000001",
  19054=>"00000100",
  19055=>"11111100",
  19056=>"11111111",
  19057=>"00000010",
  19058=>"11111110",
  19059=>"00000000",
  19060=>"00000011",
  19061=>"11111110",
  19062=>"00000001",
  19063=>"11111111",
  19064=>"11111111",
  19065=>"00000000",
  19066=>"00000000",
  19067=>"00000001",
  19068=>"11111101",
  19069=>"11111110",
  19070=>"00000000",
  19071=>"00000010",
  19072=>"11111111",
  19073=>"11111111",
  19074=>"00000000",
  19075=>"11111101",
  19076=>"00000010",
  19077=>"00000001",
  19078=>"00000011",
  19079=>"11111110",
  19080=>"11111111",
  19081=>"11111100",
  19082=>"00000000",
  19083=>"00001000",
  19084=>"00000001",
  19085=>"00000000",
  19086=>"11111101",
  19087=>"00000001",
  19088=>"11111110",
  19089=>"11111101",
  19090=>"00000000",
  19091=>"11111110",
  19092=>"00000001",
  19093=>"00000000",
  19094=>"00000000",
  19095=>"00000100",
  19096=>"00000101",
  19097=>"11111101",
  19098=>"00000010",
  19099=>"00000010",
  19100=>"00000001",
  19101=>"11111111",
  19102=>"00000010",
  19103=>"00000001",
  19104=>"00000010",
  19105=>"11111111",
  19106=>"00000100",
  19107=>"11111111",
  19108=>"11111110",
  19109=>"11111111",
  19110=>"11111111",
  19111=>"00000000",
  19112=>"00000000",
  19113=>"00000011",
  19114=>"00000011",
  19115=>"11111110",
  19116=>"11111111",
  19117=>"00000000",
  19118=>"00000010",
  19119=>"00000000",
  19120=>"00000001",
  19121=>"11111111",
  19122=>"00000001",
  19123=>"11111101",
  19124=>"00000010",
  19125=>"11111110",
  19126=>"00000011",
  19127=>"00000000",
  19128=>"00000000",
  19129=>"00000001",
  19130=>"00000001",
  19131=>"00000000",
  19132=>"11111110",
  19133=>"00000001",
  19134=>"11111110",
  19135=>"00000100",
  19136=>"11111111",
  19137=>"11111111",
  19138=>"11111101",
  19139=>"11111111",
  19140=>"00000001",
  19141=>"00000001",
  19142=>"00000010",
  19143=>"11111110",
  19144=>"00000000",
  19145=>"11111111",
  19146=>"11111101",
  19147=>"00000010",
  19148=>"00000101",
  19149=>"11111101",
  19150=>"00000000",
  19151=>"11111111",
  19152=>"00000000",
  19153=>"00000000",
  19154=>"11111111",
  19155=>"11111111",
  19156=>"00000000",
  19157=>"11111111",
  19158=>"11111110",
  19159=>"11111110",
  19160=>"11111011",
  19161=>"11111110",
  19162=>"00000010",
  19163=>"11111111",
  19164=>"00000110",
  19165=>"11111110",
  19166=>"11111110",
  19167=>"11111101",
  19168=>"00000001",
  19169=>"11111111",
  19170=>"00000000",
  19171=>"11111111",
  19172=>"11111111",
  19173=>"00000000",
  19174=>"11111111",
  19175=>"00000100",
  19176=>"00000001",
  19177=>"00000000",
  19178=>"00000000",
  19179=>"00000001",
  19180=>"00000001",
  19181=>"11111110",
  19182=>"11111101",
  19183=>"11111101",
  19184=>"00000001",
  19185=>"00000000",
  19186=>"00000000",
  19187=>"11111111",
  19188=>"00000001",
  19189=>"00000101",
  19190=>"00000000",
  19191=>"00000010",
  19192=>"00000010",
  19193=>"11111111",
  19194=>"11111111",
  19195=>"00000100",
  19196=>"00000001",
  19197=>"00000000",
  19198=>"00000010",
  19199=>"11111110",
  19200=>"00000011",
  19201=>"00000000",
  19202=>"11111111",
  19203=>"00000010",
  19204=>"00000011",
  19205=>"00000001",
  19206=>"00000010",
  19207=>"00000000",
  19208=>"11111101",
  19209=>"11111111",
  19210=>"11111111",
  19211=>"00000010",
  19212=>"00000011",
  19213=>"11111111",
  19214=>"00000100",
  19215=>"11111110",
  19216=>"11111101",
  19217=>"00000000",
  19218=>"00000000",
  19219=>"00000010",
  19220=>"00000000",
  19221=>"11111110",
  19222=>"00000011",
  19223=>"11111110",
  19224=>"11111111",
  19225=>"11111100",
  19226=>"11111110",
  19227=>"11111101",
  19228=>"11111111",
  19229=>"11111101",
  19230=>"11111101",
  19231=>"11111110",
  19232=>"00000000",
  19233=>"00000001",
  19234=>"11111111",
  19235=>"00000000",
  19236=>"11111110",
  19237=>"00000110",
  19238=>"11111111",
  19239=>"11111110",
  19240=>"11111111",
  19241=>"00000000",
  19242=>"11111110",
  19243=>"00000011",
  19244=>"11111110",
  19245=>"11111110",
  19246=>"11111110",
  19247=>"11111110",
  19248=>"11111111",
  19249=>"00000001",
  19250=>"11111110",
  19251=>"00000001",
  19252=>"00000010",
  19253=>"11111101",
  19254=>"11111110",
  19255=>"00000000",
  19256=>"11111101",
  19257=>"11111111",
  19258=>"00000001",
  19259=>"00000001",
  19260=>"00000000",
  19261=>"00000000",
  19262=>"00000011",
  19263=>"11111101",
  19264=>"11111100",
  19265=>"11111110",
  19266=>"00000001",
  19267=>"11111110",
  19268=>"11111101",
  19269=>"00000011",
  19270=>"00000011",
  19271=>"00000001",
  19272=>"00000000",
  19273=>"00000010",
  19274=>"11111111",
  19275=>"00000001",
  19276=>"00000010",
  19277=>"00000001",
  19278=>"11111101",
  19279=>"11111110",
  19280=>"11111111",
  19281=>"11111110",
  19282=>"11111110",
  19283=>"00000000",
  19284=>"11111111",
  19285=>"11111111",
  19286=>"00000001",
  19287=>"11111111",
  19288=>"00000111",
  19289=>"11111101",
  19290=>"11111111",
  19291=>"11111110",
  19292=>"00000010",
  19293=>"00000001",
  19294=>"11111111",
  19295=>"00000011",
  19296=>"11111100",
  19297=>"11111101",
  19298=>"11111110",
  19299=>"11111111",
  19300=>"00000010",
  19301=>"00000010",
  19302=>"00000001",
  19303=>"00000000",
  19304=>"00000000",
  19305=>"11111100",
  19306=>"11111110",
  19307=>"11111111",
  19308=>"00000001",
  19309=>"11111110",
  19310=>"00000100",
  19311=>"11111110",
  19312=>"00000011",
  19313=>"11111100",
  19314=>"00000000",
  19315=>"00000010",
  19316=>"00000001",
  19317=>"11111101",
  19318=>"11111111",
  19319=>"11111111",
  19320=>"11111101",
  19321=>"00000000",
  19322=>"00000010",
  19323=>"00000000",
  19324=>"11111110",
  19325=>"00000011",
  19326=>"00000000",
  19327=>"11111111",
  19328=>"00000011",
  19329=>"00000010",
  19330=>"00000000",
  19331=>"00000000",
  19332=>"00000001",
  19333=>"11111101",
  19334=>"11111110",
  19335=>"00000001",
  19336=>"11111100",
  19337=>"00000000",
  19338=>"00000010",
  19339=>"00000000",
  19340=>"00000010",
  19341=>"00000010",
  19342=>"11111111",
  19343=>"00000000",
  19344=>"00000010",
  19345=>"11111100",
  19346=>"11111110",
  19347=>"11111111",
  19348=>"11111101",
  19349=>"00000001",
  19350=>"00000000",
  19351=>"11111110",
  19352=>"11111101",
  19353=>"11111110",
  19354=>"11111101",
  19355=>"11111111",
  19356=>"11111100",
  19357=>"00000001",
  19358=>"00000000",
  19359=>"00000100",
  19360=>"00000001",
  19361=>"11111111",
  19362=>"00000000",
  19363=>"11111111",
  19364=>"11111111",
  19365=>"11111110",
  19366=>"00000001",
  19367=>"11111111",
  19368=>"00000000",
  19369=>"00000001",
  19370=>"11111110",
  19371=>"00000000",
  19372=>"00000000",
  19373=>"00000001",
  19374=>"11111101",
  19375=>"00000001",
  19376=>"00000011",
  19377=>"00000001",
  19378=>"00000011",
  19379=>"11111101",
  19380=>"11111111",
  19381=>"11111111",
  19382=>"11111110",
  19383=>"00000010",
  19384=>"11111111",
  19385=>"00000000",
  19386=>"11111101",
  19387=>"00000000",
  19388=>"11111110",
  19389=>"00000011",
  19390=>"00000000",
  19391=>"00000010",
  19392=>"11111101",
  19393=>"11111110",
  19394=>"11111111",
  19395=>"00000000",
  19396=>"11111111",
  19397=>"00000010",
  19398=>"00000010",
  19399=>"00000010",
  19400=>"00000010",
  19401=>"00000011",
  19402=>"00000000",
  19403=>"11111111",
  19404=>"00000010",
  19405=>"11111110",
  19406=>"00000001",
  19407=>"00000000",
  19408=>"00000100",
  19409=>"00000011",
  19410=>"11111111",
  19411=>"11111110",
  19412=>"11111110",
  19413=>"00000010",
  19414=>"00000000",
  19415=>"00000001",
  19416=>"11111111",
  19417=>"00000001",
  19418=>"11111111",
  19419=>"00000000",
  19420=>"00000001",
  19421=>"00000110",
  19422=>"00000000",
  19423=>"00000100",
  19424=>"11111110",
  19425=>"00000000",
  19426=>"11111111",
  19427=>"00000000",
  19428=>"00000001",
  19429=>"11111111",
  19430=>"11111110",
  19431=>"11111111",
  19432=>"11111111",
  19433=>"00000001",
  19434=>"00000010",
  19435=>"11111100",
  19436=>"00000101",
  19437=>"00000000",
  19438=>"00000000",
  19439=>"00000000",
  19440=>"11111110",
  19441=>"11111111",
  19442=>"00000011",
  19443=>"11111111",
  19444=>"11111110",
  19445=>"00000001",
  19446=>"11111100",
  19447=>"00000011",
  19448=>"11111110",
  19449=>"11111111",
  19450=>"11111110",
  19451=>"00000101",
  19452=>"00000001",
  19453=>"00000100",
  19454=>"00000001",
  19455=>"00000000",
  19456=>"00000001",
  19457=>"11111110",
  19458=>"00000100",
  19459=>"11111110",
  19460=>"11111111",
  19461=>"11111101",
  19462=>"00000001",
  19463=>"00000010",
  19464=>"00000001",
  19465=>"11111110",
  19466=>"00000011",
  19467=>"00000001",
  19468=>"00000010",
  19469=>"00000011",
  19470=>"11111111",
  19471=>"00000001",
  19472=>"00000111",
  19473=>"11111101",
  19474=>"11111111",
  19475=>"11111110",
  19476=>"00000010",
  19477=>"00000000",
  19478=>"00000101",
  19479=>"11111111",
  19480=>"00000001",
  19481=>"11111110",
  19482=>"00000011",
  19483=>"11111110",
  19484=>"11111110",
  19485=>"00000001",
  19486=>"00000000",
  19487=>"00000001",
  19488=>"11111101",
  19489=>"00000010",
  19490=>"00000011",
  19491=>"11111111",
  19492=>"00000010",
  19493=>"11111111",
  19494=>"00000000",
  19495=>"00000000",
  19496=>"00000001",
  19497=>"11111101",
  19498=>"11111111",
  19499=>"11111111",
  19500=>"00000010",
  19501=>"00000010",
  19502=>"11111111",
  19503=>"00000010",
  19504=>"11111110",
  19505=>"11111111",
  19506=>"11111110",
  19507=>"00000010",
  19508=>"00000001",
  19509=>"00000011",
  19510=>"00000010",
  19511=>"00000000",
  19512=>"11111110",
  19513=>"00000010",
  19514=>"00000001",
  19515=>"00000001",
  19516=>"00000001",
  19517=>"00000000",
  19518=>"11111110",
  19519=>"00000001",
  19520=>"11111101",
  19521=>"00000100",
  19522=>"00000001",
  19523=>"00000010",
  19524=>"00000000",
  19525=>"00000010",
  19526=>"00000011",
  19527=>"00000010",
  19528=>"11111110",
  19529=>"11111101",
  19530=>"11111110",
  19531=>"11111101",
  19532=>"00000011",
  19533=>"11111111",
  19534=>"00000001",
  19535=>"11111101",
  19536=>"00000001",
  19537=>"00000001",
  19538=>"11111100",
  19539=>"11111111",
  19540=>"00000001",
  19541=>"00000100",
  19542=>"00000010",
  19543=>"00000011",
  19544=>"00000101",
  19545=>"00000011",
  19546=>"11111110",
  19547=>"00000010",
  19548=>"11111110",
  19549=>"11111111",
  19550=>"00000000",
  19551=>"11111111",
  19552=>"11111111",
  19553=>"00000001",
  19554=>"11111110",
  19555=>"00000000",
  19556=>"00000000",
  19557=>"00000010",
  19558=>"11111110",
  19559=>"00000000",
  19560=>"00000101",
  19561=>"00000000",
  19562=>"00000010",
  19563=>"00000010",
  19564=>"11111110",
  19565=>"00000000",
  19566=>"11111101",
  19567=>"00000100",
  19568=>"00000001",
  19569=>"11111110",
  19570=>"00000000",
  19571=>"11111110",
  19572=>"11111101",
  19573=>"00000000",
  19574=>"11111110",
  19575=>"00000011",
  19576=>"11111110",
  19577=>"11111111",
  19578=>"00000000",
  19579=>"11111110",
  19580=>"00000011",
  19581=>"00000011",
  19582=>"11111110",
  19583=>"11111101",
  19584=>"00000011",
  19585=>"11111111",
  19586=>"00000000",
  19587=>"11111111",
  19588=>"11111110",
  19589=>"11111101",
  19590=>"11111101",
  19591=>"11111101",
  19592=>"00000001",
  19593=>"00000101",
  19594=>"11111110",
  19595=>"00000000",
  19596=>"11111110",
  19597=>"11111110",
  19598=>"11111111",
  19599=>"00000001",
  19600=>"11111101",
  19601=>"11111101",
  19602=>"11111110",
  19603=>"11111110",
  19604=>"00000000",
  19605=>"11111111",
  19606=>"11111101",
  19607=>"11111111",
  19608=>"00000101",
  19609=>"00000100",
  19610=>"00000000",
  19611=>"00000000",
  19612=>"00000001",
  19613=>"00000000",
  19614=>"00000010",
  19615=>"11111111",
  19616=>"11111101",
  19617=>"00000010",
  19618=>"00000101",
  19619=>"11111110",
  19620=>"00000001",
  19621=>"00000101",
  19622=>"11111110",
  19623=>"11111110",
  19624=>"00000010",
  19625=>"11111111",
  19626=>"11111101",
  19627=>"11111110",
  19628=>"00000001",
  19629=>"00000001",
  19630=>"11111101",
  19631=>"00000010",
  19632=>"00000001",
  19633=>"11111110",
  19634=>"00000011",
  19635=>"11111110",
  19636=>"11111110",
  19637=>"11111101",
  19638=>"00000000",
  19639=>"11111111",
  19640=>"00000010",
  19641=>"11111100",
  19642=>"11111101",
  19643=>"11111111",
  19644=>"00000011",
  19645=>"11111110",
  19646=>"00000010",
  19647=>"00000001",
  19648=>"00000011",
  19649=>"00000001",
  19650=>"11111110",
  19651=>"11111111",
  19652=>"00000000",
  19653=>"00000000",
  19654=>"00000000",
  19655=>"11111111",
  19656=>"00000011",
  19657=>"00000000",
  19658=>"11111110",
  19659=>"00000000",
  19660=>"00000001",
  19661=>"11111111",
  19662=>"11111111",
  19663=>"11111111",
  19664=>"11111111",
  19665=>"11111101",
  19666=>"00000000",
  19667=>"00000101",
  19668=>"00000000",
  19669=>"11111101",
  19670=>"11111101",
  19671=>"11111101",
  19672=>"11111101",
  19673=>"00000000",
  19674=>"00000000",
  19675=>"00000001",
  19676=>"00000010",
  19677=>"00000000",
  19678=>"11111111",
  19679=>"00000000",
  19680=>"00000011",
  19681=>"00000010",
  19682=>"11111111",
  19683=>"00000010",
  19684=>"00000010",
  19685=>"00000010",
  19686=>"00000011",
  19687=>"00000010",
  19688=>"00000010",
  19689=>"00000100",
  19690=>"11111111",
  19691=>"00000000",
  19692=>"11111111",
  19693=>"00000001",
  19694=>"00000010",
  19695=>"00000001",
  19696=>"11111110",
  19697=>"00000001",
  19698=>"00000000",
  19699=>"00000000",
  19700=>"11111111",
  19701=>"00000010",
  19702=>"00000000",
  19703=>"11111111",
  19704=>"11111111",
  19705=>"11111110",
  19706=>"11111110",
  19707=>"11111111",
  19708=>"11111111",
  19709=>"00000001",
  19710=>"00000000",
  19711=>"00000000",
  19712=>"11111110",
  19713=>"11111011",
  19714=>"00000100",
  19715=>"11111110",
  19716=>"00000011",
  19717=>"00000000",
  19718=>"11111101",
  19719=>"00000010",
  19720=>"00000000",
  19721=>"00000001",
  19722=>"11111110",
  19723=>"00000010",
  19724=>"00000000",
  19725=>"11111111",
  19726=>"00000000",
  19727=>"00000000",
  19728=>"00000001",
  19729=>"11111101",
  19730=>"11111111",
  19731=>"11111110",
  19732=>"11111100",
  19733=>"00000101",
  19734=>"00000100",
  19735=>"11111111",
  19736=>"00000110",
  19737=>"00000010",
  19738=>"00000010",
  19739=>"00000000",
  19740=>"00000000",
  19741=>"00000001",
  19742=>"00000100",
  19743=>"00000110",
  19744=>"00000010",
  19745=>"00000011",
  19746=>"11111110",
  19747=>"00000001",
  19748=>"11111111",
  19749=>"11111101",
  19750=>"00000101",
  19751=>"11111101",
  19752=>"00000010",
  19753=>"11111100",
  19754=>"00000011",
  19755=>"00000000",
  19756=>"11111111",
  19757=>"00000000",
  19758=>"11111101",
  19759=>"11111101",
  19760=>"00000001",
  19761=>"11111111",
  19762=>"11111110",
  19763=>"00000010",
  19764=>"11111101",
  19765=>"00000000",
  19766=>"11111110",
  19767=>"11111110",
  19768=>"00000010",
  19769=>"00000010",
  19770=>"00000001",
  19771=>"11111111",
  19772=>"00000010",
  19773=>"00000000",
  19774=>"00000000",
  19775=>"11111111",
  19776=>"00000000",
  19777=>"00000000",
  19778=>"11111101",
  19779=>"11111110",
  19780=>"00000011",
  19781=>"00000010",
  19782=>"11111101",
  19783=>"00000011",
  19784=>"00000010",
  19785=>"00000000",
  19786=>"11111110",
  19787=>"11111111",
  19788=>"00000001",
  19789=>"11111110",
  19790=>"11111111",
  19791=>"11111111",
  19792=>"00000000",
  19793=>"11111111",
  19794=>"11111101",
  19795=>"00000100",
  19796=>"11111111",
  19797=>"11111110",
  19798=>"00000101",
  19799=>"11111110",
  19800=>"11111110",
  19801=>"00000000",
  19802=>"00000001",
  19803=>"00000001",
  19804=>"11111110",
  19805=>"11111111",
  19806=>"11111101",
  19807=>"00000001",
  19808=>"00000100",
  19809=>"11111110",
  19810=>"00000010",
  19811=>"00000010",
  19812=>"11111101",
  19813=>"11111111",
  19814=>"00000001",
  19815=>"00000010",
  19816=>"11111111",
  19817=>"11111101",
  19818=>"00000010",
  19819=>"11111111",
  19820=>"11111111",
  19821=>"11111101",
  19822=>"00000001",
  19823=>"11111110",
  19824=>"00000000",
  19825=>"00000000",
  19826=>"11111100",
  19827=>"00000010",
  19828=>"00000001",
  19829=>"00000110",
  19830=>"00000010",
  19831=>"00000010",
  19832=>"00000000",
  19833=>"00000000",
  19834=>"00000010",
  19835=>"00000001",
  19836=>"00000011",
  19837=>"00000001",
  19838=>"00000000",
  19839=>"00000001",
  19840=>"00000100",
  19841=>"11111110",
  19842=>"00000010",
  19843=>"00000010",
  19844=>"00000001",
  19845=>"00000000",
  19846=>"00000000",
  19847=>"11111101",
  19848=>"00000001",
  19849=>"00000010",
  19850=>"11111111",
  19851=>"11111110",
  19852=>"00000001",
  19853=>"11111101",
  19854=>"11111110",
  19855=>"00000010",
  19856=>"00000001",
  19857=>"00000000",
  19858=>"00000010",
  19859=>"11111111",
  19860=>"11111110",
  19861=>"11111111",
  19862=>"11111111",
  19863=>"00000001",
  19864=>"11111101",
  19865=>"00000001",
  19866=>"00000000",
  19867=>"11111110",
  19868=>"00000000",
  19869=>"00000000",
  19870=>"00000011",
  19871=>"00000001",
  19872=>"00000000",
  19873=>"00000010",
  19874=>"00000000",
  19875=>"11111110",
  19876=>"11111111",
  19877=>"00000000",
  19878=>"00000001",
  19879=>"00000001",
  19880=>"00000000",
  19881=>"00000110",
  19882=>"11111101",
  19883=>"11111110",
  19884=>"00000011",
  19885=>"11111110",
  19886=>"11111111",
  19887=>"00000010",
  19888=>"00000001",
  19889=>"00000010",
  19890=>"11111110",
  19891=>"00000001",
  19892=>"00000000",
  19893=>"00000001",
  19894=>"00000011",
  19895=>"00000101",
  19896=>"00000011",
  19897=>"11111111",
  19898=>"00000001",
  19899=>"11111110",
  19900=>"00000000",
  19901=>"00000000",
  19902=>"00000001",
  19903=>"11111110",
  19904=>"00000001",
  19905=>"11111110",
  19906=>"11111111",
  19907=>"00000011",
  19908=>"11111110",
  19909=>"00000000",
  19910=>"00000000",
  19911=>"11111011",
  19912=>"00000011",
  19913=>"00000011",
  19914=>"00000001",
  19915=>"00000001",
  19916=>"11111101",
  19917=>"00000001",
  19918=>"11111110",
  19919=>"11111111",
  19920=>"00000001",
  19921=>"00000000",
  19922=>"11111111",
  19923=>"11111110",
  19924=>"11111110",
  19925=>"11111101",
  19926=>"00000010",
  19927=>"00000000",
  19928=>"00000000",
  19929=>"00000001",
  19930=>"00000001",
  19931=>"00000011",
  19932=>"11111111",
  19933=>"00000000",
  19934=>"00000010",
  19935=>"00000010",
  19936=>"00000001",
  19937=>"00000000",
  19938=>"00000001",
  19939=>"11111110",
  19940=>"11111101",
  19941=>"11111111",
  19942=>"11111101",
  19943=>"00000001",
  19944=>"11111100",
  19945=>"00000000",
  19946=>"11111110",
  19947=>"00000001",
  19948=>"11111111",
  19949=>"00000000",
  19950=>"00000001",
  19951=>"00000000",
  19952=>"11111101",
  19953=>"11111110",
  19954=>"11111110",
  19955=>"11111101",
  19956=>"00000000",
  19957=>"00000010",
  19958=>"00000000",
  19959=>"00000010",
  19960=>"00000011",
  19961=>"00000001",
  19962=>"00000010",
  19963=>"00000011",
  19964=>"00000011",
  19965=>"00000001",
  19966=>"00000010",
  19967=>"00000100",
  19968=>"11111101",
  19969=>"00000000",
  19970=>"00000000",
  19971=>"11111110",
  19972=>"00000010",
  19973=>"00000001",
  19974=>"00000010",
  19975=>"00000011",
  19976=>"11111111",
  19977=>"11111110",
  19978=>"11111110",
  19979=>"00000000",
  19980=>"00000010",
  19981=>"00000011",
  19982=>"11111110",
  19983=>"00000100",
  19984=>"11111111",
  19985=>"00000001",
  19986=>"00000010",
  19987=>"11111111",
  19988=>"11111111",
  19989=>"00000001",
  19990=>"00000001",
  19991=>"11111101",
  19992=>"11111111",
  19993=>"00000100",
  19994=>"11111101",
  19995=>"11111111",
  19996=>"11111111",
  19997=>"00000010",
  19998=>"00000010",
  19999=>"00000000",
  20000=>"11111111",
  20001=>"00000010",
  20002=>"00000000",
  20003=>"11111111",
  20004=>"11111111",
  20005=>"11111111",
  20006=>"00000000",
  20007=>"00000001",
  20008=>"00000000",
  20009=>"11111111",
  20010=>"11111101",
  20011=>"11111110",
  20012=>"00000000",
  20013=>"00000010",
  20014=>"11111110",
  20015=>"00000000",
  20016=>"11111111",
  20017=>"11111111",
  20018=>"00000000",
  20019=>"11111101",
  20020=>"00000001",
  20021=>"00000000",
  20022=>"11111110",
  20023=>"11111101",
  20024=>"00000001",
  20025=>"11111110",
  20026=>"11111111",
  20027=>"11111101",
  20028=>"11111110",
  20029=>"11111101",
  20030=>"00000000",
  20031=>"00000000",
  20032=>"00000011",
  20033=>"00000100",
  20034=>"00000100",
  20035=>"11111101",
  20036=>"11111111",
  20037=>"11111110",
  20038=>"00000010",
  20039=>"00000110",
  20040=>"00000000",
  20041=>"11111111",
  20042=>"11111110",
  20043=>"11111110",
  20044=>"11111110",
  20045=>"00000000",
  20046=>"00000010",
  20047=>"00000010",
  20048=>"00000001",
  20049=>"11111110",
  20050=>"00000010",
  20051=>"00000001",
  20052=>"00000000",
  20053=>"11111101",
  20054=>"00000001",
  20055=>"11111101",
  20056=>"11111110",
  20057=>"00000010",
  20058=>"11111111",
  20059=>"11111111",
  20060=>"11111100",
  20061=>"00000010",
  20062=>"11111101",
  20063=>"00000001",
  20064=>"00000001",
  20065=>"00000011",
  20066=>"00000010",
  20067=>"11111111",
  20068=>"11111101",
  20069=>"00000010",
  20070=>"11111110",
  20071=>"00000011",
  20072=>"11111101",
  20073=>"00000011",
  20074=>"00000010",
  20075=>"00000001",
  20076=>"00000011",
  20077=>"00000001",
  20078=>"11111110",
  20079=>"00000000",
  20080=>"00000110",
  20081=>"00000000",
  20082=>"11111110",
  20083=>"11111111",
  20084=>"00000000",
  20085=>"00000001",
  20086=>"00000001",
  20087=>"11111111",
  20088=>"00000011",
  20089=>"00000010",
  20090=>"00000010",
  20091=>"11111111",
  20092=>"00000010",
  20093=>"11111101",
  20094=>"11111110",
  20095=>"00000001",
  20096=>"00000010",
  20097=>"11111110",
  20098=>"00000000",
  20099=>"11111100",
  20100=>"11111111",
  20101=>"00000101",
  20102=>"00000010",
  20103=>"00000000",
  20104=>"11111110",
  20105=>"00000011",
  20106=>"00000001",
  20107=>"11111111",
  20108=>"00000001",
  20109=>"11111111",
  20110=>"00000100",
  20111=>"00000011",
  20112=>"11111111",
  20113=>"11111100",
  20114=>"00000100",
  20115=>"00000001",
  20116=>"00000101",
  20117=>"00000000",
  20118=>"11111110",
  20119=>"00000001",
  20120=>"11111111",
  20121=>"00000000",
  20122=>"00000001",
  20123=>"11111111",
  20124=>"11111111",
  20125=>"11111111",
  20126=>"00000100",
  20127=>"11111110",
  20128=>"00000010",
  20129=>"00000100",
  20130=>"11111111",
  20131=>"11111100",
  20132=>"00000000",
  20133=>"11111110",
  20134=>"00000000",
  20135=>"00000010",
  20136=>"11111110",
  20137=>"11111101",
  20138=>"00000000",
  20139=>"00000000",
  20140=>"00000010",
  20141=>"00000101",
  20142=>"11111110",
  20143=>"11111110",
  20144=>"00000011",
  20145=>"11111101",
  20146=>"00000010",
  20147=>"00000001",
  20148=>"00000001",
  20149=>"11111110",
  20150=>"11111111",
  20151=>"11111110",
  20152=>"11111111",
  20153=>"00000001",
  20154=>"00000010",
  20155=>"00000001",
  20156=>"11111101",
  20157=>"00000000",
  20158=>"11111101",
  20159=>"11111110",
  20160=>"11111111",
  20161=>"11111110",
  20162=>"11111110",
  20163=>"00000010",
  20164=>"00000010",
  20165=>"00000000",
  20166=>"00000001",
  20167=>"00000011",
  20168=>"00000100",
  20169=>"00000001",
  20170=>"00000011",
  20171=>"00000000",
  20172=>"00000001",
  20173=>"00000110",
  20174=>"00000001",
  20175=>"00000010",
  20176=>"11111110",
  20177=>"00000000",
  20178=>"11111111",
  20179=>"00000001",
  20180=>"00000000",
  20181=>"00000010",
  20182=>"11111111",
  20183=>"11111110",
  20184=>"11111110",
  20185=>"11111111",
  20186=>"00000011",
  20187=>"11111111",
  20188=>"11111111",
  20189=>"11111101",
  20190=>"00000000",
  20191=>"00000010",
  20192=>"11111111",
  20193=>"00000000",
  20194=>"00000100",
  20195=>"00000000",
  20196=>"11111111",
  20197=>"00000001",
  20198=>"11111111",
  20199=>"11111110",
  20200=>"00000000",
  20201=>"00000010",
  20202=>"00000011",
  20203=>"00000000",
  20204=>"00000011",
  20205=>"00000000",
  20206=>"00000011",
  20207=>"11111101",
  20208=>"11111101",
  20209=>"00000000",
  20210=>"11111110",
  20211=>"00000010",
  20212=>"11111100",
  20213=>"00000001",
  20214=>"00000011",
  20215=>"11111111",
  20216=>"00000000",
  20217=>"00000101",
  20218=>"00000011",
  20219=>"11111101",
  20220=>"00000010",
  20221=>"11111110",
  20222=>"11111101",
  20223=>"11111111",
  20224=>"00000011",
  20225=>"00000011",
  20226=>"00000000",
  20227=>"11111110",
  20228=>"11111111",
  20229=>"00000010",
  20230=>"00000000",
  20231=>"11111101",
  20232=>"00000011",
  20233=>"11111110",
  20234=>"11111111",
  20235=>"00000011",
  20236=>"00000011",
  20237=>"11111110",
  20238=>"11111101",
  20239=>"00000100",
  20240=>"00000000",
  20241=>"00000010",
  20242=>"00000010",
  20243=>"00000001",
  20244=>"00000001",
  20245=>"00000010",
  20246=>"11111110",
  20247=>"11111110",
  20248=>"00000000",
  20249=>"11111101",
  20250=>"11111110",
  20251=>"11111101",
  20252=>"11111111",
  20253=>"11111111",
  20254=>"00000000",
  20255=>"11111111",
  20256=>"11111110",
  20257=>"11111110",
  20258=>"00000000",
  20259=>"00000010",
  20260=>"11111110",
  20261=>"11111101",
  20262=>"00000010",
  20263=>"11111101",
  20264=>"11111110",
  20265=>"11111110",
  20266=>"00000101",
  20267=>"00000000",
  20268=>"00000001",
  20269=>"11111110",
  20270=>"11111110",
  20271=>"11111111",
  20272=>"11111111",
  20273=>"00000010",
  20274=>"11111101",
  20275=>"11111101",
  20276=>"00000000",
  20277=>"11111111",
  20278=>"11111110",
  20279=>"00000010",
  20280=>"00000001",
  20281=>"00000001",
  20282=>"11111101",
  20283=>"00001000",
  20284=>"11111110",
  20285=>"00000001",
  20286=>"00000000",
  20287=>"11111111",
  20288=>"00000010",
  20289=>"00000001",
  20290=>"11111111",
  20291=>"11111101",
  20292=>"00000001",
  20293=>"11111101",
  20294=>"11111101",
  20295=>"11111110",
  20296=>"00000000",
  20297=>"11111101",
  20298=>"00000001",
  20299=>"00000011",
  20300=>"11111101",
  20301=>"00000010",
  20302=>"11111100",
  20303=>"11111111",
  20304=>"00000001",
  20305=>"11111111",
  20306=>"11111111",
  20307=>"11111110",
  20308=>"00000000",
  20309=>"00000001",
  20310=>"11111110",
  20311=>"11111110",
  20312=>"11111110",
  20313=>"11111110",
  20314=>"11111101",
  20315=>"00000001",
  20316=>"00000010",
  20317=>"11111101",
  20318=>"00000000",
  20319=>"00000010",
  20320=>"11111100",
  20321=>"00000100",
  20322=>"00000001",
  20323=>"00000001",
  20324=>"11111101",
  20325=>"00000001",
  20326=>"00000010",
  20327=>"11111111",
  20328=>"00000010",
  20329=>"11111110",
  20330=>"11111110",
  20331=>"00000011",
  20332=>"11111110",
  20333=>"11111011",
  20334=>"11111110",
  20335=>"00000000",
  20336=>"11111101",
  20337=>"11111111",
  20338=>"00000010",
  20339=>"11111100",
  20340=>"11111110",
  20341=>"00000001",
  20342=>"11111111",
  20343=>"11111110",
  20344=>"11111101",
  20345=>"00000001",
  20346=>"00000000",
  20347=>"00000001",
  20348=>"00000011",
  20349=>"11111111",
  20350=>"00000010",
  20351=>"00000000",
  20352=>"11111111",
  20353=>"11111101",
  20354=>"00000001",
  20355=>"11111111",
  20356=>"11111110",
  20357=>"00000000",
  20358=>"00000000",
  20359=>"11111101",
  20360=>"00000000",
  20361=>"00000001",
  20362=>"00000010",
  20363=>"00000010",
  20364=>"00000100",
  20365=>"11111101",
  20366=>"00000010",
  20367=>"11111111",
  20368=>"00000000",
  20369=>"11111111",
  20370=>"11111111",
  20371=>"00000000",
  20372=>"11111110",
  20373=>"00000000",
  20374=>"00000001",
  20375=>"11111111",
  20376=>"11111100",
  20377=>"11111111",
  20378=>"11111111",
  20379=>"00000101",
  20380=>"00000011",
  20381=>"00000001",
  20382=>"11111111",
  20383=>"00000010",
  20384=>"11111101",
  20385=>"11111101",
  20386=>"11111110",
  20387=>"00000000",
  20388=>"00000000",
  20389=>"00000001",
  20390=>"00000011",
  20391=>"11111101",
  20392=>"00000001",
  20393=>"11111111",
  20394=>"00000000",
  20395=>"00000000",
  20396=>"11111110",
  20397=>"11111110",
  20398=>"00000010",
  20399=>"00000010",
  20400=>"00000001",
  20401=>"11111110",
  20402=>"11111111",
  20403=>"00000011",
  20404=>"00000010",
  20405=>"11111110",
  20406=>"00000000",
  20407=>"00000000",
  20408=>"11111111",
  20409=>"00000001",
  20410=>"00000000",
  20411=>"11111111",
  20412=>"00000000",
  20413=>"11111101",
  20414=>"11111111",
  20415=>"00000010",
  20416=>"11111111",
  20417=>"11111110",
  20418=>"11111111",
  20419=>"00000000",
  20420=>"11111110",
  20421=>"00000001",
  20422=>"00000000",
  20423=>"00000001",
  20424=>"11111101",
  20425=>"11111111",
  20426=>"11111111",
  20427=>"00000001",
  20428=>"00000000",
  20429=>"11111101",
  20430=>"00000001",
  20431=>"11111101",
  20432=>"11111110",
  20433=>"11111101",
  20434=>"11111101",
  20435=>"11111110",
  20436=>"11111111",
  20437=>"00000010",
  20438=>"00000001",
  20439=>"00000001",
  20440=>"11111111",
  20441=>"11111110",
  20442=>"11111110",
  20443=>"00000010",
  20444=>"11111110",
  20445=>"11111110",
  20446=>"00000010",
  20447=>"11111110",
  20448=>"11111111",
  20449=>"11111101",
  20450=>"00000011",
  20451=>"00000011",
  20452=>"00000001",
  20453=>"00000001",
  20454=>"00000011",
  20455=>"11111110",
  20456=>"00000010",
  20457=>"11111101",
  20458=>"00000000",
  20459=>"11111110",
  20460=>"11111111",
  20461=>"11111110",
  20462=>"00000100",
  20463=>"00000001",
  20464=>"11111100",
  20465=>"00000011",
  20466=>"11111111",
  20467=>"00000000",
  20468=>"11111111",
  20469=>"11111111",
  20470=>"11111101",
  20471=>"00000000",
  20472=>"00000000",
  20473=>"11111111",
  20474=>"00000100",
  20475=>"00000010",
  20476=>"00000011",
  20477=>"00000011",
  20478=>"11111111",
  20479=>"11111111",
  20480=>"00000000",
  20481=>"11111111",
  20482=>"11111110",
  20483=>"00000010",
  20484=>"00000110",
  20485=>"00000000",
  20486=>"00000000",
  20487=>"00000000",
  20488=>"00000011",
  20489=>"11111100",
  20490=>"00000010",
  20491=>"11111101",
  20492=>"11111110",
  20493=>"11111111",
  20494=>"00000001",
  20495=>"11111101",
  20496=>"11111110",
  20497=>"11111101",
  20498=>"00000000",
  20499=>"00000000",
  20500=>"00000011",
  20501=>"00000100",
  20502=>"11111111",
  20503=>"11111111",
  20504=>"11111111",
  20505=>"00000011",
  20506=>"11111111",
  20507=>"00000100",
  20508=>"11111111",
  20509=>"00000000",
  20510=>"11111110",
  20511=>"00000100",
  20512=>"00000011",
  20513=>"00000000",
  20514=>"11111111",
  20515=>"00000000",
  20516=>"11111110",
  20517=>"00000010",
  20518=>"00000011",
  20519=>"00000011",
  20520=>"00000011",
  20521=>"00000000",
  20522=>"11111100",
  20523=>"11111110",
  20524=>"11111101",
  20525=>"00000001",
  20526=>"11111111",
  20527=>"11111110",
  20528=>"00000010",
  20529=>"11111101",
  20530=>"00000010",
  20531=>"00000010",
  20532=>"00000010",
  20533=>"00000011",
  20534=>"00000010",
  20535=>"11111111",
  20536=>"00000001",
  20537=>"11111110",
  20538=>"11111111",
  20539=>"11111101",
  20540=>"00000000",
  20541=>"00000000",
  20542=>"00000101",
  20543=>"00000000",
  20544=>"00000110",
  20545=>"11111111",
  20546=>"00000001",
  20547=>"11111110",
  20548=>"11111111",
  20549=>"00000001",
  20550=>"11111101",
  20551=>"11111101",
  20552=>"11111111",
  20553=>"11111111",
  20554=>"11111111",
  20555=>"00000000",
  20556=>"00000001",
  20557=>"00000100",
  20558=>"00000010",
  20559=>"00000001",
  20560=>"00000010",
  20561=>"11111110",
  20562=>"11111110",
  20563=>"11111111",
  20564=>"11111110",
  20565=>"11111101",
  20566=>"00000010",
  20567=>"00000001",
  20568=>"11111111",
  20569=>"11111100",
  20570=>"00000001",
  20571=>"11111100",
  20572=>"00000000",
  20573=>"00000011",
  20574=>"11111111",
  20575=>"11111111",
  20576=>"11111101",
  20577=>"11111111",
  20578=>"00000010",
  20579=>"00000000",
  20580=>"00000100",
  20581=>"00000010",
  20582=>"00000000",
  20583=>"11111111",
  20584=>"00000010",
  20585=>"00000111",
  20586=>"00000000",
  20587=>"00000000",
  20588=>"11111111",
  20589=>"11111110",
  20590=>"11111111",
  20591=>"00000000",
  20592=>"00000010",
  20593=>"00000011",
  20594=>"11111101",
  20595=>"00000001",
  20596=>"00000100",
  20597=>"00000001",
  20598=>"11111111",
  20599=>"11111111",
  20600=>"00000001",
  20601=>"11111101",
  20602=>"00000001",
  20603=>"00000001",
  20604=>"00000101",
  20605=>"00000111",
  20606=>"00000010",
  20607=>"11111110",
  20608=>"11111110",
  20609=>"00000010",
  20610=>"00000000",
  20611=>"11111111",
  20612=>"11111111",
  20613=>"11111110",
  20614=>"00000001",
  20615=>"00000011",
  20616=>"11111110",
  20617=>"11111111",
  20618=>"00000001",
  20619=>"00000101",
  20620=>"00000000",
  20621=>"00000011",
  20622=>"11111101",
  20623=>"11111100",
  20624=>"00000000",
  20625=>"11111111",
  20626=>"00000001",
  20627=>"00000100",
  20628=>"11111100",
  20629=>"11111101",
  20630=>"00000110",
  20631=>"00000001",
  20632=>"11111101",
  20633=>"11111111",
  20634=>"11111111",
  20635=>"11111101",
  20636=>"00000000",
  20637=>"00000000",
  20638=>"00000000",
  20639=>"00000010",
  20640=>"00000001",
  20641=>"00000100",
  20642=>"11111101",
  20643=>"00000001",
  20644=>"11111111",
  20645=>"00000001",
  20646=>"00000010",
  20647=>"11111110",
  20648=>"11111101",
  20649=>"11111111",
  20650=>"11111110",
  20651=>"00000010",
  20652=>"11111110",
  20653=>"00000000",
  20654=>"00000010",
  20655=>"11111101",
  20656=>"00000000",
  20657=>"00000000",
  20658=>"00000001",
  20659=>"00000011",
  20660=>"00000001",
  20661=>"00000001",
  20662=>"00000000",
  20663=>"00000001",
  20664=>"11111110",
  20665=>"00000011",
  20666=>"11111101",
  20667=>"00000000",
  20668=>"11111110",
  20669=>"00000001",
  20670=>"00000000",
  20671=>"00000011",
  20672=>"00000000",
  20673=>"11111111",
  20674=>"00000001",
  20675=>"00000001",
  20676=>"11111101",
  20677=>"00000010",
  20678=>"11111101",
  20679=>"11111101",
  20680=>"11111100",
  20681=>"11111110",
  20682=>"00000010",
  20683=>"11111111",
  20684=>"11111111",
  20685=>"11111111",
  20686=>"00000000",
  20687=>"11111100",
  20688=>"00000010",
  20689=>"11111110",
  20690=>"00000010",
  20691=>"00000000",
  20692=>"00000011",
  20693=>"11111101",
  20694=>"11111110",
  20695=>"11111100",
  20696=>"11111110",
  20697=>"00000000",
  20698=>"00000010",
  20699=>"11111111",
  20700=>"00000010",
  20701=>"00000010",
  20702=>"11111111",
  20703=>"00000000",
  20704=>"11111110",
  20705=>"11111110",
  20706=>"11111111",
  20707=>"11111111",
  20708=>"00000011",
  20709=>"11111110",
  20710=>"11111110",
  20711=>"00000001",
  20712=>"11111111",
  20713=>"11111101",
  20714=>"11111111",
  20715=>"00000010",
  20716=>"00000001",
  20717=>"00000000",
  20718=>"11111110",
  20719=>"00000000",
  20720=>"00000011",
  20721=>"00000010",
  20722=>"00000001",
  20723=>"00000100",
  20724=>"11111110",
  20725=>"11111101",
  20726=>"11111101",
  20727=>"11111111",
  20728=>"11111110",
  20729=>"00000001",
  20730=>"00000100",
  20731=>"11111111",
  20732=>"00000001",
  20733=>"11111110",
  20734=>"00000011",
  20735=>"00000010",
  20736=>"00000001",
  20737=>"00000010",
  20738=>"11111101",
  20739=>"00000000",
  20740=>"11111110",
  20741=>"00000000",
  20742=>"11111110",
  20743=>"11111111",
  20744=>"00000101",
  20745=>"11111111",
  20746=>"00000000",
  20747=>"11111111",
  20748=>"11111110",
  20749=>"00000001",
  20750=>"00000010",
  20751=>"11111110",
  20752=>"00000000",
  20753=>"00000000",
  20754=>"11111110",
  20755=>"11111111",
  20756=>"11111111",
  20757=>"11111011",
  20758=>"00000011",
  20759=>"00000100",
  20760=>"00000011",
  20761=>"00000010",
  20762=>"11111110",
  20763=>"00000000",
  20764=>"11111110",
  20765=>"00000010",
  20766=>"11111111",
  20767=>"00000000",
  20768=>"00000010",
  20769=>"00000001",
  20770=>"00000101",
  20771=>"00000101",
  20772=>"11111110",
  20773=>"11111101",
  20774=>"00000000",
  20775=>"11111101",
  20776=>"00000010",
  20777=>"00000000",
  20778=>"00000000",
  20779=>"00000010",
  20780=>"00000001",
  20781=>"11111110",
  20782=>"00000010",
  20783=>"11111110",
  20784=>"11111111",
  20785=>"00000001",
  20786=>"00000100",
  20787=>"11111110",
  20788=>"00000010",
  20789=>"00000001",
  20790=>"11111101",
  20791=>"00000000",
  20792=>"00000000",
  20793=>"11111101",
  20794=>"00000011",
  20795=>"00000010",
  20796=>"11111101",
  20797=>"11111111",
  20798=>"00000000",
  20799=>"00000010",
  20800=>"00000010",
  20801=>"11111111",
  20802=>"00000010",
  20803=>"11111110",
  20804=>"00000001",
  20805=>"11111111",
  20806=>"11111110",
  20807=>"11111101",
  20808=>"00000001",
  20809=>"00000000",
  20810=>"00000011",
  20811=>"11111111",
  20812=>"00000010",
  20813=>"00000001",
  20814=>"00000000",
  20815=>"11111110",
  20816=>"11111101",
  20817=>"00000001",
  20818=>"00000000",
  20819=>"11111101",
  20820=>"11111110",
  20821=>"11111111",
  20822=>"00000000",
  20823=>"00000001",
  20824=>"00000010",
  20825=>"11111111",
  20826=>"00000000",
  20827=>"00000000",
  20828=>"00000001",
  20829=>"00000100",
  20830=>"00000000",
  20831=>"00000001",
  20832=>"00000000",
  20833=>"11111110",
  20834=>"00000100",
  20835=>"00000100",
  20836=>"00000100",
  20837=>"11111110",
  20838=>"11111100",
  20839=>"00000000",
  20840=>"00000010",
  20841=>"00000010",
  20842=>"00000010",
  20843=>"00000000",
  20844=>"11111101",
  20845=>"00000011",
  20846=>"00000010",
  20847=>"11111111",
  20848=>"00000010",
  20849=>"00000000",
  20850=>"00000000",
  20851=>"11111101",
  20852=>"11111101",
  20853=>"11111101",
  20854=>"00000010",
  20855=>"00000010",
  20856=>"00000001",
  20857=>"00000001",
  20858=>"00000000",
  20859=>"11111110",
  20860=>"00000000",
  20861=>"11111101",
  20862=>"11111111",
  20863=>"00000110",
  20864=>"00000000",
  20865=>"11111101",
  20866=>"00000010",
  20867=>"00000000",
  20868=>"11111110",
  20869=>"00000100",
  20870=>"00000110",
  20871=>"00000011",
  20872=>"00000010",
  20873=>"00000011",
  20874=>"00000011",
  20875=>"00000100",
  20876=>"11111110",
  20877=>"00000001",
  20878=>"11111111",
  20879=>"11111101",
  20880=>"11111110",
  20881=>"00000001",
  20882=>"00000000",
  20883=>"11111110",
  20884=>"00000001",
  20885=>"11111111",
  20886=>"00000010",
  20887=>"00000000",
  20888=>"00000010",
  20889=>"11111110",
  20890=>"00000001",
  20891=>"11111111",
  20892=>"11111111",
  20893=>"11111100",
  20894=>"11111111",
  20895=>"11111110",
  20896=>"11111110",
  20897=>"11111110",
  20898=>"11111111",
  20899=>"11111110",
  20900=>"11111101",
  20901=>"11111111",
  20902=>"11111110",
  20903=>"00000001",
  20904=>"11111110",
  20905=>"00000010",
  20906=>"00000000",
  20907=>"11111111",
  20908=>"00000010",
  20909=>"00000100",
  20910=>"00000001",
  20911=>"00000000",
  20912=>"11111110",
  20913=>"00001000",
  20914=>"00000000",
  20915=>"11111101",
  20916=>"11111110",
  20917=>"00000001",
  20918=>"11111111",
  20919=>"11111101",
  20920=>"00000011",
  20921=>"11111110",
  20922=>"11111111",
  20923=>"11111111",
  20924=>"11111111",
  20925=>"00000000",
  20926=>"00000001",
  20927=>"11111111",
  20928=>"00000110",
  20929=>"00000001",
  20930=>"00000010",
  20931=>"00000100",
  20932=>"11111101",
  20933=>"11111101",
  20934=>"00000010",
  20935=>"00000000",
  20936=>"11111100",
  20937=>"11111111",
  20938=>"11111101",
  20939=>"00000000",
  20940=>"11111100",
  20941=>"00000001",
  20942=>"00000110",
  20943=>"00000001",
  20944=>"00000001",
  20945=>"00000011",
  20946=>"11111111",
  20947=>"00000001",
  20948=>"11111110",
  20949=>"00000010",
  20950=>"00000101",
  20951=>"00000100",
  20952=>"11111110",
  20953=>"11111111",
  20954=>"11111111",
  20955=>"11111101",
  20956=>"00000010",
  20957=>"00000010",
  20958=>"00000001",
  20959=>"00000001",
  20960=>"00000000",
  20961=>"11111111",
  20962=>"00000000",
  20963=>"00000011",
  20964=>"00000000",
  20965=>"11111111",
  20966=>"11111111",
  20967=>"00000000",
  20968=>"00000000",
  20969=>"00000001",
  20970=>"11111100",
  20971=>"00000101",
  20972=>"11111110",
  20973=>"00000111",
  20974=>"00000000",
  20975=>"00000001",
  20976=>"00000001",
  20977=>"00000110",
  20978=>"00000000",
  20979=>"00000001",
  20980=>"00000001",
  20981=>"11111111",
  20982=>"00000000",
  20983=>"00000011",
  20984=>"11111111",
  20985=>"00000010",
  20986=>"00000100",
  20987=>"11111110",
  20988=>"00000001",
  20989=>"00000001",
  20990=>"00000011",
  20991=>"11111110",
  20992=>"11111101",
  20993=>"00000000",
  20994=>"11111101",
  20995=>"00000000",
  20996=>"00000101",
  20997=>"00000010",
  20998=>"11111101",
  20999=>"00000000",
  21000=>"00000101",
  21001=>"11111110",
  21002=>"11111111",
  21003=>"11111110",
  21004=>"11111100",
  21005=>"00000000",
  21006=>"00000010",
  21007=>"00000000",
  21008=>"11111110",
  21009=>"11111110",
  21010=>"11111101",
  21011=>"00000001",
  21012=>"00000001",
  21013=>"11111110",
  21014=>"00000000",
  21015=>"11111110",
  21016=>"00000010",
  21017=>"00000000",
  21018=>"00000000",
  21019=>"11111111",
  21020=>"11111110",
  21021=>"00000001",
  21022=>"00000001",
  21023=>"11111100",
  21024=>"11111100",
  21025=>"00000010",
  21026=>"00000000",
  21027=>"00000110",
  21028=>"11111110",
  21029=>"00000001",
  21030=>"11111111",
  21031=>"11111110",
  21032=>"00000001",
  21033=>"00000001",
  21034=>"11111110",
  21035=>"00000001",
  21036=>"11111101",
  21037=>"11111101",
  21038=>"00000010",
  21039=>"11111111",
  21040=>"11111111",
  21041=>"00000100",
  21042=>"00000000",
  21043=>"11111110",
  21044=>"00000011",
  21045=>"00000010",
  21046=>"11111110",
  21047=>"00000000",
  21048=>"00000000",
  21049=>"00000010",
  21050=>"11111111",
  21051=>"00000001",
  21052=>"11111111",
  21053=>"11111101",
  21054=>"00000011",
  21055=>"11111110",
  21056=>"00000010",
  21057=>"00000011",
  21058=>"11111111",
  21059=>"11111101",
  21060=>"00000000",
  21061=>"00000000",
  21062=>"11111110",
  21063=>"00000000",
  21064=>"11111101",
  21065=>"00000001",
  21066=>"11111101",
  21067=>"11111111",
  21068=>"11111111",
  21069=>"00000000",
  21070=>"11111111",
  21071=>"00000011",
  21072=>"11111111",
  21073=>"00000001",
  21074=>"00000011",
  21075=>"11111110",
  21076=>"00000001",
  21077=>"11111111",
  21078=>"11111101",
  21079=>"00000011",
  21080=>"00000100",
  21081=>"11111111",
  21082=>"11111111",
  21083=>"11111111",
  21084=>"11111111",
  21085=>"00000011",
  21086=>"00000000",
  21087=>"11111110",
  21088=>"00000001",
  21089=>"00000010",
  21090=>"11111110",
  21091=>"11111110",
  21092=>"11111101",
  21093=>"11111111",
  21094=>"00000001",
  21095=>"11111110",
  21096=>"00000010",
  21097=>"00000001",
  21098=>"11111111",
  21099=>"00000000",
  21100=>"11111110",
  21101=>"00000010",
  21102=>"11111110",
  21103=>"00000011",
  21104=>"00000100",
  21105=>"00000000",
  21106=>"00000010",
  21107=>"11111111",
  21108=>"00000001",
  21109=>"00000010",
  21110=>"11111110",
  21111=>"11111111",
  21112=>"11111111",
  21113=>"00000000",
  21114=>"00000101",
  21115=>"00000000",
  21116=>"11111110",
  21117=>"11111111",
  21118=>"00000000",
  21119=>"00000011",
  21120=>"11111111",
  21121=>"00000001",
  21122=>"11111101",
  21123=>"11111111",
  21124=>"11111110",
  21125=>"00000000",
  21126=>"00000100",
  21127=>"00000100",
  21128=>"11111111",
  21129=>"11111101",
  21130=>"00000000",
  21131=>"00000001",
  21132=>"00000011",
  21133=>"00000010",
  21134=>"11111110",
  21135=>"11111111",
  21136=>"11111110",
  21137=>"11111101",
  21138=>"00000001",
  21139=>"00000000",
  21140=>"00000011",
  21141=>"11111100",
  21142=>"11111101",
  21143=>"11111101",
  21144=>"11111111",
  21145=>"00000001",
  21146=>"11111111",
  21147=>"00000010",
  21148=>"11111110",
  21149=>"11111110",
  21150=>"11111111",
  21151=>"00000000",
  21152=>"00000010",
  21153=>"11111111",
  21154=>"00000101",
  21155=>"11111110",
  21156=>"11111111",
  21157=>"00000100",
  21158=>"00000101",
  21159=>"00000000",
  21160=>"00000011",
  21161=>"11111110",
  21162=>"11111111",
  21163=>"11111111",
  21164=>"11111101",
  21165=>"11111111",
  21166=>"00000010",
  21167=>"11111101",
  21168=>"11111111",
  21169=>"00000010",
  21170=>"00000000",
  21171=>"00000000",
  21172=>"00000011",
  21173=>"00000011",
  21174=>"11111111",
  21175=>"11111110",
  21176=>"00000000",
  21177=>"00000010",
  21178=>"00000011",
  21179=>"00000011",
  21180=>"11111100",
  21181=>"11111111",
  21182=>"11111110",
  21183=>"00000011",
  21184=>"11111101",
  21185=>"11111101",
  21186=>"11111101",
  21187=>"11111110",
  21188=>"00000001",
  21189=>"00000011",
  21190=>"00000011",
  21191=>"00000000",
  21192=>"11111111",
  21193=>"11111110",
  21194=>"00000101",
  21195=>"11111111",
  21196=>"00000001",
  21197=>"00000010",
  21198=>"11111111",
  21199=>"11111110",
  21200=>"00000001",
  21201=>"11111100",
  21202=>"11111111",
  21203=>"11111110",
  21204=>"00000000",
  21205=>"00000001",
  21206=>"00000001",
  21207=>"11111101",
  21208=>"00000001",
  21209=>"00000001",
  21210=>"11111110",
  21211=>"00000001",
  21212=>"11111101",
  21213=>"00000000",
  21214=>"00000000",
  21215=>"11111101",
  21216=>"00000001",
  21217=>"00000000",
  21218=>"00000000",
  21219=>"11111111",
  21220=>"00000001",
  21221=>"11111111",
  21222=>"00000010",
  21223=>"00000010",
  21224=>"00000001",
  21225=>"00000001",
  21226=>"11111111",
  21227=>"11111111",
  21228=>"00000001",
  21229=>"00000001",
  21230=>"11111110",
  21231=>"11111101",
  21232=>"00000010",
  21233=>"00000001",
  21234=>"11111111",
  21235=>"11111111",
  21236=>"11111111",
  21237=>"11111100",
  21238=>"00000001",
  21239=>"11111101",
  21240=>"00000001",
  21241=>"11111111",
  21242=>"00000001",
  21243=>"00000000",
  21244=>"11111111",
  21245=>"00000010",
  21246=>"00000011",
  21247=>"00000001",
  21248=>"11111011",
  21249=>"11111111",
  21250=>"00000000",
  21251=>"00000000",
  21252=>"00000100",
  21253=>"11111111",
  21254=>"00000011",
  21255=>"00000000",
  21256=>"00000011",
  21257=>"00000010",
  21258=>"00000001",
  21259=>"11111111",
  21260=>"00000010",
  21261=>"00000000",
  21262=>"11111111",
  21263=>"11111111",
  21264=>"00000010",
  21265=>"00000010",
  21266=>"00000011",
  21267=>"11111110",
  21268=>"00000010",
  21269=>"11111110",
  21270=>"11111111",
  21271=>"11111111",
  21272=>"11111110",
  21273=>"11111110",
  21274=>"11111111",
  21275=>"11111110",
  21276=>"00000001",
  21277=>"11111111",
  21278=>"11111101",
  21279=>"00000000",
  21280=>"00000001",
  21281=>"11111110",
  21282=>"11111110",
  21283=>"00000001",
  21284=>"00000000",
  21285=>"00000011",
  21286=>"11111100",
  21287=>"00000001",
  21288=>"00000000",
  21289=>"00000101",
  21290=>"00000010",
  21291=>"00000000",
  21292=>"11111110",
  21293=>"00000000",
  21294=>"00000010",
  21295=>"11111101",
  21296=>"11111101",
  21297=>"00000001",
  21298=>"11111111",
  21299=>"00000010",
  21300=>"00000010",
  21301=>"00000010",
  21302=>"00000001",
  21303=>"00000011",
  21304=>"11111101",
  21305=>"00000010",
  21306=>"11111110",
  21307=>"11111111",
  21308=>"00000011",
  21309=>"11111110",
  21310=>"11111110",
  21311=>"11111111",
  21312=>"00000011",
  21313=>"11111111",
  21314=>"11111110",
  21315=>"11111101",
  21316=>"11111110",
  21317=>"00000000",
  21318=>"00000001",
  21319=>"00000011",
  21320=>"11111101",
  21321=>"00000100",
  21322=>"11111110",
  21323=>"00000000",
  21324=>"11111110",
  21325=>"11111101",
  21326=>"00000001",
  21327=>"11111110",
  21328=>"00000001",
  21329=>"00000010",
  21330=>"11111110",
  21331=>"00000000",
  21332=>"00000000",
  21333=>"00000001",
  21334=>"00000000",
  21335=>"11111111",
  21336=>"00000000",
  21337=>"00000010",
  21338=>"11111110",
  21339=>"11111110",
  21340=>"00000010",
  21341=>"11111101",
  21342=>"00000010",
  21343=>"00000000",
  21344=>"00000000",
  21345=>"00000001",
  21346=>"00000010",
  21347=>"00000000",
  21348=>"00000100",
  21349=>"11111111",
  21350=>"00000001",
  21351=>"11111110",
  21352=>"11111110",
  21353=>"00000001",
  21354=>"00000000",
  21355=>"11111110",
  21356=>"00000001",
  21357=>"00000001",
  21358=>"00000000",
  21359=>"11111101",
  21360=>"11111111",
  21361=>"00000001",
  21362=>"00000010",
  21363=>"11111100",
  21364=>"11111110",
  21365=>"11111111",
  21366=>"00000010",
  21367=>"00000001",
  21368=>"00000011",
  21369=>"00000010",
  21370=>"00000000",
  21371=>"00000001",
  21372=>"00000101",
  21373=>"11111111",
  21374=>"11111111",
  21375=>"00000000",
  21376=>"11111110",
  21377=>"11111100",
  21378=>"00000010",
  21379=>"11111101",
  21380=>"00000010",
  21381=>"11111111",
  21382=>"11111101",
  21383=>"00000000",
  21384=>"00000010",
  21385=>"00000100",
  21386=>"00000011",
  21387=>"00000000",
  21388=>"11111111",
  21389=>"11111111",
  21390=>"00000001",
  21391=>"00000010",
  21392=>"11111110",
  21393=>"00000001",
  21394=>"00000101",
  21395=>"11111111",
  21396=>"00000000",
  21397=>"00000000",
  21398=>"00000011",
  21399=>"11111111",
  21400=>"11111111",
  21401=>"00000011",
  21402=>"11111101",
  21403=>"11111110",
  21404=>"00000110",
  21405=>"00000001",
  21406=>"00000011",
  21407=>"00000001",
  21408=>"11111110",
  21409=>"00000011",
  21410=>"00000010",
  21411=>"00000010",
  21412=>"11111101",
  21413=>"11111111",
  21414=>"00000000",
  21415=>"00000001",
  21416=>"00000001",
  21417=>"00000001",
  21418=>"11111110",
  21419=>"11111101",
  21420=>"00000010",
  21421=>"11111110",
  21422=>"00000100",
  21423=>"11111101",
  21424=>"11111111",
  21425=>"00000011",
  21426=>"11111111",
  21427=>"00000011",
  21428=>"00000010",
  21429=>"11111110",
  21430=>"00000000",
  21431=>"00000011",
  21432=>"00000110",
  21433=>"00000000",
  21434=>"11111110",
  21435=>"00000010",
  21436=>"00000011",
  21437=>"11111100",
  21438=>"00000001",
  21439=>"11111111",
  21440=>"00000001",
  21441=>"00000001",
  21442=>"11111111",
  21443=>"00000010",
  21444=>"00000011",
  21445=>"00000011",
  21446=>"00000010",
  21447=>"00000001",
  21448=>"11111111",
  21449=>"11111101",
  21450=>"00000001",
  21451=>"11111111",
  21452=>"11111101",
  21453=>"00000001",
  21454=>"11111110",
  21455=>"00000000",
  21456=>"00000000",
  21457=>"00000101",
  21458=>"11111111",
  21459=>"11111110",
  21460=>"11111110",
  21461=>"00000000",
  21462=>"11111101",
  21463=>"11111101",
  21464=>"11111110",
  21465=>"11111111",
  21466=>"00000001",
  21467=>"11111111",
  21468=>"11111111",
  21469=>"00000010",
  21470=>"11111111",
  21471=>"11111101",
  21472=>"11111111",
  21473=>"00000001",
  21474=>"00000010",
  21475=>"11111110",
  21476=>"11111111",
  21477=>"00000001",
  21478=>"00000010",
  21479=>"00000110",
  21480=>"00000011",
  21481=>"11111111",
  21482=>"11111101",
  21483=>"00000010",
  21484=>"00000011",
  21485=>"11111111",
  21486=>"00000011",
  21487=>"00000001",
  21488=>"11111110",
  21489=>"11111110",
  21490=>"00000100",
  21491=>"11111111",
  21492=>"00000010",
  21493=>"00000001",
  21494=>"11111101",
  21495=>"11111110",
  21496=>"11111111",
  21497=>"11111110",
  21498=>"11111110",
  21499=>"00000001",
  21500=>"00000010",
  21501=>"00000001",
  21502=>"00000100",
  21503=>"00000010",
  21504=>"11111111",
  21505=>"00000001",
  21506=>"11111110",
  21507=>"00000001",
  21508=>"11111110",
  21509=>"00000001",
  21510=>"11111111",
  21511=>"00000010",
  21512=>"11111110",
  21513=>"11111110",
  21514=>"00000010",
  21515=>"11111110",
  21516=>"00000001",
  21517=>"11111110",
  21518=>"00000000",
  21519=>"11111101",
  21520=>"00000000",
  21521=>"00000000",
  21522=>"11111111",
  21523=>"11111111",
  21524=>"11111100",
  21525=>"00000010",
  21526=>"11111111",
  21527=>"11111110",
  21528=>"00000001",
  21529=>"00000001",
  21530=>"00000000",
  21531=>"00000000",
  21532=>"00000000",
  21533=>"11111111",
  21534=>"00000000",
  21535=>"00000010",
  21536=>"00000001",
  21537=>"00000000",
  21538=>"11111110",
  21539=>"00000010",
  21540=>"11111111",
  21541=>"00000011",
  21542=>"00000010",
  21543=>"00000000",
  21544=>"11111101",
  21545=>"11111111",
  21546=>"00000010",
  21547=>"00000010",
  21548=>"00000001",
  21549=>"11111111",
  21550=>"00000011",
  21551=>"11111101",
  21552=>"00000001",
  21553=>"11111111",
  21554=>"11111111",
  21555=>"00000100",
  21556=>"11111110",
  21557=>"00000011",
  21558=>"00000001",
  21559=>"00000010",
  21560=>"11111111",
  21561=>"11111111",
  21562=>"11111111",
  21563=>"00000010",
  21564=>"00000001",
  21565=>"00000011",
  21566=>"00000000",
  21567=>"00000000",
  21568=>"00000000",
  21569=>"00000010",
  21570=>"00000000",
  21571=>"00000100",
  21572=>"00000000",
  21573=>"11111111",
  21574=>"00000001",
  21575=>"00000001",
  21576=>"00000001",
  21577=>"11111110",
  21578=>"00000000",
  21579=>"00000000",
  21580=>"00000000",
  21581=>"00000000",
  21582=>"00000000",
  21583=>"11111110",
  21584=>"00000011",
  21585=>"00000011",
  21586=>"00000010",
  21587=>"11111110",
  21588=>"11111111",
  21589=>"00000001",
  21590=>"00000101",
  21591=>"00000010",
  21592=>"11111110",
  21593=>"00000001",
  21594=>"00000001",
  21595=>"00000110",
  21596=>"11111111",
  21597=>"11111110",
  21598=>"11111111",
  21599=>"00000001",
  21600=>"00000101",
  21601=>"00000001",
  21602=>"00000000",
  21603=>"11111111",
  21604=>"11111101",
  21605=>"11111110",
  21606=>"11111101",
  21607=>"00000001",
  21608=>"11111111",
  21609=>"00000000",
  21610=>"11111110",
  21611=>"00000001",
  21612=>"11111110",
  21613=>"00000010",
  21614=>"00000001",
  21615=>"11111110",
  21616=>"00000001",
  21617=>"00000001",
  21618=>"11111101",
  21619=>"11111110",
  21620=>"11111111",
  21621=>"11111110",
  21622=>"11111101",
  21623=>"00000000",
  21624=>"00000001",
  21625=>"00000000",
  21626=>"11111110",
  21627=>"00000010",
  21628=>"00000001",
  21629=>"00000001",
  21630=>"00000000",
  21631=>"00000000",
  21632=>"00000000",
  21633=>"11111110",
  21634=>"00000010",
  21635=>"00000000",
  21636=>"11111111",
  21637=>"11111110",
  21638=>"11111111",
  21639=>"11111111",
  21640=>"00000010",
  21641=>"00000000",
  21642=>"00000000",
  21643=>"00000001",
  21644=>"00000000",
  21645=>"11111110",
  21646=>"11111110",
  21647=>"11111110",
  21648=>"00000011",
  21649=>"11111101",
  21650=>"11111111",
  21651=>"11111111",
  21652=>"11111110",
  21653=>"00000000",
  21654=>"00000100",
  21655=>"00000011",
  21656=>"11111100",
  21657=>"11111110",
  21658=>"00000000",
  21659=>"00000001",
  21660=>"00000010",
  21661=>"11111110",
  21662=>"11111111",
  21663=>"00000010",
  21664=>"11111110",
  21665=>"11111110",
  21666=>"11111101",
  21667=>"00000010",
  21668=>"11111111",
  21669=>"11111111",
  21670=>"11111110",
  21671=>"11111101",
  21672=>"00000010",
  21673=>"00000000",
  21674=>"00000010",
  21675=>"11111101",
  21676=>"00000001",
  21677=>"00000010",
  21678=>"11111110",
  21679=>"00000010",
  21680=>"11111101",
  21681=>"00000000",
  21682=>"11111111",
  21683=>"11111111",
  21684=>"00000000",
  21685=>"11111100",
  21686=>"11111110",
  21687=>"00000010",
  21688=>"11111111",
  21689=>"00000010",
  21690=>"00000000",
  21691=>"11111111",
  21692=>"00000001",
  21693=>"11111101",
  21694=>"00000010",
  21695=>"00000100",
  21696=>"00000000",
  21697=>"00000001",
  21698=>"00000001",
  21699=>"00000010",
  21700=>"11111111",
  21701=>"00000011",
  21702=>"00000011",
  21703=>"00000011",
  21704=>"11111111",
  21705=>"00000010",
  21706=>"11111110",
  21707=>"11111111",
  21708=>"00000101",
  21709=>"11111111",
  21710=>"11111111",
  21711=>"00000001",
  21712=>"00000001",
  21713=>"00000000",
  21714=>"11111110",
  21715=>"00000010",
  21716=>"00000000",
  21717=>"11111111",
  21718=>"00000000",
  21719=>"00000001",
  21720=>"00000010",
  21721=>"11111110",
  21722=>"11111110",
  21723=>"00000010",
  21724=>"11111111",
  21725=>"00000001",
  21726=>"00000000",
  21727=>"00000001",
  21728=>"00000010",
  21729=>"11111110",
  21730=>"00000001",
  21731=>"00000010",
  21732=>"11111110",
  21733=>"00000000",
  21734=>"00000100",
  21735=>"00000001",
  21736=>"11111111",
  21737=>"00000011",
  21738=>"00000011",
  21739=>"00000010",
  21740=>"11111110",
  21741=>"11111110",
  21742=>"00000010",
  21743=>"11111101",
  21744=>"00000001",
  21745=>"00000011",
  21746=>"00000010",
  21747=>"00000011",
  21748=>"11111111",
  21749=>"11111101",
  21750=>"00000010",
  21751=>"00000000",
  21752=>"11111111",
  21753=>"00000001",
  21754=>"00000010",
  21755=>"00000000",
  21756=>"00000000",
  21757=>"11111111",
  21758=>"11111101",
  21759=>"11111110",
  21760=>"00000010",
  21761=>"00000000",
  21762=>"00000100",
  21763=>"00000001",
  21764=>"00000010",
  21765=>"00000010",
  21766=>"11111111",
  21767=>"11111101",
  21768=>"00000000",
  21769=>"11111111",
  21770=>"00000010",
  21771=>"00000010",
  21772=>"00000000",
  21773=>"00000011",
  21774=>"00000010",
  21775=>"00000001",
  21776=>"00000001",
  21777=>"11111111",
  21778=>"00000010",
  21779=>"00000010",
  21780=>"00000000",
  21781=>"00000000",
  21782=>"11111101",
  21783=>"00000010",
  21784=>"11111111",
  21785=>"00000001",
  21786=>"00000000",
  21787=>"00000010",
  21788=>"11111111",
  21789=>"00000010",
  21790=>"11111110",
  21791=>"00000011",
  21792=>"11111101",
  21793=>"11111110",
  21794=>"00000000",
  21795=>"00000011",
  21796=>"00000011",
  21797=>"00000100",
  21798=>"00000011",
  21799=>"00000000",
  21800=>"11111110",
  21801=>"00000010",
  21802=>"00000100",
  21803=>"11111111",
  21804=>"00000001",
  21805=>"00000001",
  21806=>"11111111",
  21807=>"11111110",
  21808=>"11111111",
  21809=>"11111111",
  21810=>"11111101",
  21811=>"00000010",
  21812=>"00000001",
  21813=>"11111110",
  21814=>"00000010",
  21815=>"00000000",
  21816=>"00000010",
  21817=>"00000001",
  21818=>"11111101",
  21819=>"11111110",
  21820=>"00000010",
  21821=>"11111110",
  21822=>"11111110",
  21823=>"00000001",
  21824=>"11111111",
  21825=>"00000010",
  21826=>"00000001",
  21827=>"11111101",
  21828=>"00000001",
  21829=>"00000010",
  21830=>"11111101",
  21831=>"00000010",
  21832=>"00000000",
  21833=>"11111111",
  21834=>"11111111",
  21835=>"11111110",
  21836=>"11111101",
  21837=>"00000001",
  21838=>"11111110",
  21839=>"11111111",
  21840=>"11111101",
  21841=>"00000000",
  21842=>"11111101",
  21843=>"00000001",
  21844=>"00000000",
  21845=>"00000010",
  21846=>"11111101",
  21847=>"11111111",
  21848=>"11111101",
  21849=>"11111101",
  21850=>"00000001",
  21851=>"00000010",
  21852=>"00000000",
  21853=>"00000010",
  21854=>"00000001",
  21855=>"00000001",
  21856=>"00000001",
  21857=>"11111111",
  21858=>"00000000",
  21859=>"00000000",
  21860=>"11111101",
  21861=>"00000001",
  21862=>"11111101",
  21863=>"00000001",
  21864=>"11111101",
  21865=>"00000000",
  21866=>"00000010",
  21867=>"11111101",
  21868=>"11111110",
  21869=>"11111111",
  21870=>"11111110",
  21871=>"11111111",
  21872=>"00000000",
  21873=>"11111111",
  21874=>"11111110",
  21875=>"11111100",
  21876=>"11111110",
  21877=>"11111110",
  21878=>"11111111",
  21879=>"11111111",
  21880=>"11111110",
  21881=>"11111110",
  21882=>"11111110",
  21883=>"00000000",
  21884=>"00000011",
  21885=>"00000001",
  21886=>"00000010",
  21887=>"00000000",
  21888=>"00000000",
  21889=>"11111111",
  21890=>"00000010",
  21891=>"00000000",
  21892=>"11111111",
  21893=>"11111101",
  21894=>"11111111",
  21895=>"11111111",
  21896=>"00000001",
  21897=>"00000010",
  21898=>"11111110",
  21899=>"00000001",
  21900=>"11111110",
  21901=>"00000000",
  21902=>"11111110",
  21903=>"00000010",
  21904=>"00000010",
  21905=>"11111111",
  21906=>"00000010",
  21907=>"11111110",
  21908=>"00000001",
  21909=>"11111101",
  21910=>"00000000",
  21911=>"00000011",
  21912=>"11111110",
  21913=>"11111111",
  21914=>"00000010",
  21915=>"11111110",
  21916=>"11111111",
  21917=>"11111111",
  21918=>"00000001",
  21919=>"00000010",
  21920=>"00000011",
  21921=>"00000000",
  21922=>"11111110",
  21923=>"11111101",
  21924=>"00000000",
  21925=>"11111111",
  21926=>"11111111",
  21927=>"11111101",
  21928=>"11111111",
  21929=>"00000001",
  21930=>"00000100",
  21931=>"00000001",
  21932=>"11111111",
  21933=>"11111101",
  21934=>"11111111",
  21935=>"11111101",
  21936=>"11111111",
  21937=>"11111110",
  21938=>"11111110",
  21939=>"11111101",
  21940=>"11111101",
  21941=>"11111111",
  21942=>"11111101",
  21943=>"11111110",
  21944=>"00000011",
  21945=>"00000000",
  21946=>"00000000",
  21947=>"11111111",
  21948=>"00000010",
  21949=>"11111101",
  21950=>"11111110",
  21951=>"00000001",
  21952=>"00000010",
  21953=>"11111110",
  21954=>"00000001",
  21955=>"11111110",
  21956=>"00000010",
  21957=>"11111110",
  21958=>"11111101",
  21959=>"11111101",
  21960=>"00000100",
  21961=>"00000010",
  21962=>"00000001",
  21963=>"11111101",
  21964=>"11111100",
  21965=>"11111101",
  21966=>"11111110",
  21967=>"11111111",
  21968=>"11111101",
  21969=>"00000000",
  21970=>"00000000",
  21971=>"11111110",
  21972=>"00000100",
  21973=>"00000000",
  21974=>"11111111",
  21975=>"00000010",
  21976=>"11111110",
  21977=>"11111101",
  21978=>"11111101",
  21979=>"00000001",
  21980=>"11111101",
  21981=>"11111110",
  21982=>"00000010",
  21983=>"00000011",
  21984=>"11111110",
  21985=>"11111111",
  21986=>"00000010",
  21987=>"11111110",
  21988=>"00000000",
  21989=>"00000010",
  21990=>"11111110",
  21991=>"00000000",
  21992=>"00000011",
  21993=>"11111110",
  21994=>"00000000",
  21995=>"00000101",
  21996=>"11111101",
  21997=>"00000010",
  21998=>"00000000",
  21999=>"11111101",
  22000=>"11111111",
  22001=>"00000010",
  22002=>"11111111",
  22003=>"11111101",
  22004=>"00000000",
  22005=>"00000010",
  22006=>"00000011",
  22007=>"00000001",
  22008=>"00000011",
  22009=>"00000001",
  22010=>"00000000",
  22011=>"00000011",
  22012=>"00000010",
  22013=>"11111101",
  22014=>"00000010",
  22015=>"11111110",
  22016=>"00000000",
  22017=>"00000001",
  22018=>"00000000",
  22019=>"11111101",
  22020=>"00000000",
  22021=>"00000000",
  22022=>"00000000",
  22023=>"00000000",
  22024=>"00000001",
  22025=>"11111110",
  22026=>"00000000",
  22027=>"00000001",
  22028=>"00000011",
  22029=>"00000011",
  22030=>"00000010",
  22031=>"11111110",
  22032=>"00000010",
  22033=>"11111101",
  22034=>"11111111",
  22035=>"11111111",
  22036=>"00000011",
  22037=>"00000010",
  22038=>"00000010",
  22039=>"00000000",
  22040=>"00000010",
  22041=>"11111110",
  22042=>"00000000",
  22043=>"00000000",
  22044=>"11111111",
  22045=>"11111110",
  22046=>"00000001",
  22047=>"00000010",
  22048=>"00000011",
  22049=>"11111101",
  22050=>"00000011",
  22051=>"11111111",
  22052=>"00000001",
  22053=>"00000001",
  22054=>"00000011",
  22055=>"11111110",
  22056=>"00000001",
  22057=>"00000000",
  22058=>"11111100",
  22059=>"00000010",
  22060=>"11111110",
  22061=>"00000001",
  22062=>"00000001",
  22063=>"11111110",
  22064=>"00000010",
  22065=>"00000011",
  22066=>"11111111",
  22067=>"00000000",
  22068=>"00000010",
  22069=>"11111111",
  22070=>"11111101",
  22071=>"00000001",
  22072=>"00000000",
  22073=>"00000010",
  22074=>"11111110",
  22075=>"00000011",
  22076=>"11111101",
  22077=>"00000010",
  22078=>"00000001",
  22079=>"00000011",
  22080=>"00000100",
  22081=>"00000000",
  22082=>"00000000",
  22083=>"00000010",
  22084=>"11111110",
  22085=>"11111110",
  22086=>"11111110",
  22087=>"00000010",
  22088=>"11111111",
  22089=>"11111101",
  22090=>"11111111",
  22091=>"00000010",
  22092=>"00000001",
  22093=>"11111110",
  22094=>"00000010",
  22095=>"00000001",
  22096=>"11111110",
  22097=>"11111101",
  22098=>"11111110",
  22099=>"11111110",
  22100=>"00000000",
  22101=>"11111111",
  22102=>"00000001",
  22103=>"11111101",
  22104=>"11111101",
  22105=>"00000011",
  22106=>"00000010",
  22107=>"11111110",
  22108=>"00000001",
  22109=>"00000000",
  22110=>"00000010",
  22111=>"00000000",
  22112=>"11111111",
  22113=>"11111110",
  22114=>"11111111",
  22115=>"00000001",
  22116=>"11111110",
  22117=>"00000010",
  22118=>"11111111",
  22119=>"00000010",
  22120=>"11111111",
  22121=>"00000010",
  22122=>"11111111",
  22123=>"11111110",
  22124=>"00000100",
  22125=>"11111101",
  22126=>"00000100",
  22127=>"11111101",
  22128=>"11111110",
  22129=>"00000011",
  22130=>"11111101",
  22131=>"00000010",
  22132=>"11111111",
  22133=>"00000001",
  22134=>"00000001",
  22135=>"11111111",
  22136=>"00000010",
  22137=>"00000000",
  22138=>"00000000",
  22139=>"11111101",
  22140=>"00000000",
  22141=>"00000001",
  22142=>"11111101",
  22143=>"00000001",
  22144=>"00000001",
  22145=>"00000000",
  22146=>"11111111",
  22147=>"00000010",
  22148=>"00000011",
  22149=>"00000001",
  22150=>"00000000",
  22151=>"11111110",
  22152=>"11111110",
  22153=>"00000001",
  22154=>"11111111",
  22155=>"11111110",
  22156=>"00000010",
  22157=>"11111110",
  22158=>"11111111",
  22159=>"11111110",
  22160=>"11111110",
  22161=>"00000000",
  22162=>"00000101",
  22163=>"00000000",
  22164=>"11111111",
  22165=>"00000000",
  22166=>"00000011",
  22167=>"00000011",
  22168=>"11111110",
  22169=>"00000001",
  22170=>"00000010",
  22171=>"00000001",
  22172=>"11111110",
  22173=>"11111110",
  22174=>"11111111",
  22175=>"00000001",
  22176=>"00000000",
  22177=>"00000000",
  22178=>"00000001",
  22179=>"11111111",
  22180=>"11111110",
  22181=>"11111111",
  22182=>"11111111",
  22183=>"11111111",
  22184=>"11111110",
  22185=>"00000100",
  22186=>"00000001",
  22187=>"11111110",
  22188=>"11111110",
  22189=>"00000010",
  22190=>"11111111",
  22191=>"11111101",
  22192=>"11111111",
  22193=>"11111111",
  22194=>"00000010",
  22195=>"00000000",
  22196=>"00000010",
  22197=>"00000001",
  22198=>"11111110",
  22199=>"11111110",
  22200=>"11111111",
  22201=>"11111110",
  22202=>"00000001",
  22203=>"11111110",
  22204=>"11111110",
  22205=>"11111110",
  22206=>"00000101",
  22207=>"00000000",
  22208=>"00000001",
  22209=>"00000000",
  22210=>"00000001",
  22211=>"00000001",
  22212=>"00000011",
  22213=>"11111110",
  22214=>"11111110",
  22215=>"11111101",
  22216=>"11111111",
  22217=>"00000010",
  22218=>"11111110",
  22219=>"11111110",
  22220=>"00000010",
  22221=>"11111111",
  22222=>"00000000",
  22223=>"11111111",
  22224=>"00000010",
  22225=>"11111111",
  22226=>"00000011",
  22227=>"00000000",
  22228=>"00000011",
  22229=>"00000101",
  22230=>"00000010",
  22231=>"11111110",
  22232=>"11111110",
  22233=>"00000001",
  22234=>"00000000",
  22235=>"11111111",
  22236=>"00000001",
  22237=>"11111111",
  22238=>"00000011",
  22239=>"00000000",
  22240=>"11111101",
  22241=>"00000011",
  22242=>"11111110",
  22243=>"00000011",
  22244=>"11111110",
  22245=>"00000000",
  22246=>"00000010",
  22247=>"11111111",
  22248=>"00000000",
  22249=>"11111110",
  22250=>"00000000",
  22251=>"11111111",
  22252=>"00000001",
  22253=>"11111110",
  22254=>"00000100",
  22255=>"11111111",
  22256=>"00000010",
  22257=>"00000001",
  22258=>"11111110",
  22259=>"00000000",
  22260=>"00000000",
  22261=>"00000011",
  22262=>"00000001",
  22263=>"00000001",
  22264=>"00000000",
  22265=>"11111110",
  22266=>"11111111",
  22267=>"11111111",
  22268=>"00000000",
  22269=>"11111110",
  22270=>"00000001",
  22271=>"00000000",
  22272=>"00000011",
  22273=>"00000011",
  22274=>"11111111",
  22275=>"11111110",
  22276=>"11111111",
  22277=>"00000000",
  22278=>"11111111",
  22279=>"00000011",
  22280=>"00000000",
  22281=>"11111101",
  22282=>"00000000",
  22283=>"11111110",
  22284=>"11111101",
  22285=>"11111111",
  22286=>"00000010",
  22287=>"00000000",
  22288=>"00000001",
  22289=>"00000011",
  22290=>"11111110",
  22291=>"00000000",
  22292=>"00000001",
  22293=>"00000001",
  22294=>"11111110",
  22295=>"11111111",
  22296=>"00000001",
  22297=>"11111111",
  22298=>"00000010",
  22299=>"11111111",
  22300=>"00000000",
  22301=>"11111110",
  22302=>"00000000",
  22303=>"00000000",
  22304=>"11111101",
  22305=>"11111110",
  22306=>"00000000",
  22307=>"00000000",
  22308=>"00000010",
  22309=>"00000101",
  22310=>"11111110",
  22311=>"11111110",
  22312=>"00000010",
  22313=>"00000001",
  22314=>"00000010",
  22315=>"11111110",
  22316=>"11111110",
  22317=>"11111111",
  22318=>"00000001",
  22319=>"00000100",
  22320=>"11111101",
  22321=>"00000001",
  22322=>"11111110",
  22323=>"00000010",
  22324=>"00000000",
  22325=>"00000010",
  22326=>"00000011",
  22327=>"11111110",
  22328=>"11111110",
  22329=>"11111111",
  22330=>"11111111",
  22331=>"00000001",
  22332=>"11111111",
  22333=>"11111110",
  22334=>"11111110",
  22335=>"11111111",
  22336=>"00000000",
  22337=>"00000010",
  22338=>"00000011",
  22339=>"11111110",
  22340=>"00000000",
  22341=>"11111111",
  22342=>"00000000",
  22343=>"00000000",
  22344=>"11111110",
  22345=>"11111110",
  22346=>"00000001",
  22347=>"11111110",
  22348=>"11111111",
  22349=>"00000000",
  22350=>"11111101",
  22351=>"11111111",
  22352=>"11111111",
  22353=>"00000000",
  22354=>"11111111",
  22355=>"00000010",
  22356=>"11111110",
  22357=>"11111110",
  22358=>"00000010",
  22359=>"11111110",
  22360=>"00000001",
  22361=>"00000000",
  22362=>"00000011",
  22363=>"11111110",
  22364=>"00000001",
  22365=>"00000010",
  22366=>"00000100",
  22367=>"11111111",
  22368=>"00000001",
  22369=>"00000001",
  22370=>"11111111",
  22371=>"11111110",
  22372=>"00000011",
  22373=>"00000011",
  22374=>"00000011",
  22375=>"11111101",
  22376=>"11111101",
  22377=>"00000000",
  22378=>"11111110",
  22379=>"00000000",
  22380=>"11111110",
  22381=>"11111101",
  22382=>"00000011",
  22383=>"00000000",
  22384=>"00000001",
  22385=>"11111111",
  22386=>"11111110",
  22387=>"00000110",
  22388=>"00000000",
  22389=>"00000011",
  22390=>"11111101",
  22391=>"11111111",
  22392=>"11111111",
  22393=>"00000010",
  22394=>"00000000",
  22395=>"11111101",
  22396=>"00000010",
  22397=>"11111110",
  22398=>"11111111",
  22399=>"11111110",
  22400=>"00000010",
  22401=>"00000001",
  22402=>"00000000",
  22403=>"00000010",
  22404=>"00000010",
  22405=>"11111111",
  22406=>"00000010",
  22407=>"00000010",
  22408=>"00000010",
  22409=>"11111110",
  22410=>"11111110",
  22411=>"00000001",
  22412=>"11111111",
  22413=>"11111110",
  22414=>"11111111",
  22415=>"11111111",
  22416=>"00000000",
  22417=>"11111110",
  22418=>"11111100",
  22419=>"11111110",
  22420=>"11111110",
  22421=>"11111101",
  22422=>"11111111",
  22423=>"00000000",
  22424=>"00000011",
  22425=>"00000010",
  22426=>"00000001",
  22427=>"00000000",
  22428=>"11111111",
  22429=>"11111101",
  22430=>"00000001",
  22431=>"11111101",
  22432=>"00000011",
  22433=>"11111111",
  22434=>"00000100",
  22435=>"00000000",
  22436=>"00000000",
  22437=>"00000001",
  22438=>"11111110",
  22439=>"11111111",
  22440=>"00000010",
  22441=>"11111111",
  22442=>"11111101",
  22443=>"11111111",
  22444=>"00000000",
  22445=>"11111111",
  22446=>"00000000",
  22447=>"11111101",
  22448=>"00000001",
  22449=>"11111111",
  22450=>"11111101",
  22451=>"00000010",
  22452=>"00000000",
  22453=>"11111111",
  22454=>"11111111",
  22455=>"00000000",
  22456=>"11111111",
  22457=>"11111110",
  22458=>"11111111",
  22459=>"00000001",
  22460=>"11111110",
  22461=>"00000010",
  22462=>"00000001",
  22463=>"00000010",
  22464=>"11111110",
  22465=>"00000001",
  22466=>"00000000",
  22467=>"00000010",
  22468=>"11111110",
  22469=>"00000001",
  22470=>"11111101",
  22471=>"11111101",
  22472=>"11111101",
  22473=>"11111110",
  22474=>"00000000",
  22475=>"00000001",
  22476=>"11111111",
  22477=>"00000011",
  22478=>"00000000",
  22479=>"11111101",
  22480=>"11111111",
  22481=>"00000010",
  22482=>"00000011",
  22483=>"00000001",
  22484=>"11111111",
  22485=>"11111111",
  22486=>"11111111",
  22487=>"00000011",
  22488=>"11111111",
  22489=>"11111111",
  22490=>"11111111",
  22491=>"00000000",
  22492=>"11111111",
  22493=>"11111101",
  22494=>"11111111",
  22495=>"00000010",
  22496=>"00000001",
  22497=>"00000010",
  22498=>"00000000",
  22499=>"00000010",
  22500=>"00000000",
  22501=>"11111111",
  22502=>"00000010",
  22503=>"00000010",
  22504=>"00000000",
  22505=>"11111111",
  22506=>"11111110",
  22507=>"00000100",
  22508=>"00000010",
  22509=>"00000011",
  22510=>"11111101",
  22511=>"11111110",
  22512=>"00000001",
  22513=>"00000010",
  22514=>"11111101",
  22515=>"11111101",
  22516=>"11111101",
  22517=>"11111111",
  22518=>"00000101",
  22519=>"00000000",
  22520=>"00000001",
  22521=>"11111111",
  22522=>"00000011",
  22523=>"11111110",
  22524=>"11111111",
  22525=>"11111111",
  22526=>"00000011",
  22527=>"00000011",
  22528=>"11111110",
  22529=>"11111110",
  22530=>"00000001",
  22531=>"00000001",
  22532=>"00000001",
  22533=>"00000011",
  22534=>"11111110",
  22535=>"11111101",
  22536=>"00000000",
  22537=>"00000000",
  22538=>"11111101",
  22539=>"00000000",
  22540=>"11111111",
  22541=>"11111101",
  22542=>"00000001",
  22543=>"11111110",
  22544=>"00000010",
  22545=>"00000100",
  22546=>"11111111",
  22547=>"00000101",
  22548=>"11111111",
  22549=>"11111111",
  22550=>"11111110",
  22551=>"11111111",
  22552=>"00000001",
  22553=>"11111110",
  22554=>"00000000",
  22555=>"11111101",
  22556=>"11111111",
  22557=>"00000000",
  22558=>"11111101",
  22559=>"11111110",
  22560=>"00000100",
  22561=>"00000001",
  22562=>"00000010",
  22563=>"11111111",
  22564=>"11111110",
  22565=>"11111110",
  22566=>"11111111",
  22567=>"00000010",
  22568=>"00000001",
  22569=>"11111110",
  22570=>"00000010",
  22571=>"11111110",
  22572=>"00000000",
  22573=>"11111111",
  22574=>"11111111",
  22575=>"11111111",
  22576=>"11111111",
  22577=>"00000010",
  22578=>"11111111",
  22579=>"00000001",
  22580=>"11111110",
  22581=>"00000001",
  22582=>"00000100",
  22583=>"00000001",
  22584=>"00000011",
  22585=>"11111111",
  22586=>"00000010",
  22587=>"00000001",
  22588=>"11111101",
  22589=>"00000010",
  22590=>"11111110",
  22591=>"00000011",
  22592=>"00000000",
  22593=>"11111110",
  22594=>"11111110",
  22595=>"00000010",
  22596=>"00000000",
  22597=>"00000000",
  22598=>"00000000",
  22599=>"00000000",
  22600=>"00000010",
  22601=>"11111111",
  22602=>"00000001",
  22603=>"00000000",
  22604=>"00000001",
  22605=>"00000010",
  22606=>"00000010",
  22607=>"11111101",
  22608=>"00000011",
  22609=>"11111110",
  22610=>"00000001",
  22611=>"00000011",
  22612=>"00000011",
  22613=>"00000000",
  22614=>"00000000",
  22615=>"11111111",
  22616=>"11111101",
  22617=>"11111111",
  22618=>"00000000",
  22619=>"11111110",
  22620=>"11111110",
  22621=>"00000001",
  22622=>"11111100",
  22623=>"00000001",
  22624=>"11111101",
  22625=>"11111110",
  22626=>"00000010",
  22627=>"00000001",
  22628=>"00000001",
  22629=>"00000010",
  22630=>"00000011",
  22631=>"00000000",
  22632=>"11111101",
  22633=>"00000000",
  22634=>"11111101",
  22635=>"00000001",
  22636=>"11111101",
  22637=>"00000001",
  22638=>"00000001",
  22639=>"00000010",
  22640=>"11111101",
  22641=>"00000010",
  22642=>"00000010",
  22643=>"00000110",
  22644=>"11111110",
  22645=>"00000010",
  22646=>"11111111",
  22647=>"11111111",
  22648=>"00000010",
  22649=>"00000000",
  22650=>"00000011",
  22651=>"11111101",
  22652=>"11111111",
  22653=>"00000001",
  22654=>"11111110",
  22655=>"11111111",
  22656=>"00000001",
  22657=>"00000101",
  22658=>"00000110",
  22659=>"00000000",
  22660=>"00000011",
  22661=>"00000001",
  22662=>"11111111",
  22663=>"00000011",
  22664=>"11111101",
  22665=>"11111111",
  22666=>"11111111",
  22667=>"11111111",
  22668=>"11111111",
  22669=>"11111110",
  22670=>"11111111",
  22671=>"11111111",
  22672=>"00000010",
  22673=>"11111110",
  22674=>"11111111",
  22675=>"11111110",
  22676=>"00000001",
  22677=>"00000000",
  22678=>"11111111",
  22679=>"11111111",
  22680=>"11111110",
  22681=>"11111101",
  22682=>"00000001",
  22683=>"00000101",
  22684=>"00000010",
  22685=>"00000100",
  22686=>"00000010",
  22687=>"00000010",
  22688=>"00000010",
  22689=>"00000010",
  22690=>"11111111",
  22691=>"00000000",
  22692=>"00000001",
  22693=>"00000000",
  22694=>"11111101",
  22695=>"00000100",
  22696=>"11111101",
  22697=>"00000000",
  22698=>"11111110",
  22699=>"11111110",
  22700=>"00000010",
  22701=>"00000000",
  22702=>"00000011",
  22703=>"00000001",
  22704=>"00000100",
  22705=>"11111111",
  22706=>"00000100",
  22707=>"11111111",
  22708=>"00000100",
  22709=>"11111111",
  22710=>"00000100",
  22711=>"11111100",
  22712=>"11111111",
  22713=>"00000001",
  22714=>"00000000",
  22715=>"00000000",
  22716=>"11111111",
  22717=>"00000001",
  22718=>"11111101",
  22719=>"11111111",
  22720=>"00000000",
  22721=>"11111111",
  22722=>"00000001",
  22723=>"00000000",
  22724=>"00000010",
  22725=>"00000100",
  22726=>"11111101",
  22727=>"11111101",
  22728=>"11111111",
  22729=>"11111101",
  22730=>"11111111",
  22731=>"11111111",
  22732=>"00000001",
  22733=>"11111111",
  22734=>"11111110",
  22735=>"00000000",
  22736=>"11111111",
  22737=>"00000010",
  22738=>"11111110",
  22739=>"11111111",
  22740=>"11111110",
  22741=>"11111100",
  22742=>"00000000",
  22743=>"00000000",
  22744=>"00000000",
  22745=>"11111101",
  22746=>"00000010",
  22747=>"00000000",
  22748=>"00000000",
  22749=>"00000001",
  22750=>"00000010",
  22751=>"11111110",
  22752=>"11111111",
  22753=>"00000000",
  22754=>"00000000",
  22755=>"11111110",
  22756=>"00000000",
  22757=>"00000000",
  22758=>"11111111",
  22759=>"00000010",
  22760=>"00000010",
  22761=>"00000000",
  22762=>"11111111",
  22763=>"00000001",
  22764=>"00000011",
  22765=>"11111111",
  22766=>"11111111",
  22767=>"00000000",
  22768=>"11111101",
  22769=>"00000000",
  22770=>"00000001",
  22771=>"11111111",
  22772=>"00000000",
  22773=>"11111101",
  22774=>"11111101",
  22775=>"11111110",
  22776=>"11111110",
  22777=>"00000010",
  22778=>"11111110",
  22779=>"00000010",
  22780=>"00000101",
  22781=>"11111100",
  22782=>"11111101",
  22783=>"11111101",
  22784=>"11111111",
  22785=>"00000000",
  22786=>"11111110",
  22787=>"00000011",
  22788=>"11111111",
  22789=>"00000010",
  22790=>"00000011",
  22791=>"11111110",
  22792=>"11111111",
  22793=>"00000011",
  22794=>"00000100",
  22795=>"11111111",
  22796=>"11111101",
  22797=>"11111110",
  22798=>"00000001",
  22799=>"11111110",
  22800=>"00000000",
  22801=>"00000000",
  22802=>"00000000",
  22803=>"11111101",
  22804=>"00000001",
  22805=>"00000000",
  22806=>"11111110",
  22807=>"00000100",
  22808=>"00000000",
  22809=>"00000000",
  22810=>"00000001",
  22811=>"11111111",
  22812=>"00000011",
  22813=>"00000010",
  22814=>"00000000",
  22815=>"11111101",
  22816=>"11111111",
  22817=>"00000010",
  22818=>"00000010",
  22819=>"00000001",
  22820=>"00000001",
  22821=>"11111111",
  22822=>"00000010",
  22823=>"11111101",
  22824=>"00000000",
  22825=>"00000001",
  22826=>"11111111",
  22827=>"00000001",
  22828=>"00000010",
  22829=>"11111110",
  22830=>"00000010",
  22831=>"00000011",
  22832=>"00000001",
  22833=>"11111111",
  22834=>"00000010",
  22835=>"11111111",
  22836=>"00000101",
  22837=>"00000001",
  22838=>"11111111",
  22839=>"00000000",
  22840=>"00000010",
  22841=>"11111101",
  22842=>"00000011",
  22843=>"11111110",
  22844=>"00000010",
  22845=>"11111111",
  22846=>"11111111",
  22847=>"11111111",
  22848=>"11111111",
  22849=>"11111110",
  22850=>"11111110",
  22851=>"11111101",
  22852=>"00000001",
  22853=>"00000100",
  22854=>"11111101",
  22855=>"11111110",
  22856=>"00000001",
  22857=>"11111111",
  22858=>"11111111",
  22859=>"00000000",
  22860=>"00000000",
  22861=>"11111110",
  22862=>"11111110",
  22863=>"11111110",
  22864=>"00000001",
  22865=>"00000010",
  22866=>"00000100",
  22867=>"00000000",
  22868=>"00000001",
  22869=>"11111101",
  22870=>"11111110",
  22871=>"11111110",
  22872=>"11111110",
  22873=>"11111110",
  22874=>"11111111",
  22875=>"11111101",
  22876=>"00000001",
  22877=>"00000000",
  22878=>"11111111",
  22879=>"11111101",
  22880=>"00000000",
  22881=>"00000000",
  22882=>"11111101",
  22883=>"11111110",
  22884=>"00000001",
  22885=>"11111101",
  22886=>"11111110",
  22887=>"11111110",
  22888=>"00000000",
  22889=>"00000001",
  22890=>"00000010",
  22891=>"11111101",
  22892=>"00000101",
  22893=>"11111111",
  22894=>"00000000",
  22895=>"00000000",
  22896=>"00000011",
  22897=>"11111111",
  22898=>"11111111",
  22899=>"00000001",
  22900=>"11111111",
  22901=>"11111110",
  22902=>"00000011",
  22903=>"00000000",
  22904=>"11111111",
  22905=>"11111110",
  22906=>"00000000",
  22907=>"00000010",
  22908=>"00000000",
  22909=>"11111101",
  22910=>"00000010",
  22911=>"11111110",
  22912=>"00000000",
  22913=>"00000010",
  22914=>"11111111",
  22915=>"11111110",
  22916=>"11111101",
  22917=>"00000000",
  22918=>"11111111",
  22919=>"00000000",
  22920=>"11111110",
  22921=>"11111111",
  22922=>"00000001",
  22923=>"11111110",
  22924=>"11111111",
  22925=>"11111110",
  22926=>"00000010",
  22927=>"11111110",
  22928=>"00000000",
  22929=>"00000001",
  22930=>"11111101",
  22931=>"00000010",
  22932=>"11111101",
  22933=>"00000010",
  22934=>"00000000",
  22935=>"11111111",
  22936=>"11111101",
  22937=>"11111101",
  22938=>"11111110",
  22939=>"00000010",
  22940=>"11111110",
  22941=>"11111110",
  22942=>"11111101",
  22943=>"00000001",
  22944=>"11111111",
  22945=>"00000000",
  22946=>"00000010",
  22947=>"11111110",
  22948=>"11111101",
  22949=>"11111110",
  22950=>"00000001",
  22951=>"11111110",
  22952=>"00000000",
  22953=>"00000000",
  22954=>"00000000",
  22955=>"00000011",
  22956=>"00000001",
  22957=>"00000010",
  22958=>"11111110",
  22959=>"11111101",
  22960=>"11111110",
  22961=>"00000010",
  22962=>"00000011",
  22963=>"11111111",
  22964=>"11111110",
  22965=>"11111110",
  22966=>"00000001",
  22967=>"11111111",
  22968=>"00000000",
  22969=>"11111101",
  22970=>"11111110",
  22971=>"11111111",
  22972=>"00000000",
  22973=>"11111110",
  22974=>"11111101",
  22975=>"00000001",
  22976=>"00000001",
  22977=>"11111110",
  22978=>"11111101",
  22979=>"00000000",
  22980=>"00000001",
  22981=>"00000010",
  22982=>"11111101",
  22983=>"00000101",
  22984=>"11111111",
  22985=>"00000001",
  22986=>"00000101",
  22987=>"11111101",
  22988=>"11111101",
  22989=>"11111110",
  22990=>"11111101",
  22991=>"00000010",
  22992=>"00000001",
  22993=>"11111101",
  22994=>"00000001",
  22995=>"00000000",
  22996=>"11111110",
  22997=>"00000001",
  22998=>"11111101",
  22999=>"00000001",
  23000=>"00000010",
  23001=>"11111111",
  23002=>"00000011",
  23003=>"11111111",
  23004=>"00000000",
  23005=>"11111101",
  23006=>"00000010",
  23007=>"11111110",
  23008=>"11111101",
  23009=>"00000010",
  23010=>"11111101",
  23011=>"11111111",
  23012=>"00000010",
  23013=>"11111110",
  23014=>"11111111",
  23015=>"11111111",
  23016=>"00000011",
  23017=>"11111110",
  23018=>"00000010",
  23019=>"11111101",
  23020=>"00000000",
  23021=>"00000011",
  23022=>"00000001",
  23023=>"00000100",
  23024=>"00000010",
  23025=>"00000000",
  23026=>"00000000",
  23027=>"11111110",
  23028=>"11111110",
  23029=>"00000100",
  23030=>"00000001",
  23031=>"00000000",
  23032=>"11111110",
  23033=>"00000001",
  23034=>"11111101",
  23035=>"00000001",
  23036=>"00000001",
  23037=>"00000010",
  23038=>"00000010",
  23039=>"00000010",
  23040=>"00000011",
  23041=>"11111111",
  23042=>"11111110",
  23043=>"00000101",
  23044=>"00000010",
  23045=>"00000000",
  23046=>"11111101",
  23047=>"00000001",
  23048=>"00000001",
  23049=>"00000001",
  23050=>"00000001",
  23051=>"00000011",
  23052=>"00000010",
  23053=>"11111111",
  23054=>"00000001",
  23055=>"11111111",
  23056=>"00000011",
  23057=>"00000000",
  23058=>"00000001",
  23059=>"00000001",
  23060=>"11111110",
  23061=>"00000000",
  23062=>"00000001",
  23063=>"00000000",
  23064=>"11111110",
  23065=>"00000000",
  23066=>"00000001",
  23067=>"11111110",
  23068=>"00000001",
  23069=>"00000010",
  23070=>"00000011",
  23071=>"00000000",
  23072=>"11111110",
  23073=>"11111110",
  23074=>"00000000",
  23075=>"11111110",
  23076=>"00000001",
  23077=>"00000011",
  23078=>"00000000",
  23079=>"11111110",
  23080=>"00000000",
  23081=>"00000000",
  23082=>"11111110",
  23083=>"11111110",
  23084=>"00000000",
  23085=>"11111101",
  23086=>"00000010",
  23087=>"00000000",
  23088=>"11111110",
  23089=>"00000001",
  23090=>"11111111",
  23091=>"00000010",
  23092=>"11111110",
  23093=>"11111101",
  23094=>"00000000",
  23095=>"00000011",
  23096=>"00000011",
  23097=>"11111110",
  23098=>"00000001",
  23099=>"00000000",
  23100=>"11111101",
  23101=>"00000000",
  23102=>"11111101",
  23103=>"00000001",
  23104=>"00000000",
  23105=>"00000000",
  23106=>"00000000",
  23107=>"11111111",
  23108=>"11111111",
  23109=>"00000000",
  23110=>"00000011",
  23111=>"11111101",
  23112=>"00000001",
  23113=>"00000010",
  23114=>"11111110",
  23115=>"11111111",
  23116=>"00000001",
  23117=>"11111110",
  23118=>"11111101",
  23119=>"11111110",
  23120=>"00000001",
  23121=>"11111111",
  23122=>"11111110",
  23123=>"00000010",
  23124=>"00000000",
  23125=>"00000000",
  23126=>"11111111",
  23127=>"00000000",
  23128=>"00000000",
  23129=>"00000011",
  23130=>"00000000",
  23131=>"00000010",
  23132=>"00000000",
  23133=>"00000001",
  23134=>"11111111",
  23135=>"11111111",
  23136=>"11111111",
  23137=>"00000010",
  23138=>"00000001",
  23139=>"00000010",
  23140=>"00000000",
  23141=>"11111111",
  23142=>"00000010",
  23143=>"00000001",
  23144=>"11111110",
  23145=>"00000000",
  23146=>"11111111",
  23147=>"11111101",
  23148=>"11111111",
  23149=>"11111111",
  23150=>"00000000",
  23151=>"11111110",
  23152=>"00000010",
  23153=>"00000000",
  23154=>"11111101",
  23155=>"11111110",
  23156=>"11111110",
  23157=>"11111111",
  23158=>"11111111",
  23159=>"00000010",
  23160=>"11111111",
  23161=>"11111110",
  23162=>"00000001",
  23163=>"00000011",
  23164=>"00000010",
  23165=>"11111110",
  23166=>"11111101",
  23167=>"11111111",
  23168=>"00000011",
  23169=>"00000011",
  23170=>"11111110",
  23171=>"11111110",
  23172=>"11111110",
  23173=>"11111101",
  23174=>"11111101",
  23175=>"00000001",
  23176=>"00000000",
  23177=>"11111110",
  23178=>"00000001",
  23179=>"11111100",
  23180=>"00000001",
  23181=>"11111110",
  23182=>"11111110",
  23183=>"00000000",
  23184=>"00000010",
  23185=>"11111110",
  23186=>"00000010",
  23187=>"11111110",
  23188=>"00000000",
  23189=>"11111101",
  23190=>"11111101",
  23191=>"00000010",
  23192=>"11111110",
  23193=>"00000001",
  23194=>"00000000",
  23195=>"11111110",
  23196=>"00000101",
  23197=>"00000001",
  23198=>"11111111",
  23199=>"00000010",
  23200=>"00000010",
  23201=>"00000001",
  23202=>"11111101",
  23203=>"11111110",
  23204=>"00000001",
  23205=>"11111110",
  23206=>"00000001",
  23207=>"11111111",
  23208=>"00000011",
  23209=>"00000100",
  23210=>"11111111",
  23211=>"11111101",
  23212=>"00000001",
  23213=>"00000001",
  23214=>"00000001",
  23215=>"00000011",
  23216=>"00000010",
  23217=>"11111111",
  23218=>"00000010",
  23219=>"00000000",
  23220=>"11111111",
  23221=>"00000100",
  23222=>"00000000",
  23223=>"00000010",
  23224=>"00000010",
  23225=>"11111101",
  23226=>"00000001",
  23227=>"00000100",
  23228=>"00000001",
  23229=>"11111101",
  23230=>"00000000",
  23231=>"00000000",
  23232=>"00000010",
  23233=>"00000011",
  23234=>"00000011",
  23235=>"00000001",
  23236=>"00000001",
  23237=>"00000000",
  23238=>"11111101",
  23239=>"11111110",
  23240=>"11111111",
  23241=>"00000000",
  23242=>"11111111",
  23243=>"00000000",
  23244=>"11111110",
  23245=>"00000010",
  23246=>"00000010",
  23247=>"11111111",
  23248=>"11111111",
  23249=>"00000100",
  23250=>"00000001",
  23251=>"00000000",
  23252=>"00000100",
  23253=>"11111101",
  23254=>"11111111",
  23255=>"00000010",
  23256=>"11111110",
  23257=>"11111101",
  23258=>"11111111",
  23259=>"11111101",
  23260=>"11111101",
  23261=>"11111110",
  23262=>"00000000",
  23263=>"00000101",
  23264=>"00000001",
  23265=>"00000100",
  23266=>"00000000",
  23267=>"11111111",
  23268=>"11111110",
  23269=>"00000000",
  23270=>"00000000",
  23271=>"11111111",
  23272=>"11111110",
  23273=>"00000011",
  23274=>"00000001",
  23275=>"00000000",
  23276=>"00000100",
  23277=>"00000101",
  23278=>"00000001",
  23279=>"11111101",
  23280=>"00000000",
  23281=>"00000000",
  23282=>"00000011",
  23283=>"00000000",
  23284=>"00000010",
  23285=>"11111101",
  23286=>"11111111",
  23287=>"00000001",
  23288=>"11111110",
  23289=>"00000011",
  23290=>"00000001",
  23291=>"11111110",
  23292=>"00000010",
  23293=>"00000000",
  23294=>"11111111",
  23295=>"11111111",
  23296=>"11111101",
  23297=>"00000001",
  23298=>"00000110",
  23299=>"11111111",
  23300=>"11111111",
  23301=>"00000001",
  23302=>"00000011",
  23303=>"00000000",
  23304=>"00000000",
  23305=>"00000000",
  23306=>"11111101",
  23307=>"11111111",
  23308=>"11111111",
  23309=>"00000010",
  23310=>"00000001",
  23311=>"11111110",
  23312=>"11111101",
  23313=>"11111111",
  23314=>"00000001",
  23315=>"00000001",
  23316=>"00000001",
  23317=>"11111101",
  23318=>"11111111",
  23319=>"00000010",
  23320=>"00000011",
  23321=>"11111110",
  23322=>"11111110",
  23323=>"11111111",
  23324=>"00000010",
  23325=>"11111111",
  23326=>"11111101",
  23327=>"00000100",
  23328=>"00000000",
  23329=>"00000110",
  23330=>"11111110",
  23331=>"00000000",
  23332=>"00000011",
  23333=>"00000011",
  23334=>"11111111",
  23335=>"11111110",
  23336=>"00000000",
  23337=>"11111101",
  23338=>"00000011",
  23339=>"11111110",
  23340=>"00000010",
  23341=>"00000000",
  23342=>"11111110",
  23343=>"11111110",
  23344=>"11111101",
  23345=>"00000110",
  23346=>"00000100",
  23347=>"00000010",
  23348=>"00000010",
  23349=>"11111111",
  23350=>"00000000",
  23351=>"00000001",
  23352=>"00000001",
  23353=>"00000001",
  23354=>"11111111",
  23355=>"11111111",
  23356=>"11111110",
  23357=>"11111110",
  23358=>"11111111",
  23359=>"11111111",
  23360=>"11111110",
  23361=>"11111111",
  23362=>"11111101",
  23363=>"00000001",
  23364=>"00000001",
  23365=>"11111111",
  23366=>"11111101",
  23367=>"11111101",
  23368=>"00000000",
  23369=>"00000010",
  23370=>"11111101",
  23371=>"00000000",
  23372=>"11111111",
  23373=>"11111111",
  23374=>"00000001",
  23375=>"11111111",
  23376=>"11111110",
  23377=>"00000000",
  23378=>"00000000",
  23379=>"11111110",
  23380=>"00000001",
  23381=>"00000010",
  23382=>"00000001",
  23383=>"00000010",
  23384=>"11111110",
  23385=>"11111101",
  23386=>"11111101",
  23387=>"11111111",
  23388=>"11111110",
  23389=>"11111111",
  23390=>"00000011",
  23391=>"00000000",
  23392=>"00000010",
  23393=>"00000010",
  23394=>"11111110",
  23395=>"11111110",
  23396=>"11111111",
  23397=>"11111111",
  23398=>"11111110",
  23399=>"00000010",
  23400=>"11111111",
  23401=>"11111111",
  23402=>"11111111",
  23403=>"00000001",
  23404=>"00000001",
  23405=>"00000010",
  23406=>"11111101",
  23407=>"00000011",
  23408=>"11111111",
  23409=>"11111100",
  23410=>"11111110",
  23411=>"11111110",
  23412=>"00000001",
  23413=>"00000010",
  23414=>"00000001",
  23415=>"11111110",
  23416=>"00000001",
  23417=>"00000001",
  23418=>"00000000",
  23419=>"11111101",
  23420=>"11111101",
  23421=>"00000000",
  23422=>"00000000",
  23423=>"00000010",
  23424=>"00000000",
  23425=>"00000000",
  23426=>"11111101",
  23427=>"00000001",
  23428=>"11111101",
  23429=>"11111110",
  23430=>"00000000",
  23431=>"11111111",
  23432=>"11111111",
  23433=>"00000110",
  23434=>"00000010",
  23435=>"11111111",
  23436=>"00000010",
  23437=>"11111101",
  23438=>"11111101",
  23439=>"11111110",
  23440=>"11111110",
  23441=>"11111100",
  23442=>"11111110",
  23443=>"00000011",
  23444=>"00000011",
  23445=>"11111101",
  23446=>"00000101",
  23447=>"00000001",
  23448=>"00000001",
  23449=>"00000001",
  23450=>"00000001",
  23451=>"00000010",
  23452=>"11111100",
  23453=>"11111111",
  23454=>"00000011",
  23455=>"00000000",
  23456=>"11111100",
  23457=>"00000001",
  23458=>"11111110",
  23459=>"11111101",
  23460=>"00000010",
  23461=>"00000101",
  23462=>"11111111",
  23463=>"00000010",
  23464=>"00000010",
  23465=>"00000000",
  23466=>"00000011",
  23467=>"00000010",
  23468=>"11111111",
  23469=>"00000010",
  23470=>"11111101",
  23471=>"00000000",
  23472=>"00000011",
  23473=>"11111111",
  23474=>"00000000",
  23475=>"00000110",
  23476=>"11111111",
  23477=>"11111111",
  23478=>"00000001",
  23479=>"11111101",
  23480=>"00000100",
  23481=>"00000001",
  23482=>"11111101",
  23483=>"00000100",
  23484=>"00000001",
  23485=>"00000010",
  23486=>"00000000",
  23487=>"00000010",
  23488=>"00000000",
  23489=>"00000001",
  23490=>"00000001",
  23491=>"00000000",
  23492=>"00000001",
  23493=>"11111111",
  23494=>"11111101",
  23495=>"00000001",
  23496=>"00000010",
  23497=>"00000100",
  23498=>"11111111",
  23499=>"11111110",
  23500=>"00000101",
  23501=>"00000000",
  23502=>"00000001",
  23503=>"00000001",
  23504=>"00000010",
  23505=>"11111110",
  23506=>"00000100",
  23507=>"11111111",
  23508=>"00000000",
  23509=>"11111111",
  23510=>"00000011",
  23511=>"00000000",
  23512=>"00000011",
  23513=>"00000010",
  23514=>"00000000",
  23515=>"00000001",
  23516=>"00000001",
  23517=>"00000010",
  23518=>"00000000",
  23519=>"11111110",
  23520=>"00000001",
  23521=>"00000000",
  23522=>"00000001",
  23523=>"11111111",
  23524=>"00000000",
  23525=>"00000101",
  23526=>"11111101",
  23527=>"11111110",
  23528=>"00000001",
  23529=>"00000000",
  23530=>"11111101",
  23531=>"00000000",
  23532=>"00000010",
  23533=>"00000001",
  23534=>"00000000",
  23535=>"00000001",
  23536=>"11111101",
  23537=>"11111110",
  23538=>"11111110",
  23539=>"00000000",
  23540=>"00000010",
  23541=>"00000000",
  23542=>"11111110",
  23543=>"11111111",
  23544=>"11111111",
  23545=>"00000001",
  23546=>"11111101",
  23547=>"11111110",
  23548=>"11111111",
  23549=>"00000000",
  23550=>"11111110",
  23551=>"11111111",
  23552=>"00000000",
  23553=>"11111101",
  23554=>"00000001",
  23555=>"11111110",
  23556=>"00000111",
  23557=>"11111101",
  23558=>"11111110",
  23559=>"00000000",
  23560=>"00000000",
  23561=>"00000011",
  23562=>"11111110",
  23563=>"00000000",
  23564=>"11111111",
  23565=>"00000001",
  23566=>"11111100",
  23567=>"00000001",
  23568=>"11111100",
  23569=>"11111101",
  23570=>"11111110",
  23571=>"00000001",
  23572=>"00000001",
  23573=>"11111110",
  23574=>"00000000",
  23575=>"11111111",
  23576=>"00000001",
  23577=>"11111111",
  23578=>"00000000",
  23579=>"11111111",
  23580=>"11111101",
  23581=>"00000001",
  23582=>"00000011",
  23583=>"00000101",
  23584=>"00000001",
  23585=>"00000010",
  23586=>"00000001",
  23587=>"00000000",
  23588=>"00000011",
  23589=>"11111111",
  23590=>"11111111",
  23591=>"11111110",
  23592=>"00000000",
  23593=>"11111111",
  23594=>"00000010",
  23595=>"11111100",
  23596=>"00000000",
  23597=>"00000010",
  23598=>"00000000",
  23599=>"00000010",
  23600=>"11111110",
  23601=>"00000010",
  23602=>"11111110",
  23603=>"00000001",
  23604=>"00000011",
  23605=>"00000100",
  23606=>"11111110",
  23607=>"00000010",
  23608=>"00000000",
  23609=>"00000001",
  23610=>"11111111",
  23611=>"11111110",
  23612=>"11111111",
  23613=>"11111110",
  23614=>"11111101",
  23615=>"00000101",
  23616=>"11111100",
  23617=>"11111101",
  23618=>"00000000",
  23619=>"00000010",
  23620=>"11111110",
  23621=>"00000010",
  23622=>"11111100",
  23623=>"00000100",
  23624=>"00000000",
  23625=>"00000010",
  23626=>"00000100",
  23627=>"00000100",
  23628=>"00000001",
  23629=>"11111110",
  23630=>"00000010",
  23631=>"00000001",
  23632=>"11111101",
  23633=>"11111110",
  23634=>"00000010",
  23635=>"11111110",
  23636=>"11111100",
  23637=>"00000000",
  23638=>"11111100",
  23639=>"00000000",
  23640=>"11111111",
  23641=>"11111111",
  23642=>"00000011",
  23643=>"00000000",
  23644=>"00000001",
  23645=>"11111110",
  23646=>"00000010",
  23647=>"00000000",
  23648=>"11111101",
  23649=>"00000001",
  23650=>"00000001",
  23651=>"00000001",
  23652=>"11111110",
  23653=>"00000010",
  23654=>"11111110",
  23655=>"00000000",
  23656=>"11111111",
  23657=>"11111011",
  23658=>"00000000",
  23659=>"11111110",
  23660=>"00000001",
  23661=>"11111110",
  23662=>"00000010",
  23663=>"00000001",
  23664=>"00000000",
  23665=>"00000001",
  23666=>"00000001",
  23667=>"00000001",
  23668=>"00000000",
  23669=>"00000001",
  23670=>"11111100",
  23671=>"11111101",
  23672=>"11111110",
  23673=>"11111100",
  23674=>"00000100",
  23675=>"00000100",
  23676=>"11111101",
  23677=>"00000001",
  23678=>"00000000",
  23679=>"00000001",
  23680=>"11111100",
  23681=>"11111101",
  23682=>"00000010",
  23683=>"11111110",
  23684=>"00000011",
  23685=>"11111101",
  23686=>"00000010",
  23687=>"00000001",
  23688=>"11111101",
  23689=>"00000000",
  23690=>"11111111",
  23691=>"00000011",
  23692=>"00000011",
  23693=>"11111110",
  23694=>"00000010",
  23695=>"11111101",
  23696=>"00000111",
  23697=>"11111111",
  23698=>"00000001",
  23699=>"11111111",
  23700=>"11111100",
  23701=>"00000010",
  23702=>"00000010",
  23703=>"11111111",
  23704=>"00000010",
  23705=>"11111110",
  23706=>"11111110",
  23707=>"11111101",
  23708=>"11111101",
  23709=>"00000001",
  23710=>"00000001",
  23711=>"11111101",
  23712=>"00000011",
  23713=>"11111111",
  23714=>"11111110",
  23715=>"00000011",
  23716=>"00000000",
  23717=>"11111101",
  23718=>"00000010",
  23719=>"11111111",
  23720=>"11111110",
  23721=>"11111111",
  23722=>"11111110",
  23723=>"11111111",
  23724=>"11111111",
  23725=>"00000001",
  23726=>"00000000",
  23727=>"11111110",
  23728=>"00000010",
  23729=>"11111111",
  23730=>"00000000",
  23731=>"00000001",
  23732=>"00000000",
  23733=>"11111100",
  23734=>"00000000",
  23735=>"11111101",
  23736=>"11111110",
  23737=>"00000001",
  23738=>"00000000",
  23739=>"00000000",
  23740=>"11111110",
  23741=>"11111101",
  23742=>"00000000",
  23743=>"11111110",
  23744=>"11111111",
  23745=>"00000001",
  23746=>"00000010",
  23747=>"00000101",
  23748=>"00000010",
  23749=>"00000100",
  23750=>"00000000",
  23751=>"11111110",
  23752=>"00000000",
  23753=>"00000011",
  23754=>"00000000",
  23755=>"11111110",
  23756=>"00000000",
  23757=>"11111110",
  23758=>"11111110",
  23759=>"11111100",
  23760=>"00000010",
  23761=>"00000001",
  23762=>"00000010",
  23763=>"00000010",
  23764=>"00000010",
  23765=>"11111011",
  23766=>"00000000",
  23767=>"11111111",
  23768=>"00000000",
  23769=>"00000001",
  23770=>"00000001",
  23771=>"00000100",
  23772=>"00000001",
  23773=>"11111110",
  23774=>"11111110",
  23775=>"11111100",
  23776=>"00000001",
  23777=>"00000010",
  23778=>"00000010",
  23779=>"00000000",
  23780=>"00000000",
  23781=>"11111110",
  23782=>"00000011",
  23783=>"11111111",
  23784=>"00000011",
  23785=>"11111111",
  23786=>"00000000",
  23787=>"11111110",
  23788=>"00000001",
  23789=>"00000100",
  23790=>"11111110",
  23791=>"11111110",
  23792=>"11111110",
  23793=>"11111101",
  23794=>"11111110",
  23795=>"00000000",
  23796=>"11111111",
  23797=>"11111101",
  23798=>"00000000",
  23799=>"00000011",
  23800=>"00000100",
  23801=>"00000000",
  23802=>"00000000",
  23803=>"00000000",
  23804=>"00000100",
  23805=>"00000100",
  23806=>"00000001",
  23807=>"00000001",
  23808=>"00000001",
  23809=>"11111111",
  23810=>"11111100",
  23811=>"00000000",
  23812=>"00000001",
  23813=>"11111101",
  23814=>"00000011",
  23815=>"00000100",
  23816=>"00000010",
  23817=>"11111110",
  23818=>"00000100",
  23819=>"11111111",
  23820=>"00000010",
  23821=>"11111011",
  23822=>"00000001",
  23823=>"11111110",
  23824=>"11111101",
  23825=>"00000001",
  23826=>"00000000",
  23827=>"00000000",
  23828=>"00000001",
  23829=>"11111110",
  23830=>"11111111",
  23831=>"00000001",
  23832=>"00000000",
  23833=>"00000011",
  23834=>"00000000",
  23835=>"00000000",
  23836=>"00000100",
  23837=>"00000010",
  23838=>"11111101",
  23839=>"11111111",
  23840=>"11111111",
  23841=>"11111110",
  23842=>"00000010",
  23843=>"11111111",
  23844=>"11111111",
  23845=>"00000101",
  23846=>"00000010",
  23847=>"11111110",
  23848=>"00000100",
  23849=>"00000010",
  23850=>"11111111",
  23851=>"00000100",
  23852=>"00000001",
  23853=>"00000001",
  23854=>"11111110",
  23855=>"00000010",
  23856=>"11111111",
  23857=>"00000000",
  23858=>"11111111",
  23859=>"11111101",
  23860=>"00000011",
  23861=>"00000010",
  23862=>"00000010",
  23863=>"00000000",
  23864=>"00000001",
  23865=>"11111110",
  23866=>"11111110",
  23867=>"00000000",
  23868=>"11111101",
  23869=>"11111110",
  23870=>"00000110",
  23871=>"00000000",
  23872=>"00000000",
  23873=>"00000001",
  23874=>"00000100",
  23875=>"00000010",
  23876=>"00000001",
  23877=>"00000001",
  23878=>"00000101",
  23879=>"00000001",
  23880=>"11111111",
  23881=>"00000010",
  23882=>"11111111",
  23883=>"11111101",
  23884=>"11111101",
  23885=>"00000001",
  23886=>"00000011",
  23887=>"11111111",
  23888=>"11111101",
  23889=>"11111110",
  23890=>"00000010",
  23891=>"11111100",
  23892=>"00000010",
  23893=>"00000001",
  23894=>"00000000",
  23895=>"00000001",
  23896=>"00000010",
  23897=>"00000011",
  23898=>"00000010",
  23899=>"00000010",
  23900=>"00000100",
  23901=>"00000000",
  23902=>"00000001",
  23903=>"11111110",
  23904=>"00000001",
  23905=>"11111110",
  23906=>"11111110",
  23907=>"11111110",
  23908=>"11111110",
  23909=>"11111110",
  23910=>"00000001",
  23911=>"00000000",
  23912=>"00000011",
  23913=>"11111111",
  23914=>"00000000",
  23915=>"11111111",
  23916=>"00000101",
  23917=>"00000000",
  23918=>"11111100",
  23919=>"11111100",
  23920=>"00000000",
  23921=>"00000001",
  23922=>"00000000",
  23923=>"00000011",
  23924=>"11111101",
  23925=>"00000011",
  23926=>"11111110",
  23927=>"00000011",
  23928=>"00000000",
  23929=>"00000101",
  23930=>"00000010",
  23931=>"11111111",
  23932=>"00000000",
  23933=>"00000000",
  23934=>"00000001",
  23935=>"11111111",
  23936=>"00000001",
  23937=>"11111111",
  23938=>"11111110",
  23939=>"00000011",
  23940=>"00000000",
  23941=>"11111110",
  23942=>"11111111",
  23943=>"11111110",
  23944=>"00000001",
  23945=>"00000001",
  23946=>"00000001",
  23947=>"00000000",
  23948=>"11111110",
  23949=>"00000100",
  23950=>"00000001",
  23951=>"00000011",
  23952=>"00000000",
  23953=>"00000001",
  23954=>"00000000",
  23955=>"00000000",
  23956=>"11111110",
  23957=>"00000011",
  23958=>"11111111",
  23959=>"11111111",
  23960=>"00000010",
  23961=>"00000000",
  23962=>"00000000",
  23963=>"00000000",
  23964=>"00000000",
  23965=>"11111111",
  23966=>"11111110",
  23967=>"00000000",
  23968=>"00000010",
  23969=>"00000000",
  23970=>"11111111",
  23971=>"11111110",
  23972=>"00000011",
  23973=>"00000001",
  23974=>"11111110",
  23975=>"00000000",
  23976=>"11111111",
  23977=>"11111101",
  23978=>"11111101",
  23979=>"00000010",
  23980=>"00000010",
  23981=>"00000000",
  23982=>"00000010",
  23983=>"11111110",
  23984=>"11111101",
  23985=>"11111101",
  23986=>"11111100",
  23987=>"00000000",
  23988=>"00000001",
  23989=>"11111111",
  23990=>"00000000",
  23991=>"11111111",
  23992=>"00000001",
  23993=>"11111101",
  23994=>"00000001",
  23995=>"00000000",
  23996=>"00000001",
  23997=>"00000011",
  23998=>"00000010",
  23999=>"00000000",
  24000=>"11111111",
  24001=>"11111101",
  24002=>"00000000",
  24003=>"00000010",
  24004=>"00000100",
  24005=>"00000011",
  24006=>"11111110",
  24007=>"00000000",
  24008=>"11111101",
  24009=>"11111101",
  24010=>"11111111",
  24011=>"00000010",
  24012=>"00000000",
  24013=>"00000011",
  24014=>"00000000",
  24015=>"00000010",
  24016=>"11111110",
  24017=>"11111111",
  24018=>"00000001",
  24019=>"11111101",
  24020=>"00000001",
  24021=>"11111011",
  24022=>"00000001",
  24023=>"00000000",
  24024=>"11111111",
  24025=>"11111100",
  24026=>"00000010",
  24027=>"00000100",
  24028=>"11111110",
  24029=>"00000000",
  24030=>"00000000",
  24031=>"00000001",
  24032=>"00000001",
  24033=>"11111100",
  24034=>"11111110",
  24035=>"00000001",
  24036=>"11111110",
  24037=>"11111111",
  24038=>"11111111",
  24039=>"11111110",
  24040=>"00000001",
  24041=>"00000000",
  24042=>"11111110",
  24043=>"11111101",
  24044=>"00000001",
  24045=>"00000001",
  24046=>"00000010",
  24047=>"00000000",
  24048=>"00000001",
  24049=>"11111101",
  24050=>"00000001",
  24051=>"11111111",
  24052=>"11111110",
  24053=>"11111101",
  24054=>"11111100",
  24055=>"00000100",
  24056=>"11111111",
  24057=>"00000010",
  24058=>"11111111",
  24059=>"00000000",
  24060=>"11111111",
  24061=>"00000000",
  24062=>"11111110",
  24063=>"00000010",
  24064=>"00000010",
  24065=>"11111110",
  24066=>"00000000",
  24067=>"00000011",
  24068=>"00000000",
  24069=>"00000100",
  24070=>"11111011",
  24071=>"00000100",
  24072=>"11111111",
  24073=>"11111101",
  24074=>"11111110",
  24075=>"00000010",
  24076=>"00000010",
  24077=>"11111101",
  24078=>"00000010",
  24079=>"11111110",
  24080=>"00000000",
  24081=>"00000000",
  24082=>"00000011",
  24083=>"00000011",
  24084=>"00000000",
  24085=>"11111101",
  24086=>"11111110",
  24087=>"11111110",
  24088=>"00000101",
  24089=>"00000010",
  24090=>"00000001",
  24091=>"11111101",
  24092=>"11111111",
  24093=>"00000011",
  24094=>"11111110",
  24095=>"11111101",
  24096=>"00000010",
  24097=>"00000000",
  24098=>"11111111",
  24099=>"11111111",
  24100=>"00000000",
  24101=>"00000001",
  24102=>"00000000",
  24103=>"00000111",
  24104=>"11111111",
  24105=>"00000001",
  24106=>"00000001",
  24107=>"11111110",
  24108=>"11111111",
  24109=>"00000000",
  24110=>"00000000",
  24111=>"00000010",
  24112=>"00000101",
  24113=>"11111101",
  24114=>"00000000",
  24115=>"00000001",
  24116=>"11111111",
  24117=>"00000000",
  24118=>"00000011",
  24119=>"00000001",
  24120=>"11111111",
  24121=>"00000000",
  24122=>"11111111",
  24123=>"00000010",
  24124=>"11111101",
  24125=>"11111111",
  24126=>"00000100",
  24127=>"11111110",
  24128=>"11111100",
  24129=>"11111110",
  24130=>"00000000",
  24131=>"00000000",
  24132=>"00000000",
  24133=>"00000010",
  24134=>"11111110",
  24135=>"11111101",
  24136=>"11111111",
  24137=>"00000000",
  24138=>"11111110",
  24139=>"11111101",
  24140=>"00000001",
  24141=>"00000000",
  24142=>"00000100",
  24143=>"00000000",
  24144=>"00000010",
  24145=>"11111111",
  24146=>"11111110",
  24147=>"11111111",
  24148=>"11111111",
  24149=>"11111110",
  24150=>"00000001",
  24151=>"11111111",
  24152=>"00000001",
  24153=>"11111111",
  24154=>"00000010",
  24155=>"00000000",
  24156=>"11111101",
  24157=>"00000010",
  24158=>"00000000",
  24159=>"11111110",
  24160=>"11111110",
  24161=>"11111101",
  24162=>"00000000",
  24163=>"00000011",
  24164=>"11111101",
  24165=>"11111101",
  24166=>"00000011",
  24167=>"00000001",
  24168=>"11111111",
  24169=>"11111110",
  24170=>"00000010",
  24171=>"00000001",
  24172=>"00000000",
  24173=>"00000001",
  24174=>"00000001",
  24175=>"00000100",
  24176=>"11111101",
  24177=>"00000010",
  24178=>"00000011",
  24179=>"11111101",
  24180=>"00000010",
  24181=>"00000000",
  24182=>"11111111",
  24183=>"00000010",
  24184=>"11111101",
  24185=>"00000000",
  24186=>"00000010",
  24187=>"11111111",
  24188=>"11111110",
  24189=>"00000001",
  24190=>"00000010",
  24191=>"11111110",
  24192=>"00000001",
  24193=>"00000011",
  24194=>"11111101",
  24195=>"00000011",
  24196=>"11111110",
  24197=>"11111100",
  24198=>"11111111",
  24199=>"11111111",
  24200=>"11111110",
  24201=>"11111101",
  24202=>"11111111",
  24203=>"00000010",
  24204=>"00000001",
  24205=>"00000001",
  24206=>"11111111",
  24207=>"00000001",
  24208=>"11111111",
  24209=>"11111110",
  24210=>"00000011",
  24211=>"11111111",
  24212=>"00000001",
  24213=>"11111111",
  24214=>"00000001",
  24215=>"00000011",
  24216=>"00000001",
  24217=>"00000101",
  24218=>"11111101",
  24219=>"00000010",
  24220=>"00000000",
  24221=>"11111110",
  24222=>"11111101",
  24223=>"00000101",
  24224=>"11111111",
  24225=>"11111110",
  24226=>"00000001",
  24227=>"11111111",
  24228=>"11111111",
  24229=>"11111101",
  24230=>"00000001",
  24231=>"00000001",
  24232=>"11111100",
  24233=>"00000100",
  24234=>"11111110",
  24235=>"00000001",
  24236=>"00000001",
  24237=>"00000001",
  24238=>"00000001",
  24239=>"11111110",
  24240=>"11111110",
  24241=>"11111111",
  24242=>"00000010",
  24243=>"00000010",
  24244=>"11111101",
  24245=>"11111110",
  24246=>"00000001",
  24247=>"00000011",
  24248=>"11111110",
  24249=>"00000000",
  24250=>"00000000",
  24251=>"00000000",
  24252=>"11111101",
  24253=>"00000001",
  24254=>"11111111",
  24255=>"11111111",
  24256=>"00000100",
  24257=>"00000100",
  24258=>"00000011",
  24259=>"11111111",
  24260=>"00000010",
  24261=>"11111111",
  24262=>"00000000",
  24263=>"11111101",
  24264=>"00000000",
  24265=>"11111101",
  24266=>"00000000",
  24267=>"11111110",
  24268=>"00000010",
  24269=>"11111110",
  24270=>"00000000",
  24271=>"00000010",
  24272=>"11111101",
  24273=>"11111111",
  24274=>"00000010",
  24275=>"11111100",
  24276=>"00000010",
  24277=>"00000010",
  24278=>"00000001",
  24279=>"00000010",
  24280=>"00000000",
  24281=>"11111110",
  24282=>"11111111",
  24283=>"00000010",
  24284=>"11111011",
  24285=>"00000001",
  24286=>"00000011",
  24287=>"00000111",
  24288=>"00000000",
  24289=>"00000100",
  24290=>"11111101",
  24291=>"00000000",
  24292=>"11111111",
  24293=>"00000100",
  24294=>"00000000",
  24295=>"00000010",
  24296=>"00000011",
  24297=>"00000000",
  24298=>"00000000",
  24299=>"00000001",
  24300=>"00000011",
  24301=>"00000000",
  24302=>"00000011",
  24303=>"00000110",
  24304=>"11111101",
  24305=>"00000000",
  24306=>"00000010",
  24307=>"11111101",
  24308=>"11111101",
  24309=>"11111111",
  24310=>"00000100",
  24311=>"00000000",
  24312=>"11111101",
  24313=>"00000000",
  24314=>"00000010",
  24315=>"11111111",
  24316=>"11111101",
  24317=>"00000010",
  24318=>"11111101",
  24319=>"00000000",
  24320=>"00000001",
  24321=>"00000000",
  24322=>"11111101",
  24323=>"00000110",
  24324=>"11111101",
  24325=>"00000100",
  24326=>"00000001",
  24327=>"11111100",
  24328=>"11111110",
  24329=>"00000011",
  24330=>"00000001",
  24331=>"11111101",
  24332=>"00000001",
  24333=>"00000000",
  24334=>"11111110",
  24335=>"00000001",
  24336=>"00000010",
  24337=>"11111111",
  24338=>"00000000",
  24339=>"11111101",
  24340=>"00000010",
  24341=>"00000000",
  24342=>"00000000",
  24343=>"00000100",
  24344=>"11111011",
  24345=>"00000001",
  24346=>"11111111",
  24347=>"11111110",
  24348=>"11111110",
  24349=>"11111111",
  24350=>"00000000",
  24351=>"00000100",
  24352=>"00000011",
  24353=>"00000010",
  24354=>"00000000",
  24355=>"00000000",
  24356=>"00000100",
  24357=>"11111110",
  24358=>"00000001",
  24359=>"11111101",
  24360=>"00000001",
  24361=>"11111110",
  24362=>"11111111",
  24363=>"11111110",
  24364=>"00000001",
  24365=>"00000001",
  24366=>"00000011",
  24367=>"00000001",
  24368=>"00000010",
  24369=>"00000010",
  24370=>"00000011",
  24371=>"00000001",
  24372=>"11111110",
  24373=>"11111111",
  24374=>"00000001",
  24375=>"11111101",
  24376=>"11111101",
  24377=>"00000010",
  24378=>"11111110",
  24379=>"11111111",
  24380=>"11111101",
  24381=>"00000011",
  24382=>"11111110",
  24383=>"11111111",
  24384=>"00000110",
  24385=>"00000000",
  24386=>"11111110",
  24387=>"00000011",
  24388=>"00000010",
  24389=>"00000010",
  24390=>"00000001",
  24391=>"00000000",
  24392=>"11111110",
  24393=>"11111110",
  24394=>"00000001",
  24395=>"11111111",
  24396=>"00000011",
  24397=>"00000001",
  24398=>"00001000",
  24399=>"00000001",
  24400=>"11111110",
  24401=>"00000010",
  24402=>"00000010",
  24403=>"00000001",
  24404=>"11111111",
  24405=>"00000000",
  24406=>"00000000",
  24407=>"11111111",
  24408=>"11111101",
  24409=>"00000010",
  24410=>"00000010",
  24411=>"11111110",
  24412=>"00000011",
  24413=>"00000100",
  24414=>"00000011",
  24415=>"00000100",
  24416=>"00000010",
  24417=>"11111110",
  24418=>"11111110",
  24419=>"11111111",
  24420=>"11111101",
  24421=>"11111110",
  24422=>"11111100",
  24423=>"00000011",
  24424=>"11111111",
  24425=>"00000011",
  24426=>"00000010",
  24427=>"11111111",
  24428=>"00000001",
  24429=>"00000010",
  24430=>"11111110",
  24431=>"00000001",
  24432=>"00000001",
  24433=>"00000101",
  24434=>"11111110",
  24435=>"11111110",
  24436=>"11111110",
  24437=>"00000110",
  24438=>"11111111",
  24439=>"11111111",
  24440=>"11111111",
  24441=>"11111111",
  24442=>"00000100",
  24443=>"00000001",
  24444=>"11111110",
  24445=>"00000001",
  24446=>"11111101",
  24447=>"00000100",
  24448=>"00000010",
  24449=>"11111111",
  24450=>"11111111",
  24451=>"11111101",
  24452=>"00000010",
  24453=>"00000000",
  24454=>"00000000",
  24455=>"11111101",
  24456=>"11111111",
  24457=>"00000001",
  24458=>"00000001",
  24459=>"00000010",
  24460=>"11111110",
  24461=>"00000011",
  24462=>"00000001",
  24463=>"00000010",
  24464=>"00000010",
  24465=>"00000100",
  24466=>"00000010",
  24467=>"11111110",
  24468=>"00000010",
  24469=>"11111110",
  24470=>"11111111",
  24471=>"11111111",
  24472=>"00000100",
  24473=>"00000000",
  24474=>"00000001",
  24475=>"00000010",
  24476=>"00000001",
  24477=>"11111110",
  24478=>"00000011",
  24479=>"00000010",
  24480=>"00000000",
  24481=>"11111111",
  24482=>"00000001",
  24483=>"11111110",
  24484=>"00000001",
  24485=>"00000000",
  24486=>"11111111",
  24487=>"11111111",
  24488=>"00000010",
  24489=>"11111110",
  24490=>"11111111",
  24491=>"11111110",
  24492=>"11111101",
  24493=>"00000011",
  24494=>"00000011",
  24495=>"00000011",
  24496=>"00000011",
  24497=>"00000010",
  24498=>"00000100",
  24499=>"00000001",
  24500=>"11111101",
  24501=>"11111111",
  24502=>"11111101",
  24503=>"00000110",
  24504=>"00000100",
  24505=>"00000100",
  24506=>"00000011",
  24507=>"00000001",
  24508=>"00000011",
  24509=>"00000001",
  24510=>"00000000",
  24511=>"11111111",
  24512=>"11111111",
  24513=>"00000001",
  24514=>"00000010",
  24515=>"00000000",
  24516=>"11111110",
  24517=>"11111101",
  24518=>"00000000",
  24519=>"00000010",
  24520=>"11111101",
  24521=>"00000000",
  24522=>"11111110",
  24523=>"11111110",
  24524=>"00000010",
  24525=>"11111110",
  24526=>"11111101",
  24527=>"11111111",
  24528=>"00000100",
  24529=>"11111110",
  24530=>"00000011",
  24531=>"11111101",
  24532=>"00000000",
  24533=>"00000101",
  24534=>"00000011",
  24535=>"00000001",
  24536=>"00000011",
  24537=>"00000010",
  24538=>"11111101",
  24539=>"00000110",
  24540=>"00000011",
  24541=>"00000000",
  24542=>"11111111",
  24543=>"00000001",
  24544=>"11111111",
  24545=>"11111110",
  24546=>"11111100",
  24547=>"11111110",
  24548=>"11111101",
  24549=>"00000000",
  24550=>"11111110",
  24551=>"11111110",
  24552=>"11111111",
  24553=>"11111111",
  24554=>"00000100",
  24555=>"00000101",
  24556=>"11111110",
  24557=>"00000001",
  24558=>"11111100",
  24559=>"11111101",
  24560=>"00000011",
  24561=>"11111101",
  24562=>"00000001",
  24563=>"11111111",
  24564=>"11111110",
  24565=>"11111101",
  24566=>"00000101",
  24567=>"11111101",
  24568=>"00000001",
  24569=>"00000011",
  24570=>"00000101",
  24571=>"00000001",
  24572=>"00000010",
  24573=>"11111101",
  24574=>"11111101",
  24575=>"11111100",
  24576=>"11111111",
  24577=>"11111101",
  24578=>"11111111",
  24579=>"11111111",
  24580=>"00000000",
  24581=>"00000010",
  24582=>"00000010",
  24583=>"00000010",
  24584=>"00000010",
  24585=>"00000001",
  24586=>"00000000",
  24587=>"00000000",
  24588=>"00000101",
  24589=>"00000011",
  24590=>"00000001",
  24591=>"00000100",
  24592=>"00000010",
  24593=>"00000001",
  24594=>"11111110",
  24595=>"00000011",
  24596=>"00000010",
  24597=>"11111110",
  24598=>"11111111",
  24599=>"00000010",
  24600=>"11111110",
  24601=>"00000010",
  24602=>"11111100",
  24603=>"00000000",
  24604=>"11111101",
  24605=>"11111101",
  24606=>"00000001",
  24607=>"11111101",
  24608=>"11111110",
  24609=>"11111111",
  24610=>"00000000",
  24611=>"11111101",
  24612=>"00000001",
  24613=>"11111111",
  24614=>"00000101",
  24615=>"00000011",
  24616=>"00000011",
  24617=>"00000010",
  24618=>"11111110",
  24619=>"00000000",
  24620=>"11111111",
  24621=>"00000010",
  24622=>"00000001",
  24623=>"00000000",
  24624=>"00000000",
  24625=>"00000101",
  24626=>"11111110",
  24627=>"00000001",
  24628=>"00000010",
  24629=>"11111111",
  24630=>"11111110",
  24631=>"11111110",
  24632=>"11111110",
  24633=>"11111101",
  24634=>"00000010",
  24635=>"11111111",
  24636=>"00000100",
  24637=>"00000010",
  24638=>"00000001",
  24639=>"00000001",
  24640=>"11111101",
  24641=>"00000000",
  24642=>"00000010",
  24643=>"00000100",
  24644=>"00000001",
  24645=>"00000001",
  24646=>"00000000",
  24647=>"11111110",
  24648=>"11111111",
  24649=>"00000011",
  24650=>"00000001",
  24651=>"00000011",
  24652=>"00000001",
  24653=>"11111111",
  24654=>"11111101",
  24655=>"00000000",
  24656=>"11111101",
  24657=>"00000001",
  24658=>"11111100",
  24659=>"11111100",
  24660=>"00000100",
  24661=>"11111110",
  24662=>"11111110",
  24663=>"11111101",
  24664=>"11111111",
  24665=>"11111111",
  24666=>"11111110",
  24667=>"00000001",
  24668=>"11111101",
  24669=>"11111101",
  24670=>"00000001",
  24671=>"11111101",
  24672=>"11111111",
  24673=>"00000000",
  24674=>"11111110",
  24675=>"11111101",
  24676=>"11111101",
  24677=>"00000011",
  24678=>"11111110",
  24679=>"00000001",
  24680=>"00000000",
  24681=>"11111101",
  24682=>"11111111",
  24683=>"00000001",
  24684=>"00000000",
  24685=>"11111110",
  24686=>"11111101",
  24687=>"00000001",
  24688=>"00000101",
  24689=>"11111110",
  24690=>"00000001",
  24691=>"00000000",
  24692=>"11111110",
  24693=>"00000001",
  24694=>"00000001",
  24695=>"00000001",
  24696=>"00000110",
  24697=>"00000101",
  24698=>"11111111",
  24699=>"00000001",
  24700=>"00000100",
  24701=>"11111101",
  24702=>"11111101",
  24703=>"11111111",
  24704=>"00000001",
  24705=>"11111110",
  24706=>"11111110",
  24707=>"11111110",
  24708=>"11111101",
  24709=>"00000000",
  24710=>"00000010",
  24711=>"00000011",
  24712=>"00000010",
  24713=>"00000011",
  24714=>"00000000",
  24715=>"11111101",
  24716=>"11111111",
  24717=>"00000001",
  24718=>"00000011",
  24719=>"11111101",
  24720=>"11111111",
  24721=>"11111111",
  24722=>"00000001",
  24723=>"00000001",
  24724=>"11111101",
  24725=>"11111111",
  24726=>"11111110",
  24727=>"00000101",
  24728=>"11111101",
  24729=>"00000100",
  24730=>"00000000",
  24731=>"11111101",
  24732=>"00000010",
  24733=>"00000011",
  24734=>"11111111",
  24735=>"11111101",
  24736=>"11111101",
  24737=>"11111111",
  24738=>"00000100",
  24739=>"11111101",
  24740=>"11111111",
  24741=>"00000010",
  24742=>"00000100",
  24743=>"00000101",
  24744=>"00000010",
  24745=>"00000000",
  24746=>"11111101",
  24747=>"00000000",
  24748=>"00000001",
  24749=>"00000010",
  24750=>"00000100",
  24751=>"00000001",
  24752=>"11111101",
  24753=>"00000010",
  24754=>"11111110",
  24755=>"11111111",
  24756=>"00000000",
  24757=>"00000001",
  24758=>"11111110",
  24759=>"00000010",
  24760=>"00000010",
  24761=>"11111101",
  24762=>"00000101",
  24763=>"11111110",
  24764=>"11111101",
  24765=>"11111111",
  24766=>"00000000",
  24767=>"11111101",
  24768=>"00000011",
  24769=>"11111111",
  24770=>"11111111",
  24771=>"11111101",
  24772=>"00000011",
  24773=>"11111110",
  24774=>"11111101",
  24775=>"00000000",
  24776=>"00000000",
  24777=>"11111100",
  24778=>"11111111",
  24779=>"00000010",
  24780=>"00000011",
  24781=>"11111111",
  24782=>"00000001",
  24783=>"11111110",
  24784=>"00000001",
  24785=>"11111100",
  24786=>"00000000",
  24787=>"11111111",
  24788=>"00000001",
  24789=>"00000010",
  24790=>"11111110",
  24791=>"11111101",
  24792=>"00000111",
  24793=>"11111110",
  24794=>"00000010",
  24795=>"11111101",
  24796=>"00000001",
  24797=>"11111111",
  24798=>"11111101",
  24799=>"11111110",
  24800=>"00000001",
  24801=>"00000001",
  24802=>"00000000",
  24803=>"00000001",
  24804=>"11111111",
  24805=>"00000000",
  24806=>"00000011",
  24807=>"00000001",
  24808=>"00000001",
  24809=>"00000001",
  24810=>"11111101",
  24811=>"00000000",
  24812=>"00000000",
  24813=>"00000011",
  24814=>"00000010",
  24815=>"11111111",
  24816=>"11111100",
  24817=>"11111101",
  24818=>"00000000",
  24819=>"00000000",
  24820=>"11111110",
  24821=>"00000010",
  24822=>"00000001",
  24823=>"11111110",
  24824=>"11111100",
  24825=>"11111111",
  24826=>"11111110",
  24827=>"00000000",
  24828=>"11111111",
  24829=>"11111111",
  24830=>"00000010",
  24831=>"00000011",
  24832=>"11111111",
  24833=>"00000000",
  24834=>"11111110",
  24835=>"00000000",
  24836=>"00000010",
  24837=>"11111111",
  24838=>"11111111",
  24839=>"11111111",
  24840=>"00000000",
  24841=>"11111111",
  24842=>"11111100",
  24843=>"11111101",
  24844=>"00000000",
  24845=>"00000100",
  24846=>"11111111",
  24847=>"11111110",
  24848=>"11111100",
  24849=>"11111101",
  24850=>"11111111",
  24851=>"11111110",
  24852=>"00000100",
  24853=>"00000010",
  24854=>"11111101",
  24855=>"00000011",
  24856=>"11111101",
  24857=>"11111111",
  24858=>"00000010",
  24859=>"00000000",
  24860=>"11111111",
  24861=>"00000000",
  24862=>"00000000",
  24863=>"00000010",
  24864=>"00000001",
  24865=>"00000001",
  24866=>"00000000",
  24867=>"00000001",
  24868=>"00000000",
  24869=>"00000101",
  24870=>"11111101",
  24871=>"00000011",
  24872=>"11111111",
  24873=>"11111101",
  24874=>"11111101",
  24875=>"11111101",
  24876=>"00000011",
  24877=>"00000000",
  24878=>"00000010",
  24879=>"00000011",
  24880=>"00000000",
  24881=>"00000001",
  24882=>"00000010",
  24883=>"11111111",
  24884=>"00000010",
  24885=>"11111101",
  24886=>"11111111",
  24887=>"00000010",
  24888=>"11111111",
  24889=>"00000101",
  24890=>"11111111",
  24891=>"00000010",
  24892=>"00000000",
  24893=>"00000010",
  24894=>"00000000",
  24895=>"11111110",
  24896=>"00000001",
  24897=>"11111110",
  24898=>"00000010",
  24899=>"00000011",
  24900=>"11111110",
  24901=>"00000011",
  24902=>"11111111",
  24903=>"00000000",
  24904=>"11111110",
  24905=>"00000000",
  24906=>"00000001",
  24907=>"00000010",
  24908=>"11111100",
  24909=>"11111111",
  24910=>"00000010",
  24911=>"00000001",
  24912=>"00000010",
  24913=>"00000010",
  24914=>"11111101",
  24915=>"00000101",
  24916=>"11111101",
  24917=>"00000000",
  24918=>"00000011",
  24919=>"00000000",
  24920=>"11111110",
  24921=>"11111111",
  24922=>"11111110",
  24923=>"00000010",
  24924=>"11111111",
  24925=>"00000010",
  24926=>"00000101",
  24927=>"00000001",
  24928=>"11111111",
  24929=>"00000011",
  24930=>"00000000",
  24931=>"11111110",
  24932=>"00000001",
  24933=>"11111111",
  24934=>"00000010",
  24935=>"00000010",
  24936=>"11111110",
  24937=>"11111111",
  24938=>"00000001",
  24939=>"11111101",
  24940=>"00000010",
  24941=>"11111111",
  24942=>"00000101",
  24943=>"00000000",
  24944=>"00000000",
  24945=>"00000010",
  24946=>"11111110",
  24947=>"11111111",
  24948=>"11111111",
  24949=>"00000111",
  24950=>"00000100",
  24951=>"00000000",
  24952=>"11111101",
  24953=>"11111100",
  24954=>"11111111",
  24955=>"11111110",
  24956=>"11111101",
  24957=>"11111110",
  24958=>"11111110",
  24959=>"11111111",
  24960=>"00000011",
  24961=>"00000011",
  24962=>"00000000",
  24963=>"00000000",
  24964=>"11111101",
  24965=>"11111111",
  24966=>"11111110",
  24967=>"11111110",
  24968=>"00000001",
  24969=>"00000100",
  24970=>"11111111",
  24971=>"11111111",
  24972=>"00000001",
  24973=>"11111110",
  24974=>"00000011",
  24975=>"11111100",
  24976=>"00000011",
  24977=>"11111110",
  24978=>"00000001",
  24979=>"11111111",
  24980=>"11111100",
  24981=>"11111111",
  24982=>"00000010",
  24983=>"11111101",
  24984=>"00000010",
  24985=>"11111101",
  24986=>"00000010",
  24987=>"00000011",
  24988=>"11111110",
  24989=>"11111111",
  24990=>"11111111",
  24991=>"11111100",
  24992=>"11111111",
  24993=>"00000010",
  24994=>"00000000",
  24995=>"00000011",
  24996=>"11111111",
  24997=>"00000001",
  24998=>"00000001",
  24999=>"11111111",
  25000=>"00000010",
  25001=>"11111101",
  25002=>"00000001",
  25003=>"00000000",
  25004=>"11111111",
  25005=>"11111111",
  25006=>"11111111",
  25007=>"11111110",
  25008=>"11111111",
  25009=>"11111110",
  25010=>"00000000",
  25011=>"00000011",
  25012=>"00000010",
  25013=>"11111110",
  25014=>"00000110",
  25015=>"11111110",
  25016=>"11111110",
  25017=>"00000000",
  25018=>"11111110",
  25019=>"00000000",
  25020=>"11111101",
  25021=>"00000001",
  25022=>"00000001",
  25023=>"00000000",
  25024=>"11111111",
  25025=>"11111111",
  25026=>"11111100",
  25027=>"00000010",
  25028=>"11111111",
  25029=>"00000110",
  25030=>"00000011",
  25031=>"11111100",
  25032=>"00000110",
  25033=>"00000001",
  25034=>"11111111",
  25035=>"00000000",
  25036=>"00000010",
  25037=>"11111110",
  25038=>"00000000",
  25039=>"00000001",
  25040=>"11111110",
  25041=>"11111110",
  25042=>"11111111",
  25043=>"00000000",
  25044=>"11111111",
  25045=>"00000111",
  25046=>"11111101",
  25047=>"00000010",
  25048=>"11111111",
  25049=>"11111101",
  25050=>"00000000",
  25051=>"11111101",
  25052=>"00000100",
  25053=>"11111110",
  25054=>"00000001",
  25055=>"11111101",
  25056=>"00000001",
  25057=>"00000010",
  25058=>"11111110",
  25059=>"00000010",
  25060=>"00000001",
  25061=>"00000010",
  25062=>"00000001",
  25063=>"00000010",
  25064=>"11111111",
  25065=>"00000000",
  25066=>"11111101",
  25067=>"00000000",
  25068=>"00000000",
  25069=>"00000000",
  25070=>"11111110",
  25071=>"11111111",
  25072=>"00000000",
  25073=>"11111100",
  25074=>"11111111",
  25075=>"11111111",
  25076=>"11111110",
  25077=>"11111110",
  25078=>"00000011",
  25079=>"11111111",
  25080=>"00000101",
  25081=>"11111111",
  25082=>"00000001",
  25083=>"00000001",
  25084=>"00000001",
  25085=>"11111111",
  25086=>"00000001",
  25087=>"00000000",
  25088=>"00000000",
  25089=>"00000011",
  25090=>"11111101",
  25091=>"11111111",
  25092=>"00000010",
  25093=>"11111101",
  25094=>"11111100",
  25095=>"00000001",
  25096=>"11111111",
  25097=>"11111101",
  25098=>"00000010",
  25099=>"00000001",
  25100=>"00000001",
  25101=>"00000010",
  25102=>"11111101",
  25103=>"00000000",
  25104=>"11111101",
  25105=>"11111111",
  25106=>"00000001",
  25107=>"00000000",
  25108=>"00000000",
  25109=>"00000001",
  25110=>"00000001",
  25111=>"11111111",
  25112=>"11111100",
  25113=>"11111110",
  25114=>"00000010",
  25115=>"00000011",
  25116=>"00000011",
  25117=>"00000001",
  25118=>"11111111",
  25119=>"00000000",
  25120=>"00000010",
  25121=>"11111111",
  25122=>"00000010",
  25123=>"00000000",
  25124=>"00000001",
  25125=>"00000010",
  25126=>"00000011",
  25127=>"00000001",
  25128=>"00000010",
  25129=>"00000001",
  25130=>"00000001",
  25131=>"00000010",
  25132=>"00000000",
  25133=>"00000111",
  25134=>"11111111",
  25135=>"00000001",
  25136=>"11111100",
  25137=>"00000101",
  25138=>"11111101",
  25139=>"00000010",
  25140=>"11111111",
  25141=>"00000000",
  25142=>"00000001",
  25143=>"00000000",
  25144=>"00000011",
  25145=>"11111111",
  25146=>"00000000",
  25147=>"00000001",
  25148=>"11111110",
  25149=>"00000000",
  25150=>"11111110",
  25151=>"00000010",
  25152=>"11111110",
  25153=>"00000011",
  25154=>"00000001",
  25155=>"00000001",
  25156=>"00000101",
  25157=>"00000001",
  25158=>"00000011",
  25159=>"00000000",
  25160=>"11111111",
  25161=>"11111110",
  25162=>"11111111",
  25163=>"11111101",
  25164=>"00000011",
  25165=>"00000001",
  25166=>"00000100",
  25167=>"11111110",
  25168=>"00000001",
  25169=>"00000011",
  25170=>"11111110",
  25171=>"00000011",
  25172=>"11111111",
  25173=>"00000000",
  25174=>"00000001",
  25175=>"00000000",
  25176=>"11111101",
  25177=>"11111101",
  25178=>"11111111",
  25179=>"11111101",
  25180=>"00000001",
  25181=>"11111110",
  25182=>"00000001",
  25183=>"00000101",
  25184=>"11111111",
  25185=>"00000010",
  25186=>"00000010",
  25187=>"11111110",
  25188=>"11111110",
  25189=>"00000000",
  25190=>"00000011",
  25191=>"11111111",
  25192=>"00000000",
  25193=>"00000000",
  25194=>"00000001",
  25195=>"11111111",
  25196=>"00000011",
  25197=>"11111111",
  25198=>"00000000",
  25199=>"11111111",
  25200=>"00000000",
  25201=>"00000010",
  25202=>"11111111",
  25203=>"00000001",
  25204=>"00000001",
  25205=>"00000011",
  25206=>"11111110",
  25207=>"00000010",
  25208=>"11111101",
  25209=>"11111111",
  25210=>"00000001",
  25211=>"00000001",
  25212=>"00000011",
  25213=>"11111101",
  25214=>"00000010",
  25215=>"11111111",
  25216=>"00000010",
  25217=>"00000000",
  25218=>"00000010",
  25219=>"11111111",
  25220=>"00000000",
  25221=>"11111111",
  25222=>"11111111",
  25223=>"11111101",
  25224=>"00000000",
  25225=>"00000100",
  25226=>"00000001",
  25227=>"11111110",
  25228=>"11111111",
  25229=>"00000000",
  25230=>"00000001",
  25231=>"00000011",
  25232=>"11111110",
  25233=>"11111110",
  25234=>"11111110",
  25235=>"00000001",
  25236=>"11111100",
  25237=>"00000000",
  25238=>"00000001",
  25239=>"11111101",
  25240=>"11111111",
  25241=>"11111101",
  25242=>"00000011",
  25243=>"00000011",
  25244=>"00000000",
  25245=>"00000010",
  25246=>"00000000",
  25247=>"00000001",
  25248=>"11111110",
  25249=>"00000011",
  25250=>"00000001",
  25251=>"00000001",
  25252=>"00000011",
  25253=>"11111111",
  25254=>"00000010",
  25255=>"00000001",
  25256=>"11111110",
  25257=>"00000000",
  25258=>"00000000",
  25259=>"00000000",
  25260=>"11111101",
  25261=>"11111111",
  25262=>"11111110",
  25263=>"00000001",
  25264=>"00000001",
  25265=>"11111111",
  25266=>"11111110",
  25267=>"00000000",
  25268=>"11111111",
  25269=>"00000000",
  25270=>"00000001",
  25271=>"00000000",
  25272=>"00000000",
  25273=>"11111111",
  25274=>"00000000",
  25275=>"00000010",
  25276=>"11111101",
  25277=>"00000101",
  25278=>"00000010",
  25279=>"11111110",
  25280=>"00000000",
  25281=>"00000011",
  25282=>"00000101",
  25283=>"00000000",
  25284=>"00000010",
  25285=>"00000101",
  25286=>"00000011",
  25287=>"11111100",
  25288=>"11111111",
  25289=>"00000001",
  25290=>"00000000",
  25291=>"00000000",
  25292=>"11111100",
  25293=>"00000011",
  25294=>"00000100",
  25295=>"00000001",
  25296=>"00000001",
  25297=>"11111110",
  25298=>"11111101",
  25299=>"00000011",
  25300=>"00000001",
  25301=>"00000001",
  25302=>"00000000",
  25303=>"00000000",
  25304=>"00000001",
  25305=>"00000100",
  25306=>"11111111",
  25307=>"00000000",
  25308=>"00000000",
  25309=>"11111110",
  25310=>"00000000",
  25311=>"11111101",
  25312=>"00000001",
  25313=>"11111110",
  25314=>"00000000",
  25315=>"00000001",
  25316=>"11111101",
  25317=>"00000000",
  25318=>"00000010",
  25319=>"00000001",
  25320=>"11111110",
  25321=>"11111110",
  25322=>"11111110",
  25323=>"11111110",
  25324=>"11111101",
  25325=>"11111110",
  25326=>"00000000",
  25327=>"11111111",
  25328=>"11111110",
  25329=>"00000011",
  25330=>"00000000",
  25331=>"11111111",
  25332=>"00000011",
  25333=>"00000010",
  25334=>"11111110",
  25335=>"11111110",
  25336=>"00000010",
  25337=>"00000001",
  25338=>"00000000",
  25339=>"00000000",
  25340=>"00000001",
  25341=>"00000001",
  25342=>"00000011",
  25343=>"00000000",
  25344=>"11111101",
  25345=>"11111111",
  25346=>"00000010",
  25347=>"11111110",
  25348=>"00000010",
  25349=>"00000000",
  25350=>"11111110",
  25351=>"11111101",
  25352=>"00000010",
  25353=>"11111111",
  25354=>"11111110",
  25355=>"00000000",
  25356=>"11111111",
  25357=>"11111101",
  25358=>"11111110",
  25359=>"00000010",
  25360=>"00000100",
  25361=>"00000010",
  25362=>"00000011",
  25363=>"00000100",
  25364=>"00000001",
  25365=>"11111111",
  25366=>"00000000",
  25367=>"00000000",
  25368=>"00000101",
  25369=>"11111110",
  25370=>"11111110",
  25371=>"00000011",
  25372=>"11111110",
  25373=>"11111100",
  25374=>"11111110",
  25375=>"11111111",
  25376=>"11111111",
  25377=>"11111101",
  25378=>"00000001",
  25379=>"11111111",
  25380=>"00000001",
  25381=>"00000000",
  25382=>"11111111",
  25383=>"00000010",
  25384=>"00001000",
  25385=>"11111111",
  25386=>"00000000",
  25387=>"11111111",
  25388=>"00000100",
  25389=>"00000001",
  25390=>"11111101",
  25391=>"00000011",
  25392=>"00000001",
  25393=>"11111101",
  25394=>"11111101",
  25395=>"11111111",
  25396=>"00000000",
  25397=>"11111101",
  25398=>"11111101",
  25399=>"00000001",
  25400=>"11111111",
  25401=>"11111111",
  25402=>"11111101",
  25403=>"00000000",
  25404=>"11111110",
  25405=>"00000000",
  25406=>"00000001",
  25407=>"00000100",
  25408=>"11111110",
  25409=>"00000000",
  25410=>"11111101",
  25411=>"11111101",
  25412=>"11111101",
  25413=>"00000000",
  25414=>"11111111",
  25415=>"00000011",
  25416=>"00000000",
  25417=>"00000010",
  25418=>"00000000",
  25419=>"11111110",
  25420=>"00000000",
  25421=>"00000001",
  25422=>"00000000",
  25423=>"11111101",
  25424=>"00000110",
  25425=>"11111101",
  25426=>"11111111",
  25427=>"11111111",
  25428=>"11111110",
  25429=>"00000000",
  25430=>"00000011",
  25431=>"00000100",
  25432=>"11111111",
  25433=>"00000010",
  25434=>"11111101",
  25435=>"00000010",
  25436=>"11111110",
  25437=>"00000101",
  25438=>"11111111",
  25439=>"11111111",
  25440=>"11111101",
  25441=>"00000000",
  25442=>"00000001",
  25443=>"11111100",
  25444=>"11111111",
  25445=>"11111110",
  25446=>"11111101",
  25447=>"00000001",
  25448=>"00000001",
  25449=>"11111111",
  25450=>"00000001",
  25451=>"00000001",
  25452=>"11111111",
  25453=>"00000000",
  25454=>"00000001",
  25455=>"11111110",
  25456=>"00000000",
  25457=>"00000101",
  25458=>"00000000",
  25459=>"11111111",
  25460=>"11111111",
  25461=>"00000000",
  25462=>"11111110",
  25463=>"11111101",
  25464=>"00000000",
  25465=>"11111110",
  25466=>"00000010",
  25467=>"00000010",
  25468=>"00000001",
  25469=>"00000000",
  25470=>"11111101",
  25471=>"11111100",
  25472=>"11111111",
  25473=>"00000010",
  25474=>"11111111",
  25475=>"00000011",
  25476=>"00000010",
  25477=>"00000000",
  25478=>"11111111",
  25479=>"00000010",
  25480=>"00000010",
  25481=>"11111101",
  25482=>"11111111",
  25483=>"00000101",
  25484=>"00000000",
  25485=>"11111110",
  25486=>"11111101",
  25487=>"00000011",
  25488=>"11111110",
  25489=>"00000000",
  25490=>"11111111",
  25491=>"11111111",
  25492=>"11111111",
  25493=>"00000010",
  25494=>"11111111",
  25495=>"00000001",
  25496=>"00000001",
  25497=>"11111111",
  25498=>"00000001",
  25499=>"00000100",
  25500=>"11111101",
  25501=>"11111111",
  25502=>"00000011",
  25503=>"00000000",
  25504=>"11111101",
  25505=>"11111110",
  25506=>"11111111",
  25507=>"11111111",
  25508=>"11111111",
  25509=>"00000000",
  25510=>"11111110",
  25511=>"11111101",
  25512=>"00000001",
  25513=>"00000000",
  25514=>"11111101",
  25515=>"11111110",
  25516=>"00000010",
  25517=>"11111101",
  25518=>"11111110",
  25519=>"00000000",
  25520=>"00000000",
  25521=>"11111111",
  25522=>"11111011",
  25523=>"11111101",
  25524=>"11111110",
  25525=>"00000010",
  25526=>"00000000",
  25527=>"00000001",
  25528=>"00000010",
  25529=>"00000010",
  25530=>"00000000",
  25531=>"00000001",
  25532=>"00000000",
  25533=>"00000001",
  25534=>"00000000",
  25535=>"00000010",
  25536=>"00000011",
  25537=>"00000001",
  25538=>"11111110",
  25539=>"11111101",
  25540=>"11111110",
  25541=>"11111110",
  25542=>"11111110",
  25543=>"00000010",
  25544=>"00000101",
  25545=>"11111110",
  25546=>"11111100",
  25547=>"11111111",
  25548=>"11111110",
  25549=>"11111101",
  25550=>"00000101",
  25551=>"11111110",
  25552=>"00000001",
  25553=>"00000001",
  25554=>"11111101",
  25555=>"00000001",
  25556=>"11111111",
  25557=>"00000010",
  25558=>"00000000",
  25559=>"00000000",
  25560=>"00000010",
  25561=>"11111111",
  25562=>"11111101",
  25563=>"11111110",
  25564=>"11111101",
  25565=>"11111110",
  25566=>"11111110",
  25567=>"00000001",
  25568=>"00000001",
  25569=>"11111110",
  25570=>"00000010",
  25571=>"11111101",
  25572=>"00000000",
  25573=>"11111110",
  25574=>"00000001",
  25575=>"11111110",
  25576=>"11111110",
  25577=>"00000001",
  25578=>"11111110",
  25579=>"00000010",
  25580=>"11111101",
  25581=>"00000001",
  25582=>"00000010",
  25583=>"00000001",
  25584=>"11111101",
  25585=>"00000001",
  25586=>"11111110",
  25587=>"00000010",
  25588=>"00000001",
  25589=>"11111110",
  25590=>"00000010",
  25591=>"00000001",
  25592=>"11111111",
  25593=>"11111101",
  25594=>"11111100",
  25595=>"00000000",
  25596=>"00000010",
  25597=>"11111101",
  25598=>"11111110",
  25599=>"11111111",
  25600=>"00000000",
  25601=>"00000000",
  25602=>"11111111",
  25603=>"00000010",
  25604=>"11111110",
  25605=>"11111101",
  25606=>"00000010",
  25607=>"00000100",
  25608=>"11111100",
  25609=>"11111101",
  25610=>"00000000",
  25611=>"11111110",
  25612=>"11111111",
  25613=>"11111111",
  25614=>"00000110",
  25615=>"00000010",
  25616=>"11111110",
  25617=>"11111110",
  25618=>"11111110",
  25619=>"00000010",
  25620=>"00000000",
  25621=>"00000000",
  25622=>"00000001",
  25623=>"00000000",
  25624=>"00000001",
  25625=>"00000010",
  25626=>"00000000",
  25627=>"00000100",
  25628=>"00000001",
  25629=>"00000011",
  25630=>"11111111",
  25631=>"11111101",
  25632=>"11111101",
  25633=>"11111111",
  25634=>"00000100",
  25635=>"00000011",
  25636=>"00000011",
  25637=>"00000010",
  25638=>"11111111",
  25639=>"11111101",
  25640=>"00000011",
  25641=>"00000011",
  25642=>"11111110",
  25643=>"00000000",
  25644=>"11111111",
  25645=>"11111111",
  25646=>"11111111",
  25647=>"11111110",
  25648=>"00000001",
  25649=>"00000010",
  25650=>"11111110",
  25651=>"11111110",
  25652=>"00000000",
  25653=>"00000010",
  25654=>"00000010",
  25655=>"00000010",
  25656=>"00000000",
  25657=>"11111101",
  25658=>"00000100",
  25659=>"11111110",
  25660=>"00000001",
  25661=>"11111111",
  25662=>"11111110",
  25663=>"00000010",
  25664=>"00000001",
  25665=>"11111101",
  25666=>"00000000",
  25667=>"00000001",
  25668=>"00000101",
  25669=>"00000011",
  25670=>"00000101",
  25671=>"00000001",
  25672=>"00000001",
  25673=>"00000010",
  25674=>"00000010",
  25675=>"00000001",
  25676=>"11111101",
  25677=>"00000010",
  25678=>"11111110",
  25679=>"00000010",
  25680=>"00000001",
  25681=>"11111110",
  25682=>"00000101",
  25683=>"11111111",
  25684=>"00000010",
  25685=>"00000000",
  25686=>"11111101",
  25687=>"00000000",
  25688=>"00000100",
  25689=>"11111100",
  25690=>"11111111",
  25691=>"00000000",
  25692=>"11111111",
  25693=>"11111111",
  25694=>"00000000",
  25695=>"11111111",
  25696=>"00000001",
  25697=>"00000010",
  25698=>"00000110",
  25699=>"00000000",
  25700=>"00000011",
  25701=>"00000000",
  25702=>"11111111",
  25703=>"00000000",
  25704=>"00000010",
  25705=>"00000001",
  25706=>"11111111",
  25707=>"00000000",
  25708=>"00000010",
  25709=>"11111110",
  25710=>"00000010",
  25711=>"11111110",
  25712=>"11111110",
  25713=>"11111111",
  25714=>"00000010",
  25715=>"11111110",
  25716=>"11111101",
  25717=>"11111111",
  25718=>"11111111",
  25719=>"00000001",
  25720=>"11111111",
  25721=>"00000000",
  25722=>"11111110",
  25723=>"11111111",
  25724=>"11111101",
  25725=>"00000001",
  25726=>"00000010",
  25727=>"00000010",
  25728=>"00000001",
  25729=>"00000000",
  25730=>"11111110",
  25731=>"00000010",
  25732=>"11111100",
  25733=>"00000001",
  25734=>"00000011",
  25735=>"11111110",
  25736=>"11111100",
  25737=>"11111101",
  25738=>"00000011",
  25739=>"00000000",
  25740=>"11111110",
  25741=>"00000001",
  25742=>"11111101",
  25743=>"00000100",
  25744=>"00000000",
  25745=>"00000011",
  25746=>"11111110",
  25747=>"00000000",
  25748=>"11111011",
  25749=>"11111111",
  25750=>"00000001",
  25751=>"11111110",
  25752=>"11111111",
  25753=>"11111101",
  25754=>"00000010",
  25755=>"00000010",
  25756=>"11111110",
  25757=>"00000000",
  25758=>"00000000",
  25759=>"00000101",
  25760=>"11111111",
  25761=>"00000010",
  25762=>"00000000",
  25763=>"11111110",
  25764=>"00000000",
  25765=>"11111111",
  25766=>"00000100",
  25767=>"00000010",
  25768=>"00000000",
  25769=>"00000000",
  25770=>"00000001",
  25771=>"00000011",
  25772=>"11111110",
  25773=>"00000010",
  25774=>"00000000",
  25775=>"00000001",
  25776=>"00000100",
  25777=>"00000001",
  25778=>"00000001",
  25779=>"00000010",
  25780=>"11111110",
  25781=>"11111110",
  25782=>"11111100",
  25783=>"00000001",
  25784=>"11111101",
  25785=>"00000100",
  25786=>"11111101",
  25787=>"00000001",
  25788=>"11111111",
  25789=>"00000010",
  25790=>"11111111",
  25791=>"00000100",
  25792=>"00000001",
  25793=>"00000010",
  25794=>"11111110",
  25795=>"11111110",
  25796=>"11111110",
  25797=>"00000011",
  25798=>"11111110",
  25799=>"00000001",
  25800=>"00000000",
  25801=>"11111111",
  25802=>"00000000",
  25803=>"00000010",
  25804=>"00000001",
  25805=>"11111110",
  25806=>"00000001",
  25807=>"00000010",
  25808=>"00000000",
  25809=>"11111111",
  25810=>"11111111",
  25811=>"00000010",
  25812=>"00000001",
  25813=>"11111110",
  25814=>"11111111",
  25815=>"11111101",
  25816=>"00000000",
  25817=>"00000001",
  25818=>"00000000",
  25819=>"11111101",
  25820=>"11111111",
  25821=>"00000101",
  25822=>"00000010",
  25823=>"11111111",
  25824=>"00000000",
  25825=>"11111100",
  25826=>"11111110",
  25827=>"00000010",
  25828=>"11111101",
  25829=>"11111110",
  25830=>"11111111",
  25831=>"00000010",
  25832=>"00000010",
  25833=>"00000011",
  25834=>"11111111",
  25835=>"00000001",
  25836=>"11111101",
  25837=>"11111101",
  25838=>"11111101",
  25839=>"00000001",
  25840=>"00000001",
  25841=>"11111110",
  25842=>"00000001",
  25843=>"11111111",
  25844=>"00000010",
  25845=>"00000001",
  25846=>"11111110",
  25847=>"11111111",
  25848=>"11111110",
  25849=>"00000010",
  25850=>"11111110",
  25851=>"00000001",
  25852=>"00000000",
  25853=>"00000000",
  25854=>"00000000",
  25855=>"11111111",
  25856=>"00000001",
  25857=>"00000100",
  25858=>"11111110",
  25859=>"00000100",
  25860=>"11111110",
  25861=>"00000000",
  25862=>"00000000",
  25863=>"11111110",
  25864=>"11111111",
  25865=>"11111110",
  25866=>"11111111",
  25867=>"00000000",
  25868=>"11111111",
  25869=>"00000001",
  25870=>"11111111",
  25871=>"00000001",
  25872=>"00000111",
  25873=>"00000011",
  25874=>"00000001",
  25875=>"00000010",
  25876=>"00000011",
  25877=>"00000101",
  25878=>"00000000",
  25879=>"00000011",
  25880=>"00000100",
  25881=>"00000010",
  25882=>"11111111",
  25883=>"00000000",
  25884=>"11111100",
  25885=>"11111101",
  25886=>"00000100",
  25887=>"11111110",
  25888=>"00000011",
  25889=>"00000110",
  25890=>"11111111",
  25891=>"11111100",
  25892=>"00000000",
  25893=>"00000001",
  25894=>"11111101",
  25895=>"00000001",
  25896=>"00000001",
  25897=>"00000000",
  25898=>"00000001",
  25899=>"11111100",
  25900=>"00000000",
  25901=>"00000010",
  25902=>"00000010",
  25903=>"00000000",
  25904=>"00000001",
  25905=>"00000001",
  25906=>"11111110",
  25907=>"11111110",
  25908=>"11111111",
  25909=>"00000000",
  25910=>"00000010",
  25911=>"11111111",
  25912=>"00000011",
  25913=>"00000000",
  25914=>"00000001",
  25915=>"00000010",
  25916=>"00000011",
  25917=>"00000000",
  25918=>"00000000",
  25919=>"00000000",
  25920=>"00000001",
  25921=>"11111101",
  25922=>"00000000",
  25923=>"11111110",
  25924=>"11111110",
  25925=>"00000001",
  25926=>"11111101",
  25927=>"11111101",
  25928=>"11111110",
  25929=>"00000001",
  25930=>"11111110",
  25931=>"00000001",
  25932=>"00000011",
  25933=>"00000001",
  25934=>"11111101",
  25935=>"00000010",
  25936=>"11111111",
  25937=>"11111101",
  25938=>"00000000",
  25939=>"00000100",
  25940=>"00000000",
  25941=>"00000000",
  25942=>"11111110",
  25943=>"11111110",
  25944=>"00000100",
  25945=>"11111100",
  25946=>"00000000",
  25947=>"00000011",
  25948=>"00000001",
  25949=>"11111101",
  25950=>"00000010",
  25951=>"11111111",
  25952=>"11111110",
  25953=>"00000010",
  25954=>"00000001",
  25955=>"11111110",
  25956=>"11111110",
  25957=>"00000011",
  25958=>"11111100",
  25959=>"00000001",
  25960=>"00000010",
  25961=>"11111110",
  25962=>"00000000",
  25963=>"00000001",
  25964=>"11111101",
  25965=>"11111101",
  25966=>"11111101",
  25967=>"00000010",
  25968=>"00000000",
  25969=>"00000101",
  25970=>"00000000",
  25971=>"00000011",
  25972=>"11111110",
  25973=>"00000011",
  25974=>"11111111",
  25975=>"11111111",
  25976=>"00000100",
  25977=>"00000001",
  25978=>"00000010",
  25979=>"00000000",
  25980=>"00000101",
  25981=>"00000000",
  25982=>"00000001",
  25983=>"11111100",
  25984=>"11111111",
  25985=>"11111110",
  25986=>"11111110",
  25987=>"11111111",
  25988=>"11111110",
  25989=>"11111111",
  25990=>"00000011",
  25991=>"11111111",
  25992=>"00000010",
  25993=>"11111100",
  25994=>"00000000",
  25995=>"00000010",
  25996=>"11111111",
  25997=>"00000011",
  25998=>"00000000",
  25999=>"00000100",
  26000=>"00000001",
  26001=>"11111110",
  26002=>"00000001",
  26003=>"00000010",
  26004=>"00000010",
  26005=>"00000101",
  26006=>"11111101",
  26007=>"00000001",
  26008=>"00000011",
  26009=>"00000000",
  26010=>"11111111",
  26011=>"11111111",
  26012=>"00000001",
  26013=>"00000110",
  26014=>"00000010",
  26015=>"00000000",
  26016=>"00000000",
  26017=>"00000011",
  26018=>"00000011",
  26019=>"11111111",
  26020=>"11111111",
  26021=>"00000000",
  26022=>"00000000",
  26023=>"00000100",
  26024=>"00000000",
  26025=>"11111111",
  26026=>"00000010",
  26027=>"00000110",
  26028=>"11111101",
  26029=>"11111110",
  26030=>"00000001",
  26031=>"00000011",
  26032=>"00000010",
  26033=>"11111110",
  26034=>"00000000",
  26035=>"00000000",
  26036=>"00000001",
  26037=>"00000010",
  26038=>"11111110",
  26039=>"11111111",
  26040=>"11111110",
  26041=>"00000000",
  26042=>"00000001",
  26043=>"00000100",
  26044=>"11111111",
  26045=>"11111110",
  26046=>"11111110",
  26047=>"00000000",
  26048=>"11111110",
  26049=>"11111111",
  26050=>"11111100",
  26051=>"11111110",
  26052=>"11111100",
  26053=>"00000001",
  26054=>"11111110",
  26055=>"00000001",
  26056=>"00000100",
  26057=>"11111111",
  26058=>"11111111",
  26059=>"11111100",
  26060=>"00000011",
  26061=>"00000001",
  26062=>"00000000",
  26063=>"11111101",
  26064=>"00000001",
  26065=>"11111111",
  26066=>"00000010",
  26067=>"00000010",
  26068=>"11111101",
  26069=>"00000011",
  26070=>"00000010",
  26071=>"11111111",
  26072=>"11111111",
  26073=>"00000011",
  26074=>"00000000",
  26075=>"00000000",
  26076=>"00000101",
  26077=>"00000011",
  26078=>"11111101",
  26079=>"00000001",
  26080=>"00000001",
  26081=>"00000000",
  26082=>"11111111",
  26083=>"11111110",
  26084=>"00000011",
  26085=>"00000001",
  26086=>"11111110",
  26087=>"00000010",
  26088=>"00000100",
  26089=>"00000010",
  26090=>"00000001",
  26091=>"00000001",
  26092=>"11111101",
  26093=>"00000010",
  26094=>"00000010",
  26095=>"11111111",
  26096=>"11111111",
  26097=>"00000011",
  26098=>"00000001",
  26099=>"11111101",
  26100=>"00000010",
  26101=>"00000001",
  26102=>"00000010",
  26103=>"00000001",
  26104=>"00000001",
  26105=>"00000010",
  26106=>"00000000",
  26107=>"11111111",
  26108=>"00000011",
  26109=>"11111111",
  26110=>"00000010",
  26111=>"11111101",
  26112=>"00000010",
  26113=>"11111110",
  26114=>"11111111",
  26115=>"00000000",
  26116=>"11111101",
  26117=>"00000001",
  26118=>"11111111",
  26119=>"11111101",
  26120=>"11111110",
  26121=>"11111111",
  26122=>"00000010",
  26123=>"11111110",
  26124=>"11111101",
  26125=>"00000001",
  26126=>"00000111",
  26127=>"11111110",
  26128=>"11111110",
  26129=>"11111101",
  26130=>"11111111",
  26131=>"11111101",
  26132=>"00000011",
  26133=>"11111110",
  26134=>"00000100",
  26135=>"00000000",
  26136=>"11111101",
  26137=>"11111111",
  26138=>"11111101",
  26139=>"00000011",
  26140=>"00000011",
  26141=>"00000100",
  26142=>"11111101",
  26143=>"00000011",
  26144=>"11111101",
  26145=>"11111111",
  26146=>"11111111",
  26147=>"11111111",
  26148=>"00000011",
  26149=>"00000000",
  26150=>"00000000",
  26151=>"11111101",
  26152=>"00000011",
  26153=>"11111110",
  26154=>"00000000",
  26155=>"00000000",
  26156=>"00000100",
  26157=>"11111101",
  26158=>"11111101",
  26159=>"11111111",
  26160=>"00000010",
  26161=>"00000000",
  26162=>"11111111",
  26163=>"00000010",
  26164=>"00000011",
  26165=>"11111110",
  26166=>"11111110",
  26167=>"00000010",
  26168=>"00000001",
  26169=>"00000000",
  26170=>"00000001",
  26171=>"00000000",
  26172=>"00000000",
  26173=>"00000100",
  26174=>"11111110",
  26175=>"00000011",
  26176=>"11111101",
  26177=>"00000001",
  26178=>"11111110",
  26179=>"11111110",
  26180=>"11111110",
  26181=>"00000001",
  26182=>"11111111",
  26183=>"00000011",
  26184=>"00000010",
  26185=>"00000000",
  26186=>"00000101",
  26187=>"00000000",
  26188=>"00000010",
  26189=>"11111101",
  26190=>"11111101",
  26191=>"11111111",
  26192=>"00000010",
  26193=>"00000010",
  26194=>"11111101",
  26195=>"00000000",
  26196=>"00000000",
  26197=>"00000001",
  26198=>"11111110",
  26199=>"11111110",
  26200=>"00000100",
  26201=>"00000011",
  26202=>"00000011",
  26203=>"11111111",
  26204=>"00000000",
  26205=>"11111101",
  26206=>"11111111",
  26207=>"00000011",
  26208=>"00000001",
  26209=>"00000000",
  26210=>"11111101",
  26211=>"00000001",
  26212=>"11111101",
  26213=>"11111111",
  26214=>"00000010",
  26215=>"00000110",
  26216=>"00000001",
  26217=>"00000000",
  26218=>"00000010",
  26219=>"00000001",
  26220=>"00000000",
  26221=>"00000010",
  26222=>"00000100",
  26223=>"11111110",
  26224=>"11111101",
  26225=>"00000001",
  26226=>"00000011",
  26227=>"00000011",
  26228=>"11111110",
  26229=>"11111101",
  26230=>"00000010",
  26231=>"11111110",
  26232=>"11111101",
  26233=>"00000000",
  26234=>"00000000",
  26235=>"00000011",
  26236=>"00000001",
  26237=>"00000101",
  26238=>"00000000",
  26239=>"11111110",
  26240=>"11111111",
  26241=>"00000010",
  26242=>"00000100",
  26243=>"00000100",
  26244=>"00000010",
  26245=>"11111111",
  26246=>"11111110",
  26247=>"00000001",
  26248=>"11111101",
  26249=>"11111110",
  26250=>"11111111",
  26251=>"00000100",
  26252=>"00000011",
  26253=>"11111101",
  26254=>"11111111",
  26255=>"00000010",
  26256=>"00000011",
  26257=>"11111110",
  26258=>"11111111",
  26259=>"11111110",
  26260=>"11111111",
  26261=>"00000000",
  26262=>"11111101",
  26263=>"11111110",
  26264=>"00000010",
  26265=>"00000011",
  26266=>"11111101",
  26267=>"11111111",
  26268=>"00000001",
  26269=>"00000011",
  26270=>"00000001",
  26271=>"11111111",
  26272=>"11111111",
  26273=>"11111111",
  26274=>"00000001",
  26275=>"11111110",
  26276=>"11111110",
  26277=>"11111110",
  26278=>"00000011",
  26279=>"11111111",
  26280=>"11111110",
  26281=>"11111110",
  26282=>"11111110",
  26283=>"00000000",
  26284=>"11111110",
  26285=>"00000000",
  26286=>"11111111",
  26287=>"11111100",
  26288=>"00000011",
  26289=>"00000000",
  26290=>"11111110",
  26291=>"00000100",
  26292=>"00000011",
  26293=>"11111100",
  26294=>"11111111",
  26295=>"00000011",
  26296=>"11111101",
  26297=>"00000000",
  26298=>"11111111",
  26299=>"00000001",
  26300=>"11111101",
  26301=>"00000100",
  26302=>"11111110",
  26303=>"00000001",
  26304=>"00000001",
  26305=>"00000010",
  26306=>"00000001",
  26307=>"00000000",
  26308=>"11111111",
  26309=>"11111111",
  26310=>"00000001",
  26311=>"00000001",
  26312=>"00000011",
  26313=>"00000101",
  26314=>"00000010",
  26315=>"11111101",
  26316=>"11111111",
  26317=>"11111110",
  26318=>"11111110",
  26319=>"11111110",
  26320=>"00000010",
  26321=>"11111101",
  26322=>"00000001",
  26323=>"00000011",
  26324=>"11111111",
  26325=>"11111110",
  26326=>"00000001",
  26327=>"11111111",
  26328=>"00000000",
  26329=>"00000011",
  26330=>"00000000",
  26331=>"11111100",
  26332=>"00000001",
  26333=>"00000001",
  26334=>"11111110",
  26335=>"11111100",
  26336=>"00000001",
  26337=>"11111101",
  26338=>"00000000",
  26339=>"00000000",
  26340=>"00000011",
  26341=>"11111110",
  26342=>"00000011",
  26343=>"00000010",
  26344=>"00000000",
  26345=>"00000001",
  26346=>"00000000",
  26347=>"00000001",
  26348=>"00000010",
  26349=>"00000001",
  26350=>"00000011",
  26351=>"11111110",
  26352=>"00000011",
  26353=>"00000010",
  26354=>"11111111",
  26355=>"11111101",
  26356=>"00000000",
  26357=>"00000011",
  26358=>"00000010",
  26359=>"11111110",
  26360=>"00000011",
  26361=>"11111101",
  26362=>"11111110",
  26363=>"00000000",
  26364=>"00000001",
  26365=>"00000000",
  26366=>"00000001",
  26367=>"00000011",
  26368=>"00000010",
  26369=>"11111101",
  26370=>"00000000",
  26371=>"00000000",
  26372=>"11111111",
  26373=>"00000000",
  26374=>"11111110",
  26375=>"00000101",
  26376=>"11111101",
  26377=>"00000010",
  26378=>"00000000",
  26379=>"00000111",
  26380=>"11111101",
  26381=>"00000000",
  26382=>"00000010",
  26383=>"00000010",
  26384=>"00000010",
  26385=>"11111100",
  26386=>"11111100",
  26387=>"00000010",
  26388=>"11111101",
  26389=>"00000001",
  26390=>"00001000",
  26391=>"00000010",
  26392=>"00000000",
  26393=>"11111101",
  26394=>"11111110",
  26395=>"00000000",
  26396=>"00000010",
  26397=>"00000001",
  26398=>"00000000",
  26399=>"00000001",
  26400=>"00000100",
  26401=>"00000000",
  26402=>"11111111",
  26403=>"11111111",
  26404=>"11111101",
  26405=>"11111100",
  26406=>"11111110",
  26407=>"00000010",
  26408=>"00000011",
  26409=>"00000101",
  26410=>"00000000",
  26411=>"11111101",
  26412=>"11111110",
  26413=>"00000010",
  26414=>"00000100",
  26415=>"00000000",
  26416=>"00000010",
  26417=>"11111110",
  26418=>"11111111",
  26419=>"00000101",
  26420=>"00000001",
  26421=>"11111111",
  26422=>"00000011",
  26423=>"00000000",
  26424=>"00000000",
  26425=>"11111101",
  26426=>"00000010",
  26427=>"00000000",
  26428=>"00000001",
  26429=>"11111101",
  26430=>"11111110",
  26431=>"00000011",
  26432=>"00000001",
  26433=>"00000000",
  26434=>"11111101",
  26435=>"11111101",
  26436=>"00000100",
  26437=>"11111111",
  26438=>"00000011",
  26439=>"00000000",
  26440=>"11111100",
  26441=>"00000010",
  26442=>"00000000",
  26443=>"11111101",
  26444=>"00000001",
  26445=>"00000000",
  26446=>"11111101",
  26447=>"00000001",
  26448=>"00000000",
  26449=>"00000000",
  26450=>"11111111",
  26451=>"11111111",
  26452=>"00000100",
  26453=>"11111110",
  26454=>"00000001",
  26455=>"00000000",
  26456=>"00000000",
  26457=>"11111111",
  26458=>"00000010",
  26459=>"11111101",
  26460=>"00000001",
  26461=>"00000011",
  26462=>"00000100",
  26463=>"00000000",
  26464=>"11111100",
  26465=>"00000001",
  26466=>"00000001",
  26467=>"00000010",
  26468=>"11111100",
  26469=>"00000011",
  26470=>"11111110",
  26471=>"11111101",
  26472=>"11111110",
  26473=>"00000010",
  26474=>"00000000",
  26475=>"00000011",
  26476=>"11111110",
  26477=>"11111101",
  26478=>"00000000",
  26479=>"00000011",
  26480=>"11111101",
  26481=>"11111101",
  26482=>"00000010",
  26483=>"00000010",
  26484=>"00000000",
  26485=>"11111110",
  26486=>"11111110",
  26487=>"00000011",
  26488=>"00000011",
  26489=>"11111101",
  26490=>"11111110",
  26491=>"00000000",
  26492=>"00000000",
  26493=>"00000010",
  26494=>"00000001",
  26495=>"00000101",
  26496=>"00000011",
  26497=>"00000001",
  26498=>"00000010",
  26499=>"00000011",
  26500=>"00000010",
  26501=>"11111101",
  26502=>"11111101",
  26503=>"00000000",
  26504=>"00000011",
  26505=>"00000000",
  26506=>"11111111",
  26507=>"00000100",
  26508=>"11111101",
  26509=>"00000011",
  26510=>"00000001",
  26511=>"11111110",
  26512=>"11111110",
  26513=>"00000011",
  26514=>"00000100",
  26515=>"00000001",
  26516=>"00000010",
  26517=>"11111111",
  26518=>"11111111",
  26519=>"00000000",
  26520=>"11111110",
  26521=>"11111111",
  26522=>"00000110",
  26523=>"11111100",
  26524=>"00000001",
  26525=>"00000001",
  26526=>"11111011",
  26527=>"00000001",
  26528=>"00001000",
  26529=>"00000010",
  26530=>"11111111",
  26531=>"00000011",
  26532=>"00000011",
  26533=>"11111101",
  26534=>"11111110",
  26535=>"00000001",
  26536=>"00000010",
  26537=>"00000001",
  26538=>"00000010",
  26539=>"00000011",
  26540=>"00000010",
  26541=>"11111110",
  26542=>"00000011",
  26543=>"00000010",
  26544=>"00000000",
  26545=>"00000110",
  26546=>"11111101",
  26547=>"11111111",
  26548=>"00000000",
  26549=>"00000100",
  26550=>"00000100",
  26551=>"11111110",
  26552=>"11111100",
  26553=>"00000010",
  26554=>"00000011",
  26555=>"00000001",
  26556=>"00000000",
  26557=>"11111111",
  26558=>"00000011",
  26559=>"00000001",
  26560=>"00000000",
  26561=>"11111110",
  26562=>"00000001",
  26563=>"11111111",
  26564=>"00000001",
  26565=>"00000011",
  26566=>"11111100",
  26567=>"00000000",
  26568=>"00000001",
  26569=>"00000011",
  26570=>"11111111",
  26571=>"11111111",
  26572=>"00000011",
  26573=>"00000000",
  26574=>"11111110",
  26575=>"00000010",
  26576=>"00000000",
  26577=>"11111111",
  26578=>"00000011",
  26579=>"00000001",
  26580=>"11111110",
  26581=>"00000000",
  26582=>"00000010",
  26583=>"11111100",
  26584=>"00000001",
  26585=>"11111111",
  26586=>"00000110",
  26587=>"11111101",
  26588=>"11111110",
  26589=>"00000100",
  26590=>"00000101",
  26591=>"11111111",
  26592=>"11111101",
  26593=>"11111110",
  26594=>"00000010",
  26595=>"00000010",
  26596=>"11111111",
  26597=>"00000010",
  26598=>"11111100",
  26599=>"11111011",
  26600=>"00000010",
  26601=>"00000011",
  26602=>"00000001",
  26603=>"00000000",
  26604=>"00000101",
  26605=>"00000010",
  26606=>"11111101",
  26607=>"00000100",
  26608=>"11111101",
  26609=>"00000010",
  26610=>"11111110",
  26611=>"11111110",
  26612=>"00000001",
  26613=>"11111101",
  26614=>"11111101",
  26615=>"11111111",
  26616=>"00000010",
  26617=>"11111110",
  26618=>"11111101",
  26619=>"00000010",
  26620=>"11111101",
  26621=>"00000011",
  26622=>"00000000",
  26623=>"11111101",
  26624=>"11111110",
  26625=>"11111111",
  26626=>"00000010",
  26627=>"00000000",
  26628=>"11111101",
  26629=>"00000001",
  26630=>"00000001",
  26631=>"00000011",
  26632=>"11111110",
  26633=>"00000010",
  26634=>"11111111",
  26635=>"00000010",
  26636=>"00000000",
  26637=>"11111111",
  26638=>"00000010",
  26639=>"00000010",
  26640=>"11111110",
  26641=>"11111111",
  26642=>"00000001",
  26643=>"00000001",
  26644=>"00000001",
  26645=>"11111101",
  26646=>"00000010",
  26647=>"00000001",
  26648=>"11111111",
  26649=>"11111101",
  26650=>"00000000",
  26651=>"00000000",
  26652=>"00000101",
  26653=>"11111101",
  26654=>"00000000",
  26655=>"11111110",
  26656=>"11111111",
  26657=>"11111110",
  26658=>"00000101",
  26659=>"11111111",
  26660=>"11111110",
  26661=>"11111110",
  26662=>"11111111",
  26663=>"11111111",
  26664=>"11111111",
  26665=>"00000010",
  26666=>"11111110",
  26667=>"00000001",
  26668=>"00000000",
  26669=>"11111111",
  26670=>"00000000",
  26671=>"00000000",
  26672=>"00000001",
  26673=>"00000000",
  26674=>"11111111",
  26675=>"00000000",
  26676=>"11111111",
  26677=>"11111101",
  26678=>"11111111",
  26679=>"00000010",
  26680=>"11111110",
  26681=>"00000011",
  26682=>"11111110",
  26683=>"11111101",
  26684=>"11111110",
  26685=>"00000010",
  26686=>"11111111",
  26687=>"00000000",
  26688=>"11111111",
  26689=>"11111110",
  26690=>"11111101",
  26691=>"11111111",
  26692=>"11111111",
  26693=>"00000000",
  26694=>"00000001",
  26695=>"00000001",
  26696=>"00000000",
  26697=>"11111110",
  26698=>"00000000",
  26699=>"00000001",
  26700=>"11111111",
  26701=>"11111110",
  26702=>"00000000",
  26703=>"11111111",
  26704=>"00000010",
  26705=>"00000001",
  26706=>"00000011",
  26707=>"00000010",
  26708=>"00000001",
  26709=>"11111111",
  26710=>"00000011",
  26711=>"11111101",
  26712=>"11111101",
  26713=>"11111101",
  26714=>"11111111",
  26715=>"11111101",
  26716=>"11111101",
  26717=>"00000001",
  26718=>"00000010",
  26719=>"11111110",
  26720=>"00000010",
  26721=>"00000001",
  26722=>"00000000",
  26723=>"11111110",
  26724=>"11111111",
  26725=>"00000000",
  26726=>"00000100",
  26727=>"00000001",
  26728=>"00000010",
  26729=>"11111111",
  26730=>"00000011",
  26731=>"11111111",
  26732=>"00000000",
  26733=>"11111101",
  26734=>"11111111",
  26735=>"11111111",
  26736=>"00000100",
  26737=>"11111110",
  26738=>"11111111",
  26739=>"00000001",
  26740=>"11111110",
  26741=>"11111101",
  26742=>"00000101",
  26743=>"11111110",
  26744=>"11111100",
  26745=>"11111100",
  26746=>"11111110",
  26747=>"00000000",
  26748=>"00000011",
  26749=>"00000011",
  26750=>"00000000",
  26751=>"00000000",
  26752=>"00000010",
  26753=>"11111111",
  26754=>"00000000",
  26755=>"11111110",
  26756=>"00000010",
  26757=>"00000000",
  26758=>"11111101",
  26759=>"00000000",
  26760=>"11111101",
  26761=>"00000010",
  26762=>"00000010",
  26763=>"00000001",
  26764=>"11111101",
  26765=>"11111111",
  26766=>"11111111",
  26767=>"00000010",
  26768=>"00000000",
  26769=>"11111110",
  26770=>"00000001",
  26771=>"00000010",
  26772=>"00000001",
  26773=>"11111111",
  26774=>"11111111",
  26775=>"00000001",
  26776=>"11111110",
  26777=>"00000010",
  26778=>"00000000",
  26779=>"11111101",
  26780=>"00000000",
  26781=>"00000001",
  26782=>"00000000",
  26783=>"11111110",
  26784=>"11111111",
  26785=>"11111100",
  26786=>"11111110",
  26787=>"11111110",
  26788=>"00000000",
  26789=>"11111111",
  26790=>"11111101",
  26791=>"00000000",
  26792=>"11111110",
  26793=>"00000011",
  26794=>"00000001",
  26795=>"11111111",
  26796=>"00000001",
  26797=>"00000001",
  26798=>"11111101",
  26799=>"11111110",
  26800=>"11111101",
  26801=>"00000001",
  26802=>"00000010",
  26803=>"00000000",
  26804=>"11111110",
  26805=>"11111110",
  26806=>"11111111",
  26807=>"00000001",
  26808=>"00000011",
  26809=>"00000000",
  26810=>"00000100",
  26811=>"11111110",
  26812=>"00000000",
  26813=>"11111111",
  26814=>"11111111",
  26815=>"00000001",
  26816=>"11111111",
  26817=>"00000001",
  26818=>"11111101",
  26819=>"00000011",
  26820=>"11111111",
  26821=>"11111101",
  26822=>"00000000",
  26823=>"00000000",
  26824=>"11111101",
  26825=>"11111111",
  26826=>"00000001",
  26827=>"00000000",
  26828=>"00000001",
  26829=>"11111110",
  26830=>"00000000",
  26831=>"11111101",
  26832=>"00000010",
  26833=>"00000011",
  26834=>"00000001",
  26835=>"11111111",
  26836=>"00000000",
  26837=>"11111110",
  26838=>"00000011",
  26839=>"11111111",
  26840=>"00000010",
  26841=>"00000000",
  26842=>"11111111",
  26843=>"11111111",
  26844=>"00000010",
  26845=>"00000100",
  26846=>"00000000",
  26847=>"11111110",
  26848=>"00000010",
  26849=>"11111110",
  26850=>"11111110",
  26851=>"11111101",
  26852=>"11111110",
  26853=>"00000010",
  26854=>"00000001",
  26855=>"11111110",
  26856=>"11111101",
  26857=>"11111111",
  26858=>"00000001",
  26859=>"00000010",
  26860=>"00000001",
  26861=>"11111110",
  26862=>"11111101",
  26863=>"00000001",
  26864=>"00000001",
  26865=>"00000110",
  26866=>"00000001",
  26867=>"11111101",
  26868=>"00000010",
  26869=>"00000010",
  26870=>"11111111",
  26871=>"00000001",
  26872=>"00000010",
  26873=>"00000000",
  26874=>"00000110",
  26875=>"00000000",
  26876=>"11111111",
  26877=>"11111101",
  26878=>"00000001",
  26879=>"11111110",
  26880=>"11111110",
  26881=>"00000011",
  26882=>"00000010",
  26883=>"11111111",
  26884=>"00000010",
  26885=>"11111110",
  26886=>"00000001",
  26887=>"00000001",
  26888=>"00000001",
  26889=>"11111111",
  26890=>"00000100",
  26891=>"00000000",
  26892=>"00000000",
  26893=>"00000011",
  26894=>"11111101",
  26895=>"11111111",
  26896=>"00000010",
  26897=>"00000001",
  26898=>"11111110",
  26899=>"00000010",
  26900=>"00000000",
  26901=>"00000001",
  26902=>"11111110",
  26903=>"11111101",
  26904=>"11111101",
  26905=>"11111101",
  26906=>"00000000",
  26907=>"00000000",
  26908=>"11111110",
  26909=>"11111110",
  26910=>"00000001",
  26911=>"00000000",
  26912=>"11111110",
  26913=>"11111110",
  26914=>"00000010",
  26915=>"11111110",
  26916=>"11111110",
  26917=>"11111111",
  26918=>"00000100",
  26919=>"11111100",
  26920=>"00000010",
  26921=>"00000010",
  26922=>"00000000",
  26923=>"11111111",
  26924=>"00000001",
  26925=>"00000000",
  26926=>"00000000",
  26927=>"00000011",
  26928=>"00000000",
  26929=>"00000001",
  26930=>"00000001",
  26931=>"11111101",
  26932=>"11111110",
  26933=>"11111101",
  26934=>"11111110",
  26935=>"11111111",
  26936=>"11111110",
  26937=>"00000010",
  26938=>"11111101",
  26939=>"00000000",
  26940=>"00000010",
  26941=>"00000010",
  26942=>"00000001",
  26943=>"11111110",
  26944=>"11111110",
  26945=>"00000100",
  26946=>"11111111",
  26947=>"00000000",
  26948=>"11111110",
  26949=>"11111110",
  26950=>"00000101",
  26951=>"11111110",
  26952=>"11111110",
  26953=>"11111110",
  26954=>"00000000",
  26955=>"00000011",
  26956=>"00000000",
  26957=>"11111110",
  26958=>"11111110",
  26959=>"11111110",
  26960=>"11111111",
  26961=>"11111110",
  26962=>"11111111",
  26963=>"11111110",
  26964=>"00000000",
  26965=>"00000001",
  26966=>"00000010",
  26967=>"11111111",
  26968=>"11111110",
  26969=>"00000010",
  26970=>"00000001",
  26971=>"11111101",
  26972=>"00000001",
  26973=>"00000001",
  26974=>"00000000",
  26975=>"00000101",
  26976=>"11111110",
  26977=>"00000010",
  26978=>"11111111",
  26979=>"00000000",
  26980=>"11111110",
  26981=>"11111110",
  26982=>"00000011",
  26983=>"11111111",
  26984=>"11111110",
  26985=>"11111111",
  26986=>"11111111",
  26987=>"00000101",
  26988=>"11111111",
  26989=>"00000001",
  26990=>"11111101",
  26991=>"00000001",
  26992=>"00000010",
  26993=>"00000000",
  26994=>"00000010",
  26995=>"11111101",
  26996=>"11111110",
  26997=>"11111110",
  26998=>"00000000",
  26999=>"11111111",
  27000=>"11111110",
  27001=>"11111110",
  27002=>"00000000",
  27003=>"11111101",
  27004=>"11111101",
  27005=>"11111111",
  27006=>"00000010",
  27007=>"11111110",
  27008=>"00000100",
  27009=>"00000001",
  27010=>"00000011",
  27011=>"11111101",
  27012=>"00000000",
  27013=>"00000000",
  27014=>"11111111",
  27015=>"00000000",
  27016=>"00000010",
  27017=>"00000001",
  27018=>"00000101",
  27019=>"00000000",
  27020=>"00000000",
  27021=>"00000010",
  27022=>"11111101",
  27023=>"11111110",
  27024=>"00000000",
  27025=>"00000010",
  27026=>"00000000",
  27027=>"00000001",
  27028=>"11111111",
  27029=>"11111101",
  27030=>"11111110",
  27031=>"00000011",
  27032=>"11111110",
  27033=>"00000100",
  27034=>"11111100",
  27035=>"11111111",
  27036=>"00000011",
  27037=>"00000101",
  27038=>"00000001",
  27039=>"00001000",
  27040=>"11111111",
  27041=>"00000000",
  27042=>"00000101",
  27043=>"00000000",
  27044=>"00000000",
  27045=>"11111110",
  27046=>"00000001",
  27047=>"11111110",
  27048=>"11111101",
  27049=>"11111111",
  27050=>"00000001",
  27051=>"11111111",
  27052=>"11111110",
  27053=>"00000001",
  27054=>"00000001",
  27055=>"00000001",
  27056=>"00000000",
  27057=>"11111110",
  27058=>"11111110",
  27059=>"11111111",
  27060=>"11111111",
  27061=>"11111110",
  27062=>"00000000",
  27063=>"00000001",
  27064=>"11111101",
  27065=>"00000000",
  27066=>"11111110",
  27067=>"00000001",
  27068=>"00000000",
  27069=>"00000101",
  27070=>"00000011",
  27071=>"00000010",
  27072=>"11111111",
  27073=>"00000000",
  27074=>"00000000",
  27075=>"00000010",
  27076=>"00000001",
  27077=>"11111100",
  27078=>"11111110",
  27079=>"00000100",
  27080=>"11111101",
  27081=>"00000010",
  27082=>"11111111",
  27083=>"11111111",
  27084=>"00000010",
  27085=>"11111110",
  27086=>"00000010",
  27087=>"00000000",
  27088=>"11111111",
  27089=>"11111110",
  27090=>"11111100",
  27091=>"00000011",
  27092=>"00000000",
  27093=>"00000000",
  27094=>"11111111",
  27095=>"00000000",
  27096=>"00000001",
  27097=>"11111110",
  27098=>"11111111",
  27099=>"11111110",
  27100=>"11111110",
  27101=>"00000010",
  27102=>"11111101",
  27103=>"00000000",
  27104=>"11111111",
  27105=>"00000001",
  27106=>"00000001",
  27107=>"11111110",
  27108=>"00000000",
  27109=>"00000010",
  27110=>"11111101",
  27111=>"00000011",
  27112=>"00000000",
  27113=>"11111110",
  27114=>"00000000",
  27115=>"00000000",
  27116=>"00000001",
  27117=>"11111110",
  27118=>"11111110",
  27119=>"00000011",
  27120=>"00000000",
  27121=>"11111101",
  27122=>"11111111",
  27123=>"11111110",
  27124=>"00000010",
  27125=>"00000001",
  27126=>"00000000",
  27127=>"11111111",
  27128=>"11111100",
  27129=>"00000011",
  27130=>"00000001",
  27131=>"11111110",
  27132=>"00000010",
  27133=>"00000101",
  27134=>"11111101",
  27135=>"00000000",
  27136=>"00000000",
  27137=>"00000010",
  27138=>"11111111",
  27139=>"11111111",
  27140=>"00000001",
  27141=>"00000000",
  27142=>"11111110",
  27143=>"00000001",
  27144=>"00000100",
  27145=>"00000001",
  27146=>"11111111",
  27147=>"11111111",
  27148=>"00000001",
  27149=>"00000000",
  27150=>"11111111",
  27151=>"00000000",
  27152=>"00000000",
  27153=>"00000011",
  27154=>"11111111",
  27155=>"11111110",
  27156=>"11111110",
  27157=>"11111101",
  27158=>"00000010",
  27159=>"00000000",
  27160=>"11111100",
  27161=>"00000111",
  27162=>"00000010",
  27163=>"00000010",
  27164=>"00000001",
  27165=>"00000000",
  27166=>"11111111",
  27167=>"11111111",
  27168=>"11111111",
  27169=>"00000010",
  27170=>"00000001",
  27171=>"11111110",
  27172=>"00000000",
  27173=>"00000001",
  27174=>"11111101",
  27175=>"00000000",
  27176=>"11111111",
  27177=>"11111110",
  27178=>"00000101",
  27179=>"11111111",
  27180=>"00000001",
  27181=>"11111110",
  27182=>"00000000",
  27183=>"00000000",
  27184=>"00000001",
  27185=>"11111101",
  27186=>"11111101",
  27187=>"11111111",
  27188=>"11111110",
  27189=>"00000001",
  27190=>"00000000",
  27191=>"11111101",
  27192=>"00000000",
  27193=>"11111111",
  27194=>"11111101",
  27195=>"11111111",
  27196=>"00000101",
  27197=>"11111101",
  27198=>"00000001",
  27199=>"00000000",
  27200=>"11111110",
  27201=>"00000000",
  27202=>"00000001",
  27203=>"00000010",
  27204=>"11111101",
  27205=>"00000010",
  27206=>"11111111",
  27207=>"00000000",
  27208=>"11111110",
  27209=>"11111111",
  27210=>"00000000",
  27211=>"11111110",
  27212=>"00000001",
  27213=>"11111111",
  27214=>"00000001",
  27215=>"00000000",
  27216=>"11111111",
  27217=>"00000000",
  27218=>"00000011",
  27219=>"00000000",
  27220=>"00000001",
  27221=>"00000000",
  27222=>"00000000",
  27223=>"11111111",
  27224=>"00000001",
  27225=>"11111111",
  27226=>"00000001",
  27227=>"00000011",
  27228=>"00000101",
  27229=>"00000000",
  27230=>"11111110",
  27231=>"11111101",
  27232=>"00000001",
  27233=>"11111110",
  27234=>"00000001",
  27235=>"00000010",
  27236=>"00000011",
  27237=>"00000000",
  27238=>"11111111",
  27239=>"11111101",
  27240=>"00000101",
  27241=>"11111111",
  27242=>"11111111",
  27243=>"11111111",
  27244=>"00000000",
  27245=>"11111101",
  27246=>"00000001",
  27247=>"00000010",
  27248=>"00000001",
  27249=>"00000010",
  27250=>"11111111",
  27251=>"00000000",
  27252=>"11111110",
  27253=>"00000011",
  27254=>"00000010",
  27255=>"11111100",
  27256=>"00000000",
  27257=>"00000010",
  27258=>"00000001",
  27259=>"11111101",
  27260=>"11111110",
  27261=>"00000010",
  27262=>"11111110",
  27263=>"11111110",
  27264=>"11111110",
  27265=>"11111111",
  27266=>"11111101",
  27267=>"11111101",
  27268=>"00000001",
  27269=>"00000000",
  27270=>"11111110",
  27271=>"11111111",
  27272=>"00000010",
  27273=>"00000001",
  27274=>"00000001",
  27275=>"00000000",
  27276=>"00000001",
  27277=>"00000000",
  27278=>"11111111",
  27279=>"00000011",
  27280=>"11111110",
  27281=>"00000010",
  27282=>"11111101",
  27283=>"00000000",
  27284=>"00000011",
  27285=>"11111101",
  27286=>"00000001",
  27287=>"11111110",
  27288=>"00000011",
  27289=>"11111110",
  27290=>"00000000",
  27291=>"11111110",
  27292=>"11111110",
  27293=>"00000010",
  27294=>"11111111",
  27295=>"11111110",
  27296=>"11111111",
  27297=>"00000010",
  27298=>"11111110",
  27299=>"11111101",
  27300=>"11111110",
  27301=>"00000000",
  27302=>"11111110",
  27303=>"11111100",
  27304=>"11111110",
  27305=>"11111101",
  27306=>"00000001",
  27307=>"00000010",
  27308=>"00000001",
  27309=>"11111110",
  27310=>"00000001",
  27311=>"00000011",
  27312=>"11111100",
  27313=>"00000100",
  27314=>"00000000",
  27315=>"00000001",
  27316=>"00000010",
  27317=>"11111101",
  27318=>"11111101",
  27319=>"00000101",
  27320=>"11111111",
  27321=>"00000000",
  27322=>"11111110",
  27323=>"00000001",
  27324=>"00000000",
  27325=>"11111111",
  27326=>"11111111",
  27327=>"00000001",
  27328=>"11111110",
  27329=>"11111111",
  27330=>"00000100",
  27331=>"00000000",
  27332=>"00000011",
  27333=>"11111111",
  27334=>"00000000",
  27335=>"11111110",
  27336=>"00000000",
  27337=>"11111110",
  27338=>"11111101",
  27339=>"11111110",
  27340=>"11111110",
  27341=>"00000100",
  27342=>"11111110",
  27343=>"11111111",
  27344=>"11111111",
  27345=>"00000001",
  27346=>"11111110",
  27347=>"11111111",
  27348=>"00000001",
  27349=>"11111110",
  27350=>"11111111",
  27351=>"11111111",
  27352=>"00000001",
  27353=>"11111111",
  27354=>"00000010",
  27355=>"11111110",
  27356=>"11111101",
  27357=>"00000010",
  27358=>"11111111",
  27359=>"11111111",
  27360=>"11111111",
  27361=>"11111101",
  27362=>"00000011",
  27363=>"11111110",
  27364=>"00000000",
  27365=>"00000000",
  27366=>"11111110",
  27367=>"00000001",
  27368=>"00000001",
  27369=>"11111111",
  27370=>"11111101",
  27371=>"11111110",
  27372=>"11111101",
  27373=>"11111111",
  27374=>"00000000",
  27375=>"00000010",
  27376=>"11111110",
  27377=>"00000100",
  27378=>"11111101",
  27379=>"00000011",
  27380=>"00000101",
  27381=>"00000000",
  27382=>"11111101",
  27383=>"00000011",
  27384=>"00000001",
  27385=>"00000011",
  27386=>"11111110",
  27387=>"11111100",
  27388=>"00000001",
  27389=>"00000000",
  27390=>"00000001",
  27391=>"11111101",
  27392=>"11111111",
  27393=>"11111111",
  27394=>"11111110",
  27395=>"00000011",
  27396=>"00000010",
  27397=>"00000000",
  27398=>"00000001",
  27399=>"00000000",
  27400=>"11111100",
  27401=>"11111101",
  27402=>"00000010",
  27403=>"00000000",
  27404=>"00000001",
  27405=>"11111111",
  27406=>"00000001",
  27407=>"00000001",
  27408=>"11111101",
  27409=>"00000010",
  27410=>"00000000",
  27411=>"11111101",
  27412=>"11111110",
  27413=>"00000000",
  27414=>"00000010",
  27415=>"00000010",
  27416=>"00000000",
  27417=>"00000101",
  27418=>"11111101",
  27419=>"00000000",
  27420=>"11111111",
  27421=>"00000100",
  27422=>"11111111",
  27423=>"00000001",
  27424=>"00000011",
  27425=>"00000000",
  27426=>"00000001",
  27427=>"00000001",
  27428=>"11111110",
  27429=>"11111111",
  27430=>"00000001",
  27431=>"11111110",
  27432=>"00000000",
  27433=>"11111101",
  27434=>"00000000",
  27435=>"00000010",
  27436=>"00000001",
  27437=>"11111110",
  27438=>"11111111",
  27439=>"00000001",
  27440=>"00000011",
  27441=>"11111101",
  27442=>"00000110",
  27443=>"11111101",
  27444=>"00000001",
  27445=>"00000001",
  27446=>"11111110",
  27447=>"11111110",
  27448=>"00000001",
  27449=>"11111110",
  27450=>"00000000",
  27451=>"00000000",
  27452=>"00000000",
  27453=>"11111111",
  27454=>"11111111",
  27455=>"00000001",
  27456=>"00000001",
  27457=>"11111101",
  27458=>"11111111",
  27459=>"11111110",
  27460=>"00000000",
  27461=>"00000010",
  27462=>"11111110",
  27463=>"11111101",
  27464=>"11111110",
  27465=>"00000001",
  27466=>"11111111",
  27467=>"00000110",
  27468=>"11111101",
  27469=>"00000000",
  27470=>"00000000",
  27471=>"00000010",
  27472=>"00000010",
  27473=>"00000001",
  27474=>"11111101",
  27475=>"11111111",
  27476=>"00000010",
  27477=>"11111110",
  27478=>"00000010",
  27479=>"11111110",
  27480=>"11111101",
  27481=>"00000000",
  27482=>"11111101",
  27483=>"00000101",
  27484=>"00000001",
  27485=>"00000010",
  27486=>"11111111",
  27487=>"00000000",
  27488=>"00000001",
  27489=>"00000001",
  27490=>"00000000",
  27491=>"11111111",
  27492=>"11111111",
  27493=>"11111101",
  27494=>"00000001",
  27495=>"00000000",
  27496=>"00000011",
  27497=>"00000000",
  27498=>"11111111",
  27499=>"00000001",
  27500=>"11111111",
  27501=>"00000100",
  27502=>"00000011",
  27503=>"11111110",
  27504=>"11111110",
  27505=>"00000000",
  27506=>"00000000",
  27507=>"11111110",
  27508=>"11111101",
  27509=>"11111111",
  27510=>"00000001",
  27511=>"11111110",
  27512=>"00000010",
  27513=>"00000010",
  27514=>"11111110",
  27515=>"11111111",
  27516=>"00000011",
  27517=>"11111111",
  27518=>"11111111",
  27519=>"11111111",
  27520=>"11111110",
  27521=>"00000000",
  27522=>"00000001",
  27523=>"11111111",
  27524=>"00000001",
  27525=>"00000000",
  27526=>"00000011",
  27527=>"00000010",
  27528=>"11111101",
  27529=>"11111110",
  27530=>"00000000",
  27531=>"00000001",
  27532=>"11111110",
  27533=>"11111111",
  27534=>"00000100",
  27535=>"11111111",
  27536=>"11111111",
  27537=>"11111111",
  27538=>"00000010",
  27539=>"11111111",
  27540=>"00000001",
  27541=>"11111110",
  27542=>"00000000",
  27543=>"00000001",
  27544=>"11111101",
  27545=>"00000001",
  27546=>"11111101",
  27547=>"00000100",
  27548=>"11111110",
  27549=>"11111110",
  27550=>"11111111",
  27551=>"11111111",
  27552=>"00000001",
  27553=>"11111110",
  27554=>"00000010",
  27555=>"00000001",
  27556=>"00000001",
  27557=>"00000010",
  27558=>"11111101",
  27559=>"00000011",
  27560=>"11111111",
  27561=>"00000001",
  27562=>"00000000",
  27563=>"11111111",
  27564=>"11111101",
  27565=>"00000001",
  27566=>"00000001",
  27567=>"11111111",
  27568=>"00000000",
  27569=>"11111110",
  27570=>"00000011",
  27571=>"11111111",
  27572=>"11111111",
  27573=>"00000000",
  27574=>"00000010",
  27575=>"00000000",
  27576=>"11111101",
  27577=>"11111101",
  27578=>"00000000",
  27579=>"11111111",
  27580=>"11111110",
  27581=>"00000001",
  27582=>"00000001",
  27583=>"11111110",
  27584=>"11111111",
  27585=>"00000000",
  27586=>"00000001",
  27587=>"00000010",
  27588=>"00000001",
  27589=>"11111101",
  27590=>"00000001",
  27591=>"00000001",
  27592=>"00000001",
  27593=>"11111111",
  27594=>"11111101",
  27595=>"11111101",
  27596=>"00000001",
  27597=>"00000000",
  27598=>"00000001",
  27599=>"11111111",
  27600=>"11111100",
  27601=>"11111110",
  27602=>"00000010",
  27603=>"00000000",
  27604=>"00000000",
  27605=>"00000001",
  27606=>"11111111",
  27607=>"00000001",
  27608=>"00000010",
  27609=>"00000001",
  27610=>"00000001",
  27611=>"11111101",
  27612=>"00000001",
  27613=>"00000000",
  27614=>"11111110",
  27615=>"00000010",
  27616=>"11111110",
  27617=>"11111101",
  27618=>"00000000",
  27619=>"00000011",
  27620=>"11111110",
  27621=>"11111110",
  27622=>"00000101",
  27623=>"11111101",
  27624=>"00000000",
  27625=>"00000001",
  27626=>"11111110",
  27627=>"11111101",
  27628=>"00000000",
  27629=>"00000001",
  27630=>"00000001",
  27631=>"00000100",
  27632=>"00000001",
  27633=>"00000001",
  27634=>"11111110",
  27635=>"11111111",
  27636=>"11111110",
  27637=>"00000001",
  27638=>"11111101",
  27639=>"11111100",
  27640=>"11111111",
  27641=>"00000010",
  27642=>"11111110",
  27643=>"11111110",
  27644=>"11111110",
  27645=>"11111110",
  27646=>"11111101",
  27647=>"00000010",
  27648=>"11111110",
  27649=>"00000011",
  27650=>"00000011",
  27651=>"00000000",
  27652=>"00000010",
  27653=>"00000001",
  27654=>"00000000",
  27655=>"00000010",
  27656=>"00000000",
  27657=>"00000010",
  27658=>"00000001",
  27659=>"11111110",
  27660=>"00000001",
  27661=>"11111110",
  27662=>"00000011",
  27663=>"00000000",
  27664=>"00000001",
  27665=>"11111100",
  27666=>"11111101",
  27667=>"11111101",
  27668=>"00000000",
  27669=>"11111101",
  27670=>"11111101",
  27671=>"11111110",
  27672=>"11111111",
  27673=>"11111111",
  27674=>"00000001",
  27675=>"00000000",
  27676=>"00000001",
  27677=>"00000001",
  27678=>"00000010",
  27679=>"11111110",
  27680=>"11111101",
  27681=>"00000000",
  27682=>"00000010",
  27683=>"00000010",
  27684=>"11111111",
  27685=>"11111110",
  27686=>"00000000",
  27687=>"00000010",
  27688=>"11111110",
  27689=>"11111101",
  27690=>"00000010",
  27691=>"00000100",
  27692=>"00000001",
  27693=>"00000001",
  27694=>"00000000",
  27695=>"11111111",
  27696=>"00000011",
  27697=>"00000000",
  27698=>"11111111",
  27699=>"00000001",
  27700=>"00000001",
  27701=>"11111111",
  27702=>"00000000",
  27703=>"00000000",
  27704=>"00000011",
  27705=>"00000100",
  27706=>"11111110",
  27707=>"00000011",
  27708=>"00000001",
  27709=>"00000010",
  27710=>"00000001",
  27711=>"11111111",
  27712=>"11111110",
  27713=>"11111111",
  27714=>"11111110",
  27715=>"00000000",
  27716=>"00000001",
  27717=>"00000001",
  27718=>"11111101",
  27719=>"00000001",
  27720=>"00000011",
  27721=>"11111101",
  27722=>"00000011",
  27723=>"00000000",
  27724=>"00000001",
  27725=>"00000100",
  27726=>"00000001",
  27727=>"00000000",
  27728=>"11111111",
  27729=>"11111111",
  27730=>"11111100",
  27731=>"00000111",
  27732=>"00000001",
  27733=>"00000000",
  27734=>"00000011",
  27735=>"00000001",
  27736=>"00000000",
  27737=>"00000010",
  27738=>"00000000",
  27739=>"11111110",
  27740=>"00000010",
  27741=>"00000011",
  27742=>"00000000",
  27743=>"00000110",
  27744=>"11111110",
  27745=>"00000001",
  27746=>"11111101",
  27747=>"11111101",
  27748=>"00000000",
  27749=>"11111110",
  27750=>"00000011",
  27751=>"11111111",
  27752=>"00000001",
  27753=>"00000001",
  27754=>"00000001",
  27755=>"11111110",
  27756=>"00000000",
  27757=>"00000000",
  27758=>"00000001",
  27759=>"00000001",
  27760=>"00000001",
  27761=>"00000010",
  27762=>"00000101",
  27763=>"00000000",
  27764=>"11111111",
  27765=>"00000001",
  27766=>"11111110",
  27767=>"11111101",
  27768=>"11111111",
  27769=>"00000000",
  27770=>"11111110",
  27771=>"11111101",
  27772=>"00000000",
  27773=>"11111111",
  27774=>"00000011",
  27775=>"00000001",
  27776=>"11111101",
  27777=>"11111110",
  27778=>"00000010",
  27779=>"00000011",
  27780=>"11111111",
  27781=>"00000100",
  27782=>"11111111",
  27783=>"00000101",
  27784=>"11111111",
  27785=>"00000010",
  27786=>"11111100",
  27787=>"00000100",
  27788=>"00000000",
  27789=>"00000011",
  27790=>"00000001",
  27791=>"11111111",
  27792=>"11111111",
  27793=>"00000001",
  27794=>"00000001",
  27795=>"00000011",
  27796=>"11111110",
  27797=>"00000011",
  27798=>"00000100",
  27799=>"00000011",
  27800=>"00000000",
  27801=>"11111100",
  27802=>"00000000",
  27803=>"11111110",
  27804=>"00000000",
  27805=>"00000001",
  27806=>"00000011",
  27807=>"00000011",
  27808=>"00000000",
  27809=>"00000110",
  27810=>"00000010",
  27811=>"11111100",
  27812=>"00000001",
  27813=>"00000100",
  27814=>"00000000",
  27815=>"11111101",
  27816=>"00000100",
  27817=>"11111101",
  27818=>"00000010",
  27819=>"11111110",
  27820=>"00000011",
  27821=>"00000000",
  27822=>"11111111",
  27823=>"11111111",
  27824=>"11111110",
  27825=>"11111110",
  27826=>"00000001",
  27827=>"00000000",
  27828=>"11111101",
  27829=>"11111111",
  27830=>"00000010",
  27831=>"00000010",
  27832=>"11111111",
  27833=>"11111111",
  27834=>"00000000",
  27835=>"11111100",
  27836=>"00000010",
  27837=>"00000001",
  27838=>"11111110",
  27839=>"11111101",
  27840=>"00000000",
  27841=>"00000100",
  27842=>"00000000",
  27843=>"11111110",
  27844=>"00000010",
  27845=>"11111110",
  27846=>"11111110",
  27847=>"00000010",
  27848=>"00000001",
  27849=>"11111100",
  27850=>"00000000",
  27851=>"11111110",
  27852=>"00000010",
  27853=>"11111101",
  27854=>"00000010",
  27855=>"00000100",
  27856=>"11111100",
  27857=>"11111110",
  27858=>"11111111",
  27859=>"11111110",
  27860=>"00000001",
  27861=>"00000100",
  27862=>"00000100",
  27863=>"11111110",
  27864=>"11111110",
  27865=>"00000010",
  27866=>"11111110",
  27867=>"11111101",
  27868=>"11111110",
  27869=>"11111110",
  27870=>"11111111",
  27871=>"00000011",
  27872=>"11111101",
  27873=>"00000001",
  27874=>"00000000",
  27875=>"00000011",
  27876=>"11111110",
  27877=>"00000101",
  27878=>"11111110",
  27879=>"00000001",
  27880=>"00000010",
  27881=>"11111100",
  27882=>"00000011",
  27883=>"00000000",
  27884=>"11111111",
  27885=>"00000011",
  27886=>"11111111",
  27887=>"00000000",
  27888=>"00000111",
  27889=>"11111110",
  27890=>"00000010",
  27891=>"11111111",
  27892=>"11111111",
  27893=>"00000010",
  27894=>"00000010",
  27895=>"00000000",
  27896=>"11111110",
  27897=>"00000010",
  27898=>"00000001",
  27899=>"11111110",
  27900=>"11111100",
  27901=>"11111111",
  27902=>"00000001",
  27903=>"00000000",
  27904=>"00000100",
  27905=>"00000000",
  27906=>"11111101",
  27907=>"11111111",
  27908=>"11111110",
  27909=>"00000000",
  27910=>"00000010",
  27911=>"00000001",
  27912=>"00000001",
  27913=>"00000000",
  27914=>"11111110",
  27915=>"00000100",
  27916=>"11111110",
  27917=>"00000001",
  27918=>"11111111",
  27919=>"00000100",
  27920=>"00000010",
  27921=>"11111110",
  27922=>"00000000",
  27923=>"11111110",
  27924=>"00000101",
  27925=>"11111100",
  27926=>"00000011",
  27927=>"00000011",
  27928=>"00000010",
  27929=>"00000001",
  27930=>"11111101",
  27931=>"00000010",
  27932=>"00000101",
  27933=>"00000010",
  27934=>"11111101",
  27935=>"00000001",
  27936=>"11111110",
  27937=>"11111110",
  27938=>"00000100",
  27939=>"11111110",
  27940=>"00000100",
  27941=>"11111111",
  27942=>"11111011",
  27943=>"00000001",
  27944=>"00000010",
  27945=>"11111110",
  27946=>"11111111",
  27947=>"11111100",
  27948=>"00000011",
  27949=>"00000010",
  27950=>"11111101",
  27951=>"00000000",
  27952=>"00000010",
  27953=>"00000000",
  27954=>"00000011",
  27955=>"00000010",
  27956=>"00000001",
  27957=>"00000010",
  27958=>"00000010",
  27959=>"11111111",
  27960=>"00000000",
  27961=>"00000001",
  27962=>"11111111",
  27963=>"11111110",
  27964=>"11111111",
  27965=>"00000001",
  27966=>"11111101",
  27967=>"00000001",
  27968=>"00000010",
  27969=>"11111101",
  27970=>"00000001",
  27971=>"00000010",
  27972=>"00000001",
  27973=>"00000010",
  27974=>"00000000",
  27975=>"00000000",
  27976=>"11111101",
  27977=>"00000000",
  27978=>"00000011",
  27979=>"00000010",
  27980=>"00000001",
  27981=>"00000001",
  27982=>"11111111",
  27983=>"00000000",
  27984=>"11111110",
  27985=>"11111110",
  27986=>"11111101",
  27987=>"00000001",
  27988=>"00000100",
  27989=>"11111111",
  27990=>"11111110",
  27991=>"11111111",
  27992=>"11111111",
  27993=>"11111111",
  27994=>"00000001",
  27995=>"00000001",
  27996=>"11111101",
  27997=>"00000001",
  27998=>"11111111",
  27999=>"00000010",
  28000=>"00000010",
  28001=>"11111100",
  28002=>"00000000",
  28003=>"00000001",
  28004=>"00000011",
  28005=>"00000010",
  28006=>"00000100",
  28007=>"00000010",
  28008=>"00000000",
  28009=>"00000001",
  28010=>"00000000",
  28011=>"00000001",
  28012=>"11111110",
  28013=>"11111101",
  28014=>"11111111",
  28015=>"00000000",
  28016=>"11111111",
  28017=>"11111111",
  28018=>"11111111",
  28019=>"11111111",
  28020=>"00000100",
  28021=>"00000001",
  28022=>"00000001",
  28023=>"11111110",
  28024=>"00000011",
  28025=>"11111110",
  28026=>"11111100",
  28027=>"00000100",
  28028=>"11111110",
  28029=>"11111110",
  28030=>"00000001",
  28031=>"00000011",
  28032=>"11111111",
  28033=>"11111101",
  28034=>"11111111",
  28035=>"11111111",
  28036=>"00000010",
  28037=>"11111110",
  28038=>"00000101",
  28039=>"11111110",
  28040=>"00000010",
  28041=>"00000000",
  28042=>"11111101",
  28043=>"00000011",
  28044=>"00000000",
  28045=>"11111110",
  28046=>"11111111",
  28047=>"00000011",
  28048=>"00000000",
  28049=>"00000000",
  28050=>"11111110",
  28051=>"11111111",
  28052=>"00000010",
  28053=>"00000100",
  28054=>"00000000",
  28055=>"00000000",
  28056=>"00000000",
  28057=>"11111111",
  28058=>"00000001",
  28059=>"11111111",
  28060=>"00000010",
  28061=>"11111110",
  28062=>"11111110",
  28063=>"11111101",
  28064=>"00000000",
  28065=>"00000000",
  28066=>"11111110",
  28067=>"00000001",
  28068=>"00000001",
  28069=>"11111101",
  28070=>"00000001",
  28071=>"11111111",
  28072=>"00000010",
  28073=>"00000000",
  28074=>"11111111",
  28075=>"00000001",
  28076=>"00000001",
  28077=>"00000001",
  28078=>"11111110",
  28079=>"11111110",
  28080=>"11111101",
  28081=>"11111111",
  28082=>"00000010",
  28083=>"11111101",
  28084=>"00000000",
  28085=>"00000010",
  28086=>"00000010",
  28087=>"00000000",
  28088=>"11111110",
  28089=>"11111110",
  28090=>"00000010",
  28091=>"11111110",
  28092=>"00000001",
  28093=>"00000011",
  28094=>"11111111",
  28095=>"11111110",
  28096=>"11111111",
  28097=>"00000011",
  28098=>"00000000",
  28099=>"11111111",
  28100=>"00000110",
  28101=>"11111110",
  28102=>"00000100",
  28103=>"00000010",
  28104=>"00000000",
  28105=>"11111111",
  28106=>"11111101",
  28107=>"00000001",
  28108=>"11111101",
  28109=>"11111111",
  28110=>"00000011",
  28111=>"11111111",
  28112=>"00000000",
  28113=>"11111110",
  28114=>"11111111",
  28115=>"00000111",
  28116=>"11111110",
  28117=>"11111110",
  28118=>"00000000",
  28119=>"00000001",
  28120=>"11111111",
  28121=>"00000000",
  28122=>"00000001",
  28123=>"11111100",
  28124=>"11111101",
  28125=>"11111110",
  28126=>"11111110",
  28127=>"00000011",
  28128=>"00000101",
  28129=>"00000011",
  28130=>"11111101",
  28131=>"00000010",
  28132=>"00000011",
  28133=>"00000011",
  28134=>"00000000",
  28135=>"00000000",
  28136=>"11111100",
  28137=>"11111111",
  28138=>"11111110",
  28139=>"11111110",
  28140=>"00000000",
  28141=>"11111100",
  28142=>"00000010",
  28143=>"00000000",
  28144=>"00000001",
  28145=>"11111101",
  28146=>"11111111",
  28147=>"00000000",
  28148=>"11111111",
  28149=>"00000001",
  28150=>"11111111",
  28151=>"00000001",
  28152=>"00000010",
  28153=>"11111101",
  28154=>"00000100",
  28155=>"00000011",
  28156=>"11111101",
  28157=>"11111100",
  28158=>"11111111",
  28159=>"00000001",
  28160=>"00000001",
  28161=>"00000010",
  28162=>"00000000",
  28163=>"11111111",
  28164=>"00000001",
  28165=>"00000011",
  28166=>"11111100",
  28167=>"00000011",
  28168=>"11111110",
  28169=>"11111111",
  28170=>"11111110",
  28171=>"00000011",
  28172=>"00000000",
  28173=>"00000011",
  28174=>"00000001",
  28175=>"11111101",
  28176=>"11111110",
  28177=>"11111111",
  28178=>"00000010",
  28179=>"11111111",
  28180=>"00000001",
  28181=>"11111110",
  28182=>"00000000",
  28183=>"11111111",
  28184=>"11111110",
  28185=>"11111101",
  28186=>"11111101",
  28187=>"11111101",
  28188=>"11111110",
  28189=>"00000001",
  28190=>"11111101",
  28191=>"00000000",
  28192=>"00000000",
  28193=>"00000000",
  28194=>"11111111",
  28195=>"11111101",
  28196=>"11111110",
  28197=>"11111111",
  28198=>"00000001",
  28199=>"00000001",
  28200=>"00000010",
  28201=>"11111101",
  28202=>"00000010",
  28203=>"11111111",
  28204=>"00000101",
  28205=>"00000010",
  28206=>"00000000",
  28207=>"11111110",
  28208=>"00000010",
  28209=>"11111111",
  28210=>"00000001",
  28211=>"00000011",
  28212=>"11111111",
  28213=>"00000011",
  28214=>"11111110",
  28215=>"00000000",
  28216=>"00000010",
  28217=>"11111110",
  28218=>"00000011",
  28219=>"11111110",
  28220=>"00000011",
  28221=>"00000010",
  28222=>"00000011",
  28223=>"00000000",
  28224=>"11111110",
  28225=>"11111111",
  28226=>"00000000",
  28227=>"00000000",
  28228=>"00000000",
  28229=>"11111110",
  28230=>"11111110",
  28231=>"11111101",
  28232=>"11111111",
  28233=>"00000001",
  28234=>"00000010",
  28235=>"11111110",
  28236=>"00000011",
  28237=>"11111101",
  28238=>"11111110",
  28239=>"00000001",
  28240=>"00000001",
  28241=>"00000100",
  28242=>"11111111",
  28243=>"00000010",
  28244=>"00000001",
  28245=>"00000000",
  28246=>"11111111",
  28247=>"00000001",
  28248=>"00000100",
  28249=>"11111101",
  28250=>"00000001",
  28251=>"00000010",
  28252=>"00000001",
  28253=>"00000010",
  28254=>"11111111",
  28255=>"11111101",
  28256=>"00000011",
  28257=>"00000000",
  28258=>"00000000",
  28259=>"11111111",
  28260=>"00000011",
  28261=>"00000010",
  28262=>"00000001",
  28263=>"11111101",
  28264=>"00000011",
  28265=>"11111101",
  28266=>"11111111",
  28267=>"00000000",
  28268=>"11111110",
  28269=>"00000000",
  28270=>"00000101",
  28271=>"00000000",
  28272=>"00000000",
  28273=>"11111111",
  28274=>"00000100",
  28275=>"00000011",
  28276=>"00000011",
  28277=>"00000100",
  28278=>"11111111",
  28279=>"00000100",
  28280=>"11111101",
  28281=>"11111110",
  28282=>"11111111",
  28283=>"00000010",
  28284=>"00000001",
  28285=>"00000010",
  28286=>"00000100",
  28287=>"00000000",
  28288=>"11111111",
  28289=>"00000001",
  28290=>"00000011",
  28291=>"11111100",
  28292=>"11111111",
  28293=>"11111110",
  28294=>"11111110",
  28295=>"11111101",
  28296=>"00000100",
  28297=>"00000000",
  28298=>"00000000",
  28299=>"00000100",
  28300=>"11111110",
  28301=>"00000001",
  28302=>"00000001",
  28303=>"11111111",
  28304=>"00000101",
  28305=>"11111111",
  28306=>"00000001",
  28307=>"00000011",
  28308=>"11111101",
  28309=>"00000101",
  28310=>"00000001",
  28311=>"11111101",
  28312=>"11111101",
  28313=>"11111101",
  28314=>"11111110",
  28315=>"00000010",
  28316=>"00000010",
  28317=>"11111110",
  28318=>"11111101",
  28319=>"11111110",
  28320=>"00000001",
  28321=>"11111101",
  28322=>"11111110",
  28323=>"11111101",
  28324=>"00000001",
  28325=>"11111110",
  28326=>"11111110",
  28327=>"11111111",
  28328=>"00000100",
  28329=>"00000011",
  28330=>"11111111",
  28331=>"11111101",
  28332=>"11111110",
  28333=>"00000010",
  28334=>"00000001",
  28335=>"11111110",
  28336=>"11111110",
  28337=>"11111100",
  28338=>"11111101",
  28339=>"00000000",
  28340=>"11111101",
  28341=>"00000000",
  28342=>"00000010",
  28343=>"11111101",
  28344=>"00000011",
  28345=>"00000010",
  28346=>"00000100",
  28347=>"00000000",
  28348=>"00000110",
  28349=>"11111111",
  28350=>"00000100",
  28351=>"00000001",
  28352=>"00000000",
  28353=>"11111101",
  28354=>"00000001",
  28355=>"11111101",
  28356=>"00000001",
  28357=>"00000010",
  28358=>"11111111",
  28359=>"00000011",
  28360=>"00000010",
  28361=>"00000001",
  28362=>"11111111",
  28363=>"00001010",
  28364=>"11111111",
  28365=>"11111100",
  28366=>"11111101",
  28367=>"00000010",
  28368=>"11111110",
  28369=>"11111101",
  28370=>"11111110",
  28371=>"11111111",
  28372=>"00000001",
  28373=>"00000101",
  28374=>"00000000",
  28375=>"00000000",
  28376=>"00000000",
  28377=>"11111111",
  28378=>"11111111",
  28379=>"00000010",
  28380=>"00000010",
  28381=>"11111111",
  28382=>"11111111",
  28383=>"11111100",
  28384=>"11111111",
  28385=>"11111110",
  28386=>"11111100",
  28387=>"00000000",
  28388=>"00000011",
  28389=>"11111111",
  28390=>"00000110",
  28391=>"00000000",
  28392=>"00000010",
  28393=>"11111111",
  28394=>"11111110",
  28395=>"11111111",
  28396=>"00000000",
  28397=>"00000000",
  28398=>"11111110",
  28399=>"00000000",
  28400=>"00000000",
  28401=>"11111111",
  28402=>"00000100",
  28403=>"11111111",
  28404=>"11111110",
  28405=>"11111101",
  28406=>"11111101",
  28407=>"11111110",
  28408=>"00000010",
  28409=>"11111110",
  28410=>"00000010",
  28411=>"11111100",
  28412=>"00000001",
  28413=>"11111101",
  28414=>"11111111",
  28415=>"00000100",
  28416=>"11111111",
  28417=>"11111111",
  28418=>"11111111",
  28419=>"11111110",
  28420=>"00000000",
  28421=>"11111111",
  28422=>"00000010",
  28423=>"00000011",
  28424=>"00000001",
  28425=>"11111101",
  28426=>"11111110",
  28427=>"11111101",
  28428=>"00000000",
  28429=>"11111110",
  28430=>"00000010",
  28431=>"11111110",
  28432=>"00000011",
  28433=>"00000000",
  28434=>"00000001",
  28435=>"11111101",
  28436=>"00000011",
  28437=>"00000010",
  28438=>"11111101",
  28439=>"00000000",
  28440=>"11111101",
  28441=>"00000011",
  28442=>"00000000",
  28443=>"00000100",
  28444=>"00000010",
  28445=>"00000010",
  28446=>"11111110",
  28447=>"11111101",
  28448=>"11111101",
  28449=>"00000001",
  28450=>"11111111",
  28451=>"00000010",
  28452=>"11111101",
  28453=>"11111110",
  28454=>"00000000",
  28455=>"00000101",
  28456=>"11111110",
  28457=>"11111111",
  28458=>"00000001",
  28459=>"11111110",
  28460=>"00000011",
  28461=>"00000000",
  28462=>"00000000",
  28463=>"00000000",
  28464=>"11111101",
  28465=>"00000100",
  28466=>"00000001",
  28467=>"00000011",
  28468=>"00000001",
  28469=>"00000010",
  28470=>"00000000",
  28471=>"00000001",
  28472=>"00000000",
  28473=>"11111101",
  28474=>"11111111",
  28475=>"11111110",
  28476=>"00000011",
  28477=>"00000010",
  28478=>"11111110",
  28479=>"00000100",
  28480=>"11111111",
  28481=>"00000100",
  28482=>"00000001",
  28483=>"00000001",
  28484=>"00000011",
  28485=>"11111101",
  28486=>"00000010",
  28487=>"00000000",
  28488=>"00000000",
  28489=>"11111101",
  28490=>"11111111",
  28491=>"00000000",
  28492=>"00000001",
  28493=>"00000001",
  28494=>"00000010",
  28495=>"00000010",
  28496=>"00000010",
  28497=>"00000000",
  28498=>"00000010",
  28499=>"00000011",
  28500=>"11111111",
  28501=>"11111101",
  28502=>"11111110",
  28503=>"11111111",
  28504=>"11111101",
  28505=>"00000000",
  28506=>"00000010",
  28507=>"11111100",
  28508=>"11111111",
  28509=>"11111101",
  28510=>"00000011",
  28511=>"00000100",
  28512=>"00000011",
  28513=>"00000000",
  28514=>"00000011",
  28515=>"00000110",
  28516=>"11111111",
  28517=>"00000100",
  28518=>"11111101",
  28519=>"11111101",
  28520=>"11111110",
  28521=>"00000000",
  28522=>"00000000",
  28523=>"00000001",
  28524=>"11111110",
  28525=>"11111111",
  28526=>"00000000",
  28527=>"00000101",
  28528=>"00000010",
  28529=>"11111110",
  28530=>"11111111",
  28531=>"11111101",
  28532=>"11111111",
  28533=>"00000000",
  28534=>"11111111",
  28535=>"00000000",
  28536=>"11111100",
  28537=>"11111111",
  28538=>"00000000",
  28539=>"11111110",
  28540=>"11111111",
  28541=>"00000000",
  28542=>"11111111",
  28543=>"00000000",
  28544=>"11111110",
  28545=>"00000111",
  28546=>"11111110",
  28547=>"00000101",
  28548=>"00000011",
  28549=>"00000001",
  28550=>"00000001",
  28551=>"11111111",
  28552=>"00000010",
  28553=>"11111101",
  28554=>"00000100",
  28555=>"11111101",
  28556=>"11111111",
  28557=>"00000000",
  28558=>"11111100",
  28559=>"11111110",
  28560=>"00000000",
  28561=>"00000000",
  28562=>"11111101",
  28563=>"00000010",
  28564=>"00000001",
  28565=>"00000011",
  28566=>"00000000",
  28567=>"00000010",
  28568=>"11111110",
  28569=>"11111101",
  28570=>"00000001",
  28571=>"00000000",
  28572=>"11111111",
  28573=>"00000001",
  28574=>"11111101",
  28575=>"00000001",
  28576=>"00000011",
  28577=>"00000000",
  28578=>"11111011",
  28579=>"00000000",
  28580=>"00000010",
  28581=>"00000001",
  28582=>"00000001",
  28583=>"00000001",
  28584=>"00000001",
  28585=>"00000000",
  28586=>"00000011",
  28587=>"11111111",
  28588=>"00000100",
  28589=>"00000011",
  28590=>"11111111",
  28591=>"00000001",
  28592=>"11111101",
  28593=>"00000101",
  28594=>"00000000",
  28595=>"11111110",
  28596=>"00000001",
  28597=>"11111100",
  28598=>"00000011",
  28599=>"00000001",
  28600=>"11111101",
  28601=>"11111111",
  28602=>"00000011",
  28603=>"00000000",
  28604=>"00000010",
  28605=>"00000010",
  28606=>"00000011",
  28607=>"11111111",
  28608=>"00000000",
  28609=>"11111101",
  28610=>"00000010",
  28611=>"00000010",
  28612=>"00000010",
  28613=>"00000000",
  28614=>"11111101",
  28615=>"00000001",
  28616=>"11111111",
  28617=>"11111110",
  28618=>"00000011",
  28619=>"11111101",
  28620=>"11111111",
  28621=>"00000000",
  28622=>"00000001",
  28623=>"11111111",
  28624=>"00000000",
  28625=>"11111110",
  28626=>"11111111",
  28627=>"11111110",
  28628=>"11111111",
  28629=>"00000001",
  28630=>"00000010",
  28631=>"11111101",
  28632=>"00000001",
  28633=>"00000001",
  28634=>"00000010",
  28635=>"00000000",
  28636=>"00000010",
  28637=>"00000100",
  28638=>"00000011",
  28639=>"11111101",
  28640=>"00000011",
  28641=>"00000010",
  28642=>"00000000",
  28643=>"11111111",
  28644=>"00000000",
  28645=>"00000001",
  28646=>"11111110",
  28647=>"00000010",
  28648=>"00000010",
  28649=>"00000000",
  28650=>"00000010",
  28651=>"00000010",
  28652=>"00000010",
  28653=>"11111101",
  28654=>"11111101",
  28655=>"11111100",
  28656=>"11111110",
  28657=>"00000010",
  28658=>"11111110",
  28659=>"00000001",
  28660=>"11111110",
  28661=>"11111100",
  28662=>"00000000",
  28663=>"00000011",
  28664=>"00000000",
  28665=>"11111111",
  28666=>"11111110",
  28667=>"11111110",
  28668=>"00000001",
  28669=>"11111101",
  28670=>"11111110",
  28671=>"00000001",
  28672=>"00000011",
  28673=>"00000000",
  28674=>"11111110",
  28675=>"11111110",
  28676=>"11111110",
  28677=>"00000000",
  28678=>"00000010",
  28679=>"11111110",
  28680=>"00000001",
  28681=>"00000000",
  28682=>"11111110",
  28683=>"11111111",
  28684=>"00000010",
  28685=>"00000010",
  28686=>"00000000",
  28687=>"00000101",
  28688=>"11111110",
  28689=>"11111110",
  28690=>"11111111",
  28691=>"11111110",
  28692=>"00000000",
  28693=>"00000010",
  28694=>"11111110",
  28695=>"11111111",
  28696=>"11111110",
  28697=>"11111111",
  28698=>"11111101",
  28699=>"11111101",
  28700=>"00000010",
  28701=>"00000000",
  28702=>"00000001",
  28703=>"11111111",
  28704=>"11111111",
  28705=>"00000001",
  28706=>"00000001",
  28707=>"00000001",
  28708=>"11111110",
  28709=>"11111111",
  28710=>"11111101",
  28711=>"00000010",
  28712=>"00000011",
  28713=>"00000000",
  28714=>"11111110",
  28715=>"00000000",
  28716=>"00000010",
  28717=>"00000000",
  28718=>"11111111",
  28719=>"00000000",
  28720=>"11111101",
  28721=>"00000001",
  28722=>"11111101",
  28723=>"00000000",
  28724=>"00000000",
  28725=>"11111111",
  28726=>"00000001",
  28727=>"00000010",
  28728=>"00000000",
  28729=>"00000111",
  28730=>"11111101",
  28731=>"11111110",
  28732=>"00000010",
  28733=>"00000001",
  28734=>"00000010",
  28735=>"00000001",
  28736=>"11111111",
  28737=>"00000100",
  28738=>"00000010",
  28739=>"00000001",
  28740=>"11111101",
  28741=>"00000000",
  28742=>"00000010",
  28743=>"11111101",
  28744=>"00000001",
  28745=>"00000000",
  28746=>"11111111",
  28747=>"11111111",
  28748=>"11111110",
  28749=>"00000010",
  28750=>"11111101",
  28751=>"11111110",
  28752=>"11111111",
  28753=>"11111110",
  28754=>"00000010",
  28755=>"11111100",
  28756=>"00000001",
  28757=>"00000010",
  28758=>"00000010",
  28759=>"11111110",
  28760=>"00000000",
  28761=>"00000100",
  28762=>"11111111",
  28763=>"00000100",
  28764=>"00000000",
  28765=>"11111111",
  28766=>"00000011",
  28767=>"11111101",
  28768=>"00000100",
  28769=>"11111110",
  28770=>"00000010",
  28771=>"11111101",
  28772=>"00000001",
  28773=>"11111111",
  28774=>"11111110",
  28775=>"00000000",
  28776=>"11111101",
  28777=>"00000000",
  28778=>"00000110",
  28779=>"11111101",
  28780=>"00000000",
  28781=>"11111101",
  28782=>"00000000",
  28783=>"00000011",
  28784=>"11111111",
  28785=>"11111100",
  28786=>"00000010",
  28787=>"11111111",
  28788=>"11111111",
  28789=>"00000001",
  28790=>"00000000",
  28791=>"00000001",
  28792=>"00000110",
  28793=>"11111111",
  28794=>"11111111",
  28795=>"11111111",
  28796=>"00000010",
  28797=>"11111110",
  28798=>"00000011",
  28799=>"11111110",
  28800=>"00000101",
  28801=>"00000001",
  28802=>"00000000",
  28803=>"00000000",
  28804=>"11111101",
  28805=>"00000011",
  28806=>"11111111",
  28807=>"11111100",
  28808=>"11111111",
  28809=>"00000000",
  28810=>"11111101",
  28811=>"00000010",
  28812=>"11111111",
  28813=>"00000000",
  28814=>"00000011",
  28815=>"00000010",
  28816=>"00000000",
  28817=>"00000011",
  28818=>"00000011",
  28819=>"11111101",
  28820=>"00000010",
  28821=>"00000010",
  28822=>"11111111",
  28823=>"11111111",
  28824=>"00000001",
  28825=>"00000001",
  28826=>"00000101",
  28827=>"11111111",
  28828=>"00000010",
  28829=>"00000001",
  28830=>"00000010",
  28831=>"11111111",
  28832=>"00000000",
  28833=>"11111111",
  28834=>"11111101",
  28835=>"00000000",
  28836=>"11111111",
  28837=>"11111100",
  28838=>"00000011",
  28839=>"00000011",
  28840=>"00000000",
  28841=>"11111111",
  28842=>"00000011",
  28843=>"00000001",
  28844=>"00000001",
  28845=>"00000001",
  28846=>"00000011",
  28847=>"00000000",
  28848=>"11111111",
  28849=>"00000010",
  28850=>"00000000",
  28851=>"11111110",
  28852=>"11111110",
  28853=>"11111111",
  28854=>"11111111",
  28855=>"11111111",
  28856=>"00000110",
  28857=>"11111111",
  28858=>"00000001",
  28859=>"00000000",
  28860=>"00000000",
  28861=>"11111111",
  28862=>"11111101",
  28863=>"00000001",
  28864=>"00000001",
  28865=>"11111111",
  28866=>"11111110",
  28867=>"11111110",
  28868=>"11111111",
  28869=>"11111110",
  28870=>"11111101",
  28871=>"00000011",
  28872=>"00000010",
  28873=>"11111111",
  28874=>"11111111",
  28875=>"00000011",
  28876=>"00000010",
  28877=>"11111101",
  28878=>"11111110",
  28879=>"00000000",
  28880=>"00000011",
  28881=>"00000000",
  28882=>"00000000",
  28883=>"11111110",
  28884=>"11111110",
  28885=>"00000100",
  28886=>"00000000",
  28887=>"00000010",
  28888=>"11111111",
  28889=>"00000001",
  28890=>"11111111",
  28891=>"11111111",
  28892=>"11111101",
  28893=>"11111111",
  28894=>"11111111",
  28895=>"11111101",
  28896=>"11111111",
  28897=>"00000100",
  28898=>"11111110",
  28899=>"00000011",
  28900=>"11111111",
  28901=>"00000000",
  28902=>"11111111",
  28903=>"11111101",
  28904=>"00000001",
  28905=>"00000110",
  28906=>"00000000",
  28907=>"00000000",
  28908=>"11111110",
  28909=>"00000000",
  28910=>"00000011",
  28911=>"00000010",
  28912=>"11111111",
  28913=>"11111101",
  28914=>"11111110",
  28915=>"11111111",
  28916=>"00000001",
  28917=>"00000110",
  28918=>"00000000",
  28919=>"00000011",
  28920=>"11111110",
  28921=>"00000000",
  28922=>"00000011",
  28923=>"00000000",
  28924=>"11111101",
  28925=>"00000100",
  28926=>"00000100",
  28927=>"00000000",
  28928=>"00000010",
  28929=>"00000100",
  28930=>"00000010",
  28931=>"11111111",
  28932=>"11111111",
  28933=>"11111111",
  28934=>"00000000",
  28935=>"00000010",
  28936=>"11111111",
  28937=>"11111100",
  28938=>"11111111",
  28939=>"11111111",
  28940=>"00000010",
  28941=>"11111110",
  28942=>"11111111",
  28943=>"11111100",
  28944=>"00000001",
  28945=>"11111111",
  28946=>"00000000",
  28947=>"00000000",
  28948=>"11111100",
  28949=>"00000000",
  28950=>"11111101",
  28951=>"11111111",
  28952=>"11111110",
  28953=>"00000000",
  28954=>"11111101",
  28955=>"11111111",
  28956=>"11111111",
  28957=>"00000001",
  28958=>"11111101",
  28959=>"00000000",
  28960=>"00000000",
  28961=>"00000000",
  28962=>"00000010",
  28963=>"00000000",
  28964=>"00000100",
  28965=>"11111111",
  28966=>"00000000",
  28967=>"11111110",
  28968=>"11111110",
  28969=>"11111100",
  28970=>"00000000",
  28971=>"11111110",
  28972=>"00000000",
  28973=>"00000010",
  28974=>"11111100",
  28975=>"11111111",
  28976=>"00000000",
  28977=>"00000010",
  28978=>"00000000",
  28979=>"00000010",
  28980=>"11111101",
  28981=>"00000001",
  28982=>"11111110",
  28983=>"11111111",
  28984=>"11111111",
  28985=>"11111110",
  28986=>"00000010",
  28987=>"00000010",
  28988=>"00000110",
  28989=>"00000010",
  28990=>"11111111",
  28991=>"11111110",
  28992=>"00000001",
  28993=>"11111111",
  28994=>"00000000",
  28995=>"00000000",
  28996=>"00000000",
  28997=>"11111111",
  28998=>"00000011",
  28999=>"00000010",
  29000=>"00000000",
  29001=>"11111110",
  29002=>"00000001",
  29003=>"00000011",
  29004=>"00000000",
  29005=>"11111101",
  29006=>"11111111",
  29007=>"00000111",
  29008=>"00000000",
  29009=>"00000010",
  29010=>"00000000",
  29011=>"00000100",
  29012=>"11111111",
  29013=>"00000100",
  29014=>"11111101",
  29015=>"00000101",
  29016=>"00000010",
  29017=>"11111110",
  29018=>"00000000",
  29019=>"00000100",
  29020=>"11111101",
  29021=>"00000010",
  29022=>"00000101",
  29023=>"00000000",
  29024=>"11111110",
  29025=>"00000100",
  29026=>"11111110",
  29027=>"00000010",
  29028=>"11111110",
  29029=>"11111110",
  29030=>"00000011",
  29031=>"00000000",
  29032=>"11111111",
  29033=>"00000000",
  29034=>"00000000",
  29035=>"00000101",
  29036=>"00000010",
  29037=>"00000001",
  29038=>"00000110",
  29039=>"11111111",
  29040=>"00000000",
  29041=>"00000001",
  29042=>"00000010",
  29043=>"11111101",
  29044=>"00000000",
  29045=>"11111100",
  29046=>"00000011",
  29047=>"11111111",
  29048=>"11111110",
  29049=>"11111110",
  29050=>"11111100",
  29051=>"11111110",
  29052=>"00000001",
  29053=>"00000100",
  29054=>"00000010",
  29055=>"00000000",
  29056=>"11111110",
  29057=>"11111111",
  29058=>"00000010",
  29059=>"00000001",
  29060=>"11111111",
  29061=>"11111110",
  29062=>"11111110",
  29063=>"00000001",
  29064=>"00000010",
  29065=>"00000001",
  29066=>"00000001",
  29067=>"11111111",
  29068=>"00000001",
  29069=>"00000000",
  29070=>"00000001",
  29071=>"11111110",
  29072=>"11111111",
  29073=>"11111111",
  29074=>"11111111",
  29075=>"00000000",
  29076=>"00000110",
  29077=>"11111110",
  29078=>"00000010",
  29079=>"00000011",
  29080=>"00000011",
  29081=>"11111100",
  29082=>"11111111",
  29083=>"11111111",
  29084=>"11111101",
  29085=>"00000001",
  29086=>"00000010",
  29087=>"11111110",
  29088=>"11111100",
  29089=>"11111110",
  29090=>"00000000",
  29091=>"11111110",
  29092=>"11111111",
  29093=>"00000010",
  29094=>"11111111",
  29095=>"11111111",
  29096=>"00000000",
  29097=>"00000011",
  29098=>"00000000",
  29099=>"11111111",
  29100=>"11111111",
  29101=>"11111110",
  29102=>"11111111",
  29103=>"00000001",
  29104=>"00000100",
  29105=>"11111101",
  29106=>"11111110",
  29107=>"00000001",
  29108=>"11111110",
  29109=>"11111101",
  29110=>"00000000",
  29111=>"11111101",
  29112=>"11111101",
  29113=>"11111110",
  29114=>"11111110",
  29115=>"11111110",
  29116=>"11111111",
  29117=>"00000001",
  29118=>"00000100",
  29119=>"11111111",
  29120=>"11111101",
  29121=>"11111111",
  29122=>"00000011",
  29123=>"00000000",
  29124=>"11111110",
  29125=>"00000001",
  29126=>"11111111",
  29127=>"00000010",
  29128=>"00000000",
  29129=>"11111101",
  29130=>"11111111",
  29131=>"00000010",
  29132=>"00000001",
  29133=>"00000001",
  29134=>"00000000",
  29135=>"11111101",
  29136=>"00000011",
  29137=>"00000001",
  29138=>"00000001",
  29139=>"11111110",
  29140=>"00000011",
  29141=>"00000011",
  29142=>"11111110",
  29143=>"11111101",
  29144=>"11111110",
  29145=>"11111111",
  29146=>"00000000",
  29147=>"11111111",
  29148=>"11111110",
  29149=>"11111110",
  29150=>"00000010",
  29151=>"11111101",
  29152=>"00000000",
  29153=>"00000000",
  29154=>"00000011",
  29155=>"00000010",
  29156=>"11111110",
  29157=>"11111111",
  29158=>"00000010",
  29159=>"00000001",
  29160=>"00000001",
  29161=>"11111101",
  29162=>"00000001",
  29163=>"00000000",
  29164=>"00000100",
  29165=>"11111101",
  29166=>"00000001",
  29167=>"00000011",
  29168=>"00000001",
  29169=>"11111110",
  29170=>"11111110",
  29171=>"00000001",
  29172=>"11111101",
  29173=>"00000000",
  29174=>"00000100",
  29175=>"11111101",
  29176=>"00000001",
  29177=>"11111100",
  29178=>"00000000",
  29179=>"00000001",
  29180=>"00000000",
  29181=>"11111111",
  29182=>"11111110",
  29183=>"11111110",
  29184=>"00000001",
  29185=>"00000001",
  29186=>"00000100",
  29187=>"00000010",
  29188=>"11111100",
  29189=>"00000000",
  29190=>"11111111",
  29191=>"11111101",
  29192=>"00000001",
  29193=>"11111101",
  29194=>"11111110",
  29195=>"00000001",
  29196=>"11111110",
  29197=>"11111101",
  29198=>"00000000",
  29199=>"00000101",
  29200=>"11111111",
  29201=>"00000000",
  29202=>"00000000",
  29203=>"00000011",
  29204=>"00000010",
  29205=>"11111110",
  29206=>"00000001",
  29207=>"11111111",
  29208=>"00000001",
  29209=>"11111110",
  29210=>"00000001",
  29211=>"00000010",
  29212=>"00000001",
  29213=>"00000000",
  29214=>"00000010",
  29215=>"00000000",
  29216=>"00000001",
  29217=>"00000010",
  29218=>"00000000",
  29219=>"00000000",
  29220=>"00000000",
  29221=>"11111101",
  29222=>"11111101",
  29223=>"11111101",
  29224=>"11111110",
  29225=>"11111110",
  29226=>"00000011",
  29227=>"11111110",
  29228=>"00000000",
  29229=>"00000000",
  29230=>"11111100",
  29231=>"00000000",
  29232=>"11111100",
  29233=>"00000001",
  29234=>"11111111",
  29235=>"00000010",
  29236=>"00000010",
  29237=>"11111101",
  29238=>"00000001",
  29239=>"11111111",
  29240=>"00000001",
  29241=>"00000011",
  29242=>"11111111",
  29243=>"11111111",
  29244=>"00000001",
  29245=>"11111111",
  29246=>"11111101",
  29247=>"11111110",
  29248=>"00000000",
  29249=>"00000001",
  29250=>"00000001",
  29251=>"00000000",
  29252=>"00000100",
  29253=>"00000010",
  29254=>"00000011",
  29255=>"00000011",
  29256=>"11111101",
  29257=>"00000010",
  29258=>"11111101",
  29259=>"11111110",
  29260=>"11111110",
  29261=>"11111110",
  29262=>"11111110",
  29263=>"11111111",
  29264=>"00000010",
  29265=>"00000001",
  29266=>"11111110",
  29267=>"00000010",
  29268=>"11111111",
  29269=>"00000001",
  29270=>"11111111",
  29271=>"11111101",
  29272=>"00000001",
  29273=>"00000000",
  29274=>"00000000",
  29275=>"11111111",
  29276=>"00000101",
  29277=>"00000000",
  29278=>"00000000",
  29279=>"00000100",
  29280=>"11111110",
  29281=>"00000000",
  29282=>"00000100",
  29283=>"11111101",
  29284=>"00000010",
  29285=>"00000010",
  29286=>"11111110",
  29287=>"11111100",
  29288=>"11111110",
  29289=>"11111110",
  29290=>"11111110",
  29291=>"00000001",
  29292=>"00000001",
  29293=>"11111111",
  29294=>"11111100",
  29295=>"00000010",
  29296=>"00000001",
  29297=>"11111111",
  29298=>"00000000",
  29299=>"11111101",
  29300=>"00000010",
  29301=>"00000001",
  29302=>"11111110",
  29303=>"00000011",
  29304=>"00000000",
  29305=>"00000001",
  29306=>"00000100",
  29307=>"11111101",
  29308=>"00000000",
  29309=>"11111111",
  29310=>"11111111",
  29311=>"00000010",
  29312=>"00000001",
  29313=>"00000010",
  29314=>"00000000",
  29315=>"00000001",
  29316=>"11111110",
  29317=>"00000011",
  29318=>"11111111",
  29319=>"11111101",
  29320=>"00000000",
  29321=>"00000011",
  29322=>"00000001",
  29323=>"11111111",
  29324=>"11111111",
  29325=>"00000010",
  29326=>"11111111",
  29327=>"00000110",
  29328=>"11111101",
  29329=>"00000110",
  29330=>"11111110",
  29331=>"11111101",
  29332=>"00000000",
  29333=>"00000001",
  29334=>"00000010",
  29335=>"11111100",
  29336=>"11111101",
  29337=>"00000000",
  29338=>"11111110",
  29339=>"00000001",
  29340=>"11111100",
  29341=>"00000000",
  29342=>"00000100",
  29343=>"11111111",
  29344=>"00000000",
  29345=>"00000011",
  29346=>"11111110",
  29347=>"11111101",
  29348=>"00000011",
  29349=>"00000000",
  29350=>"11111101",
  29351=>"00000000",
  29352=>"00000000",
  29353=>"00000011",
  29354=>"11111101",
  29355=>"00000101",
  29356=>"00000000",
  29357=>"11111110",
  29358=>"00000010",
  29359=>"00000101",
  29360=>"00000001",
  29361=>"00000011",
  29362=>"00000010",
  29363=>"00000000",
  29364=>"11111111",
  29365=>"00000000",
  29366=>"00000000",
  29367=>"00000000",
  29368=>"11111110",
  29369=>"00000011",
  29370=>"00000000",
  29371=>"11111101",
  29372=>"00000000",
  29373=>"11111101",
  29374=>"00000011",
  29375=>"11111110",
  29376=>"00000010",
  29377=>"00000101",
  29378=>"11111111",
  29379=>"00000001",
  29380=>"00000000",
  29381=>"11111111",
  29382=>"11111111",
  29383=>"11111110",
  29384=>"11111111",
  29385=>"11111111",
  29386=>"00000100",
  29387=>"11111101",
  29388=>"00000000",
  29389=>"00000001",
  29390=>"00000001",
  29391=>"00000001",
  29392=>"00000001",
  29393=>"00000001",
  29394=>"11111110",
  29395=>"11111111",
  29396=>"11111101",
  29397=>"00000010",
  29398=>"00000001",
  29399=>"11111111",
  29400=>"00000101",
  29401=>"00000001",
  29402=>"11111111",
  29403=>"11111111",
  29404=>"11111111",
  29405=>"11111101",
  29406=>"00000001",
  29407=>"11111111",
  29408=>"00000001",
  29409=>"00000001",
  29410=>"11111111",
  29411=>"11111110",
  29412=>"11111101",
  29413=>"00000001",
  29414=>"11111111",
  29415=>"00000001",
  29416=>"11111110",
  29417=>"11111111",
  29418=>"00000000",
  29419=>"00000010",
  29420=>"00000011",
  29421=>"00000001",
  29422=>"00000000",
  29423=>"00000010",
  29424=>"11111110",
  29425=>"00000010",
  29426=>"00000010",
  29427=>"00000000",
  29428=>"00000011",
  29429=>"00000001",
  29430=>"00000011",
  29431=>"00000000",
  29432=>"00000101",
  29433=>"11111100",
  29434=>"00000010",
  29435=>"11111101",
  29436=>"11111110",
  29437=>"11111111",
  29438=>"00000001",
  29439=>"00000010",
  29440=>"11111110",
  29441=>"00000001",
  29442=>"11111111",
  29443=>"11111111",
  29444=>"11111111",
  29445=>"00000000",
  29446=>"11111110",
  29447=>"00000001",
  29448=>"00000001",
  29449=>"00000010",
  29450=>"00000001",
  29451=>"00000010",
  29452=>"00000000",
  29453=>"11111110",
  29454=>"11111110",
  29455=>"00000010",
  29456=>"11111101",
  29457=>"00000010",
  29458=>"11111110",
  29459=>"00000000",
  29460=>"11111111",
  29461=>"11111110",
  29462=>"11111111",
  29463=>"11111111",
  29464=>"00000000",
  29465=>"11111111",
  29466=>"00000000",
  29467=>"00000001",
  29468=>"00000011",
  29469=>"00000011",
  29470=>"00000000",
  29471=>"00000001",
  29472=>"00000010",
  29473=>"00000000",
  29474=>"00000000",
  29475=>"11111110",
  29476=>"11111110",
  29477=>"00000001",
  29478=>"00000001",
  29479=>"11111101",
  29480=>"00000010",
  29481=>"00000001",
  29482=>"00000000",
  29483=>"11111101",
  29484=>"00000001",
  29485=>"11111101",
  29486=>"11111100",
  29487=>"00000010",
  29488=>"11111101",
  29489=>"00000000",
  29490=>"11111111",
  29491=>"00000000",
  29492=>"00000001",
  29493=>"11111111",
  29494=>"00000000",
  29495=>"00000110",
  29496=>"00000001",
  29497=>"11111101",
  29498=>"11111111",
  29499=>"11111011",
  29500=>"11111101",
  29501=>"00000100",
  29502=>"00000011",
  29503=>"00000011",
  29504=>"11111111",
  29505=>"11111111",
  29506=>"00000110",
  29507=>"00000010",
  29508=>"11111100",
  29509=>"00000001",
  29510=>"00000100",
  29511=>"00000000",
  29512=>"00000000",
  29513=>"00000000",
  29514=>"00000100",
  29515=>"00000011",
  29516=>"00000001",
  29517=>"00000001",
  29518=>"00000000",
  29519=>"00000100",
  29520=>"11111101",
  29521=>"00000010",
  29522=>"11111111",
  29523=>"00000001",
  29524=>"00000000",
  29525=>"11111101",
  29526=>"00000010",
  29527=>"00000100",
  29528=>"11111111",
  29529=>"11111111",
  29530=>"00000011",
  29531=>"00000001",
  29532=>"11111110",
  29533=>"00000100",
  29534=>"11111110",
  29535=>"00000010",
  29536=>"11111110",
  29537=>"11111111",
  29538=>"00000001",
  29539=>"11111111",
  29540=>"00000010",
  29541=>"11111111",
  29542=>"00000010",
  29543=>"11111110",
  29544=>"11111111",
  29545=>"00000001",
  29546=>"11111110",
  29547=>"11111111",
  29548=>"00000001",
  29549=>"00000111",
  29550=>"11111101",
  29551=>"00000001",
  29552=>"00000100",
  29553=>"11111111",
  29554=>"00000001",
  29555=>"11111111",
  29556=>"00000001",
  29557=>"00000001",
  29558=>"11111110",
  29559=>"00000010",
  29560=>"00000101",
  29561=>"11111110",
  29562=>"11111111",
  29563=>"11111110",
  29564=>"11111100",
  29565=>"00000000",
  29566=>"11111101",
  29567=>"11111110",
  29568=>"00000000",
  29569=>"00000010",
  29570=>"00000010",
  29571=>"00000001",
  29572=>"11111111",
  29573=>"11111111",
  29574=>"00000010",
  29575=>"00000011",
  29576=>"11111110",
  29577=>"11111101",
  29578=>"11111110",
  29579=>"00000110",
  29580=>"00000010",
  29581=>"11111111",
  29582=>"00000000",
  29583=>"00000011",
  29584=>"00000000",
  29585=>"11111101",
  29586=>"11111111",
  29587=>"11111110",
  29588=>"00000011",
  29589=>"11111111",
  29590=>"11111110",
  29591=>"00000001",
  29592=>"00000010",
  29593=>"11111111",
  29594=>"11111101",
  29595=>"00000100",
  29596=>"00000011",
  29597=>"11111110",
  29598=>"00000000",
  29599=>"00000000",
  29600=>"11111111",
  29601=>"00000010",
  29602=>"00000010",
  29603=>"00000010",
  29604=>"11111111",
  29605=>"11111100",
  29606=>"00000011",
  29607=>"00000000",
  29608=>"11111110",
  29609=>"00000001",
  29610=>"11111110",
  29611=>"11111110",
  29612=>"00000110",
  29613=>"00000010",
  29614=>"00000100",
  29615=>"00000000",
  29616=>"11111101",
  29617=>"11111101",
  29618=>"00000010",
  29619=>"11111101",
  29620=>"00000000",
  29621=>"11111011",
  29622=>"00000010",
  29623=>"11111110",
  29624=>"11111111",
  29625=>"11111101",
  29626=>"11111110",
  29627=>"11111111",
  29628=>"11111111",
  29629=>"11111111",
  29630=>"11111110",
  29631=>"00000000",
  29632=>"11111111",
  29633=>"11111110",
  29634=>"11111110",
  29635=>"00000001",
  29636=>"11111110",
  29637=>"00000010",
  29638=>"00000000",
  29639=>"11111111",
  29640=>"00000001",
  29641=>"00000010",
  29642=>"00000000",
  29643=>"11111111",
  29644=>"00000001",
  29645=>"00000000",
  29646=>"11111101",
  29647=>"00000100",
  29648=>"00000000",
  29649=>"11111101",
  29650=>"00000011",
  29651=>"11111110",
  29652=>"11111101",
  29653=>"00000001",
  29654=>"11111111",
  29655=>"00000101",
  29656=>"00000010",
  29657=>"00000001",
  29658=>"11111101",
  29659=>"11111101",
  29660=>"11111111",
  29661=>"11111011",
  29662=>"00000000",
  29663=>"11111111",
  29664=>"00000000",
  29665=>"00000010",
  29666=>"00000000",
  29667=>"11111111",
  29668=>"00000001",
  29669=>"11111101",
  29670=>"11111111",
  29671=>"00000000",
  29672=>"11111101",
  29673=>"11111111",
  29674=>"11111101",
  29675=>"00000011",
  29676=>"00000001",
  29677=>"11111111",
  29678=>"00000001",
  29679=>"11111101",
  29680=>"11111111",
  29681=>"00000010",
  29682=>"11111101",
  29683=>"00000001",
  29684=>"00000001",
  29685=>"00000011",
  29686=>"11111100",
  29687=>"00000001",
  29688=>"00000000",
  29689=>"11111101",
  29690=>"00000100",
  29691=>"00000000",
  29692=>"11111011",
  29693=>"00000000",
  29694=>"11111111",
  29695=>"11111110",
  29696=>"00000001",
  29697=>"11111110",
  29698=>"00000010",
  29699=>"11111111",
  29700=>"11111101",
  29701=>"11111111",
  29702=>"11111110",
  29703=>"11111101",
  29704=>"00000000",
  29705=>"11111110",
  29706=>"00000010",
  29707=>"11111110",
  29708=>"00000000",
  29709=>"00000001",
  29710=>"00000001",
  29711=>"11111111",
  29712=>"00000000",
  29713=>"00000101",
  29714=>"11111111",
  29715=>"11111110",
  29716=>"00000000",
  29717=>"00000001",
  29718=>"00000010",
  29719=>"11111110",
  29720=>"00000001",
  29721=>"00000001",
  29722=>"11111100",
  29723=>"00000100",
  29724=>"11111111",
  29725=>"11111111",
  29726=>"11111110",
  29727=>"00000010",
  29728=>"00000001",
  29729=>"11111110",
  29730=>"11111101",
  29731=>"00000000",
  29732=>"00000000",
  29733=>"11111110",
  29734=>"00000000",
  29735=>"11111111",
  29736=>"00000011",
  29737=>"00000011",
  29738=>"00000000",
  29739=>"11111110",
  29740=>"11111111",
  29741=>"11111101",
  29742=>"11111111",
  29743=>"11111100",
  29744=>"00000001",
  29745=>"00000010",
  29746=>"11111111",
  29747=>"11111111",
  29748=>"00000000",
  29749=>"11111101",
  29750=>"00000001",
  29751=>"11111111",
  29752=>"00000011",
  29753=>"00000000",
  29754=>"11111110",
  29755=>"11111110",
  29756=>"11111101",
  29757=>"00000000",
  29758=>"11111101",
  29759=>"00000001",
  29760=>"00000101",
  29761=>"11111111",
  29762=>"11111111",
  29763=>"11111110",
  29764=>"00000001",
  29765=>"00000010",
  29766=>"00000000",
  29767=>"00000000",
  29768=>"00000000",
  29769=>"11111111",
  29770=>"00000001",
  29771=>"00000010",
  29772=>"11111110",
  29773=>"00000010",
  29774=>"00000011",
  29775=>"00000100",
  29776=>"00000001",
  29777=>"11111111",
  29778=>"11111110",
  29779=>"11111110",
  29780=>"00000000",
  29781=>"00000000",
  29782=>"00000000",
  29783=>"00000000",
  29784=>"00000001",
  29785=>"00000011",
  29786=>"00000001",
  29787=>"11111101",
  29788=>"11111111",
  29789=>"00000010",
  29790=>"00000001",
  29791=>"11111101",
  29792=>"11111111",
  29793=>"11111101",
  29794=>"11111111",
  29795=>"11111101",
  29796=>"00000010",
  29797=>"11111110",
  29798=>"00000000",
  29799=>"11111111",
  29800=>"11111111",
  29801=>"11111110",
  29802=>"00000001",
  29803=>"00000000",
  29804=>"11111100",
  29805=>"11111111",
  29806=>"11111110",
  29807=>"00000010",
  29808=>"00000001",
  29809=>"00000001",
  29810=>"11111101",
  29811=>"11111110",
  29812=>"11111101",
  29813=>"00000001",
  29814=>"00000010",
  29815=>"00000011",
  29816=>"00000001",
  29817=>"11111111",
  29818=>"11111101",
  29819=>"11111101",
  29820=>"00000000",
  29821=>"00000011",
  29822=>"00000001",
  29823=>"00000011",
  29824=>"00000100",
  29825=>"11111101",
  29826=>"11111101",
  29827=>"00000010",
  29828=>"11111110",
  29829=>"00000001",
  29830=>"11111110",
  29831=>"11111110",
  29832=>"00000001",
  29833=>"00000000",
  29834=>"11111110",
  29835=>"11111101",
  29836=>"11111101",
  29837=>"00000001",
  29838=>"00000010",
  29839=>"00000010",
  29840=>"11111111",
  29841=>"11111100",
  29842=>"11111101",
  29843=>"00000000",
  29844=>"00000100",
  29845=>"00000001",
  29846=>"11111111",
  29847=>"00000001",
  29848=>"11111110",
  29849=>"11111111",
  29850=>"00000100",
  29851=>"00000011",
  29852=>"00000000",
  29853=>"11111111",
  29854=>"00000001",
  29855=>"11111111",
  29856=>"11111111",
  29857=>"00000010",
  29858=>"11111110",
  29859=>"11111111",
  29860=>"00000000",
  29861=>"00000000",
  29862=>"00000010",
  29863=>"00000000",
  29864=>"11111110",
  29865=>"11111111",
  29866=>"00000001",
  29867=>"11111110",
  29868=>"11111101",
  29869=>"00000000",
  29870=>"11111100",
  29871=>"00000001",
  29872=>"00000000",
  29873=>"11111110",
  29874=>"11111110",
  29875=>"11111111",
  29876=>"00000001",
  29877=>"00000000",
  29878=>"11111110",
  29879=>"11111111",
  29880=>"11111111",
  29881=>"11111111",
  29882=>"11111101",
  29883=>"00000100",
  29884=>"00000000",
  29885=>"00000001",
  29886=>"00000000",
  29887=>"11111110",
  29888=>"00000010",
  29889=>"00000010",
  29890=>"00000010",
  29891=>"11111100",
  29892=>"00000000",
  29893=>"11111111",
  29894=>"11111111",
  29895=>"00000011",
  29896=>"00000011",
  29897=>"00000101",
  29898=>"11111110",
  29899=>"00000011",
  29900=>"11111110",
  29901=>"11111111",
  29902=>"11111111",
  29903=>"00000001",
  29904=>"11111110",
  29905=>"00000010",
  29906=>"11111111",
  29907=>"11111110",
  29908=>"11111110",
  29909=>"00000100",
  29910=>"00000000",
  29911=>"00000010",
  29912=>"00000010",
  29913=>"11111111",
  29914=>"00000001",
  29915=>"00000001",
  29916=>"11111101",
  29917=>"11111100",
  29918=>"00000011",
  29919=>"00000000",
  29920=>"11111110",
  29921=>"00000001",
  29922=>"00000001",
  29923=>"00000000",
  29924=>"11111111",
  29925=>"11111101",
  29926=>"00000000",
  29927=>"11111110",
  29928=>"11111110",
  29929=>"11111111",
  29930=>"11111101",
  29931=>"00000000",
  29932=>"11111101",
  29933=>"11111111",
  29934=>"11111111",
  29935=>"11111111",
  29936=>"11111101",
  29937=>"00000101",
  29938=>"00000001",
  29939=>"11111111",
  29940=>"00000001",
  29941=>"00000101",
  29942=>"00000011",
  29943=>"00000001",
  29944=>"00000010",
  29945=>"00000001",
  29946=>"11111100",
  29947=>"00000000",
  29948=>"00000010",
  29949=>"11111101",
  29950=>"11111111",
  29951=>"00000001",
  29952=>"00000000",
  29953=>"00000010",
  29954=>"00000010",
  29955=>"11111101",
  29956=>"11111110",
  29957=>"11111110",
  29958=>"11111111",
  29959=>"11111110",
  29960=>"00000001",
  29961=>"11111110",
  29962=>"00000011",
  29963=>"00000010",
  29964=>"00000001",
  29965=>"00000000",
  29966=>"11111111",
  29967=>"00000011",
  29968=>"11111110",
  29969=>"00000010",
  29970=>"11111101",
  29971=>"00000110",
  29972=>"00000001",
  29973=>"11111101",
  29974=>"11111110",
  29975=>"11111110",
  29976=>"00000000",
  29977=>"00000000",
  29978=>"00000010",
  29979=>"00000000",
  29980=>"11111111",
  29981=>"11111110",
  29982=>"00000000",
  29983=>"11111110",
  29984=>"11111111",
  29985=>"11111101",
  29986=>"11111111",
  29987=>"00000001",
  29988=>"11111101",
  29989=>"11111110",
  29990=>"00000010",
  29991=>"11111101",
  29992=>"00000000",
  29993=>"00000011",
  29994=>"11111110",
  29995=>"11111111",
  29996=>"11111110",
  29997=>"00000000",
  29998=>"11111111",
  29999=>"11111111",
  30000=>"00000000",
  30001=>"11111111",
  30002=>"11111110",
  30003=>"00000010",
  30004=>"11111111",
  30005=>"00000000",
  30006=>"00000010",
  30007=>"11111110",
  30008=>"11111101",
  30009=>"00000001",
  30010=>"00000010",
  30011=>"00000010",
  30012=>"00000011",
  30013=>"11111110",
  30014=>"00000001",
  30015=>"11111110",
  30016=>"11111111",
  30017=>"00000111",
  30018=>"00000000",
  30019=>"00000000",
  30020=>"11111111",
  30021=>"11111111",
  30022=>"00000111",
  30023=>"11111111",
  30024=>"11111101",
  30025=>"00000110",
  30026=>"11111111",
  30027=>"11111110",
  30028=>"00000000",
  30029=>"00000010",
  30030=>"00000000",
  30031=>"11111100",
  30032=>"11111101",
  30033=>"00000011",
  30034=>"00000000",
  30035=>"11111111",
  30036=>"11111111",
  30037=>"11111111",
  30038=>"00000010",
  30039=>"00000011",
  30040=>"11111101",
  30041=>"11111111",
  30042=>"00000011",
  30043=>"11111100",
  30044=>"00000000",
  30045=>"00000001",
  30046=>"11111111",
  30047=>"00000011",
  30048=>"00000000",
  30049=>"00000100",
  30050=>"11111111",
  30051=>"11111101",
  30052=>"11111111",
  30053=>"11111110",
  30054=>"00000000",
  30055=>"11111110",
  30056=>"11111101",
  30057=>"00000011",
  30058=>"00000000",
  30059=>"00000000",
  30060=>"00000000",
  30061=>"11111101",
  30062=>"00000010",
  30063=>"00000010",
  30064=>"00000011",
  30065=>"11111110",
  30066=>"11111110",
  30067=>"11111111",
  30068=>"00000010",
  30069=>"11111100",
  30070=>"00000001",
  30071=>"00000010",
  30072=>"00000000",
  30073=>"00000100",
  30074=>"11111110",
  30075=>"11111101",
  30076=>"00000000",
  30077=>"11111110",
  30078=>"11111111",
  30079=>"11111101",
  30080=>"11111110",
  30081=>"00000010",
  30082=>"11111110",
  30083=>"00000000",
  30084=>"00000011",
  30085=>"11111110",
  30086=>"00000010",
  30087=>"11111110",
  30088=>"11111100",
  30089=>"11111111",
  30090=>"00000001",
  30091=>"00000000",
  30092=>"00000001",
  30093=>"11111111",
  30094=>"11111111",
  30095=>"11111110",
  30096=>"00000001",
  30097=>"00000001",
  30098=>"00000011",
  30099=>"00000000",
  30100=>"00000010",
  30101=>"00000000",
  30102=>"11111111",
  30103=>"11111111",
  30104=>"00000000",
  30105=>"00000010",
  30106=>"00000000",
  30107=>"00000001",
  30108=>"00000010",
  30109=>"11111101",
  30110=>"00000010",
  30111=>"11111111",
  30112=>"00000010",
  30113=>"11111101",
  30114=>"00000000",
  30115=>"00000000",
  30116=>"11111111",
  30117=>"00000010",
  30118=>"00000011",
  30119=>"11111111",
  30120=>"00000100",
  30121=>"00000001",
  30122=>"11111101",
  30123=>"11111111",
  30124=>"11111110",
  30125=>"00000000",
  30126=>"00000011",
  30127=>"11111110",
  30128=>"11111100",
  30129=>"00000001",
  30130=>"00000000",
  30131=>"00000010",
  30132=>"11111110",
  30133=>"00000111",
  30134=>"11111110",
  30135=>"00000000",
  30136=>"11111111",
  30137=>"11111101",
  30138=>"00000001",
  30139=>"11111111",
  30140=>"11111110",
  30141=>"00000010",
  30142=>"00000001",
  30143=>"00000010",
  30144=>"00000001",
  30145=>"11111111",
  30146=>"00000010",
  30147=>"11111110",
  30148=>"00000010",
  30149=>"00000010",
  30150=>"00000100",
  30151=>"00000101",
  30152=>"11111110",
  30153=>"00000000",
  30154=>"11111111",
  30155=>"00000000",
  30156=>"00000011",
  30157=>"11111110",
  30158=>"00000000",
  30159=>"00000011",
  30160=>"00000011",
  30161=>"11111101",
  30162=>"00000001",
  30163=>"00000000",
  30164=>"11111101",
  30165=>"11111101",
  30166=>"11111100",
  30167=>"11111111",
  30168=>"11111111",
  30169=>"00000010",
  30170=>"00000000",
  30171=>"11111110",
  30172=>"11111110",
  30173=>"11111111",
  30174=>"11111111",
  30175=>"00000110",
  30176=>"11111111",
  30177=>"11111101",
  30178=>"11111100",
  30179=>"11111111",
  30180=>"00000001",
  30181=>"00000001",
  30182=>"11111101",
  30183=>"11111101",
  30184=>"11111101",
  30185=>"00000000",
  30186=>"00000000",
  30187=>"11111101",
  30188=>"00000100",
  30189=>"11111101",
  30190=>"11111101",
  30191=>"00000100",
  30192=>"11111111",
  30193=>"00000010",
  30194=>"11111101",
  30195=>"11111110",
  30196=>"00000010",
  30197=>"11111101",
  30198=>"00000000",
  30199=>"11111101",
  30200=>"00000010",
  30201=>"00000010",
  30202=>"00000000",
  30203=>"11111101",
  30204=>"00000000",
  30205=>"00000100",
  30206=>"11111101",
  30207=>"11111110",
  30208=>"00000011",
  30209=>"11111101",
  30210=>"11111111",
  30211=>"00000001",
  30212=>"00000001",
  30213=>"00000000",
  30214=>"00000001",
  30215=>"00000000",
  30216=>"11111110",
  30217=>"11111111",
  30218=>"00000001",
  30219=>"00000010",
  30220=>"00000001",
  30221=>"00000001",
  30222=>"00000000",
  30223=>"00000000",
  30224=>"00000000",
  30225=>"00000010",
  30226=>"00000011",
  30227=>"00000010",
  30228=>"00000001",
  30229=>"00000001",
  30230=>"00000001",
  30231=>"00000001",
  30232=>"11111110",
  30233=>"11111100",
  30234=>"00000000",
  30235=>"00000001",
  30236=>"11111110",
  30237=>"00000000",
  30238=>"00000001",
  30239=>"11111100",
  30240=>"00000001",
  30241=>"11111101",
  30242=>"00000001",
  30243=>"11111111",
  30244=>"00000010",
  30245=>"00000000",
  30246=>"00000011",
  30247=>"00000010",
  30248=>"00000010",
  30249=>"00000000",
  30250=>"00000110",
  30251=>"11111110",
  30252=>"11111110",
  30253=>"00000001",
  30254=>"11111100",
  30255=>"00000000",
  30256=>"11111101",
  30257=>"11111101",
  30258=>"11111110",
  30259=>"11111101",
  30260=>"00000000",
  30261=>"00000011",
  30262=>"00000001",
  30263=>"00000000",
  30264=>"11111101",
  30265=>"11111110",
  30266=>"11111101",
  30267=>"11111110",
  30268=>"00000100",
  30269=>"00000101",
  30270=>"11111111",
  30271=>"00000001",
  30272=>"11111101",
  30273=>"11111110",
  30274=>"11111101",
  30275=>"00000010",
  30276=>"00000000",
  30277=>"11111101",
  30278=>"00000010",
  30279=>"11111110",
  30280=>"00000001",
  30281=>"00000001",
  30282=>"00000000",
  30283=>"11111100",
  30284=>"11111111",
  30285=>"00000001",
  30286=>"00000000",
  30287=>"00000000",
  30288=>"00000001",
  30289=>"11111101",
  30290=>"00000001",
  30291=>"11111111",
  30292=>"11111101",
  30293=>"11111110",
  30294=>"11111110",
  30295=>"11111101",
  30296=>"11111111",
  30297=>"11111111",
  30298=>"11111111",
  30299=>"00000000",
  30300=>"11111110",
  30301=>"00000011",
  30302=>"11111110",
  30303=>"00000001",
  30304=>"00000010",
  30305=>"11111110",
  30306=>"11111111",
  30307=>"11111110",
  30308=>"00000000",
  30309=>"11111111",
  30310=>"11111100",
  30311=>"11111101",
  30312=>"00000001",
  30313=>"00000001",
  30314=>"11111110",
  30315=>"11111111",
  30316=>"00000000",
  30317=>"00000100",
  30318=>"00000001",
  30319=>"00000000",
  30320=>"11111101",
  30321=>"00000001",
  30322=>"11111101",
  30323=>"11111100",
  30324=>"00000001",
  30325=>"11111110",
  30326=>"11111101",
  30327=>"11111111",
  30328=>"11111111",
  30329=>"00000001",
  30330=>"00000011",
  30331=>"00000100",
  30332=>"11111111",
  30333=>"11111101",
  30334=>"11111101",
  30335=>"11111111",
  30336=>"11111111",
  30337=>"00000000",
  30338=>"00000010",
  30339=>"00000000",
  30340=>"00000001",
  30341=>"00000001",
  30342=>"00000100",
  30343=>"00000010",
  30344=>"00000001",
  30345=>"00000010",
  30346=>"11111110",
  30347=>"11111111",
  30348=>"00000010",
  30349=>"11111110",
  30350=>"11111110",
  30351=>"00000011",
  30352=>"00000001",
  30353=>"11111110",
  30354=>"00000011",
  30355=>"00000000",
  30356=>"00000000",
  30357=>"11111101",
  30358=>"00000010",
  30359=>"11111100",
  30360=>"00000001",
  30361=>"11111111",
  30362=>"00000010",
  30363=>"11111110",
  30364=>"00000000",
  30365=>"11111110",
  30366=>"00000001",
  30367=>"00000011",
  30368=>"00000010",
  30369=>"11111110",
  30370=>"00000001",
  30371=>"00000001",
  30372=>"00000000",
  30373=>"00000000",
  30374=>"00000001",
  30375=>"00000001",
  30376=>"11111111",
  30377=>"00000000",
  30378=>"00000000",
  30379=>"11111101",
  30380=>"00000001",
  30381=>"00000010",
  30382=>"00000010",
  30383=>"00000000",
  30384=>"00000001",
  30385=>"00000110",
  30386=>"00000010",
  30387=>"11111111",
  30388=>"00000010",
  30389=>"00000001",
  30390=>"11111111",
  30391=>"00000001",
  30392=>"11111111",
  30393=>"11111111",
  30394=>"00000010",
  30395=>"11111101",
  30396=>"11111111",
  30397=>"11111111",
  30398=>"11111101",
  30399=>"11111111",
  30400=>"00000010",
  30401=>"00000001",
  30402=>"11111110",
  30403=>"11111110",
  30404=>"11111101",
  30405=>"00000011",
  30406=>"00000010",
  30407=>"00000001",
  30408=>"11111111",
  30409=>"11111100",
  30410=>"11111111",
  30411=>"11111101",
  30412=>"00000001",
  30413=>"00000000",
  30414=>"00000000",
  30415=>"00000001",
  30416=>"11111111",
  30417=>"00000000",
  30418=>"11111101",
  30419=>"11111110",
  30420=>"11111110",
  30421=>"11111111",
  30422=>"00000010",
  30423=>"00000010",
  30424=>"00000011",
  30425=>"00000001",
  30426=>"00000001",
  30427=>"00000001",
  30428=>"11111111",
  30429=>"00000001",
  30430=>"11111110",
  30431=>"11111100",
  30432=>"00000000",
  30433=>"11111110",
  30434=>"00000001",
  30435=>"11111111",
  30436=>"11111101",
  30437=>"00000010",
  30438=>"00000010",
  30439=>"11111111",
  30440=>"00000001",
  30441=>"00000001",
  30442=>"00000000",
  30443=>"00000000",
  30444=>"00000010",
  30445=>"11111110",
  30446=>"11111110",
  30447=>"11111101",
  30448=>"11111111",
  30449=>"00000000",
  30450=>"11111110",
  30451=>"00000001",
  30452=>"00000010",
  30453=>"11111111",
  30454=>"11111111",
  30455=>"00000001",
  30456=>"11111101",
  30457=>"11111100",
  30458=>"11111111",
  30459=>"11111110",
  30460=>"00000001",
  30461=>"00000001",
  30462=>"00000000",
  30463=>"11111101",
  30464=>"11111111",
  30465=>"00000001",
  30466=>"00000000",
  30467=>"00000000",
  30468=>"00000000",
  30469=>"11111111",
  30470=>"11111101",
  30471=>"11111110",
  30472=>"00000001",
  30473=>"00000001",
  30474=>"00000010",
  30475=>"00000010",
  30476=>"11111101",
  30477=>"11111101",
  30478=>"00000001",
  30479=>"00000001",
  30480=>"00000000",
  30481=>"11111110",
  30482=>"11111110",
  30483=>"00000001",
  30484=>"00000001",
  30485=>"00000011",
  30486=>"00000000",
  30487=>"00000000",
  30488=>"00000100",
  30489=>"00000010",
  30490=>"11111100",
  30491=>"00000000",
  30492=>"11111100",
  30493=>"00000001",
  30494=>"00000010",
  30495=>"00000001",
  30496=>"11111101",
  30497=>"11111111",
  30498=>"00000000",
  30499=>"00000001",
  30500=>"00000001",
  30501=>"00000000",
  30502=>"00000010",
  30503=>"00000000",
  30504=>"00000000",
  30505=>"00000100",
  30506=>"00000000",
  30507=>"00000000",
  30508=>"00000010",
  30509=>"11111111",
  30510=>"11111100",
  30511=>"00000001",
  30512=>"00000100",
  30513=>"11111111",
  30514=>"00000010",
  30515=>"11111110",
  30516=>"11111111",
  30517=>"00000001",
  30518=>"11111110",
  30519=>"11111110",
  30520=>"00000010",
  30521=>"11111111",
  30522=>"00000010",
  30523=>"11111110",
  30524=>"00000001",
  30525=>"00000000",
  30526=>"11111110",
  30527=>"00000001",
  30528=>"00000101",
  30529=>"00000001",
  30530=>"00000000",
  30531=>"00000011",
  30532=>"11111111",
  30533=>"11111111",
  30534=>"11111110",
  30535=>"00000001",
  30536=>"11111011",
  30537=>"00000010",
  30538=>"11111110",
  30539=>"00000100",
  30540=>"11111110",
  30541=>"11111111",
  30542=>"11111111",
  30543=>"00000001",
  30544=>"00000010",
  30545=>"00000001",
  30546=>"11111110",
  30547=>"11111100",
  30548=>"11111111",
  30549=>"00000000",
  30550=>"11111111",
  30551=>"00000000",
  30552=>"00000100",
  30553=>"11111110",
  30554=>"11111110",
  30555=>"00000011",
  30556=>"00000001",
  30557=>"00000000",
  30558=>"11111111",
  30559=>"00000000",
  30560=>"11111111",
  30561=>"00000010",
  30562=>"11111111",
  30563=>"00000010",
  30564=>"11111110",
  30565=>"00000010",
  30566=>"00000000",
  30567=>"11111110",
  30568=>"00000000",
  30569=>"00000010",
  30570=>"11111110",
  30571=>"00000011",
  30572=>"00000011",
  30573=>"00000000",
  30574=>"00000101",
  30575=>"00000001",
  30576=>"00000010",
  30577=>"00000001",
  30578=>"00000010",
  30579=>"00000000",
  30580=>"11111110",
  30581=>"11111101",
  30582=>"00000010",
  30583=>"11111101",
  30584=>"11111101",
  30585=>"00000011",
  30586=>"11111111",
  30587=>"00000011",
  30588=>"00000001",
  30589=>"00000010",
  30590=>"11111111",
  30591=>"00000000",
  30592=>"00000010",
  30593=>"00000011",
  30594=>"00000000",
  30595=>"11111100",
  30596=>"00000000",
  30597=>"11111110",
  30598=>"00000000",
  30599=>"11111101",
  30600=>"11111111",
  30601=>"11111111",
  30602=>"00000001",
  30603=>"00000010",
  30604=>"11111111",
  30605=>"11111110",
  30606=>"00000011",
  30607=>"00000001",
  30608=>"00000010",
  30609=>"11111110",
  30610=>"00000010",
  30611=>"11111110",
  30612=>"11111111",
  30613=>"11111110",
  30614=>"11111110",
  30615=>"00000001",
  30616=>"11111101",
  30617=>"00000000",
  30618=>"00000000",
  30619=>"00000010",
  30620=>"00000010",
  30621=>"11111111",
  30622=>"11111111",
  30623=>"11111111",
  30624=>"11111100",
  30625=>"11111110",
  30626=>"11111111",
  30627=>"00000001",
  30628=>"11111111",
  30629=>"00000010",
  30630=>"00000100",
  30631=>"11111101",
  30632=>"11111111",
  30633=>"00000000",
  30634=>"00000001",
  30635=>"00000000",
  30636=>"00000000",
  30637=>"11111110",
  30638=>"11111110",
  30639=>"00000000",
  30640=>"00000000",
  30641=>"00000001",
  30642=>"00000100",
  30643=>"11111101",
  30644=>"00000010",
  30645=>"00000011",
  30646=>"00000010",
  30647=>"11111100",
  30648=>"00000001",
  30649=>"11111111",
  30650=>"00000001",
  30651=>"11111110",
  30652=>"00000001",
  30653=>"11111111",
  30654=>"00000000",
  30655=>"00000010",
  30656=>"00000010",
  30657=>"11111111",
  30658=>"00000000",
  30659=>"00000010",
  30660=>"11111101",
  30661=>"11111111",
  30662=>"00000011",
  30663=>"11111111",
  30664=>"00000001",
  30665=>"00000001",
  30666=>"00000010",
  30667=>"00000000",
  30668=>"00000010",
  30669=>"11111101",
  30670=>"11111110",
  30671=>"00000000",
  30672=>"00000001",
  30673=>"00000011",
  30674=>"00000000",
  30675=>"00000010",
  30676=>"00000010",
  30677=>"11111110",
  30678=>"00000010",
  30679=>"11111100",
  30680=>"00000010",
  30681=>"00000001",
  30682=>"11111111",
  30683=>"00000000",
  30684=>"11111101",
  30685=>"11111101",
  30686=>"11111110",
  30687=>"00000101",
  30688=>"11111110",
  30689=>"00000001",
  30690=>"00000000",
  30691=>"11111111",
  30692=>"11111110",
  30693=>"00000000",
  30694=>"00000010",
  30695=>"00000010",
  30696=>"11111111",
  30697=>"11111111",
  30698=>"00000000",
  30699=>"11111101",
  30700=>"00000000",
  30701=>"00000001",
  30702=>"00000000",
  30703=>"11111110",
  30704=>"00000000",
  30705=>"11111111",
  30706=>"11111101",
  30707=>"11111111",
  30708=>"00000001",
  30709=>"11111101",
  30710=>"11111111",
  30711=>"00000001",
  30712=>"00000010",
  30713=>"11111110",
  30714=>"11111110",
  30715=>"11111101",
  30716=>"11111101",
  30717=>"00000011",
  30718=>"00000000",
  30719=>"11111111",
  30720=>"11111110",
  30721=>"00000000",
  30722=>"00000001",
  30723=>"11111110",
  30724=>"11111100",
  30725=>"11111110",
  30726=>"11111110",
  30727=>"11111111",
  30728=>"00000010",
  30729=>"00000011",
  30730=>"00000001",
  30731=>"11111110",
  30732=>"11111111",
  30733=>"11111111",
  30734=>"00000001",
  30735=>"11111101",
  30736=>"00000011",
  30737=>"00000100",
  30738=>"00000010",
  30739=>"11111110",
  30740=>"11111101",
  30741=>"11111101",
  30742=>"11111101",
  30743=>"11111101",
  30744=>"11111101",
  30745=>"11111100",
  30746=>"11111101",
  30747=>"11111111",
  30748=>"00000000",
  30749=>"00000001",
  30750=>"00000010",
  30751=>"00000001",
  30752=>"11111110",
  30753=>"11111111",
  30754=>"11111101",
  30755=>"11111111",
  30756=>"00000001",
  30757=>"00000000",
  30758=>"00000000",
  30759=>"11111111",
  30760=>"11111101",
  30761=>"11111110",
  30762=>"00000010",
  30763=>"00000000",
  30764=>"00000000",
  30765=>"00000000",
  30766=>"00000001",
  30767=>"11111111",
  30768=>"11111111",
  30769=>"11111110",
  30770=>"00000001",
  30771=>"00000000",
  30772=>"11111111",
  30773=>"11111111",
  30774=>"00000000",
  30775=>"00000000",
  30776=>"00000000",
  30777=>"00000010",
  30778=>"00000010",
  30779=>"11111110",
  30780=>"11111111",
  30781=>"11111111",
  30782=>"11111101",
  30783=>"00000001",
  30784=>"00000000",
  30785=>"11111110",
  30786=>"00000001",
  30787=>"11111111",
  30788=>"00000000",
  30789=>"00000000",
  30790=>"00000011",
  30791=>"00000000",
  30792=>"00000000",
  30793=>"11111111",
  30794=>"11111110",
  30795=>"11111110",
  30796=>"00000001",
  30797=>"11111101",
  30798=>"11111110",
  30799=>"11111111",
  30800=>"11111110",
  30801=>"00000010",
  30802=>"00000011",
  30803=>"00000010",
  30804=>"11111111",
  30805=>"00000010",
  30806=>"11111101",
  30807=>"11111110",
  30808=>"11111101",
  30809=>"00000100",
  30810=>"00000000",
  30811=>"11111111",
  30812=>"00000110",
  30813=>"00000000",
  30814=>"00000001",
  30815=>"00000000",
  30816=>"00000001",
  30817=>"11111110",
  30818=>"00000010",
  30819=>"11111111",
  30820=>"00000001",
  30821=>"00000000",
  30822=>"11111101",
  30823=>"11111110",
  30824=>"11111101",
  30825=>"11111111",
  30826=>"11111111",
  30827=>"11111110",
  30828=>"00000010",
  30829=>"00000110",
  30830=>"11111111",
  30831=>"00000000",
  30832=>"00000000",
  30833=>"11111111",
  30834=>"11111101",
  30835=>"11111101",
  30836=>"11111101",
  30837=>"11111110",
  30838=>"11111111",
  30839=>"11111111",
  30840=>"00000001",
  30841=>"00000011",
  30842=>"00000001",
  30843=>"00000011",
  30844=>"00000000",
  30845=>"11111110",
  30846=>"00000000",
  30847=>"11111111",
  30848=>"11111110",
  30849=>"11111110",
  30850=>"00000010",
  30851=>"11111101",
  30852=>"11111100",
  30853=>"11111101",
  30854=>"11111111",
  30855=>"11111100",
  30856=>"00000000",
  30857=>"00000001",
  30858=>"11111111",
  30859=>"00000101",
  30860=>"11111111",
  30861=>"00000010",
  30862=>"11111110",
  30863=>"11111101",
  30864=>"00000000",
  30865=>"00000010",
  30866=>"11111111",
  30867=>"11111110",
  30868=>"00000101",
  30869=>"00000011",
  30870=>"11111110",
  30871=>"00000101",
  30872=>"00000110",
  30873=>"11111110",
  30874=>"00000001",
  30875=>"11111110",
  30876=>"00000000",
  30877=>"11111111",
  30878=>"00000010",
  30879=>"00000100",
  30880=>"00000001",
  30881=>"00000010",
  30882=>"11111100",
  30883=>"00000010",
  30884=>"11111101",
  30885=>"11111110",
  30886=>"00000100",
  30887=>"11111111",
  30888=>"11111100",
  30889=>"11111111",
  30890=>"11111111",
  30891=>"00000010",
  30892=>"00000010",
  30893=>"11111111",
  30894=>"00000000",
  30895=>"11111110",
  30896=>"11111111",
  30897=>"11111110",
  30898=>"11111110",
  30899=>"11111101",
  30900=>"00000110",
  30901=>"00000001",
  30902=>"00000011",
  30903=>"00000000",
  30904=>"11111101",
  30905=>"11111111",
  30906=>"11111110",
  30907=>"00000001",
  30908=>"00000011",
  30909=>"11111110",
  30910=>"00000001",
  30911=>"00000001",
  30912=>"11111101",
  30913=>"00000010",
  30914=>"11111111",
  30915=>"11111111",
  30916=>"11111110",
  30917=>"11111101",
  30918=>"00000001",
  30919=>"11111110",
  30920=>"11111111",
  30921=>"00000101",
  30922=>"00000001",
  30923=>"11111110",
  30924=>"00000001",
  30925=>"00000001",
  30926=>"11111111",
  30927=>"00000001",
  30928=>"00000011",
  30929=>"00000001",
  30930=>"00000000",
  30931=>"00000000",
  30932=>"00000000",
  30933=>"00000001",
  30934=>"00000001",
  30935=>"00000010",
  30936=>"00000010",
  30937=>"00000001",
  30938=>"00000000",
  30939=>"00000001",
  30940=>"00000001",
  30941=>"11111110",
  30942=>"11111110",
  30943=>"00000010",
  30944=>"11111101",
  30945=>"11111111",
  30946=>"11111101",
  30947=>"11111101",
  30948=>"00000001",
  30949=>"00000000",
  30950=>"11111110",
  30951=>"11111111",
  30952=>"11111111",
  30953=>"11111100",
  30954=>"00000000",
  30955=>"00000010",
  30956=>"00000001",
  30957=>"11111101",
  30958=>"00000000",
  30959=>"11111111",
  30960=>"00000000",
  30961=>"11111100",
  30962=>"00000010",
  30963=>"11111110",
  30964=>"11111111",
  30965=>"11111111",
  30966=>"11111101",
  30967=>"11111111",
  30968=>"00000000",
  30969=>"00000000",
  30970=>"11111110",
  30971=>"00000010",
  30972=>"00000011",
  30973=>"00000000",
  30974=>"00000001",
  30975=>"00000010",
  30976=>"11111110",
  30977=>"00000000",
  30978=>"11111110",
  30979=>"00000001",
  30980=>"11111111",
  30981=>"11111110",
  30982=>"11111101",
  30983=>"00000001",
  30984=>"11111111",
  30985=>"00000100",
  30986=>"00000001",
  30987=>"00000011",
  30988=>"00000001",
  30989=>"11111101",
  30990=>"11111110",
  30991=>"11111111",
  30992=>"11111110",
  30993=>"11111111",
  30994=>"00000010",
  30995=>"00000001",
  30996=>"00000000",
  30997=>"00000010",
  30998=>"11111101",
  30999=>"00000001",
  31000=>"11111111",
  31001=>"11111110",
  31002=>"00000000",
  31003=>"00000000",
  31004=>"00000000",
  31005=>"11111110",
  31006=>"11111111",
  31007=>"00000000",
  31008=>"11111101",
  31009=>"00000000",
  31010=>"00000001",
  31011=>"11111111",
  31012=>"00000010",
  31013=>"00000101",
  31014=>"11111101",
  31015=>"11111110",
  31016=>"00000010",
  31017=>"00000011",
  31018=>"11111101",
  31019=>"00000010",
  31020=>"00000001",
  31021=>"11111111",
  31022=>"11111101",
  31023=>"00000001",
  31024=>"11111111",
  31025=>"00000001",
  31026=>"00000000",
  31027=>"11111101",
  31028=>"00000001",
  31029=>"00000010",
  31030=>"00000000",
  31031=>"00000001",
  31032=>"00000010",
  31033=>"11111110",
  31034=>"11111101",
  31035=>"00000000",
  31036=>"11111111",
  31037=>"11111111",
  31038=>"11111101",
  31039=>"00000000",
  31040=>"00000001",
  31041=>"00000010",
  31042=>"11111101",
  31043=>"00000000",
  31044=>"00000010",
  31045=>"11111101",
  31046=>"00000011",
  31047=>"00000001",
  31048=>"00000010",
  31049=>"00000010",
  31050=>"11111100",
  31051=>"00000001",
  31052=>"00000010",
  31053=>"11111101",
  31054=>"00000001",
  31055=>"11111111",
  31056=>"11111101",
  31057=>"00000000",
  31058=>"11111111",
  31059=>"11111100",
  31060=>"00000010",
  31061=>"11111111",
  31062=>"11111111",
  31063=>"00000000",
  31064=>"00000000",
  31065=>"00000000",
  31066=>"11111110",
  31067=>"11111101",
  31068=>"00000010",
  31069=>"11111110",
  31070=>"00000001",
  31071=>"00000001",
  31072=>"11111110",
  31073=>"00000011",
  31074=>"00000000",
  31075=>"11111100",
  31076=>"00000010",
  31077=>"00000010",
  31078=>"00000001",
  31079=>"00000010",
  31080=>"00000000",
  31081=>"00000000",
  31082=>"00000010",
  31083=>"00000000",
  31084=>"00000000",
  31085=>"11111111",
  31086=>"11111101",
  31087=>"00000001",
  31088=>"00000001",
  31089=>"11111111",
  31090=>"00000011",
  31091=>"00000000",
  31092=>"00000000",
  31093=>"00000000",
  31094=>"11111110",
  31095=>"11111110",
  31096=>"00000100",
  31097=>"00000000",
  31098=>"11111101",
  31099=>"00000101",
  31100=>"00000000",
  31101=>"00000111",
  31102=>"00000000",
  31103=>"00000010",
  31104=>"00000010",
  31105=>"00000011",
  31106=>"00000010",
  31107=>"00000001",
  31108=>"00000010",
  31109=>"00000001",
  31110=>"00000010",
  31111=>"00000000",
  31112=>"00000100",
  31113=>"00000000",
  31114=>"11111111",
  31115=>"00000000",
  31116=>"00000010",
  31117=>"00000000",
  31118=>"11111111",
  31119=>"00000001",
  31120=>"00000001",
  31121=>"11111110",
  31122=>"11111111",
  31123=>"00000000",
  31124=>"11111111",
  31125=>"00000001",
  31126=>"00000000",
  31127=>"00000000",
  31128=>"11111101",
  31129=>"00000011",
  31130=>"11111111",
  31131=>"00000010",
  31132=>"00000010",
  31133=>"00000011",
  31134=>"00000000",
  31135=>"11111111",
  31136=>"00000101",
  31137=>"11111111",
  31138=>"11111110",
  31139=>"00000100",
  31140=>"00000011",
  31141=>"00000101",
  31142=>"11111111",
  31143=>"00000100",
  31144=>"00000011",
  31145=>"00000001",
  31146=>"00000000",
  31147=>"11111110",
  31148=>"11111110",
  31149=>"00000010",
  31150=>"11111101",
  31151=>"11111110",
  31152=>"00000011",
  31153=>"11111111",
  31154=>"00000000",
  31155=>"11111111",
  31156=>"11111100",
  31157=>"11111101",
  31158=>"00000000",
  31159=>"11111110",
  31160=>"00000010",
  31161=>"11111110",
  31162=>"11111101",
  31163=>"00000001",
  31164=>"11111110",
  31165=>"00000001",
  31166=>"11111111",
  31167=>"11111110",
  31168=>"11111101",
  31169=>"11111111",
  31170=>"11111100",
  31171=>"00000000",
  31172=>"11111111",
  31173=>"00000000",
  31174=>"00000010",
  31175=>"00000000",
  31176=>"00000000",
  31177=>"11111110",
  31178=>"11111110",
  31179=>"00000010",
  31180=>"11111111",
  31181=>"11111110",
  31182=>"00000001",
  31183=>"11111110",
  31184=>"00000000",
  31185=>"11111110",
  31186=>"00000010",
  31187=>"00000011",
  31188=>"11111110",
  31189=>"00000000",
  31190=>"11111101",
  31191=>"11111110",
  31192=>"00000001",
  31193=>"11111111",
  31194=>"00000010",
  31195=>"11111110",
  31196=>"00000001",
  31197=>"11111101",
  31198=>"11111110",
  31199=>"11111111",
  31200=>"11111111",
  31201=>"11111110",
  31202=>"11111110",
  31203=>"00000011",
  31204=>"00000010",
  31205=>"11111110",
  31206=>"00000100",
  31207=>"11111111",
  31208=>"00000000",
  31209=>"11111101",
  31210=>"00000011",
  31211=>"00000001",
  31212=>"11111110",
  31213=>"00000001",
  31214=>"11111110",
  31215=>"00000010",
  31216=>"00000010",
  31217=>"00000101",
  31218=>"00000001",
  31219=>"11111111",
  31220=>"11111111",
  31221=>"00000010",
  31222=>"00000000",
  31223=>"00000000",
  31224=>"11111101",
  31225=>"00000000",
  31226=>"11111110",
  31227=>"00000100",
  31228=>"00000000",
  31229=>"11111111",
  31230=>"11111101",
  31231=>"11111110",
  31232=>"00000001",
  31233=>"11111110",
  31234=>"11111111",
  31235=>"00000000",
  31236=>"11111111",
  31237=>"11111110",
  31238=>"11111100",
  31239=>"00000010",
  31240=>"11111101",
  31241=>"00000010",
  31242=>"00000000",
  31243=>"11111111",
  31244=>"00000010",
  31245=>"11111111",
  31246=>"11111111",
  31247=>"11111111",
  31248=>"00000000",
  31249=>"00000010",
  31250=>"00000010",
  31251=>"00000011",
  31252=>"00000010",
  31253=>"11111111",
  31254=>"00000010",
  31255=>"00000001",
  31256=>"00000011",
  31257=>"11111101",
  31258=>"00000010",
  31259=>"00000000",
  31260=>"00000001",
  31261=>"00000011",
  31262=>"00000001",
  31263=>"11111111",
  31264=>"11111110",
  31265=>"00000011",
  31266=>"11111101",
  31267=>"11111111",
  31268=>"00000010",
  31269=>"11111100",
  31270=>"11111110",
  31271=>"00000011",
  31272=>"11111101",
  31273=>"00000101",
  31274=>"11111110",
  31275=>"00000101",
  31276=>"11111110",
  31277=>"11111111",
  31278=>"11111110",
  31279=>"00000011",
  31280=>"11111111",
  31281=>"11111110",
  31282=>"11111111",
  31283=>"11111110",
  31284=>"00000010",
  31285=>"11111110",
  31286=>"00000010",
  31287=>"00000001",
  31288=>"11111111",
  31289=>"00000001",
  31290=>"11111110",
  31291=>"11111110",
  31292=>"00000001",
  31293=>"00000100",
  31294=>"11111111",
  31295=>"00000010",
  31296=>"00000100",
  31297=>"11111111",
  31298=>"11111101",
  31299=>"00000001",
  31300=>"00000000",
  31301=>"11111111",
  31302=>"00000001",
  31303=>"11111111",
  31304=>"11111110",
  31305=>"11111101",
  31306=>"00000000",
  31307=>"00000110",
  31308=>"11111111",
  31309=>"00000001",
  31310=>"11111111",
  31311=>"00000000",
  31312=>"11111101",
  31313=>"00000011",
  31314=>"00000001",
  31315=>"00000001",
  31316=>"11111110",
  31317=>"00000001",
  31318=>"00000000",
  31319=>"00000001",
  31320=>"11111110",
  31321=>"00000001",
  31322=>"00000000",
  31323=>"11111100",
  31324=>"00000000",
  31325=>"00000010",
  31326=>"00000001",
  31327=>"00000001",
  31328=>"11111111",
  31329=>"00000010",
  31330=>"11111111",
  31331=>"00000011",
  31332=>"11111111",
  31333=>"11111110",
  31334=>"00000000",
  31335=>"00000000",
  31336=>"11111110",
  31337=>"00000001",
  31338=>"11111110",
  31339=>"00000001",
  31340=>"00000011",
  31341=>"00000000",
  31342=>"11111110",
  31343=>"00000001",
  31344=>"11111111",
  31345=>"11111110",
  31346=>"11111111",
  31347=>"11111111",
  31348=>"00000001",
  31349=>"00000010",
  31350=>"00000100",
  31351=>"11111101",
  31352=>"00000000",
  31353=>"11111110",
  31354=>"11111110",
  31355=>"11111111",
  31356=>"11111110",
  31357=>"00000010",
  31358=>"00000101",
  31359=>"00000000",
  31360=>"00000001",
  31361=>"11111111",
  31362=>"11111111",
  31363=>"11111101",
  31364=>"00000000",
  31365=>"11111100",
  31366=>"00000000",
  31367=>"00000000",
  31368=>"00000001",
  31369=>"00000001",
  31370=>"11111110",
  31371=>"11111111",
  31372=>"00000000",
  31373=>"11111111",
  31374=>"11111111",
  31375=>"00000001",
  31376=>"11111111",
  31377=>"00000000",
  31378=>"11111111",
  31379=>"11111110",
  31380=>"00000010",
  31381=>"11111101",
  31382=>"11111111",
  31383=>"00000001",
  31384=>"00000010",
  31385=>"00000000",
  31386=>"00000000",
  31387=>"00000001",
  31388=>"11111101",
  31389=>"11111111",
  31390=>"11111110",
  31391=>"00000111",
  31392=>"00000000",
  31393=>"00000010",
  31394=>"00000000",
  31395=>"00000010",
  31396=>"00000010",
  31397=>"00000010",
  31398=>"00000001",
  31399=>"00000010",
  31400=>"00000000",
  31401=>"00000010",
  31402=>"00000011",
  31403=>"11111111",
  31404=>"00000010",
  31405=>"00000001",
  31406=>"11111110",
  31407=>"11111111",
  31408=>"11111111",
  31409=>"11111110",
  31410=>"00000000",
  31411=>"11111110",
  31412=>"00000001",
  31413=>"00000001",
  31414=>"11111111",
  31415=>"11111101",
  31416=>"11111110",
  31417=>"00000011",
  31418=>"00000010",
  31419=>"11111111",
  31420=>"11111111",
  31421=>"11111110",
  31422=>"11111110",
  31423=>"11111101",
  31424=>"11111101",
  31425=>"11111111",
  31426=>"11111100",
  31427=>"11111101",
  31428=>"11111110",
  31429=>"00000000",
  31430=>"00000010",
  31431=>"00000010",
  31432=>"11111101",
  31433=>"11111111",
  31434=>"11111101",
  31435=>"11111100",
  31436=>"00000111",
  31437=>"11111101",
  31438=>"00000000",
  31439=>"00000000",
  31440=>"00000000",
  31441=>"11111101",
  31442=>"11111111",
  31443=>"11111110",
  31444=>"00000001",
  31445=>"00000010",
  31446=>"11111111",
  31447=>"00001000",
  31448=>"00000011",
  31449=>"11111110",
  31450=>"11111110",
  31451=>"11111111",
  31452=>"00000011",
  31453=>"00000000",
  31454=>"11111111",
  31455=>"00000001",
  31456=>"11111101",
  31457=>"11111111",
  31458=>"11111111",
  31459=>"11111110",
  31460=>"00000011",
  31461=>"00000000",
  31462=>"11111100",
  31463=>"00000101",
  31464=>"00000010",
  31465=>"11111110",
  31466=>"11111110",
  31467=>"00000010",
  31468=>"11111111",
  31469=>"11111111",
  31470=>"11111110",
  31471=>"00000101",
  31472=>"00000000",
  31473=>"00000001",
  31474=>"11111110",
  31475=>"11111111",
  31476=>"00000000",
  31477=>"00000001",
  31478=>"11111111",
  31479=>"00000000",
  31480=>"00000001",
  31481=>"00000010",
  31482=>"00000001",
  31483=>"00000010",
  31484=>"11111110",
  31485=>"11111110",
  31486=>"11111101",
  31487=>"11111110",
  31488=>"00000000",
  31489=>"00000001",
  31490=>"00000000",
  31491=>"00000000",
  31492=>"11111110",
  31493=>"00000010",
  31494=>"11111110",
  31495=>"11111101",
  31496=>"00000001",
  31497=>"11111111",
  31498=>"00000001",
  31499=>"11111110",
  31500=>"00000011",
  31501=>"00000011",
  31502=>"00000000",
  31503=>"11111110",
  31504=>"00000000",
  31505=>"11111111",
  31506=>"00000000",
  31507=>"11111110",
  31508=>"00000011",
  31509=>"00000010",
  31510=>"00000001",
  31511=>"00000010",
  31512=>"00000000",
  31513=>"00000000",
  31514=>"00000000",
  31515=>"00000001",
  31516=>"00000000",
  31517=>"11111110",
  31518=>"11111100",
  31519=>"11111101",
  31520=>"11111101",
  31521=>"00000001",
  31522=>"11111111",
  31523=>"11111111",
  31524=>"11111111",
  31525=>"00000011",
  31526=>"11111111",
  31527=>"11111110",
  31528=>"00000010",
  31529=>"11111111",
  31530=>"00000010",
  31531=>"00000000",
  31532=>"11111110",
  31533=>"00000001",
  31534=>"00000100",
  31535=>"00000001",
  31536=>"11111110",
  31537=>"00000000",
  31538=>"11111100",
  31539=>"11111101",
  31540=>"00000000",
  31541=>"00000010",
  31542=>"11111110",
  31543=>"11111100",
  31544=>"11111110",
  31545=>"00000000",
  31546=>"00000001",
  31547=>"00000010",
  31548=>"00000010",
  31549=>"00000001",
  31550=>"00000010",
  31551=>"11111101",
  31552=>"00000000",
  31553=>"11111101",
  31554=>"00000000",
  31555=>"11111101",
  31556=>"00000001",
  31557=>"00000100",
  31558=>"11111111",
  31559=>"00000000",
  31560=>"11111101",
  31561=>"11111110",
  31562=>"11111111",
  31563=>"11111111",
  31564=>"11111101",
  31565=>"11111111",
  31566=>"11111110",
  31567=>"11111111",
  31568=>"00000011",
  31569=>"11111110",
  31570=>"00000001",
  31571=>"11111111",
  31572=>"00000011",
  31573=>"00000100",
  31574=>"00000000",
  31575=>"11111101",
  31576=>"00000000",
  31577=>"11111111",
  31578=>"00000011",
  31579=>"11111110",
  31580=>"11111110",
  31581=>"00000001",
  31582=>"11111110",
  31583=>"00000010",
  31584=>"11111101",
  31585=>"00000010",
  31586=>"11111101",
  31587=>"00000100",
  31588=>"00000001",
  31589=>"00000001",
  31590=>"00000000",
  31591=>"00000100",
  31592=>"00000001",
  31593=>"00000010",
  31594=>"11111111",
  31595=>"00000001",
  31596=>"11111110",
  31597=>"00000011",
  31598=>"11111101",
  31599=>"11111110",
  31600=>"00000001",
  31601=>"00000011",
  31602=>"00000001",
  31603=>"00000001",
  31604=>"00000000",
  31605=>"11111111",
  31606=>"00000010",
  31607=>"00000011",
  31608=>"00000011",
  31609=>"00000001",
  31610=>"11111111",
  31611=>"11111111",
  31612=>"00000000",
  31613=>"00000001",
  31614=>"11111101",
  31615=>"00000000",
  31616=>"11111111",
  31617=>"11111110",
  31618=>"11111111",
  31619=>"11111101",
  31620=>"00000010",
  31621=>"00000001",
  31622=>"11111110",
  31623=>"00000000",
  31624=>"00000011",
  31625=>"11111111",
  31626=>"11111111",
  31627=>"11111100",
  31628=>"00000010",
  31629=>"11111111",
  31630=>"11111110",
  31631=>"00000000",
  31632=>"11111110",
  31633=>"11111110",
  31634=>"11111110",
  31635=>"00000010",
  31636=>"00000000",
  31637=>"00000010",
  31638=>"00000001",
  31639=>"11111111",
  31640=>"00000011",
  31641=>"11111101",
  31642=>"00000000",
  31643=>"11111101",
  31644=>"00000000",
  31645=>"00000000",
  31646=>"00000001",
  31647=>"11111101",
  31648=>"00000010",
  31649=>"11111101",
  31650=>"11111110",
  31651=>"00000000",
  31652=>"00000010",
  31653=>"00000000",
  31654=>"11111101",
  31655=>"00000001",
  31656=>"00000010",
  31657=>"11111110",
  31658=>"00000010",
  31659=>"00000010",
  31660=>"00000010",
  31661=>"11111110",
  31662=>"11111111",
  31663=>"00000011",
  31664=>"11111111",
  31665=>"11111111",
  31666=>"00000001",
  31667=>"11111101",
  31668=>"00000000",
  31669=>"00000000",
  31670=>"11111111",
  31671=>"11111110",
  31672=>"00000001",
  31673=>"11111110",
  31674=>"11111110",
  31675=>"11111111",
  31676=>"00000001",
  31677=>"00000111",
  31678=>"11111111",
  31679=>"00000000",
  31680=>"11111101",
  31681=>"00000010",
  31682=>"11111110",
  31683=>"00000011",
  31684=>"11111111",
  31685=>"11111111",
  31686=>"00000101",
  31687=>"11111110",
  31688=>"00000001",
  31689=>"00000000",
  31690=>"00000011",
  31691=>"11111111",
  31692=>"00000001",
  31693=>"11111110",
  31694=>"11111111",
  31695=>"11111110",
  31696=>"00000010",
  31697=>"11111110",
  31698=>"11111101",
  31699=>"11111111",
  31700=>"00000001",
  31701=>"00000001",
  31702=>"11111110",
  31703=>"11111111",
  31704=>"00000001",
  31705=>"00000100",
  31706=>"00000000",
  31707=>"11111111",
  31708=>"00000001",
  31709=>"11111110",
  31710=>"11111100",
  31711=>"11111111",
  31712=>"00000010",
  31713=>"11111110",
  31714=>"11111111",
  31715=>"11111110",
  31716=>"00000000",
  31717=>"11111101",
  31718=>"11111110",
  31719=>"11111110",
  31720=>"00000001",
  31721=>"11111111",
  31722=>"00000100",
  31723=>"11111111",
  31724=>"00000010",
  31725=>"11111110",
  31726=>"11111111",
  31727=>"11111111",
  31728=>"00000010",
  31729=>"00000000",
  31730=>"00000100",
  31731=>"11111110",
  31732=>"11111111",
  31733=>"11111100",
  31734=>"00000010",
  31735=>"00000001",
  31736=>"00000000",
  31737=>"11111110",
  31738=>"00000001",
  31739=>"11111101",
  31740=>"11111111",
  31741=>"00000001",
  31742=>"00000000",
  31743=>"11111110",
  31744=>"00000011",
  31745=>"11111110",
  31746=>"11111110",
  31747=>"11111111",
  31748=>"00000000",
  31749=>"00000100",
  31750=>"00000000",
  31751=>"11111101",
  31752=>"00000101",
  31753=>"11111111",
  31754=>"11111111",
  31755=>"00000001",
  31756=>"00000000",
  31757=>"00000100",
  31758=>"00000000",
  31759=>"00000011",
  31760=>"00000001",
  31761=>"00000010",
  31762=>"00000110",
  31763=>"11111101",
  31764=>"11111111",
  31765=>"11111111",
  31766=>"11111101",
  31767=>"11111111",
  31768=>"00000001",
  31769=>"11111111",
  31770=>"00000001",
  31771=>"00000101",
  31772=>"00000000",
  31773=>"11111110",
  31774=>"00000100",
  31775=>"11111111",
  31776=>"11111101",
  31777=>"00000011",
  31778=>"00000011",
  31779=>"00000001",
  31780=>"11111101",
  31781=>"00000010",
  31782=>"00000001",
  31783=>"00000011",
  31784=>"11111100",
  31785=>"00000110",
  31786=>"11111111",
  31787=>"00000100",
  31788=>"00000100",
  31789=>"00000000",
  31790=>"00000000",
  31791=>"00000000",
  31792=>"11111101",
  31793=>"00000000",
  31794=>"00000010",
  31795=>"00000010",
  31796=>"11111110",
  31797=>"11111111",
  31798=>"00000001",
  31799=>"00000000",
  31800=>"11111110",
  31801=>"00000000",
  31802=>"00000001",
  31803=>"00000010",
  31804=>"11111101",
  31805=>"11111111",
  31806=>"00000010",
  31807=>"11111111",
  31808=>"00000010",
  31809=>"00000001",
  31810=>"00000011",
  31811=>"00000000",
  31812=>"11111110",
  31813=>"11111111",
  31814=>"00000100",
  31815=>"11111110",
  31816=>"11111110",
  31817=>"11111111",
  31818=>"11111110",
  31819=>"11111111",
  31820=>"00000001",
  31821=>"00000010",
  31822=>"00000010",
  31823=>"00000001",
  31824=>"11111111",
  31825=>"00000010",
  31826=>"11111111",
  31827=>"00000000",
  31828=>"11111100",
  31829=>"11111101",
  31830=>"11111111",
  31831=>"11111111",
  31832=>"11111111",
  31833=>"00000010",
  31834=>"11111110",
  31835=>"00000010",
  31836=>"11111100",
  31837=>"00000011",
  31838=>"11111100",
  31839=>"00000100",
  31840=>"11111111",
  31841=>"00000100",
  31842=>"00000010",
  31843=>"00000001",
  31844=>"11111110",
  31845=>"11111110",
  31846=>"11111101",
  31847=>"00000010",
  31848=>"00000000",
  31849=>"11111110",
  31850=>"00000011",
  31851=>"11111111",
  31852=>"11111111",
  31853=>"00000010",
  31854=>"11111111",
  31855=>"11111111",
  31856=>"11111101",
  31857=>"11111111",
  31858=>"11111111",
  31859=>"11111111",
  31860=>"00000010",
  31861=>"11111111",
  31862=>"00000011",
  31863=>"11111110",
  31864=>"11111100",
  31865=>"00000000",
  31866=>"00000010",
  31867=>"11111110",
  31868=>"11111100",
  31869=>"00000011",
  31870=>"11111101",
  31871=>"00000001",
  31872=>"00000011",
  31873=>"00000010",
  31874=>"11111101",
  31875=>"11111110",
  31876=>"11111110",
  31877=>"11111111",
  31878=>"00000000",
  31879=>"00000011",
  31880=>"00000011",
  31881=>"11111111",
  31882=>"11111110",
  31883=>"00000010",
  31884=>"11111101",
  31885=>"11111101",
  31886=>"11111111",
  31887=>"00000001",
  31888=>"00000010",
  31889=>"00000100",
  31890=>"00000010",
  31891=>"00000001",
  31892=>"00000110",
  31893=>"00000011",
  31894=>"00000001",
  31895=>"00000010",
  31896=>"00000100",
  31897=>"00000010",
  31898=>"11111110",
  31899=>"00000010",
  31900=>"00000000",
  31901=>"11111111",
  31902=>"00000000",
  31903=>"11111101",
  31904=>"00000001",
  31905=>"00000000",
  31906=>"00000000",
  31907=>"00000101",
  31908=>"00000010",
  31909=>"11111101",
  31910=>"00000000",
  31911=>"00000000",
  31912=>"11111111",
  31913=>"00000110",
  31914=>"11111110",
  31915=>"00000011",
  31916=>"11111111",
  31917=>"00000000",
  31918=>"00000011",
  31919=>"11111110",
  31920=>"00000011",
  31921=>"00000100",
  31922=>"00000000",
  31923=>"00000001",
  31924=>"00000001",
  31925=>"00000011",
  31926=>"00000000",
  31927=>"11111110",
  31928=>"11111110",
  31929=>"00000101",
  31930=>"11111110",
  31931=>"00000010",
  31932=>"00001000",
  31933=>"00000000",
  31934=>"11111110",
  31935=>"00000001",
  31936=>"11111110",
  31937=>"11111111",
  31938=>"00000000",
  31939=>"11111111",
  31940=>"00000001",
  31941=>"11111111",
  31942=>"00000001",
  31943=>"11111110",
  31944=>"11111111",
  31945=>"00000101",
  31946=>"00000011",
  31947=>"00000010",
  31948=>"00000000",
  31949=>"00000010",
  31950=>"00000001",
  31951=>"00000000",
  31952=>"00000011",
  31953=>"00000001",
  31954=>"11111110",
  31955=>"11111101",
  31956=>"11111101",
  31957=>"00000010",
  31958=>"00000000",
  31959=>"11111110",
  31960=>"00000001",
  31961=>"00000000",
  31962=>"00000010",
  31963=>"00000000",
  31964=>"11111101",
  31965=>"00000100",
  31966=>"11111110",
  31967=>"00000000",
  31968=>"00000000",
  31969=>"00000011",
  31970=>"11111111",
  31971=>"11111111",
  31972=>"11111110",
  31973=>"11111101",
  31974=>"00000000",
  31975=>"00000000",
  31976=>"00000010",
  31977=>"00000010",
  31978=>"11111110",
  31979=>"11111111",
  31980=>"11111110",
  31981=>"11111110",
  31982=>"00000001",
  31983=>"11111101",
  31984=>"00000001",
  31985=>"00000011",
  31986=>"11111110",
  31987=>"00000000",
  31988=>"00000001",
  31989=>"00000001",
  31990=>"00000010",
  31991=>"11111111",
  31992=>"11111110",
  31993=>"00000000",
  31994=>"11111110",
  31995=>"00000001",
  31996=>"11111111",
  31997=>"11111110",
  31998=>"00000101",
  31999=>"11111100",
  32000=>"11111110",
  32001=>"00000010",
  32002=>"11111100",
  32003=>"00000000",
  32004=>"11111111",
  32005=>"00000011",
  32006=>"11111100",
  32007=>"11111101",
  32008=>"11111110",
  32009=>"00000001",
  32010=>"00000000",
  32011=>"11111110",
  32012=>"11111111",
  32013=>"11111101",
  32014=>"00000000",
  32015=>"11111100",
  32016=>"11111111",
  32017=>"00000011",
  32018=>"00000000",
  32019=>"11111100",
  32020=>"00000010",
  32021=>"00000000",
  32022=>"00000001",
  32023=>"11111100",
  32024=>"11111100",
  32025=>"00000010",
  32026=>"00000001",
  32027=>"00000000",
  32028=>"11111100",
  32029=>"11111111",
  32030=>"00000010",
  32031=>"00000001",
  32032=>"00000100",
  32033=>"00000011",
  32034=>"00000000",
  32035=>"00000000",
  32036=>"00000100",
  32037=>"00000100",
  32038=>"00000010",
  32039=>"00000110",
  32040=>"11111110",
  32041=>"11111110",
  32042=>"11111111",
  32043=>"00000010",
  32044=>"00000001",
  32045=>"11111111",
  32046=>"00000010",
  32047=>"00000000",
  32048=>"11111110",
  32049=>"00000001",
  32050=>"00000001",
  32051=>"00000011",
  32052=>"00000010",
  32053=>"00000010",
  32054=>"11111110",
  32055=>"00000010",
  32056=>"11111110",
  32057=>"00000011",
  32058=>"00000000",
  32059=>"11111111",
  32060=>"11111111",
  32061=>"11111101",
  32062=>"00000001",
  32063=>"11111110",
  32064=>"00000010",
  32065=>"11111111",
  32066=>"00000000",
  32067=>"00000000",
  32068=>"11111111",
  32069=>"11111110",
  32070=>"11111101",
  32071=>"00000000",
  32072=>"00000001",
  32073=>"11111110",
  32074=>"11111110",
  32075=>"11111101",
  32076=>"00000011",
  32077=>"11111100",
  32078=>"00000011",
  32079=>"00000010",
  32080=>"11111111",
  32081=>"00000010",
  32082=>"00000001",
  32083=>"00000000",
  32084=>"11111101",
  32085=>"00000010",
  32086=>"11111101",
  32087=>"11111101",
  32088=>"11111101",
  32089=>"00000010",
  32090=>"00000001",
  32091=>"00000011",
  32092=>"00000011",
  32093=>"11111111",
  32094=>"11111101",
  32095=>"00000001",
  32096=>"00000100",
  32097=>"00000100",
  32098=>"00000000",
  32099=>"11111111",
  32100=>"00000010",
  32101=>"11111101",
  32102=>"00000110",
  32103=>"11111111",
  32104=>"11111111",
  32105=>"11111101",
  32106=>"00000000",
  32107=>"00000001",
  32108=>"11111111",
  32109=>"00000001",
  32110=>"11111110",
  32111=>"00000001",
  32112=>"11111101",
  32113=>"00000010",
  32114=>"11111100",
  32115=>"00000000",
  32116=>"00000001",
  32117=>"11111111",
  32118=>"00000000",
  32119=>"00000010",
  32120=>"11111101",
  32121=>"11111111",
  32122=>"00000110",
  32123=>"00000101",
  32124=>"00000000",
  32125=>"00000010",
  32126=>"00000001",
  32127=>"00000000",
  32128=>"11111110",
  32129=>"00000000",
  32130=>"00000010",
  32131=>"11111111",
  32132=>"11111110",
  32133=>"00000010",
  32134=>"00000000",
  32135=>"11111111",
  32136=>"00000000",
  32137=>"11111110",
  32138=>"00000010",
  32139=>"00000010",
  32140=>"00000001",
  32141=>"11111101",
  32142=>"00000001",
  32143=>"00000011",
  32144=>"11111101",
  32145=>"00000000",
  32146=>"11111011",
  32147=>"11111110",
  32148=>"00000101",
  32149=>"00000000",
  32150=>"11111110",
  32151=>"11111110",
  32152=>"00000011",
  32153=>"00000010",
  32154=>"00000100",
  32155=>"11111111",
  32156=>"11111111",
  32157=>"11111111",
  32158=>"00000011",
  32159=>"00000010",
  32160=>"00000010",
  32161=>"00000000",
  32162=>"00000101",
  32163=>"00000100",
  32164=>"00000011",
  32165=>"00000010",
  32166=>"11111110",
  32167=>"00000011",
  32168=>"00000100",
  32169=>"11111110",
  32170=>"00000010",
  32171=>"00000001",
  32172=>"11111111",
  32173=>"11111101",
  32174=>"00000011",
  32175=>"00000011",
  32176=>"00000101",
  32177=>"00000000",
  32178=>"00000010",
  32179=>"00000100",
  32180=>"11111110",
  32181=>"11111110",
  32182=>"00000010",
  32183=>"00000110",
  32184=>"11111100",
  32185=>"00000010",
  32186=>"11111111",
  32187=>"00000001",
  32188=>"11111111",
  32189=>"00000011",
  32190=>"11111111",
  32191=>"11111110",
  32192=>"00000000",
  32193=>"11111110",
  32194=>"00000000",
  32195=>"11111101",
  32196=>"11111101",
  32197=>"00000000",
  32198=>"00000010",
  32199=>"11111111",
  32200=>"00000001",
  32201=>"00000000",
  32202=>"00000010",
  32203=>"00000011",
  32204=>"00000100",
  32205=>"11111110",
  32206=>"11111110",
  32207=>"00000001",
  32208=>"00000010",
  32209=>"11111110",
  32210=>"00000000",
  32211=>"11111101",
  32212=>"00000100",
  32213=>"11111100",
  32214=>"11111101",
  32215=>"00000001",
  32216=>"11111101",
  32217=>"00000000",
  32218=>"00000000",
  32219=>"00000010",
  32220=>"11111111",
  32221=>"00000011",
  32222=>"00000001",
  32223=>"00000000",
  32224=>"11111100",
  32225=>"00000001",
  32226=>"00000011",
  32227=>"11111110",
  32228=>"00000010",
  32229=>"00000011",
  32230=>"11111111",
  32231=>"11111111",
  32232=>"00000010",
  32233=>"11111101",
  32234=>"11111110",
  32235=>"11111110",
  32236=>"11111101",
  32237=>"00000000",
  32238=>"00000010",
  32239=>"11111101",
  32240=>"11111101",
  32241=>"00000000",
  32242=>"11111111",
  32243=>"00000011",
  32244=>"00000001",
  32245=>"00000011",
  32246=>"00000001",
  32247=>"00000000",
  32248=>"11111101",
  32249=>"11111101",
  32250=>"00000000",
  32251=>"00000001",
  32252=>"00000010",
  32253=>"00000101",
  32254=>"11111110",
  32255=>"11111101",
  32256=>"00000000",
  32257=>"11111101",
  32258=>"11111111",
  32259=>"00000000",
  32260=>"11111110",
  32261=>"11111111",
  32262=>"00000110",
  32263=>"11111111",
  32264=>"11111111",
  32265=>"00000011",
  32266=>"00000001",
  32267=>"00000011",
  32268=>"00000001",
  32269=>"11111111",
  32270=>"11111100",
  32271=>"00000011",
  32272=>"00000010",
  32273=>"00000000",
  32274=>"11111110",
  32275=>"11111111",
  32276=>"00000000",
  32277=>"00000001",
  32278=>"11111110",
  32279=>"11111110",
  32280=>"00000011",
  32281=>"00000001",
  32282=>"00000100",
  32283=>"00000011",
  32284=>"11111110",
  32285=>"11111101",
  32286=>"00000010",
  32287=>"00000011",
  32288=>"00000000",
  32289=>"11111111",
  32290=>"11111111",
  32291=>"00000001",
  32292=>"11111110",
  32293=>"00000010",
  32294=>"00000010",
  32295=>"00000001",
  32296=>"00000010",
  32297=>"11111110",
  32298=>"00000000",
  32299=>"00000010",
  32300=>"00000110",
  32301=>"00000010",
  32302=>"11111110",
  32303=>"00000100",
  32304=>"00000011",
  32305=>"00000000",
  32306=>"11111101",
  32307=>"00000011",
  32308=>"00000000",
  32309=>"00000000",
  32310=>"00000000",
  32311=>"11111111",
  32312=>"00000011",
  32313=>"11111111",
  32314=>"11111110",
  32315=>"11111110",
  32316=>"11111111",
  32317=>"11111111",
  32318=>"11111101",
  32319=>"00000000",
  32320=>"00000100",
  32321=>"00000000",
  32322=>"11111110",
  32323=>"00000010",
  32324=>"11111110",
  32325=>"00000010",
  32326=>"11111110",
  32327=>"11111111",
  32328=>"00000000",
  32329=>"00000011",
  32330=>"00000101",
  32331=>"00000001",
  32332=>"00000010",
  32333=>"11111110",
  32334=>"11111100",
  32335=>"11111111",
  32336=>"00000000",
  32337=>"11111110",
  32338=>"11111111",
  32339=>"00000010",
  32340=>"00000001",
  32341=>"00000001",
  32342=>"11111111",
  32343=>"00000001",
  32344=>"11111101",
  32345=>"00000000",
  32346=>"00000001",
  32347=>"11111111",
  32348=>"00000001",
  32349=>"00000011",
  32350=>"11111100",
  32351=>"11111111",
  32352=>"11111110",
  32353=>"11111101",
  32354=>"00000100",
  32355=>"00000000",
  32356=>"11111100",
  32357=>"11111110",
  32358=>"00000001",
  32359=>"00000010",
  32360=>"00000011",
  32361=>"00000000",
  32362=>"00000001",
  32363=>"00000011",
  32364=>"00000010",
  32365=>"00000000",
  32366=>"11111110",
  32367=>"11111101",
  32368=>"00000010",
  32369=>"00000001",
  32370=>"11111111",
  32371=>"00000100",
  32372=>"11111111",
  32373=>"00000000",
  32374=>"11111110",
  32375=>"00000001",
  32376=>"11111101",
  32377=>"00000100",
  32378=>"00000010",
  32379=>"00000101",
  32380=>"00000011",
  32381=>"11111101",
  32382=>"00000000",
  32383=>"11111101",
  32384=>"11111100",
  32385=>"11111110",
  32386=>"11111111",
  32387=>"11111110",
  32388=>"11111111",
  32389=>"00000101",
  32390=>"00000001",
  32391=>"11111111",
  32392=>"11111111",
  32393=>"11111110",
  32394=>"00000011",
  32395=>"11111110",
  32396=>"11111101",
  32397=>"11111111",
  32398=>"00000001",
  32399=>"11111100",
  32400=>"00000100",
  32401=>"00000001",
  32402=>"00000011",
  32403=>"00000000",
  32404=>"11111111",
  32405=>"00000011",
  32406=>"00000010",
  32407=>"00000000",
  32408=>"00000010",
  32409=>"00000100",
  32410=>"00000000",
  32411=>"00000000",
  32412=>"00000101",
  32413=>"00000100",
  32414=>"11111111",
  32415=>"11111101",
  32416=>"00000010",
  32417=>"00000000",
  32418=>"11111110",
  32419=>"00000001",
  32420=>"00000011",
  32421=>"00000100",
  32422=>"00000001",
  32423=>"11111110",
  32424=>"11111111",
  32425=>"11111101",
  32426=>"11111111",
  32427=>"00000000",
  32428=>"00000001",
  32429=>"00000010",
  32430=>"11111101",
  32431=>"11111111",
  32432=>"00000000",
  32433=>"00000011",
  32434=>"00000010",
  32435=>"00000001",
  32436=>"00000000",
  32437=>"00000001",
  32438=>"11111110",
  32439=>"11111111",
  32440=>"00000011",
  32441=>"00000010",
  32442=>"11111101",
  32443=>"00000000",
  32444=>"00000010",
  32445=>"00000010",
  32446=>"00000000",
  32447=>"11111111",
  32448=>"11111110",
  32449=>"11111011",
  32450=>"00000000",
  32451=>"11111110",
  32452=>"00000001",
  32453=>"00000010",
  32454=>"11111111",
  32455=>"11111100",
  32456=>"11111110",
  32457=>"00000010",
  32458=>"11111111",
  32459=>"00000000",
  32460=>"00000000",
  32461=>"11111111",
  32462=>"00000011",
  32463=>"00000010",
  32464=>"11111111",
  32465=>"00000010",
  32466=>"00000010",
  32467=>"11111110",
  32468=>"11111111",
  32469=>"00000010",
  32470=>"00000000",
  32471=>"11111100",
  32472=>"00000001",
  32473=>"00000000",
  32474=>"00000001",
  32475=>"11111110",
  32476=>"00000000",
  32477=>"00000000",
  32478=>"00000010",
  32479=>"00000010",
  32480=>"00000011",
  32481=>"11111111",
  32482=>"11111111",
  32483=>"11111111",
  32484=>"11111110",
  32485=>"00000011",
  32486=>"11111101",
  32487=>"11111111",
  32488=>"00000000",
  32489=>"11111111",
  32490=>"00000101",
  32491=>"00000001",
  32492=>"11111100",
  32493=>"00000001",
  32494=>"00000000",
  32495=>"00000000",
  32496=>"00000000",
  32497=>"11111111",
  32498=>"00000000",
  32499=>"11111101",
  32500=>"11111101",
  32501=>"11111110",
  32502=>"00000000",
  32503=>"11111100",
  32504=>"00000011",
  32505=>"00000110",
  32506=>"11111111",
  32507=>"00000111",
  32508=>"00000000",
  32509=>"11111101",
  32510=>"11111101",
  32511=>"00000100",
  32512=>"00000000",
  32513=>"00000000",
  32514=>"11111111",
  32515=>"00000001",
  32516=>"00000001",
  32517=>"00000000",
  32518=>"11111101",
  32519=>"00000100",
  32520=>"11111111",
  32521=>"00000110",
  32522=>"00000010",
  32523=>"00000000",
  32524=>"00000010",
  32525=>"00000000",
  32526=>"00000010",
  32527=>"11111110",
  32528=>"00000101",
  32529=>"11111110",
  32530=>"00000010",
  32531=>"11111111",
  32532=>"11111110",
  32533=>"11111111",
  32534=>"11111111",
  32535=>"00000100",
  32536=>"11111111",
  32537=>"00000000",
  32538=>"00000011",
  32539=>"11111101",
  32540=>"00000011",
  32541=>"00000100",
  32542=>"00000101",
  32543=>"11111111",
  32544=>"00000010",
  32545=>"11111110",
  32546=>"11111101",
  32547=>"11111111",
  32548=>"11111100",
  32549=>"11111101",
  32550=>"11111100",
  32551=>"11111111",
  32552=>"00000011",
  32553=>"00000110",
  32554=>"11111111",
  32555=>"00000001",
  32556=>"11111111",
  32557=>"00000001",
  32558=>"00000010",
  32559=>"11111110",
  32560=>"11111111",
  32561=>"11111111",
  32562=>"11111111",
  32563=>"11111111",
  32564=>"00000001",
  32565=>"00000001",
  32566=>"11111110",
  32567=>"00000000",
  32568=>"00000000",
  32569=>"11111101",
  32570=>"11111110",
  32571=>"11111011",
  32572=>"00000010",
  32573=>"11111111",
  32574=>"11111111",
  32575=>"00000010",
  32576=>"00000001",
  32577=>"00000010",
  32578=>"00000011",
  32579=>"00000010",
  32580=>"11111110",
  32581=>"00000010",
  32582=>"00000011",
  32583=>"00000000",
  32584=>"11111111",
  32585=>"11111111",
  32586=>"11111101",
  32587=>"11111100",
  32588=>"00000000",
  32589=>"00000100",
  32590=>"11111111",
  32591=>"00000010",
  32592=>"11111100",
  32593=>"00000001",
  32594=>"00000001",
  32595=>"00000011",
  32596=>"00000001",
  32597=>"00000010",
  32598=>"11111100",
  32599=>"00000101",
  32600=>"00000011",
  32601=>"11111111",
  32602=>"00000101",
  32603=>"00000010",
  32604=>"00000000",
  32605=>"11111101",
  32606=>"11111111",
  32607=>"11111101",
  32608=>"00000010",
  32609=>"11111111",
  32610=>"00000001",
  32611=>"11111100",
  32612=>"00000010",
  32613=>"00000001",
  32614=>"11111111",
  32615=>"00000000",
  32616=>"11111110",
  32617=>"00000001",
  32618=>"00000001",
  32619=>"00000001",
  32620=>"11111111",
  32621=>"00000101",
  32622=>"00000000",
  32623=>"00000000",
  32624=>"00000011",
  32625=>"11111111",
  32626=>"11111111",
  32627=>"00000000",
  32628=>"00000011",
  32629=>"11111111",
  32630=>"11111101",
  32631=>"00000001",
  32632=>"00000101",
  32633=>"11111110",
  32634=>"00000000",
  32635=>"00000010",
  32636=>"11111110",
  32637=>"11111101",
  32638=>"00000010",
  32639=>"00000011",
  32640=>"11111110",
  32641=>"11111101",
  32642=>"00000010",
  32643=>"00000001",
  32644=>"11111101",
  32645=>"00000000",
  32646=>"00000010",
  32647=>"11111101",
  32648=>"00000100",
  32649=>"00000000",
  32650=>"00000010",
  32651=>"11111110",
  32652=>"11111110",
  32653=>"00000000",
  32654=>"11111111",
  32655=>"00000010",
  32656=>"00000010",
  32657=>"11111110",
  32658=>"11111111",
  32659=>"00000000",
  32660=>"00000001",
  32661=>"00000001",
  32662=>"11111111",
  32663=>"00000001",
  32664=>"00000010",
  32665=>"11111110",
  32666=>"11111110",
  32667=>"11111101",
  32668=>"11111110",
  32669=>"00000000",
  32670=>"00000100",
  32671=>"00000000",
  32672=>"11111111",
  32673=>"00000010",
  32674=>"00000011",
  32675=>"11111110",
  32676=>"11111111",
  32677=>"00000000",
  32678=>"00000000",
  32679=>"11111110",
  32680=>"00000000",
  32681=>"00000000",
  32682=>"11111111",
  32683=>"00000001",
  32684=>"11111110",
  32685=>"11111111",
  32686=>"00000010",
  32687=>"00000001",
  32688=>"00000111",
  32689=>"11111110",
  32690=>"11111111",
  32691=>"11111111",
  32692=>"00000000",
  32693=>"11111100",
  32694=>"00000011",
  32695=>"00000010",
  32696=>"11111101",
  32697=>"11111100",
  32698=>"11111111",
  32699=>"11111111",
  32700=>"00000001",
  32701=>"00000000",
  32702=>"00000001",
  32703=>"00000001",
  32704=>"11111101",
  32705=>"00000000",
  32706=>"11111110",
  32707=>"00000001",
  32708=>"00000000",
  32709=>"00000000",
  32710=>"11111101",
  32711=>"11111111",
  32712=>"00000001",
  32713=>"00000001",
  32714=>"11111110",
  32715=>"00000011",
  32716=>"11111100",
  32717=>"11111100",
  32718=>"00000001",
  32719=>"00000011",
  32720=>"11111100",
  32721=>"11111111",
  32722=>"11111110",
  32723=>"00000010",
  32724=>"11111111",
  32725=>"11111101",
  32726=>"11111111",
  32727=>"11111110",
  32728=>"11111110",
  32729=>"00000001",
  32730=>"00000001",
  32731=>"00000001",
  32732=>"11111110",
  32733=>"00000000",
  32734=>"00000000",
  32735=>"00000001",
  32736=>"00000011",
  32737=>"00000000",
  32738=>"11111110",
  32739=>"11111111",
  32740=>"11111110",
  32741=>"11111110",
  32742=>"00000001",
  32743=>"11111100",
  32744=>"00000000",
  32745=>"00000000",
  32746=>"11111100",
  32747=>"00000011",
  32748=>"00000001",
  32749=>"00000010",
  32750=>"00000010",
  32751=>"11111110",
  32752=>"00000111",
  32753=>"00000001",
  32754=>"11111101",
  32755=>"00000000",
  32756=>"00000001",
  32757=>"11111110",
  32758=>"00000010",
  32759=>"00000100",
  32760=>"11111111",
  32761=>"11111111",
  32762=>"00000001",
  32763=>"11111111",
  32764=>"00000110",
  32765=>"11111111",
  32766=>"00000010",
  32767=>"00000000",
  32768=>"00000011",
  32769=>"00000010",
  32770=>"00000010",
  32771=>"11111110",
  32772=>"11111111",
  32773=>"11111110",
  32774=>"11111111",
  32775=>"11111111",
  32776=>"11111110",
  32777=>"11111110",
  32778=>"00000011",
  32779=>"11111110",
  32780=>"00000011",
  32781=>"00000010",
  32782=>"11111101",
  32783=>"00000010",
  32784=>"11111110",
  32785=>"11111111",
  32786=>"00000010",
  32787=>"00000011",
  32788=>"00000010",
  32789=>"00000100",
  32790=>"00000001",
  32791=>"00000010",
  32792=>"11111111",
  32793=>"11111111",
  32794=>"11111101",
  32795=>"00000011",
  32796=>"00000001",
  32797=>"00000010",
  32798=>"11111111",
  32799=>"00000001",
  32800=>"00000001",
  32801=>"11111110",
  32802=>"00000010",
  32803=>"11111101",
  32804=>"00000000",
  32805=>"11111111",
  32806=>"11111110",
  32807=>"00000000",
  32808=>"11111110",
  32809=>"11111101",
  32810=>"00000001",
  32811=>"00000001",
  32812=>"00000000",
  32813=>"00000001",
  32814=>"11111111",
  32815=>"00000001",
  32816=>"00000011",
  32817=>"00000000",
  32818=>"00000001",
  32819=>"11111111",
  32820=>"11111111",
  32821=>"11111111",
  32822=>"11111111",
  32823=>"00000001",
  32824=>"00000010",
  32825=>"11111110",
  32826=>"00000000",
  32827=>"00000011",
  32828=>"11111101",
  32829=>"00000010",
  32830=>"11111111",
  32831=>"00000010",
  32832=>"11111111",
  32833=>"11111110",
  32834=>"00000010",
  32835=>"00000000",
  32836=>"11111111",
  32837=>"11111101",
  32838=>"11111101",
  32839=>"00000010",
  32840=>"11111110",
  32841=>"00000001",
  32842=>"00000010",
  32843=>"00000001",
  32844=>"00000010",
  32845=>"11111111",
  32846=>"00000000",
  32847=>"00000000",
  32848=>"00000010",
  32849=>"11111111",
  32850=>"00000010",
  32851=>"11111110",
  32852=>"00000000",
  32853=>"11111101",
  32854=>"00000010",
  32855=>"00000000",
  32856=>"11111111",
  32857=>"00000000",
  32858=>"11111101",
  32859=>"00000001",
  32860=>"11111111",
  32861=>"00000000",
  32862=>"00000001",
  32863=>"00000000",
  32864=>"00000011",
  32865=>"11111111",
  32866=>"00000011",
  32867=>"00000010",
  32868=>"11111111",
  32869=>"11111101",
  32870=>"11111111",
  32871=>"00000001",
  32872=>"00000001",
  32873=>"11111111",
  32874=>"11111110",
  32875=>"00000000",
  32876=>"00000001",
  32877=>"00000001",
  32878=>"00000001",
  32879=>"11111111",
  32880=>"00000010",
  32881=>"00000010",
  32882=>"00000010",
  32883=>"11111111",
  32884=>"00000100",
  32885=>"11111110",
  32886=>"00000001",
  32887=>"11111111",
  32888=>"00000000",
  32889=>"00000101",
  32890=>"00000010",
  32891=>"00000010",
  32892=>"11111111",
  32893=>"11111111",
  32894=>"11111111",
  32895=>"00000001",
  32896=>"00000010",
  32897=>"11111111",
  32898=>"00000010",
  32899=>"00000001",
  32900=>"11111110",
  32901=>"11111111",
  32902=>"11111111",
  32903=>"11111101",
  32904=>"00000010",
  32905=>"00000000",
  32906=>"11111111",
  32907=>"00000000",
  32908=>"00000000",
  32909=>"11111111",
  32910=>"00000001",
  32911=>"11111110",
  32912=>"00000010",
  32913=>"00000000",
  32914=>"00000001",
  32915=>"00000010",
  32916=>"00000001",
  32917=>"11111110",
  32918=>"11111111",
  32919=>"11111110",
  32920=>"11111110",
  32921=>"11111110",
  32922=>"11111110",
  32923=>"00000000",
  32924=>"00000000",
  32925=>"11111111",
  32926=>"00000000",
  32927=>"11111101",
  32928=>"00000001",
  32929=>"11111111",
  32930=>"00000100",
  32931=>"11111110",
  32932=>"00000001",
  32933=>"11111111",
  32934=>"11111111",
  32935=>"11111111",
  32936=>"00000110",
  32937=>"00000010",
  32938=>"00000001",
  32939=>"11111110",
  32940=>"11111110",
  32941=>"00000001",
  32942=>"11111110",
  32943=>"11111101",
  32944=>"00000011",
  32945=>"00000001",
  32946=>"00000100",
  32947=>"11111111",
  32948=>"11111101",
  32949=>"11111110",
  32950=>"11111111",
  32951=>"11111111",
  32952=>"11111111",
  32953=>"00000000",
  32954=>"11111101",
  32955=>"00000010",
  32956=>"00000010",
  32957=>"00000001",
  32958=>"00000010",
  32959=>"00000000",
  32960=>"00000010",
  32961=>"00000010",
  32962=>"00000100",
  32963=>"11111111",
  32964=>"11111111",
  32965=>"11111110",
  32966=>"00000001",
  32967=>"11111110",
  32968=>"00000010",
  32969=>"00000001",
  32970=>"00000010",
  32971=>"11111101",
  32972=>"11111111",
  32973=>"00000001",
  32974=>"11111110",
  32975=>"11111110",
  32976=>"00000000",
  32977=>"11111101",
  32978=>"00000000",
  32979=>"00000001",
  32980=>"00000000",
  32981=>"00000010",
  32982=>"00000010",
  32983=>"00000000",
  32984=>"11111111",
  32985=>"11111110",
  32986=>"00000000",
  32987=>"11111111",
  32988=>"00000001",
  32989=>"11111111",
  32990=>"11111110",
  32991=>"00000010",
  32992=>"11111111",
  32993=>"11111110",
  32994=>"11111110",
  32995=>"00000001",
  32996=>"11111110",
  32997=>"00000011",
  32998=>"00000010",
  32999=>"11111110",
  33000=>"00000000",
  33001=>"11111111",
  33002=>"11111110",
  33003=>"00000010",
  33004=>"00000001",
  33005=>"11111111",
  33006=>"00000010",
  33007=>"11111111",
  33008=>"00000000",
  33009=>"11111111",
  33010=>"00000010",
  33011=>"00000000",
  33012=>"11111111",
  33013=>"00000000",
  33014=>"11111110",
  33015=>"00000001",
  33016=>"00000001",
  33017=>"00000001",
  33018=>"11111101",
  33019=>"00000000",
  33020=>"11111101",
  33021=>"11111111",
  33022=>"11111101",
  33023=>"00000001",
  33024=>"00000000",
  33025=>"11111111",
  33026=>"11111101",
  33027=>"00000001",
  33028=>"11111110",
  33029=>"00000001",
  33030=>"00000010",
  33031=>"00000010",
  33032=>"11111101",
  33033=>"11111101",
  33034=>"00000001",
  33035=>"00000100",
  33036=>"00000000",
  33037=>"00000001",
  33038=>"11111101",
  33039=>"00000010",
  33040=>"11111101",
  33041=>"00000010",
  33042=>"00000001",
  33043=>"11111110",
  33044=>"00000000",
  33045=>"00000001",
  33046=>"11111110",
  33047=>"11111110",
  33048=>"00000000",
  33049=>"11111111",
  33050=>"00000001",
  33051=>"00000010",
  33052=>"00000000",
  33053=>"00000001",
  33054=>"11111111",
  33055=>"11111110",
  33056=>"00000011",
  33057=>"00000000",
  33058=>"00000010",
  33059=>"11111110",
  33060=>"11111101",
  33061=>"00000001",
  33062=>"11111101",
  33063=>"11111110",
  33064=>"00000010",
  33065=>"00000010",
  33066=>"11111101",
  33067=>"00000000",
  33068=>"00000000",
  33069=>"11111110",
  33070=>"11111111",
  33071=>"11111111",
  33072=>"00000001",
  33073=>"00000100",
  33074=>"00000001",
  33075=>"11111111",
  33076=>"00000010",
  33077=>"11111101",
  33078=>"00000000",
  33079=>"00000000",
  33080=>"11111111",
  33081=>"11111111",
  33082=>"11111110",
  33083=>"11111101",
  33084=>"11111110",
  33085=>"11111111",
  33086=>"11111111",
  33087=>"11111110",
  33088=>"00000001",
  33089=>"11111101",
  33090=>"11111110",
  33091=>"00000100",
  33092=>"00000010",
  33093=>"11111110",
  33094=>"11111100",
  33095=>"00000101",
  33096=>"00000000",
  33097=>"11111101",
  33098=>"11111111",
  33099=>"00000000",
  33100=>"11111110",
  33101=>"00000001",
  33102=>"00000011",
  33103=>"00000011",
  33104=>"00000011",
  33105=>"00000010",
  33106=>"11111110",
  33107=>"11111111",
  33108=>"00000010",
  33109=>"00000001",
  33110=>"00000100",
  33111=>"11111110",
  33112=>"11111101",
  33113=>"00000100",
  33114=>"11111111",
  33115=>"11111111",
  33116=>"11111111",
  33117=>"00000000",
  33118=>"11111111",
  33119=>"11111101",
  33120=>"00000001",
  33121=>"00000000",
  33122=>"00000010",
  33123=>"00000011",
  33124=>"00000011",
  33125=>"00000011",
  33126=>"11111111",
  33127=>"11111110",
  33128=>"11111101",
  33129=>"11111110",
  33130=>"00000000",
  33131=>"11111110",
  33132=>"00000010",
  33133=>"11111111",
  33134=>"11111101",
  33135=>"00000000",
  33136=>"11111111",
  33137=>"11111111",
  33138=>"11111110",
  33139=>"11111111",
  33140=>"11111111",
  33141=>"00000011",
  33142=>"11111111",
  33143=>"11111111",
  33144=>"00000100",
  33145=>"00000000",
  33146=>"00000101",
  33147=>"11111110",
  33148=>"11111111",
  33149=>"11111101",
  33150=>"11111111",
  33151=>"00000010",
  33152=>"00000001",
  33153=>"11111110",
  33154=>"00000001",
  33155=>"00000001",
  33156=>"11111110",
  33157=>"11111110",
  33158=>"00000010",
  33159=>"11111111",
  33160=>"11111111",
  33161=>"00000001",
  33162=>"00000000",
  33163=>"11111110",
  33164=>"00000001",
  33165=>"00000000",
  33166=>"00000001",
  33167=>"11111100",
  33168=>"00000010",
  33169=>"00000100",
  33170=>"11111110",
  33171=>"11111110",
  33172=>"00000001",
  33173=>"00000001",
  33174=>"00000001",
  33175=>"00000000",
  33176=>"11111110",
  33177=>"11111110",
  33178=>"00000100",
  33179=>"00000001",
  33180=>"11111110",
  33181=>"11111111",
  33182=>"00000000",
  33183=>"11111101",
  33184=>"11111111",
  33185=>"11111111",
  33186=>"00000010",
  33187=>"00000101",
  33188=>"00000000",
  33189=>"00000001",
  33190=>"00000011",
  33191=>"00000010",
  33192=>"00000000",
  33193=>"00000000",
  33194=>"00000011",
  33195=>"00000001",
  33196=>"00000010",
  33197=>"00000000",
  33198=>"11111111",
  33199=>"00000001",
  33200=>"11111111",
  33201=>"00000100",
  33202=>"11111101",
  33203=>"11111101",
  33204=>"11111111",
  33205=>"00000000",
  33206=>"00000000",
  33207=>"00000001",
  33208=>"00000010",
  33209=>"00000010",
  33210=>"11111111",
  33211=>"11111111",
  33212=>"00000001",
  33213=>"00000001",
  33214=>"11111101",
  33215=>"11111101",
  33216=>"11111101",
  33217=>"00000011",
  33218=>"00000000",
  33219=>"00000000",
  33220=>"00000000",
  33221=>"00000001",
  33222=>"11111111",
  33223=>"11111110",
  33224=>"11111101",
  33225=>"11111101",
  33226=>"00000001",
  33227=>"00000010",
  33228=>"00000000",
  33229=>"11111111",
  33230=>"00000001",
  33231=>"00000011",
  33232=>"00000100",
  33233=>"00000010",
  33234=>"11111110",
  33235=>"11111110",
  33236=>"11111111",
  33237=>"00000011",
  33238=>"11111101",
  33239=>"11111111",
  33240=>"11111111",
  33241=>"11111111",
  33242=>"00000000",
  33243=>"00000001",
  33244=>"11111110",
  33245=>"00000010",
  33246=>"00000011",
  33247=>"11111110",
  33248=>"00000100",
  33249=>"00000001",
  33250=>"00000011",
  33251=>"11111110",
  33252=>"11111110",
  33253=>"11111111",
  33254=>"11111111",
  33255=>"11111111",
  33256=>"11111110",
  33257=>"11111110",
  33258=>"11111110",
  33259=>"00000100",
  33260=>"11111110",
  33261=>"00000011",
  33262=>"00000001",
  33263=>"11111110",
  33264=>"00000010",
  33265=>"00000001",
  33266=>"00000000",
  33267=>"11111101",
  33268=>"00000000",
  33269=>"00000000",
  33270=>"00000000",
  33271=>"00000000",
  33272=>"00000010",
  33273=>"11111101",
  33274=>"00000000",
  33275=>"00000000",
  33276=>"00000001",
  33277=>"11111110",
  33278=>"00000000",
  33279=>"00000000",
  33280=>"00000010",
  33281=>"00000000",
  33282=>"00000000",
  33283=>"11111111",
  33284=>"00000000",
  33285=>"11111101",
  33286=>"00000000",
  33287=>"00000010",
  33288=>"11111110",
  33289=>"00000011",
  33290=>"00000000",
  33291=>"00000000",
  33292=>"00000000",
  33293=>"11111111",
  33294=>"00000000",
  33295=>"11111110",
  33296=>"11111101",
  33297=>"11111101",
  33298=>"11111111",
  33299=>"00000000",
  33300=>"00000000",
  33301=>"11111101",
  33302=>"11111110",
  33303=>"00000001",
  33304=>"11111101",
  33305=>"00000000",
  33306=>"00000001",
  33307=>"00000010",
  33308=>"00000010",
  33309=>"11111111",
  33310=>"11111111",
  33311=>"00000100",
  33312=>"00000010",
  33313=>"00000100",
  33314=>"00000100",
  33315=>"11111111",
  33316=>"00000011",
  33317=>"00000000",
  33318=>"11111110",
  33319=>"11111101",
  33320=>"11111101",
  33321=>"00000010",
  33322=>"00000010",
  33323=>"00000001",
  33324=>"00000011",
  33325=>"11111111",
  33326=>"00000011",
  33327=>"00000010",
  33328=>"11111110",
  33329=>"00000000",
  33330=>"00000000",
  33331=>"11111110",
  33332=>"11111111",
  33333=>"00000000",
  33334=>"00000000",
  33335=>"00000000",
  33336=>"11111110",
  33337=>"00000000",
  33338=>"11111111",
  33339=>"11111110",
  33340=>"00000010",
  33341=>"11111110",
  33342=>"00000100",
  33343=>"00000010",
  33344=>"11111111",
  33345=>"00000011",
  33346=>"00000000",
  33347=>"11111110",
  33348=>"11111111",
  33349=>"00000000",
  33350=>"11111111",
  33351=>"00000000",
  33352=>"11111110",
  33353=>"00000010",
  33354=>"11111110",
  33355=>"00000101",
  33356=>"11111110",
  33357=>"11111101",
  33358=>"00000101",
  33359=>"00000000",
  33360=>"00000000",
  33361=>"00000000",
  33362=>"11111111",
  33363=>"00000011",
  33364=>"11111110",
  33365=>"11111110",
  33366=>"00000000",
  33367=>"11111110",
  33368=>"00000000",
  33369=>"00000001",
  33370=>"00000000",
  33371=>"00000000",
  33372=>"11111110",
  33373=>"00000000",
  33374=>"00000001",
  33375=>"00000000",
  33376=>"00000000",
  33377=>"00000001",
  33378=>"00000001",
  33379=>"00000010",
  33380=>"11111110",
  33381=>"11111110",
  33382=>"11111111",
  33383=>"11111111",
  33384=>"11111110",
  33385=>"11111111",
  33386=>"00000000",
  33387=>"11111110",
  33388=>"00000000",
  33389=>"11111110",
  33390=>"00000001",
  33391=>"00000110",
  33392=>"00000000",
  33393=>"11111101",
  33394=>"00000010",
  33395=>"00000010",
  33396=>"11111111",
  33397=>"11111111",
  33398=>"00000111",
  33399=>"00000011",
  33400=>"11111101",
  33401=>"00000000",
  33402=>"11111110",
  33403=>"11111110",
  33404=>"00000010",
  33405=>"00000001",
  33406=>"00000000",
  33407=>"11111110",
  33408=>"00000000",
  33409=>"11111111",
  33410=>"11111101",
  33411=>"00000001",
  33412=>"00000010",
  33413=>"11111110",
  33414=>"11111101",
  33415=>"00000010",
  33416=>"00000100",
  33417=>"11111110",
  33418=>"00000011",
  33419=>"11111110",
  33420=>"00000001",
  33421=>"00000000",
  33422=>"11111101",
  33423=>"11111111",
  33424=>"00000000",
  33425=>"00000010",
  33426=>"11111101",
  33427=>"00000010",
  33428=>"00000000",
  33429=>"11111101",
  33430=>"11111111",
  33431=>"11111111",
  33432=>"11111111",
  33433=>"00000001",
  33434=>"00000000",
  33435=>"11111110",
  33436=>"00000001",
  33437=>"11111110",
  33438=>"00000000",
  33439=>"11111101",
  33440=>"00000001",
  33441=>"00000001",
  33442=>"00000001",
  33443=>"11111111",
  33444=>"00000010",
  33445=>"00000001",
  33446=>"11111110",
  33447=>"00000000",
  33448=>"11111110",
  33449=>"00000001",
  33450=>"00000000",
  33451=>"00000010",
  33452=>"00000010",
  33453=>"00000010",
  33454=>"11111110",
  33455=>"11111111",
  33456=>"00000000",
  33457=>"11111111",
  33458=>"00000011",
  33459=>"00000010",
  33460=>"11111110",
  33461=>"00000000",
  33462=>"11111110",
  33463=>"00000000",
  33464=>"11111111",
  33465=>"00000010",
  33466=>"00000011",
  33467=>"00000010",
  33468=>"00000010",
  33469=>"11111110",
  33470=>"11111110",
  33471=>"00000001",
  33472=>"00000010",
  33473=>"00000001",
  33474=>"00000010",
  33475=>"00000001",
  33476=>"00000000",
  33477=>"00000101",
  33478=>"11111111",
  33479=>"00000001",
  33480=>"00000011",
  33481=>"11111101",
  33482=>"11111111",
  33483=>"11111111",
  33484=>"00000001",
  33485=>"00000010",
  33486=>"00000010",
  33487=>"11111111",
  33488=>"00000010",
  33489=>"00000010",
  33490=>"11111111",
  33491=>"11111110",
  33492=>"11111110",
  33493=>"11111110",
  33494=>"00000001",
  33495=>"00000010",
  33496=>"11111100",
  33497=>"00000000",
  33498=>"00000001",
  33499=>"00000010",
  33500=>"00000100",
  33501=>"00000001",
  33502=>"00000000",
  33503=>"00000010",
  33504=>"11111111",
  33505=>"11111111",
  33506=>"00000001",
  33507=>"00000011",
  33508=>"00000010",
  33509=>"11111111",
  33510=>"00000010",
  33511=>"00000000",
  33512=>"11111110",
  33513=>"11111111",
  33514=>"11111111",
  33515=>"00000011",
  33516=>"11111101",
  33517=>"00000000",
  33518=>"11111110",
  33519=>"00000001",
  33520=>"00000000",
  33521=>"11111111",
  33522=>"11111101",
  33523=>"00000010",
  33524=>"00000000",
  33525=>"00000001",
  33526=>"11111111",
  33527=>"00000001",
  33528=>"00000000",
  33529=>"00000010",
  33530=>"00000000",
  33531=>"11111111",
  33532=>"00000000",
  33533=>"11111110",
  33534=>"11111110",
  33535=>"11111110",
  33536=>"00000000",
  33537=>"00000101",
  33538=>"00000011",
  33539=>"11111110",
  33540=>"00000011",
  33541=>"00000001",
  33542=>"00000000",
  33543=>"11111111",
  33544=>"00000100",
  33545=>"00000001",
  33546=>"00000010",
  33547=>"00000011",
  33548=>"00000000",
  33549=>"11111101",
  33550=>"00000001",
  33551=>"00000010",
  33552=>"00000000",
  33553=>"00000011",
  33554=>"00000001",
  33555=>"11111110",
  33556=>"00000001",
  33557=>"00000110",
  33558=>"00000001",
  33559=>"11111101",
  33560=>"00000001",
  33561=>"11111110",
  33562=>"11111110",
  33563=>"00000000",
  33564=>"00000000",
  33565=>"00000000",
  33566=>"00000011",
  33567=>"11111110",
  33568=>"11111111",
  33569=>"00000000",
  33570=>"00000000",
  33571=>"00000000",
  33572=>"11111110",
  33573=>"11111101",
  33574=>"00000010",
  33575=>"00000000",
  33576=>"00000011",
  33577=>"00000000",
  33578=>"11111111",
  33579=>"00000000",
  33580=>"00000001",
  33581=>"11111110",
  33582=>"11111111",
  33583=>"11111111",
  33584=>"11111110",
  33585=>"00000010",
  33586=>"11111110",
  33587=>"00000011",
  33588=>"00000010",
  33589=>"00000100",
  33590=>"00000010",
  33591=>"00000010",
  33592=>"11111111",
  33593=>"00000000",
  33594=>"00000000",
  33595=>"00000011",
  33596=>"00000010",
  33597=>"11111101",
  33598=>"00000101",
  33599=>"11111110",
  33600=>"00000000",
  33601=>"00000000",
  33602=>"00000001",
  33603=>"00000001",
  33604=>"00000011",
  33605=>"11111110",
  33606=>"11111101",
  33607=>"00000001",
  33608=>"00000000",
  33609=>"11111111",
  33610=>"00000101",
  33611=>"11111111",
  33612=>"00000001",
  33613=>"00000000",
  33614=>"11111111",
  33615=>"00000010",
  33616=>"11111111",
  33617=>"00000010",
  33618=>"00000000",
  33619=>"11111111",
  33620=>"00000001",
  33621=>"11111111",
  33622=>"11111101",
  33623=>"11111101",
  33624=>"00000000",
  33625=>"00000001",
  33626=>"00000000",
  33627=>"11111111",
  33628=>"00000000",
  33629=>"00000010",
  33630=>"00000000",
  33631=>"11111101",
  33632=>"11111101",
  33633=>"11111111",
  33634=>"00000011",
  33635=>"00000001",
  33636=>"00000000",
  33637=>"11111111",
  33638=>"11111111",
  33639=>"11111111",
  33640=>"00000001",
  33641=>"11111110",
  33642=>"00000011",
  33643=>"00000011",
  33644=>"00000001",
  33645=>"11111110",
  33646=>"00000000",
  33647=>"00000010",
  33648=>"00000011",
  33649=>"11111101",
  33650=>"11111110",
  33651=>"00000001",
  33652=>"00000000",
  33653=>"11111110",
  33654=>"00000001",
  33655=>"11111110",
  33656=>"00000000",
  33657=>"00000000",
  33658=>"00000010",
  33659=>"11111110",
  33660=>"11111111",
  33661=>"00000010",
  33662=>"11111110",
  33663=>"00000010",
  33664=>"00000010",
  33665=>"11111101",
  33666=>"11111111",
  33667=>"00000001",
  33668=>"11111110",
  33669=>"00000010",
  33670=>"00000001",
  33671=>"00000001",
  33672=>"11111110",
  33673=>"11111111",
  33674=>"00000001",
  33675=>"11111101",
  33676=>"00000000",
  33677=>"11111111",
  33678=>"00000110",
  33679=>"00000000",
  33680=>"00000000",
  33681=>"11111111",
  33682=>"11111110",
  33683=>"11111110",
  33684=>"11111111",
  33685=>"00000010",
  33686=>"11111110",
  33687=>"00000100",
  33688=>"11111111",
  33689=>"00000010",
  33690=>"00000011",
  33691=>"00000000",
  33692=>"11111111",
  33693=>"11111110",
  33694=>"11111111",
  33695=>"11111111",
  33696=>"11111111",
  33697=>"00000010",
  33698=>"00000000",
  33699=>"00000000",
  33700=>"00000001",
  33701=>"11111111",
  33702=>"11111111",
  33703=>"11111101",
  33704=>"00000001",
  33705=>"00000001",
  33706=>"11111101",
  33707=>"11111111",
  33708=>"11111110",
  33709=>"11111101",
  33710=>"00000001",
  33711=>"00000000",
  33712=>"11111101",
  33713=>"00000001",
  33714=>"11111111",
  33715=>"11111111",
  33716=>"00000011",
  33717=>"00000001",
  33718=>"00000001",
  33719=>"11111110",
  33720=>"00000010",
  33721=>"11111111",
  33722=>"11111101",
  33723=>"11111110",
  33724=>"11111111",
  33725=>"11111111",
  33726=>"00000000",
  33727=>"00000001",
  33728=>"11111110",
  33729=>"11111101",
  33730=>"11111110",
  33731=>"00000010",
  33732=>"00000000",
  33733=>"00000001",
  33734=>"00000101",
  33735=>"11111111",
  33736=>"11111101",
  33737=>"00000011",
  33738=>"00000000",
  33739=>"11111101",
  33740=>"11111101",
  33741=>"11111110",
  33742=>"00000001",
  33743=>"11111110",
  33744=>"11111110",
  33745=>"11111101",
  33746=>"00000000",
  33747=>"00000010",
  33748=>"00000001",
  33749=>"00000100",
  33750=>"11111110",
  33751=>"11111111",
  33752=>"11111101",
  33753=>"11111111",
  33754=>"00000000",
  33755=>"00000000",
  33756=>"00000011",
  33757=>"00000011",
  33758=>"11111110",
  33759=>"11111110",
  33760=>"11111111",
  33761=>"00000000",
  33762=>"11111101",
  33763=>"00000000",
  33764=>"00000001",
  33765=>"00000011",
  33766=>"00000000",
  33767=>"00000011",
  33768=>"00000010",
  33769=>"11111110",
  33770=>"00000100",
  33771=>"11111101",
  33772=>"11111111",
  33773=>"00000000",
  33774=>"11111101",
  33775=>"00000000",
  33776=>"00000000",
  33777=>"00000001",
  33778=>"00000000",
  33779=>"11111111",
  33780=>"11111111",
  33781=>"00000001",
  33782=>"00000010",
  33783=>"00000000",
  33784=>"11111111",
  33785=>"11111110",
  33786=>"11111111",
  33787=>"00000010",
  33788=>"11111100",
  33789=>"11111111",
  33790=>"00000110",
  33791=>"11111101",
  33792=>"00000011",
  33793=>"11111110",
  33794=>"00000001",
  33795=>"00000010",
  33796=>"11111100",
  33797=>"11111110",
  33798=>"00000001",
  33799=>"11111101",
  33800=>"11111111",
  33801=>"00000011",
  33802=>"11111101",
  33803=>"00000011",
  33804=>"11111111",
  33805=>"11111110",
  33806=>"00000001",
  33807=>"00000011",
  33808=>"00000100",
  33809=>"00000001",
  33810=>"00000010",
  33811=>"11111111",
  33812=>"00000001",
  33813=>"00000000",
  33814=>"00000101",
  33815=>"00000010",
  33816=>"00000001",
  33817=>"11111101",
  33818=>"00000001",
  33819=>"00000000",
  33820=>"00000000",
  33821=>"00000001",
  33822=>"00000001",
  33823=>"11111111",
  33824=>"00000011",
  33825=>"00000000",
  33826=>"11111111",
  33827=>"00000001",
  33828=>"00000001",
  33829=>"00000001",
  33830=>"00000011",
  33831=>"00000000",
  33832=>"00000001",
  33833=>"00000000",
  33834=>"11111110",
  33835=>"00000001",
  33836=>"00000001",
  33837=>"00000001",
  33838=>"00000000",
  33839=>"00000010",
  33840=>"00000000",
  33841=>"11111111",
  33842=>"11111110",
  33843=>"11111110",
  33844=>"11111110",
  33845=>"11111101",
  33846=>"00000010",
  33847=>"00000100",
  33848=>"11111111",
  33849=>"00000001",
  33850=>"00000001",
  33851=>"00000001",
  33852=>"11111111",
  33853=>"00000000",
  33854=>"11111111",
  33855=>"11111101",
  33856=>"11111100",
  33857=>"00000001",
  33858=>"00000011",
  33859=>"00000010",
  33860=>"00000010",
  33861=>"00000000",
  33862=>"11111101",
  33863=>"11111101",
  33864=>"00000000",
  33865=>"00000000",
  33866=>"00000001",
  33867=>"11111110",
  33868=>"00000110",
  33869=>"11111110",
  33870=>"00000001",
  33871=>"00000000",
  33872=>"00000000",
  33873=>"00000010",
  33874=>"00000011",
  33875=>"00000000",
  33876=>"00000100",
  33877=>"00000010",
  33878=>"00000000",
  33879=>"11111110",
  33880=>"11111110",
  33881=>"11111110",
  33882=>"11111110",
  33883=>"00000000",
  33884=>"00000001",
  33885=>"00000000",
  33886=>"00000010",
  33887=>"00000001",
  33888=>"11111110",
  33889=>"11111111",
  33890=>"00000000",
  33891=>"00000001",
  33892=>"00000001",
  33893=>"00000010",
  33894=>"00000010",
  33895=>"11111101",
  33896=>"11111101",
  33897=>"00000001",
  33898=>"11111110",
  33899=>"11111110",
  33900=>"11111100",
  33901=>"00000010",
  33902=>"00000010",
  33903=>"00000001",
  33904=>"00000010",
  33905=>"11111110",
  33906=>"00000001",
  33907=>"00000001",
  33908=>"00000001",
  33909=>"00000000",
  33910=>"00000110",
  33911=>"00000010",
  33912=>"00000001",
  33913=>"11111111",
  33914=>"11111111",
  33915=>"00000000",
  33916=>"00000010",
  33917=>"11111110",
  33918=>"00000000",
  33919=>"00000100",
  33920=>"00000000",
  33921=>"11111110",
  33922=>"00000000",
  33923=>"00000000",
  33924=>"11111110",
  33925=>"00000000",
  33926=>"00000001",
  33927=>"11111110",
  33928=>"11111110",
  33929=>"00000000",
  33930=>"00000001",
  33931=>"11111111",
  33932=>"11111111",
  33933=>"00000010",
  33934=>"11111110",
  33935=>"11111111",
  33936=>"00000001",
  33937=>"00000000",
  33938=>"00000011",
  33939=>"00000000",
  33940=>"00000011",
  33941=>"00000001",
  33942=>"11111110",
  33943=>"00000000",
  33944=>"11111111",
  33945=>"00000011",
  33946=>"11111101",
  33947=>"00000001",
  33948=>"11111110",
  33949=>"00000000",
  33950=>"00000001",
  33951=>"00000001",
  33952=>"00000000",
  33953=>"11111111",
  33954=>"11111111",
  33955=>"00000001",
  33956=>"00000011",
  33957=>"00000010",
  33958=>"11111101",
  33959=>"11111111",
  33960=>"11111111",
  33961=>"11111111",
  33962=>"00000011",
  33963=>"00000010",
  33964=>"00000001",
  33965=>"00000001",
  33966=>"11111110",
  33967=>"11111110",
  33968=>"00000001",
  33969=>"11111101",
  33970=>"00000000",
  33971=>"00000000",
  33972=>"11111101",
  33973=>"00000111",
  33974=>"11111101",
  33975=>"11111110",
  33976=>"00000010",
  33977=>"11111101",
  33978=>"00000011",
  33979=>"00000001",
  33980=>"11111111",
  33981=>"00000000",
  33982=>"00000001",
  33983=>"11111111",
  33984=>"00000010",
  33985=>"00000010",
  33986=>"00000000",
  33987=>"00000001",
  33988=>"00000000",
  33989=>"11111111",
  33990=>"11111110",
  33991=>"00000011",
  33992=>"00000100",
  33993=>"00000010",
  33994=>"00000001",
  33995=>"11111100",
  33996=>"11111111",
  33997=>"00000010",
  33998=>"11111111",
  33999=>"11111110",
  34000=>"00000001",
  34001=>"00000010",
  34002=>"00000001",
  34003=>"00000010",
  34004=>"00000001",
  34005=>"00000000",
  34006=>"00000010",
  34007=>"00000100",
  34008=>"00000011",
  34009=>"00000001",
  34010=>"00000000",
  34011=>"11111111",
  34012=>"11111111",
  34013=>"11111110",
  34014=>"00000110",
  34015=>"11111110",
  34016=>"11111110",
  34017=>"11111110",
  34018=>"11111110",
  34019=>"00000001",
  34020=>"00000000",
  34021=>"11111110",
  34022=>"00000000",
  34023=>"00000000",
  34024=>"11111110",
  34025=>"11111111",
  34026=>"00000001",
  34027=>"00000010",
  34028=>"11111110",
  34029=>"00000010",
  34030=>"11111110",
  34031=>"11111101",
  34032=>"00000001",
  34033=>"00000001",
  34034=>"00000001",
  34035=>"11111111",
  34036=>"00000000",
  34037=>"00000001",
  34038=>"00000010",
  34039=>"00000000",
  34040=>"00000000",
  34041=>"00000000",
  34042=>"11111111",
  34043=>"11111110",
  34044=>"00000001",
  34045=>"11111100",
  34046=>"11111111",
  34047=>"00000001",
  34048=>"11111111",
  34049=>"11111111",
  34050=>"00000001",
  34051=>"00000010",
  34052=>"00000001",
  34053=>"11111101",
  34054=>"00000000",
  34055=>"00000001",
  34056=>"00000000",
  34057=>"00000000",
  34058=>"00000010",
  34059=>"00000000",
  34060=>"11111111",
  34061=>"11111101",
  34062=>"00000010",
  34063=>"00000110",
  34064=>"00000011",
  34065=>"00000000",
  34066=>"11111110",
  34067=>"00000001",
  34068=>"11111111",
  34069=>"00000000",
  34070=>"11111111",
  34071=>"11111101",
  34072=>"00000001",
  34073=>"11111111",
  34074=>"11111110",
  34075=>"00000000",
  34076=>"11111111",
  34077=>"11111111",
  34078=>"11111111",
  34079=>"00000001",
  34080=>"00000011",
  34081=>"00000011",
  34082=>"00000001",
  34083=>"11111111",
  34084=>"11111101",
  34085=>"11111110",
  34086=>"00000000",
  34087=>"11111111",
  34088=>"11111111",
  34089=>"11111110",
  34090=>"11111110",
  34091=>"00000001",
  34092=>"11111111",
  34093=>"00000010",
  34094=>"00000010",
  34095=>"00000001",
  34096=>"00000001",
  34097=>"11111110",
  34098=>"11111101",
  34099=>"00000010",
  34100=>"11111111",
  34101=>"11111110",
  34102=>"00000010",
  34103=>"11111111",
  34104=>"00000000",
  34105=>"11111101",
  34106=>"00000010",
  34107=>"11111110",
  34108=>"11111111",
  34109=>"11111111",
  34110=>"00000010",
  34111=>"11111110",
  34112=>"11111111",
  34113=>"00000001",
  34114=>"00000000",
  34115=>"11111111",
  34116=>"00000010",
  34117=>"11111110",
  34118=>"00000001",
  34119=>"11111111",
  34120=>"00000011",
  34121=>"11111100",
  34122=>"11111101",
  34123=>"00000010",
  34124=>"00000001",
  34125=>"00000001",
  34126=>"11111110",
  34127=>"11111111",
  34128=>"00000101",
  34129=>"11111101",
  34130=>"11111111",
  34131=>"00000001",
  34132=>"00000000",
  34133=>"00000000",
  34134=>"00000001",
  34135=>"11111111",
  34136=>"11111111",
  34137=>"00000010",
  34138=>"11111111",
  34139=>"00000011",
  34140=>"00000010",
  34141=>"11111111",
  34142=>"00000011",
  34143=>"11111111",
  34144=>"00000001",
  34145=>"11111111",
  34146=>"00000000",
  34147=>"00000001",
  34148=>"00000001",
  34149=>"00000000",
  34150=>"11111101",
  34151=>"11111111",
  34152=>"11111111",
  34153=>"11111111",
  34154=>"11111110",
  34155=>"11111110",
  34156=>"11111101",
  34157=>"11111101",
  34158=>"00000110",
  34159=>"11111101",
  34160=>"11111111",
  34161=>"11111110",
  34162=>"11111111",
  34163=>"00000001",
  34164=>"00000001",
  34165=>"11111101",
  34166=>"11111110",
  34167=>"00000010",
  34168=>"00000001",
  34169=>"11111111",
  34170=>"00000000",
  34171=>"00000001",
  34172=>"00000000",
  34173=>"00000001",
  34174=>"00000100",
  34175=>"00000000",
  34176=>"11111111",
  34177=>"11111111",
  34178=>"11111111",
  34179=>"11111101",
  34180=>"00000010",
  34181=>"11111111",
  34182=>"11111110",
  34183=>"11111111",
  34184=>"00000001",
  34185=>"00000001",
  34186=>"00000100",
  34187=>"00000010",
  34188=>"00000001",
  34189=>"00000000",
  34190=>"00000011",
  34191=>"00000000",
  34192=>"00000010",
  34193=>"11111111",
  34194=>"00000011",
  34195=>"11111111",
  34196=>"11111111",
  34197=>"00000000",
  34198=>"11111110",
  34199=>"11111111",
  34200=>"11111101",
  34201=>"00000001",
  34202=>"11111101",
  34203=>"00000001",
  34204=>"00000001",
  34205=>"00000100",
  34206=>"11111111",
  34207=>"00000010",
  34208=>"11111111",
  34209=>"00000001",
  34210=>"00000100",
  34211=>"11111110",
  34212=>"11111111",
  34213=>"11111110",
  34214=>"00000100",
  34215=>"00000001",
  34216=>"11111111",
  34217=>"00000000",
  34218=>"00000010",
  34219=>"00000010",
  34220=>"11111101",
  34221=>"00000000",
  34222=>"00000000",
  34223=>"00000010",
  34224=>"11111110",
  34225=>"11111110",
  34226=>"11111110",
  34227=>"00000010",
  34228=>"00000011",
  34229=>"11111111",
  34230=>"00000100",
  34231=>"11111111",
  34232=>"11111111",
  34233=>"00000001",
  34234=>"00000001",
  34235=>"00000000",
  34236=>"00000010",
  34237=>"11111110",
  34238=>"11111111",
  34239=>"00000000",
  34240=>"00000010",
  34241=>"11111101",
  34242=>"00000001",
  34243=>"11111101",
  34244=>"11111101",
  34245=>"11111111",
  34246=>"11111101",
  34247=>"11111111",
  34248=>"00000001",
  34249=>"00000101",
  34250=>"11111111",
  34251=>"00000010",
  34252=>"00000011",
  34253=>"11111110",
  34254=>"00000001",
  34255=>"00000000",
  34256=>"11111111",
  34257=>"00000011",
  34258=>"11111101",
  34259=>"11111110",
  34260=>"11111111",
  34261=>"11111101",
  34262=>"11111111",
  34263=>"00000000",
  34264=>"00000010",
  34265=>"11111101",
  34266=>"11111110",
  34267=>"00000001",
  34268=>"11111110",
  34269=>"11111111",
  34270=>"11111101",
  34271=>"11111110",
  34272=>"11111111",
  34273=>"00000001",
  34274=>"00000001",
  34275=>"00000001",
  34276=>"00000011",
  34277=>"00000000",
  34278=>"11111110",
  34279=>"00000001",
  34280=>"00000000",
  34281=>"00000001",
  34282=>"11111111",
  34283=>"11111110",
  34284=>"00000001",
  34285=>"11111110",
  34286=>"00000001",
  34287=>"11111111",
  34288=>"11111110",
  34289=>"11111110",
  34290=>"11111111",
  34291=>"00000000",
  34292=>"11111101",
  34293=>"00000001",
  34294=>"11111101",
  34295=>"00000001",
  34296=>"00000100",
  34297=>"11111111",
  34298=>"00000001",
  34299=>"11111110",
  34300=>"00000010",
  34301=>"00000000",
  34302=>"11111111",
  34303=>"00000000",
  34304=>"00000000",
  34305=>"11111110",
  34306=>"00000010",
  34307=>"11111111",
  34308=>"00000001",
  34309=>"11111101",
  34310=>"11111110",
  34311=>"00000010",
  34312=>"00000001",
  34313=>"00000011",
  34314=>"00000010",
  34315=>"11111111",
  34316=>"00000001",
  34317=>"00000010",
  34318=>"00000000",
  34319=>"11111111",
  34320=>"00000011",
  34321=>"00000001",
  34322=>"00000000",
  34323=>"00000001",
  34324=>"00000000",
  34325=>"00000010",
  34326=>"00000010",
  34327=>"00000000",
  34328=>"11111101",
  34329=>"00000001",
  34330=>"00000000",
  34331=>"00000001",
  34332=>"11111110",
  34333=>"11111110",
  34334=>"11111101",
  34335=>"00000001",
  34336=>"11111110",
  34337=>"00000011",
  34338=>"11111101",
  34339=>"11111110",
  34340=>"11111101",
  34341=>"11111110",
  34342=>"00000001",
  34343=>"00000001",
  34344=>"00000010",
  34345=>"00000000",
  34346=>"11111110",
  34347=>"00000000",
  34348=>"11111110",
  34349=>"00000010",
  34350=>"00000000",
  34351=>"11111101",
  34352=>"00000001",
  34353=>"11111111",
  34354=>"00000011",
  34355=>"11111111",
  34356=>"11111110",
  34357=>"00000011",
  34358=>"11111111",
  34359=>"11111110",
  34360=>"11111110",
  34361=>"00000001",
  34362=>"11111101",
  34363=>"00000000",
  34364=>"11111100",
  34365=>"11111101",
  34366=>"11111110",
  34367=>"11111111",
  34368=>"11111101",
  34369=>"00000001",
  34370=>"00000000",
  34371=>"11111110",
  34372=>"00000011",
  34373=>"11111111",
  34374=>"00000001",
  34375=>"11111111",
  34376=>"00000010",
  34377=>"11111101",
  34378=>"11111110",
  34379=>"11111110",
  34380=>"00000011",
  34381=>"11111111",
  34382=>"11111111",
  34383=>"00000001",
  34384=>"00000010",
  34385=>"00000000",
  34386=>"11111111",
  34387=>"11111110",
  34388=>"11111101",
  34389=>"11111110",
  34390=>"11111111",
  34391=>"11111111",
  34392=>"00000010",
  34393=>"00000000",
  34394=>"00000010",
  34395=>"00000101",
  34396=>"00000010",
  34397=>"11111111",
  34398=>"00000010",
  34399=>"00000001",
  34400=>"00000000",
  34401=>"00000011",
  34402=>"00000001",
  34403=>"11111110",
  34404=>"11111111",
  34405=>"11111110",
  34406=>"00000010",
  34407=>"11111101",
  34408=>"00000010",
  34409=>"11111101",
  34410=>"00000000",
  34411=>"00000000",
  34412=>"11111111",
  34413=>"00000100",
  34414=>"11111101",
  34415=>"11111100",
  34416=>"11111101",
  34417=>"11111110",
  34418=>"11111101",
  34419=>"11111101",
  34420=>"00000000",
  34421=>"11111111",
  34422=>"11111111",
  34423=>"11111111",
  34424=>"00000010",
  34425=>"11111111",
  34426=>"11111111",
  34427=>"11111111",
  34428=>"00000001",
  34429=>"00000001",
  34430=>"11111101",
  34431=>"11111111",
  34432=>"00000001",
  34433=>"00000000",
  34434=>"00000000",
  34435=>"11111101",
  34436=>"11111110",
  34437=>"11111110",
  34438=>"11111111",
  34439=>"00000001",
  34440=>"00000000",
  34441=>"00000010",
  34442=>"00000011",
  34443=>"00000000",
  34444=>"00000000",
  34445=>"11111110",
  34446=>"00000010",
  34447=>"00000000",
  34448=>"11111111",
  34449=>"00000110",
  34450=>"00000000",
  34451=>"00000010",
  34452=>"11111101",
  34453=>"11111101",
  34454=>"00000000",
  34455=>"11111110",
  34456=>"00000000",
  34457=>"00000010",
  34458=>"00000101",
  34459=>"00000000",
  34460=>"00000001",
  34461=>"00000010",
  34462=>"00000101",
  34463=>"00000000",
  34464=>"00000000",
  34465=>"11111110",
  34466=>"00000000",
  34467=>"00000000",
  34468=>"00000010",
  34469=>"11111101",
  34470=>"11111110",
  34471=>"11111110",
  34472=>"00000010",
  34473=>"11111111",
  34474=>"11111110",
  34475=>"00000010",
  34476=>"00000001",
  34477=>"00000010",
  34478=>"11111110",
  34479=>"00000010",
  34480=>"00000010",
  34481=>"00000011",
  34482=>"00000001",
  34483=>"11111101",
  34484=>"11111101",
  34485=>"11111101",
  34486=>"11111111",
  34487=>"00000001",
  34488=>"00000010",
  34489=>"11111110",
  34490=>"00000011",
  34491=>"00000010",
  34492=>"00000100",
  34493=>"00000000",
  34494=>"00000000",
  34495=>"00000000",
  34496=>"00000010",
  34497=>"11111110",
  34498=>"11111110",
  34499=>"00000001",
  34500=>"11111110",
  34501=>"00000101",
  34502=>"00000010",
  34503=>"11111111",
  34504=>"11111110",
  34505=>"00000010",
  34506=>"00000000",
  34507=>"00000000",
  34508=>"00000001",
  34509=>"00000100",
  34510=>"11111111",
  34511=>"00000000",
  34512=>"00000001",
  34513=>"11111101",
  34514=>"00000000",
  34515=>"00000100",
  34516=>"11111110",
  34517=>"00000001",
  34518=>"11111111",
  34519=>"11111100",
  34520=>"00000111",
  34521=>"11111111",
  34522=>"00000010",
  34523=>"00000010",
  34524=>"00000010",
  34525=>"11111110",
  34526=>"00000000",
  34527=>"00000010",
  34528=>"11111110",
  34529=>"00000001",
  34530=>"00000010",
  34531=>"11111111",
  34532=>"00000010",
  34533=>"00000000",
  34534=>"11111111",
  34535=>"00000010",
  34536=>"11111111",
  34537=>"11111101",
  34538=>"11111110",
  34539=>"00000000",
  34540=>"00000010",
  34541=>"00000000",
  34542=>"00000000",
  34543=>"00000010",
  34544=>"00000001",
  34545=>"11111110",
  34546=>"11111110",
  34547=>"00000010",
  34548=>"11111101",
  34549=>"00000001",
  34550=>"00000010",
  34551=>"11111110",
  34552=>"11111100",
  34553=>"00000001",
  34554=>"11111110",
  34555=>"11111101",
  34556=>"00000010",
  34557=>"00000000",
  34558=>"11111101",
  34559=>"00000011",
  34560=>"11111111",
  34561=>"00000000",
  34562=>"11111110",
  34563=>"11111111",
  34564=>"11111101",
  34565=>"00000001",
  34566=>"11111101",
  34567=>"00000000",
  34568=>"00000011",
  34569=>"11111111",
  34570=>"00000010",
  34571=>"00000010",
  34572=>"11111110",
  34573=>"00000000",
  34574=>"11111111",
  34575=>"00000011",
  34576=>"00000011",
  34577=>"00000001",
  34578=>"00000001",
  34579=>"00000100",
  34580=>"00000000",
  34581=>"00000000",
  34582=>"11111110",
  34583=>"00000001",
  34584=>"11111111",
  34585=>"11111101",
  34586=>"00000000",
  34587=>"11111110",
  34588=>"00000011",
  34589=>"11111111",
  34590=>"11111110",
  34591=>"11111111",
  34592=>"11111110",
  34593=>"00000000",
  34594=>"00000011",
  34595=>"00000000",
  34596=>"11111110",
  34597=>"00000001",
  34598=>"11111101",
  34599=>"11111101",
  34600=>"00000000",
  34601=>"00000001",
  34602=>"11111100",
  34603=>"11111111",
  34604=>"00000001",
  34605=>"00000000",
  34606=>"11111110",
  34607=>"00000000",
  34608=>"11111111",
  34609=>"11111101",
  34610=>"00000000",
  34611=>"00000001",
  34612=>"00000001",
  34613=>"11111110",
  34614=>"00000000",
  34615=>"11111101",
  34616=>"11111111",
  34617=>"11111110",
  34618=>"00000000",
  34619=>"11111111",
  34620=>"00000010",
  34621=>"00000010",
  34622=>"00000010",
  34623=>"11111110",
  34624=>"11111101",
  34625=>"00000000",
  34626=>"00000000",
  34627=>"00000000",
  34628=>"11111111",
  34629=>"00000001",
  34630=>"00000000",
  34631=>"00000001",
  34632=>"00000100",
  34633=>"00000001",
  34634=>"11111101",
  34635=>"11111111",
  34636=>"11111111",
  34637=>"11111111",
  34638=>"00000000",
  34639=>"00000010",
  34640=>"11111111",
  34641=>"11111110",
  34642=>"00000000",
  34643=>"11111101",
  34644=>"11111111",
  34645=>"11111101",
  34646=>"11111111",
  34647=>"11111110",
  34648=>"11111110",
  34649=>"00000001",
  34650=>"11111111",
  34651=>"11111111",
  34652=>"11111111",
  34653=>"11111111",
  34654=>"11111101",
  34655=>"00000000",
  34656=>"00000010",
  34657=>"00000100",
  34658=>"11111110",
  34659=>"11111111",
  34660=>"00000001",
  34661=>"00000001",
  34662=>"00000010",
  34663=>"11111110",
  34664=>"00000001",
  34665=>"00000011",
  34666=>"00000000",
  34667=>"00000010",
  34668=>"11111111",
  34669=>"11111100",
  34670=>"00000000",
  34671=>"00000000",
  34672=>"11111101",
  34673=>"11111111",
  34674=>"00000001",
  34675=>"00000000",
  34676=>"00000001",
  34677=>"11111101",
  34678=>"00000000",
  34679=>"00000000",
  34680=>"00000010",
  34681=>"11111110",
  34682=>"00000001",
  34683=>"11111111",
  34684=>"00000001",
  34685=>"00000001",
  34686=>"00000110",
  34687=>"11111101",
  34688=>"11111111",
  34689=>"00000110",
  34690=>"00000000",
  34691=>"00000001",
  34692=>"00000001",
  34693=>"11111111",
  34694=>"00000011",
  34695=>"11111111",
  34696=>"11111111",
  34697=>"11111111",
  34698=>"11111111",
  34699=>"00000010",
  34700=>"11111111",
  34701=>"11111111",
  34702=>"00000000",
  34703=>"00000001",
  34704=>"11111111",
  34705=>"11111110",
  34706=>"11111110",
  34707=>"00000001",
  34708=>"11111110",
  34709=>"00000001",
  34710=>"11111111",
  34711=>"11111110",
  34712=>"00000001",
  34713=>"00000010",
  34714=>"00000001",
  34715=>"11111110",
  34716=>"00000000",
  34717=>"11111111",
  34718=>"11111111",
  34719=>"11111101",
  34720=>"11111101",
  34721=>"00000010",
  34722=>"00000010",
  34723=>"11111110",
  34724=>"11111111",
  34725=>"00000011",
  34726=>"00000001",
  34727=>"00000001",
  34728=>"11111111",
  34729=>"00000001",
  34730=>"00000000",
  34731=>"00000010",
  34732=>"00000010",
  34733=>"00000001",
  34734=>"00000000",
  34735=>"11111110",
  34736=>"11111110",
  34737=>"00000000",
  34738=>"00000110",
  34739=>"00000001",
  34740=>"00000000",
  34741=>"00000010",
  34742=>"00000001",
  34743=>"11111110",
  34744=>"11111110",
  34745=>"11111111",
  34746=>"00000000",
  34747=>"00000010",
  34748=>"00000000",
  34749=>"11111101",
  34750=>"11111101",
  34751=>"00000010",
  34752=>"00000100",
  34753=>"11111101",
  34754=>"00000010",
  34755=>"11111110",
  34756=>"00000010",
  34757=>"11111111",
  34758=>"11111101",
  34759=>"11111111",
  34760=>"00000000",
  34761=>"00000000",
  34762=>"11111101",
  34763=>"11111101",
  34764=>"11111111",
  34765=>"00000001",
  34766=>"00000001",
  34767=>"00000001",
  34768=>"11111111",
  34769=>"11111111",
  34770=>"11111110",
  34771=>"00000011",
  34772=>"00000001",
  34773=>"11111110",
  34774=>"11111111",
  34775=>"00000011",
  34776=>"00000000",
  34777=>"11111101",
  34778=>"00000010",
  34779=>"11111101",
  34780=>"11111110",
  34781=>"00000001",
  34782=>"11111101",
  34783=>"00000011",
  34784=>"00000001",
  34785=>"11111101",
  34786=>"11111111",
  34787=>"00000011",
  34788=>"00000001",
  34789=>"11111111",
  34790=>"11111110",
  34791=>"00000001",
  34792=>"00000001",
  34793=>"11111110",
  34794=>"11111101",
  34795=>"11111110",
  34796=>"11111101",
  34797=>"00000001",
  34798=>"11111101",
  34799=>"00000001",
  34800=>"00000010",
  34801=>"00000000",
  34802=>"11111111",
  34803=>"00000000",
  34804=>"00000001",
  34805=>"00000100",
  34806=>"00000000",
  34807=>"11111110",
  34808=>"00000001",
  34809=>"00000000",
  34810=>"11111110",
  34811=>"00000001",
  34812=>"11111110",
  34813=>"11111111",
  34814=>"00000001",
  34815=>"11111111",
  34816=>"00000000",
  34817=>"00000000",
  34818=>"11111110",
  34819=>"11111110",
  34820=>"11111111",
  34821=>"00000000",
  34822=>"11111110",
  34823=>"00000000",
  34824=>"00000001",
  34825=>"11111101",
  34826=>"00000001",
  34827=>"00000001",
  34828=>"00000010",
  34829=>"00000011",
  34830=>"11111011",
  34831=>"00000001",
  34832=>"11111110",
  34833=>"11111110",
  34834=>"11111110",
  34835=>"11111101",
  34836=>"11111101",
  34837=>"00000010",
  34838=>"11111111",
  34839=>"00000010",
  34840=>"11111110",
  34841=>"00000010",
  34842=>"00000101",
  34843=>"00000010",
  34844=>"11111111",
  34845=>"00000001",
  34846=>"00000010",
  34847=>"00000100",
  34848=>"00000000",
  34849=>"11111101",
  34850=>"00000010",
  34851=>"00000100",
  34852=>"11111110",
  34853=>"11111100",
  34854=>"11111110",
  34855=>"00000011",
  34856=>"11111011",
  34857=>"00000100",
  34858=>"00000001",
  34859=>"00000010",
  34860=>"00000010",
  34861=>"00000000",
  34862=>"11111110",
  34863=>"11111101",
  34864=>"00000011",
  34865=>"00000000",
  34866=>"11111110",
  34867=>"11111101",
  34868=>"11111111",
  34869=>"00000000",
  34870=>"00000010",
  34871=>"00000001",
  34872=>"11111101",
  34873=>"00000000",
  34874=>"11111111",
  34875=>"11111110",
  34876=>"11111110",
  34877=>"11111110",
  34878=>"11111110",
  34879=>"00000010",
  34880=>"11111110",
  34881=>"11111100",
  34882=>"00000000",
  34883=>"00000001",
  34884=>"11111110",
  34885=>"00000100",
  34886=>"00000000",
  34887=>"11111110",
  34888=>"00000010",
  34889=>"11111110",
  34890=>"11111101",
  34891=>"00000000",
  34892=>"00000001",
  34893=>"00000000",
  34894=>"00000010",
  34895=>"00000000",
  34896=>"00000011",
  34897=>"00000011",
  34898=>"00000100",
  34899=>"11111101",
  34900=>"00000001",
  34901=>"00000001",
  34902=>"11111101",
  34903=>"00000001",
  34904=>"00000010",
  34905=>"11111110",
  34906=>"00000100",
  34907=>"00000000",
  34908=>"00000001",
  34909=>"11111101",
  34910=>"11111111",
  34911=>"00000110",
  34912=>"11111100",
  34913=>"11111100",
  34914=>"00000001",
  34915=>"11111110",
  34916=>"11111100",
  34917=>"00000010",
  34918=>"00000000",
  34919=>"00000010",
  34920=>"00000011",
  34921=>"11111111",
  34922=>"00000000",
  34923=>"00000001",
  34924=>"00000100",
  34925=>"11111101",
  34926=>"00000000",
  34927=>"00000010",
  34928=>"11111101",
  34929=>"11111110",
  34930=>"11111101",
  34931=>"11111111",
  34932=>"00000010",
  34933=>"11111111",
  34934=>"11111101",
  34935=>"11111110",
  34936=>"00000001",
  34937=>"11111101",
  34938=>"00000001",
  34939=>"11111111",
  34940=>"11111101",
  34941=>"11111110",
  34942=>"11111111",
  34943=>"11111111",
  34944=>"11111101",
  34945=>"00000010",
  34946=>"11111111",
  34947=>"11111110",
  34948=>"00000011",
  34949=>"00000010",
  34950=>"11111110",
  34951=>"00000100",
  34952=>"11111101",
  34953=>"11111111",
  34954=>"00000000",
  34955=>"11111011",
  34956=>"00000001",
  34957=>"00000001",
  34958=>"00000010",
  34959=>"00000010",
  34960=>"00000011",
  34961=>"11111101",
  34962=>"11111111",
  34963=>"00000001",
  34964=>"11111101",
  34965=>"11111110",
  34966=>"00000100",
  34967=>"11111101",
  34968=>"00000000",
  34969=>"00000010",
  34970=>"00000000",
  34971=>"00000010",
  34972=>"00000010",
  34973=>"11111100",
  34974=>"00000001",
  34975=>"11111100",
  34976=>"00000101",
  34977=>"11111111",
  34978=>"11111110",
  34979=>"00000011",
  34980=>"11111110",
  34981=>"11111111",
  34982=>"00000101",
  34983=>"11111111",
  34984=>"00000011",
  34985=>"11111111",
  34986=>"00000000",
  34987=>"11111111",
  34988=>"11111101",
  34989=>"00000000",
  34990=>"11111111",
  34991=>"00000100",
  34992=>"11111110",
  34993=>"11111111",
  34994=>"11111111",
  34995=>"00000011",
  34996=>"11111100",
  34997=>"11111110",
  34998=>"00000100",
  34999=>"11111111",
  35000=>"11111101",
  35001=>"11111110",
  35002=>"00000000",
  35003=>"00000001",
  35004=>"00000001",
  35005=>"11111111",
  35006=>"00000011",
  35007=>"00000001",
  35008=>"00000001",
  35009=>"11111110",
  35010=>"11111111",
  35011=>"00000010",
  35012=>"00000000",
  35013=>"11111111",
  35014=>"00000000",
  35015=>"00000001",
  35016=>"00000001",
  35017=>"11111100",
  35018=>"11111110",
  35019=>"00000000",
  35020=>"00000000",
  35021=>"00000000",
  35022=>"00000001",
  35023=>"00000110",
  35024=>"00000101",
  35025=>"11111111",
  35026=>"00000001",
  35027=>"00000011",
  35028=>"00000001",
  35029=>"00000000",
  35030=>"00000001",
  35031=>"00000010",
  35032=>"11111101",
  35033=>"00000011",
  35034=>"11111111",
  35035=>"11111111",
  35036=>"11111100",
  35037=>"00000100",
  35038=>"11111110",
  35039=>"00000100",
  35040=>"00000000",
  35041=>"00000000",
  35042=>"00000001",
  35043=>"11111101",
  35044=>"00000010",
  35045=>"00000000",
  35046=>"00000000",
  35047=>"11111111",
  35048=>"11111110",
  35049=>"00000011",
  35050=>"11111101",
  35051=>"00000010",
  35052=>"11111110",
  35053=>"00000010",
  35054=>"00000000",
  35055=>"11111110",
  35056=>"00000100",
  35057=>"11111110",
  35058=>"11111110",
  35059=>"00000010",
  35060=>"00000011",
  35061=>"00000010",
  35062=>"11111111",
  35063=>"00000010",
  35064=>"11111111",
  35065=>"00000011",
  35066=>"00000000",
  35067=>"00000010",
  35068=>"11111101",
  35069=>"00000011",
  35070=>"00000001",
  35071=>"00000001",
  35072=>"00000000",
  35073=>"11111110",
  35074=>"11111101",
  35075=>"00000000",
  35076=>"00000001",
  35077=>"00000011",
  35078=>"00000011",
  35079=>"00000011",
  35080=>"00000000",
  35081=>"11111101",
  35082=>"00000000",
  35083=>"00000010",
  35084=>"00000010",
  35085=>"00000001",
  35086=>"00000010",
  35087=>"00000010",
  35088=>"00000001",
  35089=>"00000110",
  35090=>"00000000",
  35091=>"00000000",
  35092=>"00000011",
  35093=>"00000010",
  35094=>"00000000",
  35095=>"00000001",
  35096=>"00000001",
  35097=>"11111111",
  35098=>"00000001",
  35099=>"00000010",
  35100=>"11111101",
  35101=>"00000001",
  35102=>"00000011",
  35103=>"00000000",
  35104=>"00000001",
  35105=>"00000001",
  35106=>"11111110",
  35107=>"11111111",
  35108=>"11111110",
  35109=>"11111101",
  35110=>"11111111",
  35111=>"00000100",
  35112=>"11111110",
  35113=>"11111110",
  35114=>"00000001",
  35115=>"00000010",
  35116=>"00000000",
  35117=>"11111111",
  35118=>"00000100",
  35119=>"11111110",
  35120=>"11111111",
  35121=>"11111110",
  35122=>"00000010",
  35123=>"00000011",
  35124=>"00000101",
  35125=>"00000001",
  35126=>"11111101",
  35127=>"00000000",
  35128=>"11111111",
  35129=>"11111100",
  35130=>"00000000",
  35131=>"00000011",
  35132=>"00000001",
  35133=>"11111110",
  35134=>"11111110",
  35135=>"00000000",
  35136=>"00000010",
  35137=>"11111110",
  35138=>"00000010",
  35139=>"11111110",
  35140=>"00000000",
  35141=>"11111110",
  35142=>"00000000",
  35143=>"00000000",
  35144=>"00000000",
  35145=>"00000001",
  35146=>"00000100",
  35147=>"11111110",
  35148=>"11111101",
  35149=>"00000000",
  35150=>"00000000",
  35151=>"00000000",
  35152=>"11111111",
  35153=>"11111110",
  35154=>"11111111",
  35155=>"11111111",
  35156=>"00000010",
  35157=>"11111111",
  35158=>"11111101",
  35159=>"11111110",
  35160=>"00000000",
  35161=>"00000000",
  35162=>"00000001",
  35163=>"00000000",
  35164=>"00000000",
  35165=>"00000010",
  35166=>"00000001",
  35167=>"00000000",
  35168=>"11111110",
  35169=>"00000000",
  35170=>"00000001",
  35171=>"00000000",
  35172=>"11111101",
  35173=>"11111101",
  35174=>"11111111",
  35175=>"00000001",
  35176=>"00000100",
  35177=>"00000010",
  35178=>"00000010",
  35179=>"00000100",
  35180=>"11111110",
  35181=>"11111110",
  35182=>"11111110",
  35183=>"00000010",
  35184=>"00000000",
  35185=>"00000000",
  35186=>"00000000",
  35187=>"11111111",
  35188=>"11111110",
  35189=>"11111111",
  35190=>"11111110",
  35191=>"00000010",
  35192=>"00000001",
  35193=>"11111101",
  35194=>"11111101",
  35195=>"00000001",
  35196=>"11111101",
  35197=>"00000100",
  35198=>"11111110",
  35199=>"11111111",
  35200=>"11111110",
  35201=>"00000011",
  35202=>"11111101",
  35203=>"00000001",
  35204=>"00000010",
  35205=>"11111111",
  35206=>"11111111",
  35207=>"00000011",
  35208=>"11111101",
  35209=>"11111101",
  35210=>"00000000",
  35211=>"11111111",
  35212=>"11111111",
  35213=>"00000010",
  35214=>"11111101",
  35215=>"00000110",
  35216=>"00000001",
  35217=>"11111111",
  35218=>"11111110",
  35219=>"00000010",
  35220=>"00000100",
  35221=>"00000000",
  35222=>"00000001",
  35223=>"00000001",
  35224=>"00000001",
  35225=>"00000010",
  35226=>"11111110",
  35227=>"00000001",
  35228=>"00000001",
  35229=>"11111101",
  35230=>"11111101",
  35231=>"11111101",
  35232=>"11111101",
  35233=>"11111110",
  35234=>"00000001",
  35235=>"11111101",
  35236=>"00000000",
  35237=>"00000011",
  35238=>"00000000",
  35239=>"00000011",
  35240=>"00000010",
  35241=>"11111111",
  35242=>"11111110",
  35243=>"11111110",
  35244=>"11111111",
  35245=>"00000000",
  35246=>"11111101",
  35247=>"00000011",
  35248=>"00000101",
  35249=>"11111110",
  35250=>"00000010",
  35251=>"00000010",
  35252=>"00000010",
  35253=>"11111111",
  35254=>"11111110",
  35255=>"11111111",
  35256=>"00000000",
  35257=>"00000000",
  35258=>"00000010",
  35259=>"11111111",
  35260=>"00000001",
  35261=>"00000011",
  35262=>"11111110",
  35263=>"00000010",
  35264=>"11111011",
  35265=>"00000101",
  35266=>"00000101",
  35267=>"11111111",
  35268=>"00000000",
  35269=>"00000000",
  35270=>"00000001",
  35271=>"00000000",
  35272=>"11111110",
  35273=>"00000000",
  35274=>"00000011",
  35275=>"00000000",
  35276=>"00000000",
  35277=>"11111101",
  35278=>"00000000",
  35279=>"11111111",
  35280=>"11111111",
  35281=>"11111110",
  35282=>"11111110",
  35283=>"11111101",
  35284=>"00000010",
  35285=>"11111110",
  35286=>"11111110",
  35287=>"11111111",
  35288=>"00000011",
  35289=>"11111101",
  35290=>"11111110",
  35291=>"11111111",
  35292=>"00000101",
  35293=>"00000000",
  35294=>"00000001",
  35295=>"11111011",
  35296=>"11111111",
  35297=>"00000000",
  35298=>"00000001",
  35299=>"00000001",
  35300=>"11111101",
  35301=>"11111101",
  35302=>"11111111",
  35303=>"11111110",
  35304=>"00000010",
  35305=>"00000001",
  35306=>"11111111",
  35307=>"11111101",
  35308=>"11111111",
  35309=>"00000000",
  35310=>"11111111",
  35311=>"00000010",
  35312=>"00000100",
  35313=>"00000000",
  35314=>"00000011",
  35315=>"00000010",
  35316=>"00000010",
  35317=>"11111111",
  35318=>"00000011",
  35319=>"00000100",
  35320=>"11111110",
  35321=>"11111111",
  35322=>"00000000",
  35323=>"11111110",
  35324=>"00000010",
  35325=>"00000100",
  35326=>"11111111",
  35327=>"11111101",
  35328=>"11111111",
  35329=>"00000110",
  35330=>"00000011",
  35331=>"11111111",
  35332=>"11111100",
  35333=>"00000001",
  35334=>"00000001",
  35335=>"00000011",
  35336=>"00000011",
  35337=>"00000100",
  35338=>"11111110",
  35339=>"00000000",
  35340=>"00000010",
  35341=>"00000010",
  35342=>"11111110",
  35343=>"00000100",
  35344=>"11111110",
  35345=>"00000000",
  35346=>"00000001",
  35347=>"11111101",
  35348=>"00000010",
  35349=>"00000000",
  35350=>"11111101",
  35351=>"00000010",
  35352=>"00000001",
  35353=>"00000000",
  35354=>"11111101",
  35355=>"11111111",
  35356=>"00000001",
  35357=>"00000001",
  35358=>"00000001",
  35359=>"00000011",
  35360=>"00000000",
  35361=>"00000000",
  35362=>"11111110",
  35363=>"11111111",
  35364=>"11111101",
  35365=>"00000001",
  35366=>"11111111",
  35367=>"11111101",
  35368=>"00000011",
  35369=>"00000000",
  35370=>"00000001",
  35371=>"00000001",
  35372=>"11111110",
  35373=>"11111101",
  35374=>"11111110",
  35375=>"00000000",
  35376=>"00000011",
  35377=>"11111100",
  35378=>"00000001",
  35379=>"11111110",
  35380=>"11111111",
  35381=>"00000110",
  35382=>"11111111",
  35383=>"11111111",
  35384=>"11111111",
  35385=>"00000000",
  35386=>"00000011",
  35387=>"00000010",
  35388=>"11111110",
  35389=>"00000000",
  35390=>"00000011",
  35391=>"00000000",
  35392=>"11111100",
  35393=>"11111101",
  35394=>"11111110",
  35395=>"11111110",
  35396=>"11111101",
  35397=>"00000000",
  35398=>"11111101",
  35399=>"11111101",
  35400=>"11111111",
  35401=>"00000010",
  35402=>"00000101",
  35403=>"00000011",
  35404=>"00000011",
  35405=>"00000001",
  35406=>"11111110",
  35407=>"00000000",
  35408=>"11111111",
  35409=>"00000010",
  35410=>"00000000",
  35411=>"00000010",
  35412=>"00000000",
  35413=>"00000001",
  35414=>"11111111",
  35415=>"11111100",
  35416=>"11111110",
  35417=>"11111101",
  35418=>"00000010",
  35419=>"11111110",
  35420=>"00000011",
  35421=>"00000001",
  35422=>"00000010",
  35423=>"00000001",
  35424=>"11111101",
  35425=>"00000100",
  35426=>"00000100",
  35427=>"11111101",
  35428=>"00000001",
  35429=>"11111101",
  35430=>"11111110",
  35431=>"11111101",
  35432=>"00000010",
  35433=>"11111101",
  35434=>"00000010",
  35435=>"00000011",
  35436=>"00000000",
  35437=>"11111111",
  35438=>"00000010",
  35439=>"00000010",
  35440=>"11111101",
  35441=>"11111111",
  35442=>"11111111",
  35443=>"00000011",
  35444=>"11111100",
  35445=>"00000010",
  35446=>"00000100",
  35447=>"11111110",
  35448=>"00000100",
  35449=>"00000010",
  35450=>"11111101",
  35451=>"00000000",
  35452=>"00000000",
  35453=>"11111110",
  35454=>"00000010",
  35455=>"00000001",
  35456=>"11111101",
  35457=>"11111111",
  35458=>"00000101",
  35459=>"00000111",
  35460=>"11111101",
  35461=>"00000000",
  35462=>"11111110",
  35463=>"11111101",
  35464=>"00000000",
  35465=>"00000101",
  35466=>"00000001",
  35467=>"00000010",
  35468=>"11111101",
  35469=>"00000000",
  35470=>"00000001",
  35471=>"11111110",
  35472=>"00000011",
  35473=>"11111111",
  35474=>"11111100",
  35475=>"00000010",
  35476=>"11111110",
  35477=>"11111101",
  35478=>"11111101",
  35479=>"11111101",
  35480=>"00000001",
  35481=>"11111111",
  35482=>"00000000",
  35483=>"00000000",
  35484=>"11111111",
  35485=>"00000011",
  35486=>"11111101",
  35487=>"00000000",
  35488=>"11111101",
  35489=>"11111101",
  35490=>"11111111",
  35491=>"11111111",
  35492=>"11111111",
  35493=>"00000000",
  35494=>"11111111",
  35495=>"00000001",
  35496=>"11111111",
  35497=>"00000001",
  35498=>"00000011",
  35499=>"00000000",
  35500=>"00000000",
  35501=>"00000001",
  35502=>"00000010",
  35503=>"00000000",
  35504=>"00000101",
  35505=>"00000100",
  35506=>"11111111",
  35507=>"11111101",
  35508=>"00000010",
  35509=>"00000010",
  35510=>"11111110",
  35511=>"00000100",
  35512=>"00000011",
  35513=>"00000001",
  35514=>"11111111",
  35515=>"11111111",
  35516=>"00000011",
  35517=>"00000000",
  35518=>"11111100",
  35519=>"00000001",
  35520=>"00000000",
  35521=>"11111111",
  35522=>"11111101",
  35523=>"11111101",
  35524=>"11111101",
  35525=>"11111101",
  35526=>"00000011",
  35527=>"00000000",
  35528=>"11111111",
  35529=>"00000010",
  35530=>"11111101",
  35531=>"00000001",
  35532=>"11111111",
  35533=>"00000000",
  35534=>"11111101",
  35535=>"11111101",
  35536=>"00000010",
  35537=>"11111111",
  35538=>"00000000",
  35539=>"00000110",
  35540=>"00000001",
  35541=>"11111110",
  35542=>"00000000",
  35543=>"00000000",
  35544=>"11111100",
  35545=>"00000001",
  35546=>"11111110",
  35547=>"00000001",
  35548=>"11111111",
  35549=>"11111110",
  35550=>"00000001",
  35551=>"00000101",
  35552=>"00000001",
  35553=>"11111111",
  35554=>"00000010",
  35555=>"00000001",
  35556=>"00000010",
  35557=>"00000001",
  35558=>"11111111",
  35559=>"11111100",
  35560=>"00000001",
  35561=>"00000000",
  35562=>"00000011",
  35563=>"11111101",
  35564=>"11111110",
  35565=>"00000010",
  35566=>"11111110",
  35567=>"11111101",
  35568=>"11111111",
  35569=>"00000000",
  35570=>"00000011",
  35571=>"11111111",
  35572=>"00000101",
  35573=>"00000010",
  35574=>"11111100",
  35575=>"00000011",
  35576=>"00000001",
  35577=>"11111101",
  35578=>"11111111",
  35579=>"00000101",
  35580=>"11111111",
  35581=>"11111101",
  35582=>"00000011",
  35583=>"11111110",
  35584=>"11111111",
  35585=>"00000001",
  35586=>"11111101",
  35587=>"11111111",
  35588=>"00000000",
  35589=>"11111111",
  35590=>"11111111",
  35591=>"11111110",
  35592=>"00000111",
  35593=>"00000000",
  35594=>"00000000",
  35595=>"11111101",
  35596=>"11111110",
  35597=>"00000000",
  35598=>"11111110",
  35599=>"00000001",
  35600=>"00000001",
  35601=>"11111110",
  35602=>"00000010",
  35603=>"00000001",
  35604=>"00000001",
  35605=>"00000001",
  35606=>"00000001",
  35607=>"11111100",
  35608=>"11111101",
  35609=>"11111111",
  35610=>"00000011",
  35611=>"00000001",
  35612=>"11111101",
  35613=>"11111111",
  35614=>"00000110",
  35615=>"00000000",
  35616=>"11111101",
  35617=>"00000010",
  35618=>"11111101",
  35619=>"00000010",
  35620=>"11111111",
  35621=>"11111110",
  35622=>"11111110",
  35623=>"00000010",
  35624=>"11111111",
  35625=>"11111101",
  35626=>"11111111",
  35627=>"00000010",
  35628=>"00000001",
  35629=>"00000010",
  35630=>"00000001",
  35631=>"00000001",
  35632=>"00000011",
  35633=>"00000001",
  35634=>"00000000",
  35635=>"00000001",
  35636=>"00000000",
  35637=>"11111101",
  35638=>"00000000",
  35639=>"00000010",
  35640=>"11111110",
  35641=>"00000000",
  35642=>"11111111",
  35643=>"11111111",
  35644=>"00000011",
  35645=>"11111110",
  35646=>"11111110",
  35647=>"11111111",
  35648=>"11111101",
  35649=>"11111110",
  35650=>"11111100",
  35651=>"11111111",
  35652=>"00000000",
  35653=>"11111100",
  35654=>"00000100",
  35655=>"11111110",
  35656=>"00000001",
  35657=>"11111110",
  35658=>"11111110",
  35659=>"11111101",
  35660=>"00000011",
  35661=>"00000010",
  35662=>"11111110",
  35663=>"00000001",
  35664=>"00000000",
  35665=>"00000000",
  35666=>"11111110",
  35667=>"11111100",
  35668=>"00000010",
  35669=>"00000001",
  35670=>"00000011",
  35671=>"00000010",
  35672=>"11111101",
  35673=>"11111110",
  35674=>"11111111",
  35675=>"11111110",
  35676=>"11111111",
  35677=>"00000010",
  35678=>"11111111",
  35679=>"11111111",
  35680=>"00000100",
  35681=>"00000000",
  35682=>"00000001",
  35683=>"11111111",
  35684=>"00000010",
  35685=>"00000000",
  35686=>"00000001",
  35687=>"11111100",
  35688=>"00000001",
  35689=>"11111100",
  35690=>"11111111",
  35691=>"00000000",
  35692=>"00000010",
  35693=>"00000001",
  35694=>"11111111",
  35695=>"11111111",
  35696=>"00000010",
  35697=>"00000010",
  35698=>"00000000",
  35699=>"00000001",
  35700=>"00000001",
  35701=>"00000000",
  35702=>"00000000",
  35703=>"11111101",
  35704=>"00000010",
  35705=>"11111101",
  35706=>"11111111",
  35707=>"00000010",
  35708=>"00000000",
  35709=>"00000010",
  35710=>"11111110",
  35711=>"00000000",
  35712=>"00000000",
  35713=>"00000100",
  35714=>"00000011",
  35715=>"11111100",
  35716=>"00000000",
  35717=>"00000001",
  35718=>"11111110",
  35719=>"11111110",
  35720=>"00000110",
  35721=>"11111111",
  35722=>"00000010",
  35723=>"00000000",
  35724=>"00000001",
  35725=>"00000000",
  35726=>"11111101",
  35727=>"00000010",
  35728=>"11111101",
  35729=>"00000011",
  35730=>"00000001",
  35731=>"00000001",
  35732=>"11111111",
  35733=>"00000111",
  35734=>"00000001",
  35735=>"00000010",
  35736=>"00000010",
  35737=>"11111111",
  35738=>"00000001",
  35739=>"00000000",
  35740=>"11111110",
  35741=>"00000101",
  35742=>"11111100",
  35743=>"00000001",
  35744=>"00000011",
  35745=>"11111110",
  35746=>"00000110",
  35747=>"00000000",
  35748=>"00000100",
  35749=>"11111101",
  35750=>"00000010",
  35751=>"00000100",
  35752=>"00000001",
  35753=>"00000001",
  35754=>"00000000",
  35755=>"00000000",
  35756=>"00000010",
  35757=>"11111111",
  35758=>"11111110",
  35759=>"00000011",
  35760=>"11111110",
  35761=>"00000000",
  35762=>"00000001",
  35763=>"11111111",
  35764=>"00000000",
  35765=>"00000100",
  35766=>"11111101",
  35767=>"00000000",
  35768=>"11111110",
  35769=>"00000001",
  35770=>"11111101",
  35771=>"11111110",
  35772=>"00000011",
  35773=>"11111110",
  35774=>"11111110",
  35775=>"00000001",
  35776=>"00000000",
  35777=>"00000010",
  35778=>"11111111",
  35779=>"11111111",
  35780=>"11111101",
  35781=>"11111101",
  35782=>"00000100",
  35783=>"00000001",
  35784=>"11111111",
  35785=>"11111110",
  35786=>"11111110",
  35787=>"00000000",
  35788=>"00000001",
  35789=>"11111111",
  35790=>"11111111",
  35791=>"00000100",
  35792=>"00000001",
  35793=>"11111110",
  35794=>"00000000",
  35795=>"00000001",
  35796=>"11111110",
  35797=>"00000000",
  35798=>"00000010",
  35799=>"11111101",
  35800=>"11111111",
  35801=>"11111101",
  35802=>"00000000",
  35803=>"11111111",
  35804=>"11111111",
  35805=>"00000001",
  35806=>"11111111",
  35807=>"00000001",
  35808=>"00000001",
  35809=>"00000000",
  35810=>"00000011",
  35811=>"00000001",
  35812=>"00000000",
  35813=>"00000100",
  35814=>"11111110",
  35815=>"11111110",
  35816=>"00000000",
  35817=>"11111111",
  35818=>"00000001",
  35819=>"00000100",
  35820=>"00000000",
  35821=>"00000010",
  35822=>"00000011",
  35823=>"00000000",
  35824=>"11111110",
  35825=>"11111111",
  35826=>"00000010",
  35827=>"11111101",
  35828=>"00000001",
  35829=>"00000100",
  35830=>"00000000",
  35831=>"11111101",
  35832=>"00000001",
  35833=>"00000011",
  35834=>"11111111",
  35835=>"11111101",
  35836=>"00000000",
  35837=>"00000000",
  35838=>"00000001",
  35839=>"00000101",
  35840=>"11111110",
  35841=>"00000001",
  35842=>"00000000",
  35843=>"00000010",
  35844=>"00000000",
  35845=>"00000011",
  35846=>"00000001",
  35847=>"00000010",
  35848=>"00000010",
  35849=>"11111110",
  35850=>"00000011",
  35851=>"00000000",
  35852=>"11111111",
  35853=>"00000001",
  35854=>"00000100",
  35855=>"11111111",
  35856=>"11111110",
  35857=>"00000001",
  35858=>"00000000",
  35859=>"00000110",
  35860=>"11111110",
  35861=>"00000010",
  35862=>"11111101",
  35863=>"11111110",
  35864=>"00000100",
  35865=>"11111111",
  35866=>"11111111",
  35867=>"11111101",
  35868=>"11111111",
  35869=>"11111101",
  35870=>"11111101",
  35871=>"11111111",
  35872=>"00000100",
  35873=>"00000000",
  35874=>"11111111",
  35875=>"00000000",
  35876=>"11111111",
  35877=>"11111101",
  35878=>"00000000",
  35879=>"11111111",
  35880=>"00000000",
  35881=>"11111110",
  35882=>"00000001",
  35883=>"00000001",
  35884=>"11111110",
  35885=>"00000000",
  35886=>"11111110",
  35887=>"11111110",
  35888=>"11111111",
  35889=>"00000010",
  35890=>"00000010",
  35891=>"00000001",
  35892=>"00000011",
  35893=>"11111111",
  35894=>"00000011",
  35895=>"00000001",
  35896=>"00000011",
  35897=>"11111110",
  35898=>"00000010",
  35899=>"11111110",
  35900=>"11111111",
  35901=>"00000010",
  35902=>"00000010",
  35903=>"11111110",
  35904=>"00000000",
  35905=>"11111110",
  35906=>"00000010",
  35907=>"00000010",
  35908=>"11111111",
  35909=>"00000000",
  35910=>"11111101",
  35911=>"00000110",
  35912=>"00000101",
  35913=>"00000001",
  35914=>"00000001",
  35915=>"11111110",
  35916=>"11111111",
  35917=>"00000011",
  35918=>"00000000",
  35919=>"00000000",
  35920=>"00000011",
  35921=>"00000001",
  35922=>"11111110",
  35923=>"00000100",
  35924=>"11111110",
  35925=>"11111111",
  35926=>"00000000",
  35927=>"11111101",
  35928=>"00000000",
  35929=>"11111111",
  35930=>"00000000",
  35931=>"00000011",
  35932=>"11111111",
  35933=>"11111101",
  35934=>"11111110",
  35935=>"11111100",
  35936=>"11111110",
  35937=>"11111110",
  35938=>"00000000",
  35939=>"00000010",
  35940=>"00000001",
  35941=>"00000010",
  35942=>"00000000",
  35943=>"00000001",
  35944=>"00000010",
  35945=>"00000101",
  35946=>"11111100",
  35947=>"11111110",
  35948=>"00000010",
  35949=>"00000001",
  35950=>"00000001",
  35951=>"00000010",
  35952=>"00000000",
  35953=>"11111110",
  35954=>"00000000",
  35955=>"00000011",
  35956=>"11111111",
  35957=>"11111111",
  35958=>"00000001",
  35959=>"11111110",
  35960=>"00000001",
  35961=>"00000000",
  35962=>"00000110",
  35963=>"11111111",
  35964=>"00000001",
  35965=>"11111110",
  35966=>"11111111",
  35967=>"11111110",
  35968=>"11111110",
  35969=>"11111111",
  35970=>"00000011",
  35971=>"11111110",
  35972=>"00000000",
  35973=>"00000010",
  35974=>"00000011",
  35975=>"00000011",
  35976=>"00000010",
  35977=>"00000011",
  35978=>"00000101",
  35979=>"00000001",
  35980=>"00000011",
  35981=>"00000000",
  35982=>"00000001",
  35983=>"00000010",
  35984=>"00000010",
  35985=>"11111101",
  35986=>"00000000",
  35987=>"11111111",
  35988=>"11111111",
  35989=>"00000100",
  35990=>"11111111",
  35991=>"11111111",
  35992=>"00000010",
  35993=>"11111110",
  35994=>"00000001",
  35995=>"00000011",
  35996=>"00000000",
  35997=>"11111101",
  35998=>"00000001",
  35999=>"11111111",
  36000=>"11111110",
  36001=>"11111101",
  36002=>"11111101",
  36003=>"11111101",
  36004=>"00000011",
  36005=>"11111101",
  36006=>"11111100",
  36007=>"00000000",
  36008=>"11111101",
  36009=>"11111101",
  36010=>"11111111",
  36011=>"00000001",
  36012=>"00000010",
  36013=>"00000011",
  36014=>"00000100",
  36015=>"00000000",
  36016=>"11111110",
  36017=>"00000010",
  36018=>"00000100",
  36019=>"00000001",
  36020=>"00000100",
  36021=>"11111111",
  36022=>"11111110",
  36023=>"00000110",
  36024=>"00000000",
  36025=>"00000001",
  36026=>"11111110",
  36027=>"11111110",
  36028=>"00000000",
  36029=>"00000010",
  36030=>"11111110",
  36031=>"00000011",
  36032=>"00000010",
  36033=>"00000000",
  36034=>"11111110",
  36035=>"00000100",
  36036=>"00000000",
  36037=>"11111111",
  36038=>"00000001",
  36039=>"00000000",
  36040=>"11111110",
  36041=>"11111100",
  36042=>"11111110",
  36043=>"00000010",
  36044=>"11111100",
  36045=>"00000001",
  36046=>"00000001",
  36047=>"11111110",
  36048=>"00000000",
  36049=>"00000000",
  36050=>"00000010",
  36051=>"11111111",
  36052=>"00000010",
  36053=>"00000100",
  36054=>"11111101",
  36055=>"00000010",
  36056=>"00000001",
  36057=>"11111111",
  36058=>"00000010",
  36059=>"00000101",
  36060=>"11111110",
  36061=>"11111101",
  36062=>"11111111",
  36063=>"11111100",
  36064=>"00000011",
  36065=>"00000001",
  36066=>"00000010",
  36067=>"11111110",
  36068=>"00000110",
  36069=>"11111111",
  36070=>"00000110",
  36071=>"11111110",
  36072=>"00000000",
  36073=>"11111101",
  36074=>"11111110",
  36075=>"00000000",
  36076=>"00000010",
  36077=>"00000001",
  36078=>"00000010",
  36079=>"00000001",
  36080=>"11111110",
  36081=>"00000000",
  36082=>"11111101",
  36083=>"11111110",
  36084=>"00000000",
  36085=>"11111101",
  36086=>"00000001",
  36087=>"11111111",
  36088=>"00000001",
  36089=>"00000001",
  36090=>"00000100",
  36091=>"00000001",
  36092=>"00000100",
  36093=>"11111110",
  36094=>"00000000",
  36095=>"00000001",
  36096=>"00000001",
  36097=>"00000000",
  36098=>"00000100",
  36099=>"00000010",
  36100=>"11111101",
  36101=>"00000010",
  36102=>"00000010",
  36103=>"00000001",
  36104=>"00000010",
  36105=>"00000010",
  36106=>"11111111",
  36107=>"00000001",
  36108=>"00000000",
  36109=>"00000000",
  36110=>"11111110",
  36111=>"00000011",
  36112=>"11111111",
  36113=>"11111101",
  36114=>"00000011",
  36115=>"11111110",
  36116=>"11111110",
  36117=>"00000000",
  36118=>"11111111",
  36119=>"00000011",
  36120=>"11111111",
  36121=>"11111110",
  36122=>"00000001",
  36123=>"00000010",
  36124=>"00000100",
  36125=>"00000000",
  36126=>"11111111",
  36127=>"11111110",
  36128=>"11111101",
  36129=>"11111101",
  36130=>"00000011",
  36131=>"11111101",
  36132=>"00000010",
  36133=>"00000010",
  36134=>"00000000",
  36135=>"00000000",
  36136=>"00000100",
  36137=>"00000001",
  36138=>"11111101",
  36139=>"00000000",
  36140=>"11111111",
  36141=>"11111110",
  36142=>"11111100",
  36143=>"00000001",
  36144=>"11111110",
  36145=>"00000010",
  36146=>"00000010",
  36147=>"00000001",
  36148=>"00000000",
  36149=>"11111110",
  36150=>"00000000",
  36151=>"00000001",
  36152=>"00000001",
  36153=>"11111111",
  36154=>"00000001",
  36155=>"00000010",
  36156=>"00000000",
  36157=>"00000011",
  36158=>"11111111",
  36159=>"00000010",
  36160=>"11111110",
  36161=>"11111110",
  36162=>"00000011",
  36163=>"00000010",
  36164=>"11111101",
  36165=>"00000000",
  36166=>"11111110",
  36167=>"00000000",
  36168=>"11111110",
  36169=>"11111111",
  36170=>"00000101",
  36171=>"00000000",
  36172=>"11111111",
  36173=>"00000100",
  36174=>"11111111",
  36175=>"00000001",
  36176=>"00000100",
  36177=>"11111110",
  36178=>"00000001",
  36179=>"11111111",
  36180=>"11111110",
  36181=>"11111110",
  36182=>"11111101",
  36183=>"00000001",
  36184=>"11111111",
  36185=>"00000000",
  36186=>"00000001",
  36187=>"11111110",
  36188=>"00000001",
  36189=>"00000011",
  36190=>"11111101",
  36191=>"00000010",
  36192=>"11111110",
  36193=>"11111100",
  36194=>"00000010",
  36195=>"11111111",
  36196=>"00000010",
  36197=>"00000001",
  36198=>"11111100",
  36199=>"00000001",
  36200=>"11111110",
  36201=>"00000010",
  36202=>"11111111",
  36203=>"00000000",
  36204=>"00000001",
  36205=>"00000010",
  36206=>"00000000",
  36207=>"00000010",
  36208=>"00000001",
  36209=>"11111101",
  36210=>"11111110",
  36211=>"00000001",
  36212=>"11111110",
  36213=>"11111101",
  36214=>"00000000",
  36215=>"00000000",
  36216=>"00000011",
  36217=>"11111111",
  36218=>"00000001",
  36219=>"11111111",
  36220=>"11111110",
  36221=>"11111101",
  36222=>"11111110",
  36223=>"11111111",
  36224=>"11111111",
  36225=>"00000011",
  36226=>"00000001",
  36227=>"00000001",
  36228=>"00000011",
  36229=>"00000001",
  36230=>"00000010",
  36231=>"00000010",
  36232=>"00000001",
  36233=>"11111100",
  36234=>"11111111",
  36235=>"00000010",
  36236=>"00000001",
  36237=>"11111110",
  36238=>"11111101",
  36239=>"11111101",
  36240=>"11111111",
  36241=>"11111111",
  36242=>"11111101",
  36243=>"00000000",
  36244=>"00000000",
  36245=>"00000000",
  36246=>"11111110",
  36247=>"11111110",
  36248=>"00000001",
  36249=>"11111110",
  36250=>"00000000",
  36251=>"11111110",
  36252=>"11111110",
  36253=>"00000001",
  36254=>"00000000",
  36255=>"11111111",
  36256=>"00000000",
  36257=>"00000000",
  36258=>"11111110",
  36259=>"11111110",
  36260=>"11111111",
  36261=>"00000010",
  36262=>"11111110",
  36263=>"00000001",
  36264=>"00000100",
  36265=>"00000000",
  36266=>"11111110",
  36267=>"11111111",
  36268=>"00000100",
  36269=>"00000100",
  36270=>"00000011",
  36271=>"00000010",
  36272=>"11111110",
  36273=>"00000001",
  36274=>"00000001",
  36275=>"00000001",
  36276=>"11111110",
  36277=>"11111111",
  36278=>"11111100",
  36279=>"11111101",
  36280=>"00000000",
  36281=>"00000001",
  36282=>"11111110",
  36283=>"00000001",
  36284=>"00000001",
  36285=>"00000000",
  36286=>"00000101",
  36287=>"11111111",
  36288=>"11111101",
  36289=>"11111110",
  36290=>"00000001",
  36291=>"11111101",
  36292=>"11111101",
  36293=>"00000001",
  36294=>"11111101",
  36295=>"11111101",
  36296=>"11111111",
  36297=>"11111111",
  36298=>"00000000",
  36299=>"11111110",
  36300=>"11111110",
  36301=>"11111111",
  36302=>"11111101",
  36303=>"00000011",
  36304=>"11111101",
  36305=>"00000010",
  36306=>"11111101",
  36307=>"11111110",
  36308=>"11111101",
  36309=>"11111111",
  36310=>"00000000",
  36311=>"00000001",
  36312=>"00000010",
  36313=>"11111111",
  36314=>"11111110",
  36315=>"00000100",
  36316=>"11111110",
  36317=>"11111110",
  36318=>"00000010",
  36319=>"11111111",
  36320=>"11111111",
  36321=>"00000000",
  36322=>"00000000",
  36323=>"00000000",
  36324=>"11111111",
  36325=>"00000000",
  36326=>"00000101",
  36327=>"00000001",
  36328=>"11111101",
  36329=>"11111111",
  36330=>"00000100",
  36331=>"11111111",
  36332=>"00000001",
  36333=>"11111101",
  36334=>"00000001",
  36335=>"00000001",
  36336=>"00000001",
  36337=>"00000010",
  36338=>"00000010",
  36339=>"00000101",
  36340=>"00000010",
  36341=>"00000001",
  36342=>"11111111",
  36343=>"00000010",
  36344=>"11111101",
  36345=>"00000010",
  36346=>"00000000",
  36347=>"11111111",
  36348=>"00000001",
  36349=>"00000001",
  36350=>"00000100",
  36351=>"11111111",
  36352=>"11111110",
  36353=>"11111111",
  36354=>"00000001",
  36355=>"00000000",
  36356=>"11111110",
  36357=>"11111111",
  36358=>"00000001",
  36359=>"11111101",
  36360=>"00000010",
  36361=>"11111110",
  36362=>"00000000",
  36363=>"11111111",
  36364=>"11111111",
  36365=>"11111110",
  36366=>"00000100",
  36367=>"11111110",
  36368=>"11111101",
  36369=>"00000100",
  36370=>"00000101",
  36371=>"11111101",
  36372=>"11111101",
  36373=>"00000000",
  36374=>"00000011",
  36375=>"11111110",
  36376=>"00000100",
  36377=>"00000000",
  36378=>"00000001",
  36379=>"00000001",
  36380=>"00000100",
  36381=>"00000001",
  36382=>"00000011",
  36383=>"00000010",
  36384=>"00001000",
  36385=>"00000001",
  36386=>"11111111",
  36387=>"00000010",
  36388=>"11111111",
  36389=>"00000100",
  36390=>"00000010",
  36391=>"00000101",
  36392=>"00000100",
  36393=>"00000000",
  36394=>"11111110",
  36395=>"11111101",
  36396=>"00000000",
  36397=>"11111110",
  36398=>"00000001",
  36399=>"00000000",
  36400=>"11111100",
  36401=>"00000000",
  36402=>"00000001",
  36403=>"11111110",
  36404=>"00000011",
  36405=>"00000001",
  36406=>"11111111",
  36407=>"00000001",
  36408=>"11111101",
  36409=>"11111110",
  36410=>"00000000",
  36411=>"11111110",
  36412=>"00000000",
  36413=>"11111110",
  36414=>"00000011",
  36415=>"00000000",
  36416=>"11111101",
  36417=>"11111110",
  36418=>"11111101",
  36419=>"00000000",
  36420=>"00000010",
  36421=>"11111110",
  36422=>"11111111",
  36423=>"00000011",
  36424=>"00000010",
  36425=>"00000001",
  36426=>"11111100",
  36427=>"11111111",
  36428=>"00000001",
  36429=>"00000000",
  36430=>"11111101",
  36431=>"00000010",
  36432=>"00000001",
  36433=>"00000010",
  36434=>"11111111",
  36435=>"00000000",
  36436=>"00000000",
  36437=>"00000001",
  36438=>"11111110",
  36439=>"00000001",
  36440=>"00000000",
  36441=>"00000101",
  36442=>"00000011",
  36443=>"11111111",
  36444=>"11111110",
  36445=>"00000001",
  36446=>"00000001",
  36447=>"11111111",
  36448=>"11111111",
  36449=>"11111110",
  36450=>"00000001",
  36451=>"11111101",
  36452=>"00000000",
  36453=>"11111110",
  36454=>"00000010",
  36455=>"11111101",
  36456=>"00000010",
  36457=>"00000100",
  36458=>"11111111",
  36459=>"00000010",
  36460=>"11111111",
  36461=>"00000000",
  36462=>"00000001",
  36463=>"11111111",
  36464=>"00000000",
  36465=>"00000001",
  36466=>"00000001",
  36467=>"11111101",
  36468=>"11111111",
  36469=>"00000101",
  36470=>"00000001",
  36471=>"11111100",
  36472=>"00000010",
  36473=>"00000001",
  36474=>"00000000",
  36475=>"11111111",
  36476=>"00000001",
  36477=>"11111111",
  36478=>"11111110",
  36479=>"00000011",
  36480=>"00000000",
  36481=>"00000000",
  36482=>"11111101",
  36483=>"00000011",
  36484=>"00000011",
  36485=>"11111101",
  36486=>"00000010",
  36487=>"00000010",
  36488=>"11111101",
  36489=>"11111111",
  36490=>"11111111",
  36491=>"11111111",
  36492=>"00000010",
  36493=>"11111111",
  36494=>"00000001",
  36495=>"11111110",
  36496=>"00000011",
  36497=>"11111111",
  36498=>"11111110",
  36499=>"11111111",
  36500=>"11111110",
  36501=>"11111110",
  36502=>"11111111",
  36503=>"11111110",
  36504=>"00000001",
  36505=>"00000101",
  36506=>"11111110",
  36507=>"00000000",
  36508=>"11111101",
  36509=>"00000010",
  36510=>"11111111",
  36511=>"00000000",
  36512=>"11111110",
  36513=>"11111111",
  36514=>"00000000",
  36515=>"00000001",
  36516=>"00000001",
  36517=>"11111110",
  36518=>"00000000",
  36519=>"00000011",
  36520=>"00000000",
  36521=>"11111111",
  36522=>"11111101",
  36523=>"11111110",
  36524=>"11111110",
  36525=>"00000001",
  36526=>"00000000",
  36527=>"11111101",
  36528=>"11111101",
  36529=>"00000010",
  36530=>"00000000",
  36531=>"00000001",
  36532=>"00000011",
  36533=>"00000010",
  36534=>"00000000",
  36535=>"00000001",
  36536=>"00000001",
  36537=>"00000001",
  36538=>"11111111",
  36539=>"00000011",
  36540=>"00000000",
  36541=>"00000001",
  36542=>"11111100",
  36543=>"00000000",
  36544=>"00000000",
  36545=>"11111111",
  36546=>"00000000",
  36547=>"00000101",
  36548=>"00000001",
  36549=>"11111101",
  36550=>"00000000",
  36551=>"00000001",
  36552=>"11111110",
  36553=>"00000010",
  36554=>"11111110",
  36555=>"00000000",
  36556=>"00000000",
  36557=>"00000001",
  36558=>"00000000",
  36559=>"00000001",
  36560=>"11111111",
  36561=>"00000011",
  36562=>"11111101",
  36563=>"11111101",
  36564=>"00000010",
  36565=>"00000000",
  36566=>"00000010",
  36567=>"11111111",
  36568=>"11111110",
  36569=>"11111101",
  36570=>"00000001",
  36571=>"00000011",
  36572=>"00000001",
  36573=>"00000010",
  36574=>"00000001",
  36575=>"11111100",
  36576=>"00000010",
  36577=>"00000011",
  36578=>"00000100",
  36579=>"11111110",
  36580=>"11111100",
  36581=>"00000010",
  36582=>"11111101",
  36583=>"11111110",
  36584=>"11111111",
  36585=>"00000001",
  36586=>"00000000",
  36587=>"00000010",
  36588=>"11111101",
  36589=>"00000001",
  36590=>"00000001",
  36591=>"00000001",
  36592=>"11111110",
  36593=>"11111111",
  36594=>"00000010",
  36595=>"00000001",
  36596=>"11111110",
  36597=>"11111101",
  36598=>"11111101",
  36599=>"00000000",
  36600=>"11111110",
  36601=>"00000011",
  36602=>"11111101",
  36603=>"11111101",
  36604=>"11111111",
  36605=>"00000011",
  36606=>"11111101",
  36607=>"11111111",
  36608=>"11111110",
  36609=>"11111101",
  36610=>"00000011",
  36611=>"00000001",
  36612=>"00000011",
  36613=>"11111110",
  36614=>"00000010",
  36615=>"11111101",
  36616=>"11111111",
  36617=>"11111111",
  36618=>"00000010",
  36619=>"11111111",
  36620=>"00000000",
  36621=>"00000000",
  36622=>"00000101",
  36623=>"11111110",
  36624=>"00000010",
  36625=>"00000000",
  36626=>"11111101",
  36627=>"11111101",
  36628=>"00000001",
  36629=>"11111101",
  36630=>"11111111",
  36631=>"00000011",
  36632=>"00000100",
  36633=>"00000000",
  36634=>"00000100",
  36635=>"11111111",
  36636=>"11111100",
  36637=>"11111110",
  36638=>"00000001",
  36639=>"11111111",
  36640=>"11111101",
  36641=>"00000100",
  36642=>"00000001",
  36643=>"00000001",
  36644=>"00000011",
  36645=>"11111111",
  36646=>"00000011",
  36647=>"00000000",
  36648=>"00000001",
  36649=>"00000100",
  36650=>"00000001",
  36651=>"00000000",
  36652=>"11111110",
  36653=>"00000010",
  36654=>"00000000",
  36655=>"11111110",
  36656=>"00000000",
  36657=>"11111111",
  36658=>"11111111",
  36659=>"11111101",
  36660=>"00000001",
  36661=>"00000110",
  36662=>"11111101",
  36663=>"11111111",
  36664=>"11111111",
  36665=>"11111110",
  36666=>"00000010",
  36667=>"11111110",
  36668=>"11111101",
  36669=>"00000000",
  36670=>"00000001",
  36671=>"11111110",
  36672=>"11111110",
  36673=>"11111111",
  36674=>"11111101",
  36675=>"11111111",
  36676=>"00000010",
  36677=>"00000011",
  36678=>"11111111",
  36679=>"00000000",
  36680=>"00000010",
  36681=>"00000000",
  36682=>"11111101",
  36683=>"11111101",
  36684=>"00000010",
  36685=>"00000000",
  36686=>"00000000",
  36687=>"00000100",
  36688=>"11111110",
  36689=>"00000010",
  36690=>"11111101",
  36691=>"00000001",
  36692=>"11111111",
  36693=>"11111110",
  36694=>"11111110",
  36695=>"00000010",
  36696=>"11111101",
  36697=>"11111110",
  36698=>"11111110",
  36699=>"11111110",
  36700=>"00000001",
  36701=>"00000010",
  36702=>"00000000",
  36703=>"11111101",
  36704=>"00000001",
  36705=>"11111111",
  36706=>"00000010",
  36707=>"11111101",
  36708=>"11111111",
  36709=>"11111101",
  36710=>"00000011",
  36711=>"00000100",
  36712=>"00000010",
  36713=>"00000011",
  36714=>"11111101",
  36715=>"11111110",
  36716=>"11111110",
  36717=>"11111111",
  36718=>"11111110",
  36719=>"11111111",
  36720=>"11111101",
  36721=>"11111111",
  36722=>"11111110",
  36723=>"00000010",
  36724=>"11111111",
  36725=>"00000000",
  36726=>"00000001",
  36727=>"11111111",
  36728=>"11111111",
  36729=>"00000001",
  36730=>"11111111",
  36731=>"11111111",
  36732=>"00000001",
  36733=>"00000011",
  36734=>"00000000",
  36735=>"00000100",
  36736=>"11111110",
  36737=>"00000000",
  36738=>"11111101",
  36739=>"11111111",
  36740=>"00000001",
  36741=>"00000001",
  36742=>"00000000",
  36743=>"11111111",
  36744=>"11111111",
  36745=>"11111110",
  36746=>"00000001",
  36747=>"00000000",
  36748=>"00000100",
  36749=>"00000011",
  36750=>"11111101",
  36751=>"00000010",
  36752=>"11111111",
  36753=>"11111101",
  36754=>"11111111",
  36755=>"00000001",
  36756=>"00000011",
  36757=>"00000001",
  36758=>"00000111",
  36759=>"11111111",
  36760=>"00000010",
  36761=>"11111111",
  36762=>"00000000",
  36763=>"11111101",
  36764=>"00000000",
  36765=>"00000010",
  36766=>"00000100",
  36767=>"11111111",
  36768=>"00000000",
  36769=>"00000011",
  36770=>"00000001",
  36771=>"11111111",
  36772=>"00000001",
  36773=>"11111111",
  36774=>"00000000",
  36775=>"11111110",
  36776=>"00000001",
  36777=>"11111111",
  36778=>"00000011",
  36779=>"11111111",
  36780=>"11111111",
  36781=>"00000010",
  36782=>"11111111",
  36783=>"00000000",
  36784=>"11111101",
  36785=>"00000010",
  36786=>"11111100",
  36787=>"00000000",
  36788=>"00000001",
  36789=>"00000010",
  36790=>"00000001",
  36791=>"11111110",
  36792=>"11111110",
  36793=>"00000000",
  36794=>"11111110",
  36795=>"00000001",
  36796=>"11111111",
  36797=>"11111101",
  36798=>"11111110",
  36799=>"00000001",
  36800=>"11111101",
  36801=>"00000100",
  36802=>"11111110",
  36803=>"00000001",
  36804=>"11111110",
  36805=>"00000010",
  36806=>"11111100",
  36807=>"00000001",
  36808=>"00000010",
  36809=>"00000011",
  36810=>"11111110",
  36811=>"00000110",
  36812=>"00000001",
  36813=>"00000011",
  36814=>"11111111",
  36815=>"11111111",
  36816=>"11111111",
  36817=>"11111111",
  36818=>"11111101",
  36819=>"11111111",
  36820=>"11111111",
  36821=>"11111110",
  36822=>"00000011",
  36823=>"00000001",
  36824=>"00000000",
  36825=>"00000011",
  36826=>"11111111",
  36827=>"00000110",
  36828=>"11111110",
  36829=>"11111111",
  36830=>"00000010",
  36831=>"11111110",
  36832=>"11111111",
  36833=>"00000101",
  36834=>"11111111",
  36835=>"00000000",
  36836=>"00000100",
  36837=>"11111111",
  36838=>"00000010",
  36839=>"11111101",
  36840=>"11111101",
  36841=>"00000000",
  36842=>"00000010",
  36843=>"00000001",
  36844=>"11111110",
  36845=>"11111110",
  36846=>"11111101",
  36847=>"00000010",
  36848=>"00000001",
  36849=>"00000000",
  36850=>"11111111",
  36851=>"00000001",
  36852=>"00000011",
  36853=>"00000011",
  36854=>"00000001",
  36855=>"11111111",
  36856=>"00000001",
  36857=>"00000011",
  36858=>"11111111",
  36859=>"00000010",
  36860=>"11111101",
  36861=>"11111101",
  36862=>"11111101",
  36863=>"00000100",
  36864=>"00000010",
  36865=>"11111111",
  36866=>"00000000",
  36867=>"00000001",
  36868=>"00000000",
  36869=>"00000100",
  36870=>"00000011",
  36871=>"00000001",
  36872=>"00000100",
  36873=>"00000011",
  36874=>"00000000",
  36875=>"00000010",
  36876=>"11111110",
  36877=>"11111111",
  36878=>"00000000",
  36879=>"00000010",
  36880=>"11111101",
  36881=>"00000010",
  36882=>"00000010",
  36883=>"00000010",
  36884=>"00000001",
  36885=>"11111111",
  36886=>"00000000",
  36887=>"11111111",
  36888=>"11111111",
  36889=>"00000100",
  36890=>"00000011",
  36891=>"00000001",
  36892=>"00000011",
  36893=>"11111110",
  36894=>"00000010",
  36895=>"00000010",
  36896=>"11111111",
  36897=>"11111110",
  36898=>"00000001",
  36899=>"11111110",
  36900=>"11111111",
  36901=>"00000001",
  36902=>"00000001",
  36903=>"00000010",
  36904=>"11111111",
  36905=>"11111111",
  36906=>"00000011",
  36907=>"00000000",
  36908=>"00000000",
  36909=>"11111111",
  36910=>"00000000",
  36911=>"00000001",
  36912=>"00000011",
  36913=>"11111110",
  36914=>"00000011",
  36915=>"00000000",
  36916=>"11111111",
  36917=>"11111110",
  36918=>"00000001",
  36919=>"00000001",
  36920=>"00000100",
  36921=>"00000000",
  36922=>"00000000",
  36923=>"00000000",
  36924=>"00000001",
  36925=>"11111111",
  36926=>"00000011",
  36927=>"11111110",
  36928=>"11111111",
  36929=>"11111110",
  36930=>"00000000",
  36931=>"00000001",
  36932=>"00000010",
  36933=>"11111110",
  36934=>"11111111",
  36935=>"11111111",
  36936=>"11111111",
  36937=>"00000010",
  36938=>"00000010",
  36939=>"00000001",
  36940=>"11111110",
  36941=>"11111111",
  36942=>"11111111",
  36943=>"11111111",
  36944=>"00000000",
  36945=>"00000001",
  36946=>"11111111",
  36947=>"00000010",
  36948=>"00000010",
  36949=>"11111101",
  36950=>"00000000",
  36951=>"00000100",
  36952=>"00000010",
  36953=>"00000001",
  36954=>"00000010",
  36955=>"00000000",
  36956=>"00000010",
  36957=>"00000000",
  36958=>"00000000",
  36959=>"11111110",
  36960=>"00000010",
  36961=>"00000101",
  36962=>"00000011",
  36963=>"00000001",
  36964=>"11111110",
  36965=>"00000000",
  36966=>"00000101",
  36967=>"00000000",
  36968=>"11111110",
  36969=>"00000001",
  36970=>"00000001",
  36971=>"00000000",
  36972=>"11111101",
  36973=>"11111110",
  36974=>"00000000",
  36975=>"00000000",
  36976=>"11111101",
  36977=>"11111101",
  36978=>"11111111",
  36979=>"00000100",
  36980=>"11111111",
  36981=>"00000001",
  36982=>"00000001",
  36983=>"00000001",
  36984=>"00000001",
  36985=>"00000000",
  36986=>"11111101",
  36987=>"00000010",
  36988=>"00000001",
  36989=>"00000010",
  36990=>"11111110",
  36991=>"00000000",
  36992=>"00000001",
  36993=>"11111110",
  36994=>"11111110",
  36995=>"00000110",
  36996=>"00000001",
  36997=>"00000011",
  36998=>"11111110",
  36999=>"00000001",
  37000=>"00000110",
  37001=>"11111101",
  37002=>"00000000",
  37003=>"11111101",
  37004=>"11111110",
  37005=>"00000010",
  37006=>"00000010",
  37007=>"11111110",
  37008=>"00000010",
  37009=>"11111111",
  37010=>"11111110",
  37011=>"11111110",
  37012=>"11111100",
  37013=>"00000010",
  37014=>"00000001",
  37015=>"00000010",
  37016=>"11111101",
  37017=>"11111101",
  37018=>"11111111",
  37019=>"00000001",
  37020=>"11111111",
  37021=>"11111111",
  37022=>"11111110",
  37023=>"00000010",
  37024=>"00000001",
  37025=>"11111110",
  37026=>"00000001",
  37027=>"00000100",
  37028=>"00000000",
  37029=>"00000011",
  37030=>"00000001",
  37031=>"11111110",
  37032=>"00000011",
  37033=>"00000001",
  37034=>"11111111",
  37035=>"11111101",
  37036=>"11111111",
  37037=>"11111101",
  37038=>"11111110",
  37039=>"11111111",
  37040=>"11111111",
  37041=>"11111111",
  37042=>"11111111",
  37043=>"00000000",
  37044=>"11111110",
  37045=>"00000000",
  37046=>"00000100",
  37047=>"11111111",
  37048=>"11111111",
  37049=>"00000000",
  37050=>"11111111",
  37051=>"00000010",
  37052=>"11111111",
  37053=>"00000000",
  37054=>"00000000",
  37055=>"11111101",
  37056=>"00000010",
  37057=>"11111101",
  37058=>"00000010",
  37059=>"11111101",
  37060=>"00000010",
  37061=>"11111111",
  37062=>"00000000",
  37063=>"00000001",
  37064=>"11111110",
  37065=>"00000011",
  37066=>"00000001",
  37067=>"00000001",
  37068=>"00000010",
  37069=>"11111110",
  37070=>"00000100",
  37071=>"11111101",
  37072=>"11111111",
  37073=>"11111111",
  37074=>"00000000",
  37075=>"00000010",
  37076=>"00000001",
  37077=>"11111110",
  37078=>"11111101",
  37079=>"00000001",
  37080=>"00000100",
  37081=>"00000000",
  37082=>"11111111",
  37083=>"00000000",
  37084=>"00000101",
  37085=>"00000000",
  37086=>"00000001",
  37087=>"00000010",
  37088=>"00000001",
  37089=>"11111111",
  37090=>"11111101",
  37091=>"00000000",
  37092=>"00000010",
  37093=>"00000010",
  37094=>"11111110",
  37095=>"00000011",
  37096=>"00000000",
  37097=>"11111101",
  37098=>"00000010",
  37099=>"11111111",
  37100=>"11111111",
  37101=>"00000001",
  37102=>"00000000",
  37103=>"00000001",
  37104=>"00000010",
  37105=>"00000010",
  37106=>"00000001",
  37107=>"00000000",
  37108=>"11111111",
  37109=>"11111110",
  37110=>"11111110",
  37111=>"00000011",
  37112=>"00000000",
  37113=>"00000000",
  37114=>"00000000",
  37115=>"00000001",
  37116=>"11111110",
  37117=>"11111101",
  37118=>"11111110",
  37119=>"00000100",
  37120=>"00000000",
  37121=>"11111111",
  37122=>"11111111",
  37123=>"11111111",
  37124=>"00000010",
  37125=>"00000010",
  37126=>"00000000",
  37127=>"11111111",
  37128=>"00000010",
  37129=>"00000100",
  37130=>"11111111",
  37131=>"11111101",
  37132=>"00000000",
  37133=>"00000011",
  37134=>"00000001",
  37135=>"11111110",
  37136=>"11111111",
  37137=>"11111101",
  37138=>"11111111",
  37139=>"00000001",
  37140=>"11111111",
  37141=>"00000000",
  37142=>"00000000",
  37143=>"11111110",
  37144=>"11111110",
  37145=>"11111110",
  37146=>"00000001",
  37147=>"00000000",
  37148=>"11111101",
  37149=>"00000011",
  37150=>"11111111",
  37151=>"00000001",
  37152=>"11111111",
  37153=>"00000001",
  37154=>"00000010",
  37155=>"11111110",
  37156=>"00000000",
  37157=>"11111110",
  37158=>"11111110",
  37159=>"11111101",
  37160=>"11111110",
  37161=>"00000000",
  37162=>"00000001",
  37163=>"11111111",
  37164=>"11111111",
  37165=>"11111110",
  37166=>"00000001",
  37167=>"00000010",
  37168=>"11111110",
  37169=>"11111110",
  37170=>"11111110",
  37171=>"11111111",
  37172=>"00000010",
  37173=>"11111100",
  37174=>"00000001",
  37175=>"00000010",
  37176=>"11111110",
  37177=>"00000000",
  37178=>"11111111",
  37179=>"11111101",
  37180=>"11111101",
  37181=>"00000100",
  37182=>"00000100",
  37183=>"00000001",
  37184=>"00000000",
  37185=>"00000001",
  37186=>"00000001",
  37187=>"00000010",
  37188=>"00000011",
  37189=>"00000101",
  37190=>"11111101",
  37191=>"11111110",
  37192=>"00000000",
  37193=>"00000010",
  37194=>"00000000",
  37195=>"00000011",
  37196=>"00000001",
  37197=>"00000000",
  37198=>"00000001",
  37199=>"00000000",
  37200=>"00000000",
  37201=>"00000011",
  37202=>"00000000",
  37203=>"11111101",
  37204=>"00000101",
  37205=>"00000010",
  37206=>"11111110",
  37207=>"11111101",
  37208=>"11111110",
  37209=>"00000001",
  37210=>"00000000",
  37211=>"11111110",
  37212=>"11111111",
  37213=>"00000011",
  37214=>"00000001",
  37215=>"00000000",
  37216=>"00000010",
  37217=>"11111110",
  37218=>"00000000",
  37219=>"00000001",
  37220=>"11111111",
  37221=>"00000010",
  37222=>"00000000",
  37223=>"00000010",
  37224=>"11111110",
  37225=>"11111111",
  37226=>"00000001",
  37227=>"00000001",
  37228=>"00000000",
  37229=>"11111111",
  37230=>"11111110",
  37231=>"00000011",
  37232=>"00000000",
  37233=>"00000010",
  37234=>"11111110",
  37235=>"11111111",
  37236=>"00000000",
  37237=>"11111110",
  37238=>"11111110",
  37239=>"00000000",
  37240=>"00000000",
  37241=>"11111111",
  37242=>"00000010",
  37243=>"00000000",
  37244=>"11111111",
  37245=>"11111111",
  37246=>"11111110",
  37247=>"00000010",
  37248=>"00000100",
  37249=>"00000001",
  37250=>"00000000",
  37251=>"11111111",
  37252=>"11111110",
  37253=>"11111101",
  37254=>"11111111",
  37255=>"00000000",
  37256=>"11111111",
  37257=>"11111110",
  37258=>"11111101",
  37259=>"00000010",
  37260=>"11111111",
  37261=>"00000010",
  37262=>"00000110",
  37263=>"00000001",
  37264=>"11111111",
  37265=>"11111110",
  37266=>"00000001",
  37267=>"00000001",
  37268=>"11111101",
  37269=>"00000011",
  37270=>"11111111",
  37271=>"00000010",
  37272=>"11111111",
  37273=>"00000001",
  37274=>"00000000",
  37275=>"00000000",
  37276=>"11111111",
  37277=>"00000001",
  37278=>"00000000",
  37279=>"11111111",
  37280=>"11111110",
  37281=>"00000011",
  37282=>"00000000",
  37283=>"11111111",
  37284=>"11111101",
  37285=>"00000011",
  37286=>"00000000",
  37287=>"11111110",
  37288=>"11111011",
  37289=>"00000000",
  37290=>"00000000",
  37291=>"11111111",
  37292=>"11111110",
  37293=>"11111110",
  37294=>"00000011",
  37295=>"00000000",
  37296=>"11111110",
  37297=>"00000001",
  37298=>"11111111",
  37299=>"11111111",
  37300=>"00000000",
  37301=>"11111110",
  37302=>"11111110",
  37303=>"00000001",
  37304=>"00000010",
  37305=>"00000101",
  37306=>"00000000",
  37307=>"11111111",
  37308=>"00000000",
  37309=>"11111101",
  37310=>"00000000",
  37311=>"00000001",
  37312=>"00000111",
  37313=>"11111101",
  37314=>"00000001",
  37315=>"11111101",
  37316=>"11111111",
  37317=>"11111110",
  37318=>"11111111",
  37319=>"11111110",
  37320=>"00000010",
  37321=>"00000000",
  37322=>"00000001",
  37323=>"11111110",
  37324=>"00000001",
  37325=>"00000000",
  37326=>"00000000",
  37327=>"11111100",
  37328=>"11111110",
  37329=>"00000001",
  37330=>"00000001",
  37331=>"00000000",
  37332=>"00000010",
  37333=>"00000001",
  37334=>"11111110",
  37335=>"00000001",
  37336=>"00000010",
  37337=>"00000001",
  37338=>"00000011",
  37339=>"11111101",
  37340=>"00000100",
  37341=>"00000000",
  37342=>"00000011",
  37343=>"00000010",
  37344=>"00000001",
  37345=>"00000000",
  37346=>"00000010",
  37347=>"11111110",
  37348=>"00000010",
  37349=>"11111110",
  37350=>"11111110",
  37351=>"00000010",
  37352=>"00000010",
  37353=>"00000011",
  37354=>"00000100",
  37355=>"00000000",
  37356=>"11111111",
  37357=>"11111111",
  37358=>"00000001",
  37359=>"11111111",
  37360=>"00000001",
  37361=>"11111101",
  37362=>"00000010",
  37363=>"11111111",
  37364=>"00000011",
  37365=>"11111101",
  37366=>"00000010",
  37367=>"11111111",
  37368=>"11111100",
  37369=>"00000000",
  37370=>"00000001",
  37371=>"00000010",
  37372=>"11111110",
  37373=>"11111110",
  37374=>"00000000",
  37375=>"00000011",
  37376=>"11111110",
  37377=>"11111111",
  37378=>"00000010",
  37379=>"00000011",
  37380=>"11111110",
  37381=>"00000000",
  37382=>"00000001",
  37383=>"11111110",
  37384=>"00000000",
  37385=>"11111111",
  37386=>"00000001",
  37387=>"00000010",
  37388=>"00000010",
  37389=>"11111111",
  37390=>"11111111",
  37391=>"00000000",
  37392=>"11111111",
  37393=>"11111110",
  37394=>"00000001",
  37395=>"11111101",
  37396=>"11111111",
  37397=>"00000010",
  37398=>"00000001",
  37399=>"11111111",
  37400=>"11111111",
  37401=>"11111110",
  37402=>"11111110",
  37403=>"00000000",
  37404=>"00000001",
  37405=>"00000010",
  37406=>"00000000",
  37407=>"00000010",
  37408=>"00000011",
  37409=>"11111110",
  37410=>"00000001",
  37411=>"11111110",
  37412=>"00000000",
  37413=>"11111111",
  37414=>"00000000",
  37415=>"00000011",
  37416=>"00000100",
  37417=>"11111101",
  37418=>"11111110",
  37419=>"00000010",
  37420=>"11111101",
  37421=>"00000000",
  37422=>"11111101",
  37423=>"00000000",
  37424=>"00000100",
  37425=>"00000011",
  37426=>"00000010",
  37427=>"11111110",
  37428=>"11111111",
  37429=>"11111101",
  37430=>"11111111",
  37431=>"00000010",
  37432=>"11111111",
  37433=>"00000000",
  37434=>"11111111",
  37435=>"11111101",
  37436=>"11111110",
  37437=>"00000001",
  37438=>"00000001",
  37439=>"11111111",
  37440=>"00000001",
  37441=>"00000000",
  37442=>"00000000",
  37443=>"11111101",
  37444=>"00000011",
  37445=>"00000100",
  37446=>"00000100",
  37447=>"00000010",
  37448=>"00000100",
  37449=>"11111110",
  37450=>"00000001",
  37451=>"11111101",
  37452=>"00000001",
  37453=>"00000101",
  37454=>"00000011",
  37455=>"00000001",
  37456=>"00000001",
  37457=>"11111101",
  37458=>"00000001",
  37459=>"11111110",
  37460=>"11111110",
  37461=>"11111110",
  37462=>"00000011",
  37463=>"00000001",
  37464=>"00000011",
  37465=>"11111110",
  37466=>"00000001",
  37467=>"00000011",
  37468=>"00000000",
  37469=>"11111110",
  37470=>"11111101",
  37471=>"11111110",
  37472=>"00000010",
  37473=>"11111111",
  37474=>"11111111",
  37475=>"00000101",
  37476=>"00000001",
  37477=>"11111110",
  37478=>"00000010",
  37479=>"11111110",
  37480=>"11111111",
  37481=>"11111110",
  37482=>"00000000",
  37483=>"11111110",
  37484=>"00000010",
  37485=>"00000011",
  37486=>"00000011",
  37487=>"00000001",
  37488=>"11111101",
  37489=>"11111111",
  37490=>"00000011",
  37491=>"11111110",
  37492=>"00000010",
  37493=>"00000001",
  37494=>"00000001",
  37495=>"11111110",
  37496=>"00000011",
  37497=>"11111111",
  37498=>"11111110",
  37499=>"11111111",
  37500=>"00000001",
  37501=>"00000000",
  37502=>"00000001",
  37503=>"00000001",
  37504=>"00000011",
  37505=>"11111110",
  37506=>"11111111",
  37507=>"00000000",
  37508=>"11111110",
  37509=>"00000001",
  37510=>"11111110",
  37511=>"00000000",
  37512=>"11111111",
  37513=>"00000010",
  37514=>"00000100",
  37515=>"11111110",
  37516=>"00000010",
  37517=>"00000001",
  37518=>"00000010",
  37519=>"00000001",
  37520=>"11111101",
  37521=>"11111111",
  37522=>"11111110",
  37523=>"00000010",
  37524=>"11111110",
  37525=>"00000101",
  37526=>"11111110",
  37527=>"11111100",
  37528=>"11111111",
  37529=>"11111110",
  37530=>"00000000",
  37531=>"00000011",
  37532=>"00000001",
  37533=>"11111111",
  37534=>"11111111",
  37535=>"00000001",
  37536=>"00000000",
  37537=>"00000001",
  37538=>"00000001",
  37539=>"00000101",
  37540=>"00000001",
  37541=>"11111110",
  37542=>"11111111",
  37543=>"00000011",
  37544=>"00000011",
  37545=>"11111101",
  37546=>"11111101",
  37547=>"00000000",
  37548=>"00000001",
  37549=>"00000010",
  37550=>"00000001",
  37551=>"00000001",
  37552=>"11111111",
  37553=>"11111111",
  37554=>"00000001",
  37555=>"00000000",
  37556=>"00000000",
  37557=>"00000010",
  37558=>"00000001",
  37559=>"00000011",
  37560=>"11111110",
  37561=>"11111110",
  37562=>"00000010",
  37563=>"00000010",
  37564=>"00000001",
  37565=>"11111111",
  37566=>"00000000",
  37567=>"11111111",
  37568=>"11111101",
  37569=>"11111101",
  37570=>"00000010",
  37571=>"00000001",
  37572=>"11111110",
  37573=>"11111101",
  37574=>"00000010",
  37575=>"11111101",
  37576=>"11111111",
  37577=>"00000100",
  37578=>"00000010",
  37579=>"00000011",
  37580=>"00000010",
  37581=>"11111101",
  37582=>"00000010",
  37583=>"11111110",
  37584=>"00000010",
  37585=>"00000000",
  37586=>"00000010",
  37587=>"11111110",
  37588=>"00000101",
  37589=>"11111111",
  37590=>"11111111",
  37591=>"11111101",
  37592=>"00000000",
  37593=>"11111110",
  37594=>"00000010",
  37595=>"11111101",
  37596=>"11111110",
  37597=>"11111111",
  37598=>"11111101",
  37599=>"00000000",
  37600=>"00000000",
  37601=>"00000011",
  37602=>"11111111",
  37603=>"00000011",
  37604=>"11111110",
  37605=>"11111110",
  37606=>"00000011",
  37607=>"11111111",
  37608=>"11111111",
  37609=>"00000001",
  37610=>"11111110",
  37611=>"11111110",
  37612=>"00000001",
  37613=>"11111101",
  37614=>"00000000",
  37615=>"11111110",
  37616=>"00000000",
  37617=>"11111110",
  37618=>"00000000",
  37619=>"00000000",
  37620=>"11111111",
  37621=>"00000001",
  37622=>"11111111",
  37623=>"00000010",
  37624=>"00000001",
  37625=>"11111110",
  37626=>"00000010",
  37627=>"11111110",
  37628=>"00000001",
  37629=>"00000001",
  37630=>"00000011",
  37631=>"00000010",
  37632=>"00000011",
  37633=>"00000000",
  37634=>"00000001",
  37635=>"00000010",
  37636=>"00000001",
  37637=>"11111111",
  37638=>"11111111",
  37639=>"00000010",
  37640=>"00000001",
  37641=>"00000001",
  37642=>"00000011",
  37643=>"11111110",
  37644=>"00000001",
  37645=>"00000000",
  37646=>"11111111",
  37647=>"11111110",
  37648=>"11111110",
  37649=>"11111110",
  37650=>"00000001",
  37651=>"00000001",
  37652=>"00000011",
  37653=>"00000001",
  37654=>"11111110",
  37655=>"00000011",
  37656=>"11111101",
  37657=>"11111110",
  37658=>"11111101",
  37659=>"00000001",
  37660=>"11111110",
  37661=>"11111101",
  37662=>"00000000",
  37663=>"00000011",
  37664=>"00000010",
  37665=>"11111111",
  37666=>"00000010",
  37667=>"11111111",
  37668=>"00000001",
  37669=>"11111100",
  37670=>"11111110",
  37671=>"11111110",
  37672=>"00000000",
  37673=>"11111101",
  37674=>"11111111",
  37675=>"11111111",
  37676=>"11111111",
  37677=>"00000010",
  37678=>"00000000",
  37679=>"00000010",
  37680=>"11111101",
  37681=>"00000001",
  37682=>"11111110",
  37683=>"00000110",
  37684=>"00000011",
  37685=>"11111111",
  37686=>"00000011",
  37687=>"00000010",
  37688=>"00000011",
  37689=>"11111110",
  37690=>"00000010",
  37691=>"00000100",
  37692=>"11111111",
  37693=>"11111111",
  37694=>"00000011",
  37695=>"00000010",
  37696=>"00000000",
  37697=>"00000010",
  37698=>"11111101",
  37699=>"00000100",
  37700=>"00000011",
  37701=>"11111110",
  37702=>"11111100",
  37703=>"00000010",
  37704=>"00000001",
  37705=>"00000000",
  37706=>"11111101",
  37707=>"00000001",
  37708=>"00000000",
  37709=>"00000000",
  37710=>"00000001",
  37711=>"00000000",
  37712=>"00000000",
  37713=>"00000000",
  37714=>"00000001",
  37715=>"11111110",
  37716=>"11111110",
  37717=>"11111111",
  37718=>"11111110",
  37719=>"00000011",
  37720=>"11111110",
  37721=>"00000010",
  37722=>"00000010",
  37723=>"00000000",
  37724=>"00000011",
  37725=>"00000000",
  37726=>"11111111",
  37727=>"11111111",
  37728=>"00000000",
  37729=>"00000000",
  37730=>"11111110",
  37731=>"00000000",
  37732=>"00000010",
  37733=>"11111110",
  37734=>"11111110",
  37735=>"11111111",
  37736=>"00000001",
  37737=>"11111101",
  37738=>"11111101",
  37739=>"11111111",
  37740=>"00000001",
  37741=>"11111110",
  37742=>"00000001",
  37743=>"11111110",
  37744=>"11111110",
  37745=>"11111110",
  37746=>"11111111",
  37747=>"00000001",
  37748=>"00000000",
  37749=>"00000000",
  37750=>"00000000",
  37751=>"00000011",
  37752=>"11111110",
  37753=>"11111110",
  37754=>"00000001",
  37755=>"00000010",
  37756=>"11111101",
  37757=>"00000010",
  37758=>"11111111",
  37759=>"00000010",
  37760=>"00000000",
  37761=>"11111110",
  37762=>"11111110",
  37763=>"11111101",
  37764=>"00000000",
  37765=>"11111111",
  37766=>"00000000",
  37767=>"00000000",
  37768=>"11111111",
  37769=>"00000000",
  37770=>"00000010",
  37771=>"11111100",
  37772=>"11111101",
  37773=>"11111111",
  37774=>"11111110",
  37775=>"11111110",
  37776=>"00000001",
  37777=>"00000000",
  37778=>"11111110",
  37779=>"11111111",
  37780=>"00000011",
  37781=>"00000000",
  37782=>"11111101",
  37783=>"00000011",
  37784=>"00000011",
  37785=>"00000000",
  37786=>"00000001",
  37787=>"00000010",
  37788=>"11111111",
  37789=>"11111110",
  37790=>"00000000",
  37791=>"00000010",
  37792=>"00000000",
  37793=>"00000001",
  37794=>"11111100",
  37795=>"00000011",
  37796=>"00000100",
  37797=>"00000000",
  37798=>"11111101",
  37799=>"00000000",
  37800=>"11111110",
  37801=>"00000010",
  37802=>"00000010",
  37803=>"11111110",
  37804=>"11111101",
  37805=>"00000100",
  37806=>"11111110",
  37807=>"00000010",
  37808=>"00000010",
  37809=>"00000000",
  37810=>"00000001",
  37811=>"11111111",
  37812=>"11111111",
  37813=>"00000010",
  37814=>"00000000",
  37815=>"11111110",
  37816=>"00000001",
  37817=>"11111111",
  37818=>"11111111",
  37819=>"00000011",
  37820=>"11111111",
  37821=>"00000001",
  37822=>"00000001",
  37823=>"00000010",
  37824=>"11111110",
  37825=>"00000010",
  37826=>"00000001",
  37827=>"11111110",
  37828=>"00000000",
  37829=>"00000011",
  37830=>"00000001",
  37831=>"00000000",
  37832=>"00000000",
  37833=>"00000000",
  37834=>"00000000",
  37835=>"00000001",
  37836=>"11111111",
  37837=>"00000001",
  37838=>"11111110",
  37839=>"00000010",
  37840=>"00000000",
  37841=>"11111110",
  37842=>"11111111",
  37843=>"00000000",
  37844=>"11111110",
  37845=>"00000001",
  37846=>"00000010",
  37847=>"00000010",
  37848=>"00000100",
  37849=>"00000011",
  37850=>"00000001",
  37851=>"11111110",
  37852=>"00000000",
  37853=>"11111101",
  37854=>"00000100",
  37855=>"00000001",
  37856=>"11111101",
  37857=>"00000001",
  37858=>"00000100",
  37859=>"11111111",
  37860=>"11111111",
  37861=>"00000000",
  37862=>"00000001",
  37863=>"00000011",
  37864=>"11111110",
  37865=>"00000000",
  37866=>"00000000",
  37867=>"11111111",
  37868=>"11111101",
  37869=>"00000010",
  37870=>"11111111",
  37871=>"00000000",
  37872=>"11111101",
  37873=>"00000001",
  37874=>"00000010",
  37875=>"11111111",
  37876=>"11111111",
  37877=>"00000011",
  37878=>"00000011",
  37879=>"11111110",
  37880=>"00000010",
  37881=>"00000000",
  37882=>"11111111",
  37883=>"11111111",
  37884=>"00000000",
  37885=>"11111111",
  37886=>"00000011",
  37887=>"00000000",
  37888=>"00000010",
  37889=>"00000001",
  37890=>"00000010",
  37891=>"11111111",
  37892=>"00000001",
  37893=>"00000001",
  37894=>"11111111",
  37895=>"00000001",
  37896=>"11111110",
  37897=>"00000001",
  37898=>"11111111",
  37899=>"11111110",
  37900=>"00000001",
  37901=>"00000000",
  37902=>"00000000",
  37903=>"00000001",
  37904=>"11111111",
  37905=>"00000000",
  37906=>"11111111",
  37907=>"00000000",
  37908=>"11111111",
  37909=>"00000001",
  37910=>"00000000",
  37911=>"00000001",
  37912=>"00000000",
  37913=>"00000001",
  37914=>"11111111",
  37915=>"00000001",
  37916=>"11111111",
  37917=>"11111111",
  37918=>"00000000",
  37919=>"11111111",
  37920=>"11111110",
  37921=>"00000000",
  37922=>"00000001",
  37923=>"00000001",
  37924=>"11111111",
  37925=>"11111111",
  37926=>"00000000",
  37927=>"11111111",
  37928=>"00000001",
  37929=>"00000001",
  37930=>"11111111",
  37931=>"00000001",
  37932=>"11111111",
  37933=>"00000001",
  37934=>"00000000",
  37935=>"00000000",
  37936=>"11111111",
  37937=>"00000001",
  37938=>"00000010",
  37939=>"00000000",
  37940=>"00000001",
  37941=>"00000000",
  37942=>"00000000",
  37943=>"00000010",
  37944=>"00000000",
  37945=>"00000001",
  37946=>"00000001",
  37947=>"00000001",
  37948=>"00000001",
  37949=>"11111111",
  37950=>"11111111",
  37951=>"00000001",
  37952=>"00000001",
  37953=>"00000001",
  37954=>"00000001",
  37955=>"00000010",
  37956=>"00000001",
  37957=>"11111111",
  37958=>"11111111",
  37959=>"00000001",
  37960=>"11111111",
  37961=>"00000000",
  37962=>"00000000",
  37963=>"00000000",
  37964=>"11111111",
  37965=>"11111111",
  37966=>"11111110",
  37967=>"00000000",
  37968=>"11111110",
  37969=>"00000010",
  37970=>"11111110",
  37971=>"00000001",
  37972=>"00000000",
  37973=>"00000000",
  37974=>"00000001",
  37975=>"00000001",
  37976=>"11111111",
  37977=>"00000000",
  37978=>"00000000",
  37979=>"00000010",
  37980=>"00000010",
  37981=>"00000001",
  37982=>"00000001",
  37983=>"00000001",
  37984=>"00000000",
  37985=>"00000001",
  37986=>"00000001",
  37987=>"11111111",
  37988=>"00000001",
  37989=>"00000001",
  37990=>"11111111",
  37991=>"00000010",
  37992=>"11111111",
  37993=>"00000000",
  37994=>"00000000",
  37995=>"00000000",
  37996=>"11111111",
  37997=>"00000000",
  37998=>"11111111",
  37999=>"11111110",
  38000=>"00000000",
  38001=>"11111111",
  38002=>"00000001",
  38003=>"00000010",
  38004=>"00000000",
  38005=>"00000001",
  38006=>"00000001",
  38007=>"00000001",
  38008=>"00000000",
  38009=>"00000000",
  38010=>"00000001",
  38011=>"11111111",
  38012=>"11111111",
  38013=>"00000000",
  38014=>"11111110",
  38015=>"00000000",
  38016=>"11111111",
  38017=>"00000001",
  38018=>"00000001",
  38019=>"11111110",
  38020=>"00000001",
  38021=>"00000001",
  38022=>"00000010",
  38023=>"00000001",
  38024=>"00000001",
  38025=>"00000000",
  38026=>"00000000",
  38027=>"00000001",
  38028=>"00000001",
  38029=>"00000001",
  38030=>"00000001",
  38031=>"11111111",
  38032=>"00000010",
  38033=>"00000000",
  38034=>"11111111",
  38035=>"00000000",
  38036=>"11111111",
  38037=>"11111111",
  38038=>"00000000",
  38039=>"00000001",
  38040=>"00000000",
  38041=>"11111111",
  38042=>"00000001",
  38043=>"00000000",
  38044=>"00000001",
  38045=>"00000001",
  38046=>"11111110",
  38047=>"00000001",
  38048=>"00000001",
  38049=>"00000001",
  38050=>"00000010",
  38051=>"11111111",
  38052=>"00000001",
  38053=>"00000001",
  38054=>"11111111",
  38055=>"11111111",
  38056=>"11111111",
  38057=>"00000000",
  38058=>"11111110",
  38059=>"11111111",
  38060=>"11111111",
  38061=>"00000001",
  38062=>"00000000",
  38063=>"11111111",
  38064=>"00000000",
  38065=>"00000001",
  38066=>"00000000",
  38067=>"00000010",
  38068=>"00000001",
  38069=>"11111111",
  38070=>"00000000",
  38071=>"11111111",
  38072=>"00000000",
  38073=>"11111111",
  38074=>"00000001",
  38075=>"11111110",
  38076=>"11111111",
  38077=>"00000001",
  38078=>"00000010",
  38079=>"00000001",
  38080=>"00000000",
  38081=>"00000010",
  38082=>"11111111",
  38083=>"11111111",
  38084=>"00000010",
  38085=>"11111111",
  38086=>"00000000",
  38087=>"00000000",
  38088=>"00000001",
  38089=>"00000001",
  38090=>"11111111",
  38091=>"11111110",
  38092=>"00000001",
  38093=>"00000010",
  38094=>"11111111",
  38095=>"11111111",
  38096=>"00000000",
  38097=>"00000010",
  38098=>"11111110",
  38099=>"00000000",
  38100=>"00000010",
  38101=>"00000000",
  38102=>"00000000",
  38103=>"11111111",
  38104=>"00000001",
  38105=>"00000000",
  38106=>"11111111",
  38107=>"00000000",
  38108=>"11111110",
  38109=>"11111111",
  38110=>"11111111",
  38111=>"00000001",
  38112=>"11111111",
  38113=>"00000000",
  38114=>"00000010",
  38115=>"11111110",
  38116=>"00000001",
  38117=>"00000000",
  38118=>"00000000",
  38119=>"00000000",
  38120=>"11111111",
  38121=>"00000000",
  38122=>"00000000",
  38123=>"11111110",
  38124=>"00000001",
  38125=>"00000001",
  38126=>"11111111",
  38127=>"11111111",
  38128=>"00000001",
  38129=>"11111111",
  38130=>"00000001",
  38131=>"00000000",
  38132=>"00000001",
  38133=>"00000000",
  38134=>"00000001",
  38135=>"00000001",
  38136=>"00000001",
  38137=>"00000010",
  38138=>"11111111",
  38139=>"00000001",
  38140=>"11111111",
  38141=>"00000000",
  38142=>"00000000",
  38143=>"11111111",
  38144=>"00000001",
  38145=>"00000000",
  38146=>"11111111",
  38147=>"11111111",
  38148=>"00000010",
  38149=>"00000000",
  38150=>"00000001",
  38151=>"00000000",
  38152=>"11111111",
  38153=>"00000000",
  38154=>"00000000",
  38155=>"00000010",
  38156=>"11111110",
  38157=>"00000000",
  38158=>"11111111",
  38159=>"00000001",
  38160=>"00000001",
  38161=>"11111110",
  38162=>"11111111",
  38163=>"00000001",
  38164=>"00000000",
  38165=>"00000010",
  38166=>"00000000",
  38167=>"11111110",
  38168=>"00000001",
  38169=>"00000000",
  38170=>"00000010",
  38171=>"11111110",
  38172=>"11111111",
  38173=>"00000000",
  38174=>"00000000",
  38175=>"00000001",
  38176=>"00000000",
  38177=>"00000001",
  38178=>"11111111",
  38179=>"00000000",
  38180=>"11111111",
  38181=>"00000001",
  38182=>"11111110",
  38183=>"00000000",
  38184=>"11111111",
  38185=>"00000000",
  38186=>"11111111",
  38187=>"11111111",
  38188=>"11111110",
  38189=>"00000001",
  38190=>"00000001",
  38191=>"00000001",
  38192=>"00000001",
  38193=>"11111111",
  38194=>"00000000",
  38195=>"11111110",
  38196=>"11111111",
  38197=>"11111111",
  38198=>"11111111",
  38199=>"11111110",
  38200=>"00000001",
  38201=>"11111110",
  38202=>"11111111",
  38203=>"00000001",
  38204=>"00000000",
  38205=>"00000001",
  38206=>"00000000",
  38207=>"11111110",
  38208=>"11111111",
  38209=>"00000001",
  38210=>"00000000",
  38211=>"00000000",
  38212=>"00000001",
  38213=>"00000001",
  38214=>"00000010",
  38215=>"00000001",
  38216=>"11111111",
  38217=>"11111111",
  38218=>"11111111",
  38219=>"11111111",
  38220=>"00000000",
  38221=>"11111110",
  38222=>"11111111",
  38223=>"00000000",
  38224=>"11111111",
  38225=>"00000001",
  38226=>"00000000",
  38227=>"11111111",
  38228=>"00000001",
  38229=>"00000000",
  38230=>"11111111",
  38231=>"00000000",
  38232=>"00000000",
  38233=>"00000000",
  38234=>"11111111",
  38235=>"11111111",
  38236=>"11111111",
  38237=>"00000001",
  38238=>"11111111",
  38239=>"00000000",
  38240=>"00000000",
  38241=>"00000001",
  38242=>"00000001",
  38243=>"11111111",
  38244=>"00000001",
  38245=>"00000000",
  38246=>"11111110",
  38247=>"00000001",
  38248=>"00000001",
  38249=>"11111111",
  38250=>"11111111",
  38251=>"00000000",
  38252=>"11111111",
  38253=>"11111111",
  38254=>"00000001",
  38255=>"11111111",
  38256=>"00000010",
  38257=>"11111111",
  38258=>"00000001",
  38259=>"00000000",
  38260=>"00000001",
  38261=>"00000001",
  38262=>"11111111",
  38263=>"00000000",
  38264=>"00000000",
  38265=>"11111111",
  38266=>"00000001",
  38267=>"00000001",
  38268=>"11111111",
  38269=>"00000001",
  38270=>"00000010",
  38271=>"00000001",
  38272=>"00000001",
  38273=>"00000001",
  38274=>"00000010",
  38275=>"11111111",
  38276=>"00000000",
  38277=>"00000001",
  38278=>"11111111",
  38279=>"11111111",
  38280=>"11111111",
  38281=>"00000000",
  38282=>"00000001",
  38283=>"11111111",
  38284=>"00000001",
  38285=>"00000001",
  38286=>"00000001",
  38287=>"00000000",
  38288=>"11111110",
  38289=>"11111111",
  38290=>"11111111",
  38291=>"00000001",
  38292=>"11111111",
  38293=>"11111111",
  38294=>"00000001",
  38295=>"00000001",
  38296=>"00000001",
  38297=>"00000000",
  38298=>"00000000",
  38299=>"00000010",
  38300=>"11111111",
  38301=>"11111111",
  38302=>"00000000",
  38303=>"11111110",
  38304=>"11111111",
  38305=>"00000000",
  38306=>"00000000",
  38307=>"00000000",
  38308=>"00000000",
  38309=>"00000001",
  38310=>"00000001",
  38311=>"00000000",
  38312=>"11111111",
  38313=>"00000000",
  38314=>"11111111",
  38315=>"00000001",
  38316=>"11111111",
  38317=>"00000001",
  38318=>"00000000",
  38319=>"00000000",
  38320=>"00000001",
  38321=>"00000000",
  38322=>"11111111",
  38323=>"11111111",
  38324=>"00000001",
  38325=>"11111111",
  38326=>"00000001",
  38327=>"00000000",
  38328=>"11111111",
  38329=>"00000010",
  38330=>"00000000",
  38331=>"00000001",
  38332=>"11111111",
  38333=>"11111110",
  38334=>"00000001",
  38335=>"11111111",
  38336=>"00000001",
  38337=>"11111111",
  38338=>"00000001",
  38339=>"11111111",
  38340=>"00000010",
  38341=>"00000000",
  38342=>"11111110",
  38343=>"11111111",
  38344=>"11111111",
  38345=>"11111110",
  38346=>"11111111",
  38347=>"00000000",
  38348=>"00000001",
  38349=>"00000000",
  38350=>"00000001",
  38351=>"00000001",
  38352=>"00000001",
  38353=>"11111111",
  38354=>"00000001",
  38355=>"00000001",
  38356=>"11111111",
  38357=>"00000000",
  38358=>"11111111",
  38359=>"00000000",
  38360=>"00000000",
  38361=>"00000001",
  38362=>"11111111",
  38363=>"00000001",
  38364=>"00000001",
  38365=>"00000010",
  38366=>"11111110",
  38367=>"00000000",
  38368=>"11111111",
  38369=>"00000010",
  38370=>"00000010",
  38371=>"11111110",
  38372=>"00000000",
  38373=>"00000001",
  38374=>"11111111",
  38375=>"00000000",
  38376=>"00000001",
  38377=>"11111111",
  38378=>"11111111",
  38379=>"00000000",
  38380=>"00000000",
  38381=>"00000001",
  38382=>"00000000",
  38383=>"00000001",
  38384=>"11111111",
  38385=>"00000000",
  38386=>"00000000",
  38387=>"00000000",
  38388=>"00000001",
  38389=>"00000001",
  38390=>"11111111",
  38391=>"00000000",
  38392=>"00000000",
  38393=>"00000000",
  38394=>"11111111",
  38395=>"11111111",
  38396=>"00000000",
  38397=>"00000000",
  38398=>"00000010",
  38399=>"00000001",
  38400=>"11111111",
  38401=>"00000001",
  38402=>"00000000",
  38403=>"00000000",
  38404=>"00000001",
  38405=>"11111110",
  38406=>"11111111",
  38407=>"00000001",
  38408=>"11111111",
  38409=>"11111111",
  38410=>"00000000",
  38411=>"11111110",
  38412=>"11111111",
  38413=>"00000001",
  38414=>"00000001",
  38415=>"00000000",
  38416=>"11111111",
  38417=>"11111111",
  38418=>"11111110",
  38419=>"11111111",
  38420=>"00000001",
  38421=>"11111111",
  38422=>"00000000",
  38423=>"11111111",
  38424=>"00000001",
  38425=>"00000001",
  38426=>"00000000",
  38427=>"11111110",
  38428=>"11111111",
  38429=>"00000000",
  38430=>"00000010",
  38431=>"11111111",
  38432=>"00000000",
  38433=>"00000000",
  38434=>"11111110",
  38435=>"00000001",
  38436=>"00000001",
  38437=>"11111111",
  38438=>"00000001",
  38439=>"11111111",
  38440=>"00000000",
  38441=>"11111111",
  38442=>"11111111",
  38443=>"00000000",
  38444=>"00000001",
  38445=>"00000001",
  38446=>"11111111",
  38447=>"11111111",
  38448=>"11111111",
  38449=>"11111110",
  38450=>"11111111",
  38451=>"00000010",
  38452=>"11111111",
  38453=>"00000001",
  38454=>"11111111",
  38455=>"11111111",
  38456=>"00000000",
  38457=>"00000001",
  38458=>"11111111",
  38459=>"00000001",
  38460=>"11111111",
  38461=>"11111111",
  38462=>"11111111",
  38463=>"00000000",
  38464=>"00000010",
  38465=>"11111111",
  38466=>"00000000",
  38467=>"00000000",
  38468=>"00000000",
  38469=>"00000010",
  38470=>"00000001",
  38471=>"00000010",
  38472=>"00000010",
  38473=>"00000001",
  38474=>"00000001",
  38475=>"00000001",
  38476=>"00000001",
  38477=>"00000001",
  38478=>"00000001",
  38479=>"00000010",
  38480=>"00000010",
  38481=>"11111111",
  38482=>"00000001",
  38483=>"11111111",
  38484=>"00000001",
  38485=>"00000001",
  38486=>"00000000",
  38487=>"11111111",
  38488=>"00000000",
  38489=>"00000001",
  38490=>"11111111",
  38491=>"00000001",
  38492=>"11111111",
  38493=>"00000000",
  38494=>"00000000",
  38495=>"00000010",
  38496=>"00000000",
  38497=>"00000000",
  38498=>"00000000",
  38499=>"11111111",
  38500=>"00000000",
  38501=>"11111111",
  38502=>"11111111",
  38503=>"00000000",
  38504=>"11111111",
  38505=>"00000001",
  38506=>"11111111",
  38507=>"00000010",
  38508=>"00000000",
  38509=>"00000000",
  38510=>"00000001",
  38511=>"00000001",
  38512=>"00000000",
  38513=>"00000001",
  38514=>"11111110",
  38515=>"00000000",
  38516=>"00000000",
  38517=>"00000000",
  38518=>"00000001",
  38519=>"11111111",
  38520=>"11111111",
  38521=>"11111111",
  38522=>"00000001",
  38523=>"11111111",
  38524=>"00000000",
  38525=>"11111110",
  38526=>"11111111",
  38527=>"00000000",
  38528=>"00000001",
  38529=>"00000001",
  38530=>"00000000",
  38531=>"00000000",
  38532=>"00000001",
  38533=>"00000010",
  38534=>"00000001",
  38535=>"11111110",
  38536=>"00000001",
  38537=>"11111111",
  38538=>"11111110",
  38539=>"11111111",
  38540=>"00000001",
  38541=>"00000001",
  38542=>"11111111",
  38543=>"11111111",
  38544=>"00000000",
  38545=>"11111111",
  38546=>"00000001",
  38547=>"00000010",
  38548=>"00000001",
  38549=>"00000000",
  38550=>"00000001",
  38551=>"00000001",
  38552=>"00000001",
  38553=>"00000001",
  38554=>"11111111",
  38555=>"00000000",
  38556=>"00000001",
  38557=>"00000000",
  38558=>"00000001",
  38559=>"00000000",
  38560=>"11111110",
  38561=>"00000000",
  38562=>"00000001",
  38563=>"11111110",
  38564=>"00000000",
  38565=>"00000000",
  38566=>"11111110",
  38567=>"11111111",
  38568=>"11111111",
  38569=>"11111111",
  38570=>"00000000",
  38571=>"00000001",
  38572=>"11111110",
  38573=>"00000001",
  38574=>"11111110",
  38575=>"00000001",
  38576=>"00000001",
  38577=>"00000001",
  38578=>"11111111",
  38579=>"00000001",
  38580=>"11111111",
  38581=>"00000001",
  38582=>"00000000",
  38583=>"00000000",
  38584=>"00000000",
  38585=>"00000001",
  38586=>"00000001",
  38587=>"11111111",
  38588=>"11111111",
  38589=>"00000001",
  38590=>"00000001",
  38591=>"11111111",
  38592=>"11111110",
  38593=>"00000001",
  38594=>"11111111",
  38595=>"00000000",
  38596=>"00000000",
  38597=>"11111111",
  38598=>"00000001",
  38599=>"00000000",
  38600=>"00000001",
  38601=>"00000000",
  38602=>"11111111",
  38603=>"00000001",
  38604=>"11111111",
  38605=>"00000000",
  38606=>"00000000",
  38607=>"11111111",
  38608=>"11111111",
  38609=>"00000001",
  38610=>"00000001",
  38611=>"00000001",
  38612=>"11111111",
  38613=>"11111111",
  38614=>"00000010",
  38615=>"00000000",
  38616=>"00000001",
  38617=>"00000000",
  38618=>"00000001",
  38619=>"11111110",
  38620=>"11111111",
  38621=>"00000001",
  38622=>"11111111",
  38623=>"00000000",
  38624=>"11111111",
  38625=>"00000000",
  38626=>"11111111",
  38627=>"00000001",
  38628=>"00000001",
  38629=>"00000001",
  38630=>"11111111",
  38631=>"00000000",
  38632=>"11111111",
  38633=>"00000000",
  38634=>"11111111",
  38635=>"00000000",
  38636=>"00000001",
  38637=>"00000000",
  38638=>"00000000",
  38639=>"11111111",
  38640=>"00000000",
  38641=>"11111111",
  38642=>"00000001",
  38643=>"00000001",
  38644=>"00000000",
  38645=>"00000001",
  38646=>"00000000",
  38647=>"00000000",
  38648=>"00000001",
  38649=>"11111111",
  38650=>"00000000",
  38651=>"00000001",
  38652=>"11111110",
  38653=>"00000001",
  38654=>"00000000",
  38655=>"00000000",
  38656=>"00000000",
  38657=>"11111111",
  38658=>"11111111",
  38659=>"11111111",
  38660=>"11111111",
  38661=>"00000000",
  38662=>"00000000",
  38663=>"00000000",
  38664=>"11111111",
  38665=>"00000001",
  38666=>"00000001",
  38667=>"11111110",
  38668=>"00000000",
  38669=>"11111111",
  38670=>"11111111",
  38671=>"00000001",
  38672=>"00000000",
  38673=>"11111110",
  38674=>"00000000",
  38675=>"11111110",
  38676=>"00000010",
  38677=>"11111110",
  38678=>"00000000",
  38679=>"00000000",
  38680=>"00000000",
  38681=>"00000000",
  38682=>"00000000",
  38683=>"00000000",
  38684=>"11111111",
  38685=>"00000000",
  38686=>"00000001",
  38687=>"00000000",
  38688=>"00000010",
  38689=>"00000010",
  38690=>"00000001",
  38691=>"11111110",
  38692=>"00000000",
  38693=>"11111111",
  38694=>"00000000",
  38695=>"00000000",
  38696=>"00000000",
  38697=>"11111111",
  38698=>"00000000",
  38699=>"00000001",
  38700=>"00000000",
  38701=>"00000000",
  38702=>"00000001",
  38703=>"11111111",
  38704=>"00000001",
  38705=>"11111111",
  38706=>"11111111",
  38707=>"00000001",
  38708=>"00000000",
  38709=>"00000010",
  38710=>"11111110",
  38711=>"00000000",
  38712=>"11111111",
  38713=>"11111111",
  38714=>"11111110",
  38715=>"11111111",
  38716=>"00000001",
  38717=>"00000001",
  38718=>"00000000",
  38719=>"00000001",
  38720=>"00000001",
  38721=>"11111111",
  38722=>"00000010",
  38723=>"11111111",
  38724=>"00000000",
  38725=>"11111111",
  38726=>"00000001",
  38727=>"11111111",
  38728=>"00000001",
  38729=>"11111111",
  38730=>"00000010",
  38731=>"11111111",
  38732=>"00000001",
  38733=>"00000000",
  38734=>"00000000",
  38735=>"00000000",
  38736=>"00000001",
  38737=>"00000000",
  38738=>"00000000",
  38739=>"11111111",
  38740=>"00000000",
  38741=>"00000000",
  38742=>"00000001",
  38743=>"00000000",
  38744=>"00000001",
  38745=>"00000010",
  38746=>"00000000",
  38747=>"00000000",
  38748=>"00000001",
  38749=>"11111111",
  38750=>"11111111",
  38751=>"00000001",
  38752=>"00000000",
  38753=>"11111111",
  38754=>"00000010",
  38755=>"11111111",
  38756=>"00000000",
  38757=>"00000000",
  38758=>"11111111",
  38759=>"11111110",
  38760=>"00000001",
  38761=>"00000001",
  38762=>"11111111",
  38763=>"00000001",
  38764=>"11111111",
  38765=>"00000001",
  38766=>"00000000",
  38767=>"11111111",
  38768=>"11111111",
  38769=>"00000001",
  38770=>"11111111",
  38771=>"00000001",
  38772=>"11111111",
  38773=>"11111111",
  38774=>"11111110",
  38775=>"00000001",
  38776=>"11111110",
  38777=>"00000001",
  38778=>"11111111",
  38779=>"00000001",
  38780=>"00000001",
  38781=>"00000000",
  38782=>"00000000",
  38783=>"11111111",
  38784=>"00000001",
  38785=>"11111111",
  38786=>"11111111",
  38787=>"11111110",
  38788=>"00000001",
  38789=>"11111111",
  38790=>"11111111",
  38791=>"00000000",
  38792=>"11111111",
  38793=>"00000000",
  38794=>"11111111",
  38795=>"11111111",
  38796=>"11111111",
  38797=>"00000001",
  38798=>"00000000",
  38799=>"00000000",
  38800=>"00000001",
  38801=>"00000001",
  38802=>"00000000",
  38803=>"00000001",
  38804=>"00000010",
  38805=>"00000000",
  38806=>"00000001",
  38807=>"00000010",
  38808=>"11111111",
  38809=>"00000001",
  38810=>"00000001",
  38811=>"00000001",
  38812=>"00000000",
  38813=>"11111111",
  38814=>"11111111",
  38815=>"11111110",
  38816=>"00000000",
  38817=>"11111111",
  38818=>"11111111",
  38819=>"11111111",
  38820=>"00000000",
  38821=>"11111111",
  38822=>"11111110",
  38823=>"00000000",
  38824=>"00000001",
  38825=>"00000000",
  38826=>"00000010",
  38827=>"11111110",
  38828=>"11111111",
  38829=>"00000000",
  38830=>"00000000",
  38831=>"00000001",
  38832=>"00000000",
  38833=>"00000001",
  38834=>"00000000",
  38835=>"11111111",
  38836=>"11111111",
  38837=>"11111111",
  38838=>"11111111",
  38839=>"00000000",
  38840=>"00000001",
  38841=>"11111111",
  38842=>"11111111",
  38843=>"00000000",
  38844=>"11111111",
  38845=>"00000000",
  38846=>"00000000",
  38847=>"00000010",
  38848=>"00000000",
  38849=>"00000000",
  38850=>"11111111",
  38851=>"00000010",
  38852=>"00000001",
  38853=>"11111111",
  38854=>"00000000",
  38855=>"00000000",
  38856=>"00000000",
  38857=>"11111111",
  38858=>"00000001",
  38859=>"11111110",
  38860=>"00000001",
  38861=>"11111111",
  38862=>"00000001",
  38863=>"11111111",
  38864=>"11111110",
  38865=>"11111111",
  38866=>"00000000",
  38867=>"11111111",
  38868=>"00000000",
  38869=>"00000001",
  38870=>"00000001",
  38871=>"00000000",
  38872=>"00000010",
  38873=>"00000010",
  38874=>"00000000",
  38875=>"11111111",
  38876=>"11111111",
  38877=>"11111110",
  38878=>"11111111",
  38879=>"00000001",
  38880=>"00000000",
  38881=>"00000000",
  38882=>"00000001",
  38883=>"11111111",
  38884=>"00000001",
  38885=>"11111111",
  38886=>"00000001",
  38887=>"00000000",
  38888=>"00000000",
  38889=>"00000000",
  38890=>"00000000",
  38891=>"00000000",
  38892=>"00000000",
  38893=>"11111111",
  38894=>"00000000",
  38895=>"00000000",
  38896=>"00000000",
  38897=>"11111111",
  38898=>"00000001",
  38899=>"11111110",
  38900=>"00000001",
  38901=>"00000001",
  38902=>"00000000",
  38903=>"00000001",
  38904=>"00000000",
  38905=>"11111110",
  38906=>"11111111",
  38907=>"00000001",
  38908=>"11111111",
  38909=>"00000000",
  38910=>"00000000",
  38911=>"00000001",
  38912=>"00000001",
  38913=>"11111111",
  38914=>"00000001",
  38915=>"11111111",
  38916=>"00000000",
  38917=>"00000001",
  38918=>"00000010",
  38919=>"00000010",
  38920=>"00000000",
  38921=>"11111111",
  38922=>"00000000",
  38923=>"00000010",
  38924=>"00000000",
  38925=>"00000001",
  38926=>"11111111",
  38927=>"00000000",
  38928=>"11111111",
  38929=>"00000000",
  38930=>"00000000",
  38931=>"11111110",
  38932=>"00000001",
  38933=>"00000001",
  38934=>"00000001",
  38935=>"11111110",
  38936=>"00000001",
  38937=>"11111110",
  38938=>"11111111",
  38939=>"00000010",
  38940=>"00000000",
  38941=>"00000000",
  38942=>"00000001",
  38943=>"11111110",
  38944=>"00000001",
  38945=>"00000001",
  38946=>"00000000",
  38947=>"11111111",
  38948=>"11111111",
  38949=>"00000000",
  38950=>"11111110",
  38951=>"00000001",
  38952=>"00000001",
  38953=>"00000000",
  38954=>"00000000",
  38955=>"00000000",
  38956=>"00000000",
  38957=>"00000001",
  38958=>"00000010",
  38959=>"00000000",
  38960=>"11111111",
  38961=>"00000000",
  38962=>"00000000",
  38963=>"11111110",
  38964=>"11111110",
  38965=>"00000000",
  38966=>"11111111",
  38967=>"00000001",
  38968=>"11111111",
  38969=>"00000000",
  38970=>"00000010",
  38971=>"00000001",
  38972=>"00000001",
  38973=>"00000001",
  38974=>"00000001",
  38975=>"00000000",
  38976=>"11111111",
  38977=>"11111111",
  38978=>"00000001",
  38979=>"00000010",
  38980=>"00000001",
  38981=>"00000001",
  38982=>"00000000",
  38983=>"11111111",
  38984=>"11111110",
  38985=>"11111110",
  38986=>"00000001",
  38987=>"00000000",
  38988=>"11111110",
  38989=>"00000001",
  38990=>"11111110",
  38991=>"11111111",
  38992=>"11111110",
  38993=>"00000000",
  38994=>"11111111",
  38995=>"11111111",
  38996=>"00000001",
  38997=>"00000000",
  38998=>"11111111",
  38999=>"11111111",
  39000=>"00000010",
  39001=>"11111111",
  39002=>"00000010",
  39003=>"00000001",
  39004=>"00000001",
  39005=>"00000001",
  39006=>"00000000",
  39007=>"11111111",
  39008=>"11111111",
  39009=>"00000010",
  39010=>"00000001",
  39011=>"00000001",
  39012=>"00000001",
  39013=>"00000000",
  39014=>"11111110",
  39015=>"11111110",
  39016=>"00000000",
  39017=>"11111110",
  39018=>"00000000",
  39019=>"00000001",
  39020=>"00000001",
  39021=>"00000000",
  39022=>"00000001",
  39023=>"00000001",
  39024=>"11111111",
  39025=>"11111111",
  39026=>"11111110",
  39027=>"00000001",
  39028=>"00000010",
  39029=>"11111111",
  39030=>"11111110",
  39031=>"00000001",
  39032=>"00000000",
  39033=>"11111110",
  39034=>"00000000",
  39035=>"11111111",
  39036=>"00000010",
  39037=>"00000001",
  39038=>"11111111",
  39039=>"00000010",
  39040=>"00000001",
  39041=>"11111111",
  39042=>"00000000",
  39043=>"00000000",
  39044=>"00000000",
  39045=>"00000001",
  39046=>"00000000",
  39047=>"11111111",
  39048=>"00000001",
  39049=>"11111111",
  39050=>"00000001",
  39051=>"00000001",
  39052=>"00000001",
  39053=>"00000000",
  39054=>"00000000",
  39055=>"00000010",
  39056=>"11111111",
  39057=>"00000000",
  39058=>"00000001",
  39059=>"11111111",
  39060=>"00000010",
  39061=>"00000001",
  39062=>"00000001",
  39063=>"00000000",
  39064=>"00000010",
  39065=>"00000000",
  39066=>"00000000",
  39067=>"00000000",
  39068=>"11111111",
  39069=>"00000000",
  39070=>"00000000",
  39071=>"00000010",
  39072=>"00000010",
  39073=>"00000000",
  39074=>"00000000",
  39075=>"00000000",
  39076=>"11111111",
  39077=>"11111111",
  39078=>"00000001",
  39079=>"11111111",
  39080=>"00000000",
  39081=>"00000010",
  39082=>"00000000",
  39083=>"11111111",
  39084=>"00000000",
  39085=>"11111111",
  39086=>"00000001",
  39087=>"00000001",
  39088=>"11111110",
  39089=>"00000000",
  39090=>"00000010",
  39091=>"00000010",
  39092=>"00000000",
  39093=>"00000000",
  39094=>"11111111",
  39095=>"00000000",
  39096=>"11111111",
  39097=>"00000001",
  39098=>"11111111",
  39099=>"11111111",
  39100=>"11111111",
  39101=>"11111110",
  39102=>"00000000",
  39103=>"00000000",
  39104=>"00000000",
  39105=>"00000010",
  39106=>"00000001",
  39107=>"00000000",
  39108=>"11111110",
  39109=>"00000000",
  39110=>"00000000",
  39111=>"00000000",
  39112=>"11111111",
  39113=>"00000000",
  39114=>"00000001",
  39115=>"00000010",
  39116=>"00000010",
  39117=>"00000000",
  39118=>"00000001",
  39119=>"00000010",
  39120=>"11111111",
  39121=>"00000001",
  39122=>"00000001",
  39123=>"00000010",
  39124=>"11111111",
  39125=>"00000001",
  39126=>"00000000",
  39127=>"00000000",
  39128=>"00000001",
  39129=>"11111110",
  39130=>"00000001",
  39131=>"11111111",
  39132=>"11111111",
  39133=>"11111111",
  39134=>"00000000",
  39135=>"00000001",
  39136=>"11111111",
  39137=>"00000000",
  39138=>"11111111",
  39139=>"11111111",
  39140=>"11111110",
  39141=>"00000010",
  39142=>"00000001",
  39143=>"00000000",
  39144=>"00000000",
  39145=>"11111111",
  39146=>"00000000",
  39147=>"11111111",
  39148=>"00000010",
  39149=>"11111111",
  39150=>"11111111",
  39151=>"11111110",
  39152=>"00000010",
  39153=>"00000001",
  39154=>"11111110",
  39155=>"11111111",
  39156=>"00000001",
  39157=>"00000001",
  39158=>"00000010",
  39159=>"00000000",
  39160=>"00000001",
  39161=>"00000001",
  39162=>"00000000",
  39163=>"00000010",
  39164=>"00000001",
  39165=>"00000010",
  39166=>"00000000",
  39167=>"11111111",
  39168=>"11111111",
  39169=>"00000001",
  39170=>"00000000",
  39171=>"11111111",
  39172=>"00000001",
  39173=>"00000010",
  39174=>"00000001",
  39175=>"11111111",
  39176=>"00000000",
  39177=>"11111111",
  39178=>"00000000",
  39179=>"11111110",
  39180=>"00000001",
  39181=>"00000000",
  39182=>"11111111",
  39183=>"00000000",
  39184=>"00000000",
  39185=>"00000000",
  39186=>"00000001",
  39187=>"00000001",
  39188=>"11111111",
  39189=>"00000000",
  39190=>"11111111",
  39191=>"00000001",
  39192=>"11111111",
  39193=>"00000001",
  39194=>"00000001",
  39195=>"11111110",
  39196=>"00000000",
  39197=>"00000000",
  39198=>"11111111",
  39199=>"00000001",
  39200=>"00000001",
  39201=>"00000000",
  39202=>"11111111",
  39203=>"00000001",
  39204=>"11111111",
  39205=>"00000000",
  39206=>"00000001",
  39207=>"00000000",
  39208=>"00000001",
  39209=>"11111110",
  39210=>"00000000",
  39211=>"11111111",
  39212=>"00000000",
  39213=>"00000010",
  39214=>"00000001",
  39215=>"00000001",
  39216=>"11111111",
  39217=>"00000000",
  39218=>"00000000",
  39219=>"00000000",
  39220=>"11111111",
  39221=>"11111110",
  39222=>"11111111",
  39223=>"00000000",
  39224=>"00000001",
  39225=>"11111111",
  39226=>"00000000",
  39227=>"00000000",
  39228=>"11111111",
  39229=>"00000001",
  39230=>"11111111",
  39231=>"11111111",
  39232=>"11111111",
  39233=>"00000001",
  39234=>"00000001",
  39235=>"00000001",
  39236=>"00000010",
  39237=>"00000001",
  39238=>"11111111",
  39239=>"00000000",
  39240=>"00000001",
  39241=>"00000010",
  39242=>"00000010",
  39243=>"11111111",
  39244=>"00000001",
  39245=>"00000001",
  39246=>"00000010",
  39247=>"11111110",
  39248=>"00000001",
  39249=>"00000000",
  39250=>"11111111",
  39251=>"00000010",
  39252=>"00000001",
  39253=>"00000000",
  39254=>"11111111",
  39255=>"00000000",
  39256=>"00000001",
  39257=>"11111111",
  39258=>"00000010",
  39259=>"00000010",
  39260=>"00000001",
  39261=>"11111111",
  39262=>"11111111",
  39263=>"11111111",
  39264=>"11111110",
  39265=>"11111111",
  39266=>"00000001",
  39267=>"11111111",
  39268=>"00000001",
  39269=>"00000010",
  39270=>"00000000",
  39271=>"00000000",
  39272=>"00000010",
  39273=>"00000001",
  39274=>"00000010",
  39275=>"00000000",
  39276=>"11111111",
  39277=>"00000001",
  39278=>"00000000",
  39279=>"00000001",
  39280=>"00000000",
  39281=>"11111110",
  39282=>"00000000",
  39283=>"11111111",
  39284=>"00000000",
  39285=>"00000001",
  39286=>"00000000",
  39287=>"00000000",
  39288=>"00000001",
  39289=>"00000000",
  39290=>"11111111",
  39291=>"00000001",
  39292=>"00000001",
  39293=>"00000000",
  39294=>"00000010",
  39295=>"00000001",
  39296=>"00000001",
  39297=>"00000000",
  39298=>"00000001",
  39299=>"00000000",
  39300=>"00000000",
  39301=>"00000000",
  39302=>"11111110",
  39303=>"11111111",
  39304=>"00000010",
  39305=>"00000001",
  39306=>"11111110",
  39307=>"00000000",
  39308=>"00000001",
  39309=>"00000001",
  39310=>"00000001",
  39311=>"00000000",
  39312=>"00000001",
  39313=>"00000000",
  39314=>"11111111",
  39315=>"11111111",
  39316=>"00000000",
  39317=>"11111111",
  39318=>"00000001",
  39319=>"11111111",
  39320=>"00000000",
  39321=>"11111111",
  39322=>"00000010",
  39323=>"11111111",
  39324=>"00000000",
  39325=>"00000001",
  39326=>"11111111",
  39327=>"11111111",
  39328=>"11111111",
  39329=>"00000010",
  39330=>"00000000",
  39331=>"00000001",
  39332=>"00000000",
  39333=>"00000001",
  39334=>"11111111",
  39335=>"00000000",
  39336=>"00000001",
  39337=>"11111111",
  39338=>"00000000",
  39339=>"11111111",
  39340=>"00000001",
  39341=>"11111111",
  39342=>"00000001",
  39343=>"00000000",
  39344=>"00000001",
  39345=>"11111111",
  39346=>"11111101",
  39347=>"11111111",
  39348=>"11111111",
  39349=>"00000001",
  39350=>"11111111",
  39351=>"00000001",
  39352=>"00000001",
  39353=>"11111111",
  39354=>"00000010",
  39355=>"11111111",
  39356=>"00000010",
  39357=>"11111111",
  39358=>"00000000",
  39359=>"11111111",
  39360=>"11111110",
  39361=>"11111111",
  39362=>"11111110",
  39363=>"11111111",
  39364=>"00000001",
  39365=>"11111110",
  39366=>"00000001",
  39367=>"00000000",
  39368=>"11111111",
  39369=>"11111111",
  39370=>"00000001",
  39371=>"11111110",
  39372=>"00000000",
  39373=>"11111111",
  39374=>"00000001",
  39375=>"00000000",
  39376=>"00000000",
  39377=>"00000001",
  39378=>"00000000",
  39379=>"00000001",
  39380=>"00000001",
  39381=>"11111110",
  39382=>"00000000",
  39383=>"11111111",
  39384=>"00000000",
  39385=>"00000000",
  39386=>"00000001",
  39387=>"11111111",
  39388=>"00000000",
  39389=>"11111111",
  39390=>"00000000",
  39391=>"11111111",
  39392=>"11111111",
  39393=>"00000001",
  39394=>"00000001",
  39395=>"11111101",
  39396=>"11111111",
  39397=>"11111111",
  39398=>"11111111",
  39399=>"00000010",
  39400=>"00000001",
  39401=>"11111110",
  39402=>"11111110",
  39403=>"11111111",
  39404=>"11111111",
  39405=>"00000001",
  39406=>"00000001",
  39407=>"00000001",
  39408=>"00000000",
  39409=>"00000000",
  39410=>"00000000",
  39411=>"11111111",
  39412=>"00000000",
  39413=>"00000001",
  39414=>"00000000",
  39415=>"00000001",
  39416=>"11111110",
  39417=>"11111110",
  39418=>"11111111",
  39419=>"00000000",
  39420=>"11111111",
  39421=>"00000000",
  39422=>"00000010",
  39423=>"00000000",
  39424=>"11111110",
  39425=>"00000001",
  39426=>"00000000",
  39427=>"00000000",
  39428=>"11111111",
  39429=>"00000001",
  39430=>"00000000",
  39431=>"00000001",
  39432=>"00000010",
  39433=>"00000001",
  39434=>"11111111",
  39435=>"00000000",
  39436=>"00000001",
  39437=>"11111111",
  39438=>"11111111",
  39439=>"11111111",
  39440=>"11111111",
  39441=>"00000001",
  39442=>"11111111",
  39443=>"00000010",
  39444=>"00000000",
  39445=>"00000001",
  39446=>"00000001",
  39447=>"00000001",
  39448=>"00000010",
  39449=>"00000001",
  39450=>"11111111",
  39451=>"11111111",
  39452=>"00000000",
  39453=>"11111111",
  39454=>"00000001",
  39455=>"11111111",
  39456=>"00000001",
  39457=>"11111111",
  39458=>"11111110",
  39459=>"11111110",
  39460=>"11111111",
  39461=>"00000001",
  39462=>"00000001",
  39463=>"11111111",
  39464=>"00000000",
  39465=>"11111111",
  39466=>"00000000",
  39467=>"11111111",
  39468=>"11111111",
  39469=>"00000001",
  39470=>"11111111",
  39471=>"00000000",
  39472=>"00000000",
  39473=>"00000001",
  39474=>"00000000",
  39475=>"11111110",
  39476=>"11111111",
  39477=>"11111111",
  39478=>"00000001",
  39479=>"11111111",
  39480=>"11111110",
  39481=>"11111111",
  39482=>"11111111",
  39483=>"11111111",
  39484=>"00000000",
  39485=>"11111110",
  39486=>"00000000",
  39487=>"11111111",
  39488=>"00000000",
  39489=>"00000000",
  39490=>"11111111",
  39491=>"00000000",
  39492=>"00000000",
  39493=>"11111111",
  39494=>"00000001",
  39495=>"00000010",
  39496=>"11111111",
  39497=>"00000000",
  39498=>"11111111",
  39499=>"00000000",
  39500=>"00000000",
  39501=>"00000000",
  39502=>"00000010",
  39503=>"00000010",
  39504=>"11111111",
  39505=>"11111111",
  39506=>"11111110",
  39507=>"11111111",
  39508=>"00000001",
  39509=>"11111110",
  39510=>"00000000",
  39511=>"00000001",
  39512=>"11111111",
  39513=>"00000010",
  39514=>"11111110",
  39515=>"00000000",
  39516=>"11111110",
  39517=>"00000001",
  39518=>"00000000",
  39519=>"00000000",
  39520=>"00000000",
  39521=>"00000001",
  39522=>"11111111",
  39523=>"00000010",
  39524=>"00000010",
  39525=>"11111111",
  39526=>"00000001",
  39527=>"11111111",
  39528=>"00000001",
  39529=>"00000010",
  39530=>"00000001",
  39531=>"11111110",
  39532=>"00000000",
  39533=>"00000000",
  39534=>"00000001",
  39535=>"00000000",
  39536=>"11111111",
  39537=>"00000010",
  39538=>"00000010",
  39539=>"00000010",
  39540=>"11111101",
  39541=>"00000000",
  39542=>"00000001",
  39543=>"11111111",
  39544=>"00000000",
  39545=>"00000010",
  39546=>"00000001",
  39547=>"00000000",
  39548=>"00000001",
  39549=>"00000000",
  39550=>"11111111",
  39551=>"00000000",
  39552=>"00000000",
  39553=>"11111111",
  39554=>"11111111",
  39555=>"11111111",
  39556=>"11111111",
  39557=>"11111111",
  39558=>"00000000",
  39559=>"11111111",
  39560=>"11111110",
  39561=>"11111111",
  39562=>"11111111",
  39563=>"00000000",
  39564=>"00000001",
  39565=>"11111110",
  39566=>"11111110",
  39567=>"11111110",
  39568=>"11111110",
  39569=>"00000001",
  39570=>"11111111",
  39571=>"11111110",
  39572=>"00000000",
  39573=>"00000001",
  39574=>"11111111",
  39575=>"00000010",
  39576=>"00000001",
  39577=>"11111110",
  39578=>"00000000",
  39579=>"00000001",
  39580=>"00000000",
  39581=>"00000001",
  39582=>"00000001",
  39583=>"00000001",
  39584=>"11111110",
  39585=>"11111110",
  39586=>"11111110",
  39587=>"00000000",
  39588=>"11111111",
  39589=>"00000001",
  39590=>"00000001",
  39591=>"00000000",
  39592=>"11111111",
  39593=>"00000000",
  39594=>"11111110",
  39595=>"11111110",
  39596=>"00000001",
  39597=>"11111110",
  39598=>"11111111",
  39599=>"00000001",
  39600=>"11111111",
  39601=>"11111111",
  39602=>"00000010",
  39603=>"00000000",
  39604=>"00000001",
  39605=>"11111111",
  39606=>"00000000",
  39607=>"00000001",
  39608=>"11111111",
  39609=>"11111110",
  39610=>"11111110",
  39611=>"00000001",
  39612=>"00000000",
  39613=>"11111111",
  39614=>"00000001",
  39615=>"00000001",
  39616=>"11111111",
  39617=>"00000010",
  39618=>"11111111",
  39619=>"00000000",
  39620=>"00000001",
  39621=>"00000010",
  39622=>"00000001",
  39623=>"00000010",
  39624=>"00000001",
  39625=>"00000001",
  39626=>"00000010",
  39627=>"11111111",
  39628=>"11111110",
  39629=>"00000010",
  39630=>"11111110",
  39631=>"11111111",
  39632=>"11111110",
  39633=>"11111111",
  39634=>"00000000",
  39635=>"00000010",
  39636=>"11111111",
  39637=>"11111111",
  39638=>"00000000",
  39639=>"00000000",
  39640=>"11111111",
  39641=>"00000001",
  39642=>"11111110",
  39643=>"00000010",
  39644=>"00000001",
  39645=>"00000001",
  39646=>"00000001",
  39647=>"00000010",
  39648=>"00000001",
  39649=>"00000010",
  39650=>"11111111",
  39651=>"00000000",
  39652=>"00000001",
  39653=>"00000000",
  39654=>"00000000",
  39655=>"00000000",
  39656=>"11111111",
  39657=>"11111111",
  39658=>"00000001",
  39659=>"11111111",
  39660=>"00000000",
  39661=>"11111101",
  39662=>"00000000",
  39663=>"00000000",
  39664=>"11111111",
  39665=>"11111111",
  39666=>"11111111",
  39667=>"11111111",
  39668=>"11111111",
  39669=>"00000001",
  39670=>"00000001",
  39671=>"11111111",
  39672=>"00000000",
  39673=>"00000001",
  39674=>"11111111",
  39675=>"11111111",
  39676=>"11111111",
  39677=>"00000001",
  39678=>"11111111",
  39679=>"00000001",
  39680=>"00000001",
  39681=>"00000000",
  39682=>"11111111",
  39683=>"00000000",
  39684=>"00000010",
  39685=>"00000001",
  39686=>"11111110",
  39687=>"11111111",
  39688=>"11111111",
  39689=>"00000010",
  39690=>"00000001",
  39691=>"00000000",
  39692=>"00000001",
  39693=>"11111111",
  39694=>"00000001",
  39695=>"00000010",
  39696=>"11111111",
  39697=>"11111111",
  39698=>"11111111",
  39699=>"11111111",
  39700=>"00000001",
  39701=>"00000001",
  39702=>"00000000",
  39703=>"11111111",
  39704=>"11111111",
  39705=>"00000000",
  39706=>"00000000",
  39707=>"00000001",
  39708=>"11111111",
  39709=>"00000001",
  39710=>"00000000",
  39711=>"00000000",
  39712=>"11111111",
  39713=>"11111110",
  39714=>"00000001",
  39715=>"11111111",
  39716=>"00000010",
  39717=>"00000010",
  39718=>"00000000",
  39719=>"11111110",
  39720=>"00000001",
  39721=>"00000000",
  39722=>"00000000",
  39723=>"00000001",
  39724=>"00000000",
  39725=>"11111111",
  39726=>"00000000",
  39727=>"00000001",
  39728=>"00000000",
  39729=>"00000001",
  39730=>"00000001",
  39731=>"00000000",
  39732=>"00000000",
  39733=>"11111111",
  39734=>"00000001",
  39735=>"00000010",
  39736=>"00000001",
  39737=>"11111111",
  39738=>"00000000",
  39739=>"11111111",
  39740=>"11111111",
  39741=>"11111111",
  39742=>"00000000",
  39743=>"00000000",
  39744=>"11111111",
  39745=>"00000000",
  39746=>"00000001",
  39747=>"11111111",
  39748=>"11111111",
  39749=>"00000000",
  39750=>"11111111",
  39751=>"00000001",
  39752=>"00000001",
  39753=>"00000000",
  39754=>"00000000",
  39755=>"11111111",
  39756=>"11111110",
  39757=>"11111111",
  39758=>"00000001",
  39759=>"00000000",
  39760=>"00000001",
  39761=>"00000001",
  39762=>"11111111",
  39763=>"00000000",
  39764=>"11111110",
  39765=>"00000001",
  39766=>"11111111",
  39767=>"00000001",
  39768=>"11111110",
  39769=>"00000001",
  39770=>"00000000",
  39771=>"11111111",
  39772=>"11111111",
  39773=>"00000001",
  39774=>"00000000",
  39775=>"00000000",
  39776=>"11111110",
  39777=>"00000000",
  39778=>"00000000",
  39779=>"11111111",
  39780=>"00000001",
  39781=>"00000001",
  39782=>"11111110",
  39783=>"11111111",
  39784=>"11111111",
  39785=>"00000001",
  39786=>"00000000",
  39787=>"00000000",
  39788=>"00000001",
  39789=>"00000000",
  39790=>"11111111",
  39791=>"00000001",
  39792=>"11111111",
  39793=>"11111111",
  39794=>"11111110",
  39795=>"11111111",
  39796=>"00000001",
  39797=>"00000000",
  39798=>"11111111",
  39799=>"11111110",
  39800=>"00000000",
  39801=>"00000000",
  39802=>"11111111",
  39803=>"11111111",
  39804=>"11111111",
  39805=>"00000001",
  39806=>"00000000",
  39807=>"00000000",
  39808=>"11111110",
  39809=>"00000000",
  39810=>"00000000",
  39811=>"00000001",
  39812=>"00000010",
  39813=>"00000001",
  39814=>"11111110",
  39815=>"00000000",
  39816=>"11111111",
  39817=>"00000001",
  39818=>"00000001",
  39819=>"11111111",
  39820=>"11111111",
  39821=>"00000000",
  39822=>"00000001",
  39823=>"11111111",
  39824=>"00000010",
  39825=>"00000010",
  39826=>"00000000",
  39827=>"00000001",
  39828=>"11111111",
  39829=>"00000001",
  39830=>"00000001",
  39831=>"00000000",
  39832=>"11111110",
  39833=>"11111110",
  39834=>"11111111",
  39835=>"00000000",
  39836=>"00000010",
  39837=>"00000001",
  39838=>"00000000",
  39839=>"11111111",
  39840=>"11111111",
  39841=>"00000010",
  39842=>"00000010",
  39843=>"11111111",
  39844=>"00000000",
  39845=>"11111110",
  39846=>"11111111",
  39847=>"00000001",
  39848=>"00000010",
  39849=>"11111111",
  39850=>"00000001",
  39851=>"11111110",
  39852=>"00000001",
  39853=>"00000000",
  39854=>"00000000",
  39855=>"00000001",
  39856=>"00000001",
  39857=>"00000000",
  39858=>"00000000",
  39859=>"11111110",
  39860=>"00000000",
  39861=>"11111111",
  39862=>"00000000",
  39863=>"00000000",
  39864=>"11111111",
  39865=>"00000001",
  39866=>"00000010",
  39867=>"11111110",
  39868=>"00000001",
  39869=>"00000000",
  39870=>"11111111",
  39871=>"00000001",
  39872=>"00000000",
  39873=>"11111110",
  39874=>"00000001",
  39875=>"11111110",
  39876=>"11111111",
  39877=>"00000000",
  39878=>"00000001",
  39879=>"11111110",
  39880=>"11111111",
  39881=>"00000001",
  39882=>"11111110",
  39883=>"11111111",
  39884=>"00000001",
  39885=>"00000000",
  39886=>"00000001",
  39887=>"11111111",
  39888=>"11111101",
  39889=>"00000000",
  39890=>"11111111",
  39891=>"00000001",
  39892=>"00000001",
  39893=>"00000001",
  39894=>"00000000",
  39895=>"11111111",
  39896=>"00000001",
  39897=>"00000000",
  39898=>"11111111",
  39899=>"00000000",
  39900=>"00000001",
  39901=>"00000000",
  39902=>"11111111",
  39903=>"00000000",
  39904=>"00000000",
  39905=>"11111110",
  39906=>"11111111",
  39907=>"00000001",
  39908=>"00000000",
  39909=>"00000000",
  39910=>"00000001",
  39911=>"00000001",
  39912=>"11111110",
  39913=>"00000001",
  39914=>"11111111",
  39915=>"00000000",
  39916=>"11111111",
  39917=>"11111110",
  39918=>"00000010",
  39919=>"00000001",
  39920=>"00000000",
  39921=>"11111110",
  39922=>"00000000",
  39923=>"11111111",
  39924=>"00000010",
  39925=>"00000001",
  39926=>"11111111",
  39927=>"00000001",
  39928=>"11111111",
  39929=>"11111111",
  39930=>"11111111",
  39931=>"11111111",
  39932=>"00000001",
  39933=>"00000000",
  39934=>"00000000",
  39935=>"11111111",
  39936=>"00000000",
  39937=>"00000000",
  39938=>"00000000",
  39939=>"00000000",
  39940=>"00000000",
  39941=>"00000000",
  39942=>"00000000",
  39943=>"00000000",
  39944=>"00000000",
  39945=>"00000000",
  39946=>"00000000",
  39947=>"00000000",
  39948=>"00000000",
  39949=>"00000000",
  39950=>"00000000",
  39951=>"00000000",
  39952=>"00000000",
  39953=>"00000000",
  39954=>"00000000",
  39955=>"00000000",
  39956=>"00000000",
  39957=>"00000000",
  39958=>"00000000",
  39959=>"00000000",
  39960=>"00000000",
  39961=>"00000000",
  39962=>"00000000",
  39963=>"00000000",
  39964=>"00000000",
  39965=>"00000000",
  39966=>"00000000",
  39967=>"00000000",
  39968=>"00000000",
  39969=>"00000000",
  39970=>"00000000",
  39971=>"00000000",
  39972=>"00000000",
  39973=>"00000000",
  39974=>"00000000",
  39975=>"00000000",
  39976=>"00000000",
  39977=>"00000000",
  39978=>"00000000",
  39979=>"00000000",
  39980=>"00000001",
  39981=>"00000000",
  39982=>"00000000",
  39983=>"00000000",
  39984=>"00000000",
  39985=>"00000000",
  39986=>"00000000",
  39987=>"00000000",
  39988=>"00000000",
  39989=>"00000000",
  39990=>"00000000",
  39991=>"00000000",
  39992=>"00000000",
  39993=>"00000000",
  39994=>"00000000",
  39995=>"00000000",
  39996=>"00000000",
  39997=>"00000000",
  39998=>"00000000",
  39999=>"00000000",
  40000=>"00000000",
  40001=>"00000000",
  40002=>"00000000",
  40003=>"00000000",
  40004=>"00000000",
  40005=>"00000000",
  40006=>"00000000",
  40007=>"00000000",
  40008=>"00000000",
  40009=>"00000000",
  40010=>"00000000",
  40011=>"00000000",
  40012=>"00000000",
  40013=>"00000000",
  40014=>"00000000",
  40015=>"00000000",
  40016=>"00000000",
  40017=>"00000000",
  40018=>"00000000",
  40019=>"00000000",
  40020=>"00000000",
  40021=>"00000000",
  40022=>"00000000",
  40023=>"00000000",
  40024=>"00000000",
  40025=>"00000000",
  40026=>"00000000",
  40027=>"00000000",
  40028=>"00000000",
  40029=>"00000000",
  40030=>"00000000",
  40031=>"00000000",
  40032=>"00000000",
  40033=>"00000000",
  40034=>"00000000",
  40035=>"00000000",
  40036=>"00000000",
  40037=>"00000000",
  40038=>"00000000",
  40039=>"00000000",
  40040=>"00000000",
  40041=>"00000000",
  40042=>"00000000",
  40043=>"00000000",
  40044=>"00000000",
  40045=>"00000000",
  40046=>"00000000",
  40047=>"00000000",
  40048=>"00000000",
  40049=>"00000000",
  40050=>"00000000",
  40051=>"00000000",
  40052=>"00000000",
  40053=>"00000000",
  40054=>"00000000",
  40055=>"00000000",
  40056=>"00000000",
  40057=>"00000000",
  40058=>"00000000",
  40059=>"00000000",
  40060=>"00000000",
  40061=>"00000000",
  40062=>"00000000",
  40063=>"00000000",
  40064=>"00000000",
  40065=>"00000000",
  40066=>"00000000",
  40067=>"00000000",
  40068=>"00000000",
  40069=>"00000000",
  40070=>"00000000",
  40071=>"00000000",
  40072=>"00000000",
  40073=>"00000000",
  40074=>"00000000",
  40075=>"00000000",
  40076=>"00000000",
  40077=>"00000000",
  40078=>"00000000",
  40079=>"00000000",
  40080=>"00000000",
  40081=>"00000000",
  40082=>"00000000",
  40083=>"00000000",
  40084=>"00000000",
  40085=>"00000000",
  40086=>"00000000",
  40087=>"00000000",
  40088=>"00000000",
  40089=>"00000000",
  40090=>"00000000",
  40091=>"00000000",
  40092=>"00000000",
  40093=>"00000000",
  40094=>"00000000",
  40095=>"00000000",
  40096=>"00000000",
  40097=>"00000000",
  40098=>"00000000",
  40099=>"00000000",
  40100=>"00000001",
  40101=>"00000000",
  40102=>"00000000",
  40103=>"00000000",
  40104=>"00000000",
  40105=>"00000000",
  40106=>"00000000",
  40107=>"00000000",
  40108=>"00000000",
  40109=>"00000000",
  40110=>"00000000",
  40111=>"00000000",
  40112=>"00000000",
  40113=>"00000000",
  40114=>"00000000",
  40115=>"00000000",
  40116=>"00000000",
  40117=>"00000000",
  40118=>"00000000",
  40119=>"00000000",
  40120=>"00000000",
  40121=>"00000000",
  40122=>"00000000",
  40123=>"00000000",
  40124=>"00000000",
  40125=>"11111111",
  40126=>"00000000",
  40127=>"00000000",
  40128=>"00000000",
  40129=>"00000001",
  40130=>"00000000",
  40131=>"00000000",
  40132=>"00000000",
  40133=>"00000000",
  40134=>"00000000",
  40135=>"00000000",
  40136=>"00000000",
  40137=>"00000000",
  40138=>"00000000",
  40139=>"00000000",
  40140=>"00000000",
  40141=>"00000000",
  40142=>"00000000",
  40143=>"00000000",
  40144=>"00000000",
  40145=>"00000000",
  40146=>"00000001",
  40147=>"00000000",
  40148=>"00000000",
  40149=>"00000000",
  40150=>"00000000",
  40151=>"00000000",
  40152=>"00000000",
  40153=>"00000000",
  40154=>"00000000",
  40155=>"00000000",
  40156=>"00000000",
  40157=>"00000000",
  40158=>"00000000",
  40159=>"00000000",
  40160=>"00000000",
  40161=>"00000000",
  40162=>"00000000",
  40163=>"00000000",
  40164=>"00000000",
  40165=>"00000000",
  40166=>"00000000",
  40167=>"00000000",
  40168=>"00000000",
  40169=>"00000000",
  40170=>"00000000",
  40171=>"00000000",
  40172=>"00000000",
  40173=>"00000000",
  40174=>"00000000",
  40175=>"11111111",
  40176=>"00000000",
  40177=>"00000000",
  40178=>"00000000",
  40179=>"00000000",
  40180=>"00000000",
  40181=>"00000000",
  40182=>"00000000",
  40183=>"00000000",
  40184=>"00000000",
  40185=>"00000000",
  40186=>"00000000",
  40187=>"00000000",
  40188=>"00000000",
  40189=>"00000000",
  40190=>"00000000",
  40191=>"00000000",
  40192=>"00000000",
  40193=>"00000000",
  40194=>"00000000",
  40195=>"00000000",
  40196=>"00000000",
  40197=>"00000000",
  40198=>"00000000",
  40199=>"00000000",
  40200=>"00000000",
  40201=>"00000000",
  40202=>"00000000",
  40203=>"00000000",
  40204=>"00000000",
  40205=>"00000000",
  40206=>"00000000",
  40207=>"00000000",
  40208=>"00000000",
  40209=>"00000000",
  40210=>"00000000",
  40211=>"00000000",
  40212=>"00000000",
  40213=>"00000000",
  40214=>"00000000",
  40215=>"00000000",
  40216=>"00000000",
  40217=>"00000000",
  40218=>"00000000",
  40219=>"11111111",
  40220=>"00000000",
  40221=>"00000000",
  40222=>"00000000",
  40223=>"00000000",
  40224=>"00000000",
  40225=>"00000000",
  40226=>"00000000",
  40227=>"00000000",
  40228=>"00000000",
  40229=>"00000000",
  40230=>"00000000",
  40231=>"00000000",
  40232=>"00000000",
  40233=>"00000000",
  40234=>"00000000",
  40235=>"00000000",
  40236=>"00000000",
  40237=>"00000000",
  40238=>"00000000",
  40239=>"00000000",
  40240=>"00000000",
  40241=>"00000000",
  40242=>"11111111",
  40243=>"00000000",
  40244=>"00000000",
  40245=>"00000000",
  40246=>"00000000",
  40247=>"00000000",
  40248=>"00000000",
  40249=>"00000000",
  40250=>"11111111",
  40251=>"00000000",
  40252=>"00000000",
  40253=>"00000000",
  40254=>"00000000",
  40255=>"00000000",
  40256=>"00000000",
  40257=>"00000000",
  40258=>"00000000",
  40259=>"00000000",
  40260=>"00000000",
  40261=>"00000000",
  40262=>"00000000",
  40263=>"00000000",
  40264=>"00000000",
  40265=>"00000000",
  40266=>"00000000",
  40267=>"00000000",
  40268=>"00000000",
  40269=>"00000000",
  40270=>"00000000",
  40271=>"00000000",
  40272=>"00000000",
  40273=>"00000000",
  40274=>"00000000",
  40275=>"00000000",
  40276=>"00000000",
  40277=>"00000000",
  40278=>"00000000",
  40279=>"00000000",
  40280=>"00000000",
  40281=>"00000000",
  40282=>"00000000",
  40283=>"00000000",
  40284=>"00000000",
  40285=>"00000000",
  40286=>"00000000",
  40287=>"00000000",
  40288=>"00000000",
  40289=>"00000000",
  40290=>"00000000",
  40291=>"00000000",
  40292=>"00000000",
  40293=>"00000000",
  40294=>"11111111",
  40295=>"00000000",
  40296=>"00000000",
  40297=>"00000000",
  40298=>"00000000",
  40299=>"00000000",
  40300=>"00000000",
  40301=>"00000000",
  40302=>"00000000",
  40303=>"00000000",
  40304=>"00000000",
  40305=>"00000000",
  40306=>"00000000",
  40307=>"00000000",
  40308=>"00000000",
  40309=>"00000000",
  40310=>"00000000",
  40311=>"00000000",
  40312=>"00000000",
  40313=>"00000000",
  40314=>"00000000",
  40315=>"00000000",
  40316=>"00000000",
  40317=>"00000000",
  40318=>"00000000",
  40319=>"00000000",
  40320=>"00000000",
  40321=>"00000000",
  40322=>"00000000",
  40323=>"00000000",
  40324=>"00000000",
  40325=>"00000000",
  40326=>"00000000",
  40327=>"00000000",
  40328=>"00000000",
  40329=>"00000000",
  40330=>"00000000",
  40331=>"00000000",
  40332=>"00000000",
  40333=>"00000000",
  40334=>"00000000",
  40335=>"00000000",
  40336=>"00000000",
  40337=>"00000000",
  40338=>"00000000",
  40339=>"00000000",
  40340=>"00000000",
  40341=>"00000000",
  40342=>"00000000",
  40343=>"00000000",
  40344=>"00000000",
  40345=>"00000000",
  40346=>"00000000",
  40347=>"00000000",
  40348=>"00000000",
  40349=>"00000000",
  40350=>"00000000",
  40351=>"00000000",
  40352=>"00000000",
  40353=>"00000000",
  40354=>"00000000",
  40355=>"00000000",
  40356=>"00000000",
  40357=>"00000000",
  40358=>"00000000",
  40359=>"00000000",
  40360=>"00000000",
  40361=>"00000000",
  40362=>"00000000",
  40363=>"00000000",
  40364=>"00000000",
  40365=>"00000000",
  40366=>"00000000",
  40367=>"00000000",
  40368=>"00000000",
  40369=>"00000000",
  40370=>"00000000",
  40371=>"00000000",
  40372=>"00000000",
  40373=>"00000000",
  40374=>"00000000",
  40375=>"00000000",
  40376=>"00000000",
  40377=>"00000000",
  40378=>"00000000",
  40379=>"00000000",
  40380=>"00000000",
  40381=>"00000000",
  40382=>"00000000",
  40383=>"00000000",
  40384=>"00000000",
  40385=>"00000000",
  40386=>"00000000",
  40387=>"00000000",
  40388=>"00000000",
  40389=>"00000000",
  40390=>"00000000",
  40391=>"00000000",
  40392=>"00000000",
  40393=>"00000000",
  40394=>"00000000",
  40395=>"00000000",
  40396=>"00000000",
  40397=>"00000000",
  40398=>"00000000",
  40399=>"00000000",
  40400=>"00000000",
  40401=>"00000000",
  40402=>"00000000",
  40403=>"00000000",
  40404=>"00000000",
  40405=>"00000000",
  40406=>"00000000",
  40407=>"00000000",
  40408=>"00000000",
  40409=>"00000000",
  40410=>"00000000",
  40411=>"00000000",
  40412=>"00000000",
  40413=>"00000000",
  40414=>"00000000",
  40415=>"00000000",
  40416=>"00000000",
  40417=>"00000000",
  40418=>"00000000",
  40419=>"00000000",
  40420=>"00000000",
  40421=>"00000000",
  40422=>"00000000",
  40423=>"00000000",
  40424=>"00000000",
  40425=>"00000000",
  40426=>"00000000",
  40427=>"00000000",
  40428=>"11111111",
  40429=>"00000000",
  40430=>"00000000",
  40431=>"00000000",
  40432=>"00000000",
  40433=>"00000000",
  40434=>"00000000",
  40435=>"00000000",
  40436=>"00000000",
  40437=>"00000000",
  40438=>"00000000",
  40439=>"00000000",
  40440=>"00000000",
  40441=>"00000000",
  40442=>"00000000",
  40443=>"00000000",
  40444=>"00000000",
  40445=>"00000000",
  40446=>"00000000",
  40447=>"00000000",
  40448=>"00000001",
  40449=>"00000000",
  40450=>"00000000",
  40451=>"00000000",
  40452=>"00000000",
  40453=>"00000000",
  40454=>"00000000",
  40455=>"00000000",
  40456=>"00000000",
  40457=>"00000000",
  40458=>"00000000",
  40459=>"00000000",
  40460=>"00000000",
  40461=>"00000000",
  40462=>"00000000",
  40463=>"00000000",
  40464=>"00000000",
  40465=>"00000000",
  40466=>"00000000",
  40467=>"00000000",
  40468=>"00000000",
  40469=>"00000000",
  40470=>"00000000",
  40471=>"00000000",
  40472=>"00000000",
  40473=>"00000000",
  40474=>"00000000",
  40475=>"00000000",
  40476=>"00000000",
  40477=>"00000000",
  40478=>"00000000",
  40479=>"00000000",
  40480=>"00000000",
  40481=>"00000000",
  40482=>"00000000",
  40483=>"00000000",
  40484=>"00000000",
  40485=>"00000000",
  40486=>"00000000",
  40487=>"00000000",
  40488=>"00000000",
  40489=>"00000000",
  40490=>"00000000",
  40491=>"00000000",
  40492=>"00000000",
  40493=>"00000000",
  40494=>"00000000",
  40495=>"00000000",
  40496=>"00000000",
  40497=>"00000000",
  40498=>"00000000",
  40499=>"00000000",
  40500=>"00000000",
  40501=>"00000000",
  40502=>"00000000",
  40503=>"00000000",
  40504=>"00000000",
  40505=>"00000000",
  40506=>"00000000",
  40507=>"00000000",
  40508=>"00000000",
  40509=>"00000000",
  40510=>"00000000",
  40511=>"00000000",
  40512=>"00000000",
  40513=>"00000000",
  40514=>"00000000",
  40515=>"00000000",
  40516=>"00000000",
  40517=>"00000000",
  40518=>"00000000",
  40519=>"00000000",
  40520=>"00000000",
  40521=>"00000000",
  40522=>"00000000",
  40523=>"00000000",
  40524=>"00000000",
  40525=>"00000000",
  40526=>"00000000",
  40527=>"00000000",
  40528=>"00000000",
  40529=>"00000000",
  40530=>"00000000",
  40531=>"00000000",
  40532=>"00000000",
  40533=>"00000000",
  40534=>"00000000",
  40535=>"00000000",
  40536=>"00000000",
  40537=>"00000000",
  40538=>"00000000",
  40539=>"00000000",
  40540=>"00000000",
  40541=>"00000000",
  40542=>"00000000",
  40543=>"00000000",
  40544=>"00000000",
  40545=>"00000000",
  40546=>"00000000",
  40547=>"00000000",
  40548=>"00000000",
  40549=>"00000000",
  40550=>"00000000",
  40551=>"00000000",
  40552=>"00000000",
  40553=>"00000000",
  40554=>"00000000",
  40555=>"00000000",
  40556=>"00000000",
  40557=>"00000000",
  40558=>"00000000",
  40559=>"00000000",
  40560=>"00000000",
  40561=>"00000000",
  40562=>"00000000",
  40563=>"00000000",
  40564=>"00000000",
  40565=>"00000000",
  40566=>"00000000",
  40567=>"00000000",
  40568=>"00000000",
  40569=>"00000000",
  40570=>"00000000",
  40571=>"00000000",
  40572=>"00000000",
  40573=>"00000000",
  40574=>"00000000",
  40575=>"00000000",
  40576=>"00000000",
  40577=>"00000000",
  40578=>"00000000",
  40579=>"00000000",
  40580=>"00000000",
  40581=>"00000000",
  40582=>"00000000",
  40583=>"00000000",
  40584=>"00000000",
  40585=>"00000000",
  40586=>"00000000",
  40587=>"00000000",
  40588=>"00000000",
  40589=>"00000001",
  40590=>"00000000",
  40591=>"00000000",
  40592=>"00000000",
  40593=>"00000000",
  40594=>"00000000",
  40595=>"00000000",
  40596=>"00000000",
  40597=>"00000000",
  40598=>"00000000",
  40599=>"00000000",
  40600=>"00000000",
  40601=>"00000000",
  40602=>"00000000",
  40603=>"00000001",
  40604=>"00000000",
  40605=>"00000000",
  40606=>"00000000",
  40607=>"00000000",
  40608=>"00000000",
  40609=>"00000000",
  40610=>"00000000",
  40611=>"00000000",
  40612=>"00000000",
  40613=>"00000000",
  40614=>"00000000",
  40615=>"00000000",
  40616=>"00000000",
  40617=>"00000000",
  40618=>"00000000",
  40619=>"00000000",
  40620=>"00000000",
  40621=>"00000000",
  40622=>"00000000",
  40623=>"00000000",
  40624=>"00000000",
  40625=>"00000000",
  40626=>"00000000",
  40627=>"00000000",
  40628=>"00000000",
  40629=>"00000000",
  40630=>"00000000",
  40631=>"00000000",
  40632=>"00000000",
  40633=>"00000000",
  40634=>"00000001",
  40635=>"00000000",
  40636=>"00000000",
  40637=>"00000000",
  40638=>"00000000",
  40639=>"00000000",
  40640=>"00000000",
  40641=>"00000000",
  40642=>"00000000",
  40643=>"00000000",
  40644=>"00000000",
  40645=>"00000000",
  40646=>"00000000",
  40647=>"00000000",
  40648=>"00000000",
  40649=>"00000000",
  40650=>"00000000",
  40651=>"00000000",
  40652=>"00000000",
  40653=>"00000000",
  40654=>"00000000",
  40655=>"00000000",
  40656=>"00000000",
  40657=>"00000000",
  40658=>"00000000",
  40659=>"00000000",
  40660=>"00000000",
  40661=>"00000000",
  40662=>"00000000",
  40663=>"00000000",
  40664=>"00000000",
  40665=>"00000000",
  40666=>"00000000",
  40667=>"00000000",
  40668=>"00000000",
  40669=>"11111111",
  40670=>"00000000",
  40671=>"00000000",
  40672=>"00000000",
  40673=>"00000000",
  40674=>"00000000",
  40675=>"00000000",
  40676=>"00000000",
  40677=>"00000000",
  40678=>"00000000",
  40679=>"00000000",
  40680=>"00000000",
  40681=>"00000000",
  40682=>"00000000",
  40683=>"00000000",
  40684=>"00000000",
  40685=>"00000000",
  40686=>"00000000",
  40687=>"00000000",
  40688=>"00000000",
  40689=>"00000000",
  40690=>"00000000",
  40691=>"00000000",
  40692=>"00000000",
  40693=>"00000000",
  40694=>"00000000",
  40695=>"00000000",
  40696=>"00000000",
  40697=>"00000000",
  40698=>"00000000",
  40699=>"00000000",
  40700=>"00000000",
  40701=>"00000000",
  40702=>"00000000",
  40703=>"00000000",
  40704=>"00000000",
  40705=>"00000000",
  40706=>"00000000",
  40707=>"00000000",
  40708=>"00000000",
  40709=>"00000000",
  40710=>"00000000",
  40711=>"00000000",
  40712=>"00000000",
  40713=>"00000000",
  40714=>"00000000",
  40715=>"00000000",
  40716=>"00000000",
  40717=>"00000000",
  40718=>"00000000",
  40719=>"00000000",
  40720=>"00000000",
  40721=>"00000000",
  40722=>"00000000",
  40723=>"00000000",
  40724=>"00000000",
  40725=>"00000000",
  40726=>"00000000",
  40727=>"00000000",
  40728=>"00000000",
  40729=>"00000000",
  40730=>"00000000",
  40731=>"00000000",
  40732=>"00000000",
  40733=>"00000000",
  40734=>"00000000",
  40735=>"00000000",
  40736=>"00000000",
  40737=>"00000000",
  40738=>"00000000",
  40739=>"00000000",
  40740=>"00000000",
  40741=>"00000000",
  40742=>"00000000",
  40743=>"00000000",
  40744=>"00000000",
  40745=>"00000000",
  40746=>"00000000",
  40747=>"00000000",
  40748=>"00000000",
  40749=>"00000000",
  40750=>"00000000",
  40751=>"00000000",
  40752=>"00000000",
  40753=>"00000000",
  40754=>"00000000",
  40755=>"00000000",
  40756=>"00000000",
  40757=>"00000000",
  40758=>"00000000",
  40759=>"00000000",
  40760=>"00000000",
  40761=>"00000000",
  40762=>"00000000",
  40763=>"00000000",
  40764=>"00000000",
  40765=>"00000000",
  40766=>"00000000",
  40767=>"00000000",
  40768=>"00000000",
  40769=>"00000000",
  40770=>"00000000",
  40771=>"00000000",
  40772=>"00000000",
  40773=>"00000000",
  40774=>"00000000",
  40775=>"00000000",
  40776=>"00000000",
  40777=>"00000000",
  40778=>"00000000",
  40779=>"00000000",
  40780=>"00000000",
  40781=>"00000000",
  40782=>"00000000",
  40783=>"00000000",
  40784=>"00000000",
  40785=>"00000000",
  40786=>"00000000",
  40787=>"00000000",
  40788=>"00000000",
  40789=>"00000000",
  40790=>"00000000",
  40791=>"00000000",
  40792=>"00000000",
  40793=>"00000000",
  40794=>"00000000",
  40795=>"00000000",
  40796=>"00000000",
  40797=>"00000000",
  40798=>"00000000",
  40799=>"00000000",
  40800=>"00000000",
  40801=>"00000000",
  40802=>"00000000",
  40803=>"00000000",
  40804=>"00000000",
  40805=>"00000000",
  40806=>"00000000",
  40807=>"00000000",
  40808=>"00000000",
  40809=>"00000000",
  40810=>"00000000",
  40811=>"00000000",
  40812=>"00000000",
  40813=>"00000000",
  40814=>"00000000",
  40815=>"00000000",
  40816=>"00000000",
  40817=>"00000000",
  40818=>"00000001",
  40819=>"00000000",
  40820=>"00000000",
  40821=>"00000000",
  40822=>"00000000",
  40823=>"00000000",
  40824=>"00000000",
  40825=>"00000000",
  40826=>"00000000",
  40827=>"00000000",
  40828=>"00000000",
  40829=>"00000000",
  40830=>"00000000",
  40831=>"00000000",
  40832=>"00000000",
  40833=>"00000000",
  40834=>"00000000",
  40835=>"00000000",
  40836=>"00000000",
  40837=>"00000000",
  40838=>"00000000",
  40839=>"00000000",
  40840=>"00000000",
  40841=>"00000000",
  40842=>"00000001",
  40843=>"00000000",
  40844=>"00000000",
  40845=>"00000000",
  40846=>"00000000",
  40847=>"00000000",
  40848=>"00000000",
  40849=>"00000000",
  40850=>"00000000",
  40851=>"00000000",
  40852=>"00000000",
  40853=>"00000000",
  40854=>"00000000",
  40855=>"00000000",
  40856=>"00000000",
  40857=>"00000000",
  40858=>"00000000",
  40859=>"00000000",
  40860=>"00000000",
  40861=>"00000000",
  40862=>"00000000",
  40863=>"00000000",
  40864=>"00000000",
  40865=>"00000000",
  40866=>"00000000",
  40867=>"00000000",
  40868=>"00000000",
  40869=>"00000000",
  40870=>"00000000",
  40871=>"00000000",
  40872=>"00000000",
  40873=>"00000000",
  40874=>"00000000",
  40875=>"00000000",
  40876=>"00000000",
  40877=>"00000000",
  40878=>"00000000",
  40879=>"00000000",
  40880=>"00000000",
  40881=>"00000000",
  40882=>"00000000",
  40883=>"00000000",
  40884=>"00000000",
  40885=>"00000000",
  40886=>"00000000",
  40887=>"00000000",
  40888=>"00000000",
  40889=>"00000000",
  40890=>"00000000",
  40891=>"00000000",
  40892=>"00000000",
  40893=>"00000000",
  40894=>"00000000",
  40895=>"00000000",
  40896=>"00000000",
  40897=>"00000000",
  40898=>"00000000",
  40899=>"00000000",
  40900=>"00000000",
  40901=>"00000000",
  40902=>"00000000",
  40903=>"11111111",
  40904=>"00000000",
  40905=>"00000000",
  40906=>"00000000",
  40907=>"00000000",
  40908=>"00000000",
  40909=>"00000000",
  40910=>"00000000",
  40911=>"00000000",
  40912=>"00000001",
  40913=>"00000000",
  40914=>"00000000",
  40915=>"00000000",
  40916=>"00000000",
  40917=>"00000000",
  40918=>"00000000",
  40919=>"00000000",
  40920=>"00000000",
  40921=>"00000000",
  40922=>"00000000",
  40923=>"00000000",
  40924=>"00000000",
  40925=>"00000000",
  40926=>"00000000",
  40927=>"00000000",
  40928=>"00000000",
  40929=>"00000000",
  40930=>"00000001",
  40931=>"00000000",
  40932=>"00000000",
  40933=>"00000000",
  40934=>"00000000",
  40935=>"00000000",
  40936=>"00000000",
  40937=>"00000000",
  40938=>"00000000",
  40939=>"00000000",
  40940=>"00000000",
  40941=>"00000000",
  40942=>"00000000",
  40943=>"00000000",
  40944=>"00000000",
  40945=>"00000000",
  40946=>"00000000",
  40947=>"00000000",
  40948=>"00000000",
  40949=>"00000000",
  40950=>"00000000",
  40951=>"00000000",
  40952=>"00000000",
  40953=>"00000000",
  40954=>"00000000",
  40955=>"00000000",
  40956=>"00000000",
  40957=>"00000000",
  40958=>"00000000",
  40959=>"00000000",
  40960=>"00000000",
  40961=>"00000000",
  40962=>"00000000",
  40963=>"00000000",
  40964=>"00000000",
  40965=>"00000000",
  40966=>"00000000",
  40967=>"00000000",
  40968=>"00000000",
  40969=>"00000000",
  40970=>"00000000",
  40971=>"00000000",
  40972=>"00000000",
  40973=>"00000000",
  40974=>"00000000",
  40975=>"00000000",
  40976=>"00000000",
  40977=>"00000000",
  40978=>"00000000",
  40979=>"00000000",
  40980=>"00000000",
  40981=>"00000000",
  40982=>"00000000",
  40983=>"00000001",
  40984=>"00000000",
  40985=>"00000000",
  40986=>"00000000",
  40987=>"00000000",
  40988=>"00000000",
  40989=>"00000000",
  40990=>"00000000",
  40991=>"00000000",
  40992=>"00000000",
  40993=>"00000000",
  40994=>"00000000",
  40995=>"00000000",
  40996=>"00000000",
  40997=>"00000000",
  40998=>"00000000",
  40999=>"00000000",
  41000=>"00000000",
  41001=>"00000000",
  41002=>"00000000",
  41003=>"00000000",
  41004=>"00000000",
  41005=>"00000000",
  41006=>"00000000",
  41007=>"00000000",
  41008=>"00000000",
  41009=>"00000000",
  41010=>"00000000",
  41011=>"00000000",
  41012=>"00000001",
  41013=>"00000000",
  41014=>"00000000",
  41015=>"00000000",
  41016=>"00000000",
  41017=>"00000000",
  41018=>"00000000",
  41019=>"00000000",
  41020=>"00000000",
  41021=>"00000000",
  41022=>"00000000",
  41023=>"00000000",
  41024=>"00000000",
  41025=>"11111111",
  41026=>"00000001",
  41027=>"00000000",
  41028=>"00000000",
  41029=>"00000000",
  41030=>"00000000",
  41031=>"00000001",
  41032=>"00000000",
  41033=>"00000000",
  41034=>"00000000",
  41035=>"00000000",
  41036=>"00000000",
  41037=>"00000000",
  41038=>"00000000",
  41039=>"00000000",
  41040=>"00000000",
  41041=>"00000000",
  41042=>"00000000",
  41043=>"00000000",
  41044=>"00000000",
  41045=>"00000000",
  41046=>"00000000",
  41047=>"00000001",
  41048=>"00000000",
  41049=>"00000000",
  41050=>"00000000",
  41051=>"00000000",
  41052=>"00000000",
  41053=>"00000000",
  41054=>"00000000",
  41055=>"00000000",
  41056=>"00000000",
  41057=>"00000000",
  41058=>"00000000",
  41059=>"00000000",
  41060=>"00000000",
  41061=>"00000000",
  41062=>"00000000",
  41063=>"00000000",
  41064=>"11111111",
  41065=>"00000000",
  41066=>"00000000",
  41067=>"00000000",
  41068=>"00000000",
  41069=>"00000000",
  41070=>"00000000",
  41071=>"00000000",
  41072=>"00000000",
  41073=>"00000000",
  41074=>"00000000",
  41075=>"00000000",
  41076=>"00000000",
  41077=>"00000000",
  41078=>"00000000",
  41079=>"00000000",
  41080=>"00000000",
  41081=>"00000000",
  41082=>"00000000",
  41083=>"00000000",
  41084=>"00000000",
  41085=>"11111111",
  41086=>"00000000",
  41087=>"00000000",
  41088=>"00000000",
  41089=>"00000000",
  41090=>"00000000",
  41091=>"00000000",
  41092=>"00000000",
  41093=>"00000001",
  41094=>"00000000",
  41095=>"11111111",
  41096=>"00000000",
  41097=>"00000000",
  41098=>"00000000",
  41099=>"00000000",
  41100=>"00000000",
  41101=>"00000000",
  41102=>"00000000",
  41103=>"00000000",
  41104=>"00000000",
  41105=>"00000000",
  41106=>"00000000",
  41107=>"00000000",
  41108=>"00000000",
  41109=>"00000000",
  41110=>"00000000",
  41111=>"00000000",
  41112=>"00000000",
  41113=>"00000000",
  41114=>"00000000",
  41115=>"00000000",
  41116=>"11111111",
  41117=>"00000000",
  41118=>"00000000",
  41119=>"00000000",
  41120=>"00000000",
  41121=>"00000000",
  41122=>"00000000",
  41123=>"00000000",
  41124=>"00000000",
  41125=>"00000000",
  41126=>"00000000",
  41127=>"00000000",
  41128=>"00000000",
  41129=>"00000000",
  41130=>"00000000",
  41131=>"00000000",
  41132=>"00000000",
  41133=>"00000000",
  41134=>"00000000",
  41135=>"00000000",
  41136=>"00000000",
  41137=>"00000000",
  41138=>"00000000",
  41139=>"00000000",
  41140=>"00000000",
  41141=>"00000000",
  41142=>"00000000",
  41143=>"00000000",
  41144=>"00000000",
  41145=>"00000000",
  41146=>"00000000",
  41147=>"00000000",
  41148=>"00000000",
  41149=>"11111111",
  41150=>"00000000",
  41151=>"00000000",
  41152=>"00000001",
  41153=>"00000000",
  41154=>"00000000",
  41155=>"00000000",
  41156=>"00000000",
  41157=>"00000000",
  41158=>"00000000",
  41159=>"00000000",
  41160=>"00000000",
  41161=>"00000000",
  41162=>"00000000",
  41163=>"00000000",
  41164=>"00000000",
  41165=>"00000000",
  41166=>"00000000",
  41167=>"00000000",
  41168=>"00000000",
  41169=>"00000000",
  41170=>"00000000",
  41171=>"00000000",
  41172=>"11111111",
  41173=>"00000000",
  41174=>"00000000",
  41175=>"00000000",
  41176=>"00000000",
  41177=>"00000000",
  41178=>"00000000",
  41179=>"00000000",
  41180=>"00000000",
  41181=>"00000000",
  41182=>"00000000",
  41183=>"00000000",
  41184=>"00000000",
  41185=>"00000000",
  41186=>"00000000",
  41187=>"00000000",
  41188=>"00000000",
  41189=>"00000000",
  41190=>"00000000",
  41191=>"00000000",
  41192=>"00000000",
  41193=>"00000000",
  41194=>"00000000",
  41195=>"00000001",
  41196=>"00000000",
  41197=>"00000000",
  41198=>"00000000",
  41199=>"00000010",
  41200=>"00000000",
  41201=>"00000000",
  41202=>"00000000",
  41203=>"00000000",
  41204=>"00000000",
  41205=>"00000000",
  41206=>"00000000",
  41207=>"00000000",
  41208=>"00000000",
  41209=>"00000000",
  41210=>"00000000",
  41211=>"00000000",
  41212=>"00000000",
  41213=>"00000000",
  41214=>"00000000",
  41215=>"11111111",
  41216=>"00000000",
  41217=>"00000000",
  41218=>"00000000",
  41219=>"00000000",
  41220=>"00000000",
  41221=>"00000000",
  41222=>"00000000",
  41223=>"00000000",
  41224=>"00000000",
  41225=>"00000000",
  41226=>"00000000",
  41227=>"11111111",
  41228=>"00000000",
  41229=>"00000000",
  41230=>"00000000",
  41231=>"00000000",
  41232=>"00000000",
  41233=>"11111111",
  41234=>"00000000",
  41235=>"00000000",
  41236=>"00000000",
  41237=>"00000000",
  41238=>"00000000",
  41239=>"00000000",
  41240=>"00000000",
  41241=>"00000000",
  41242=>"00000000",
  41243=>"00000001",
  41244=>"00000000",
  41245=>"00000000",
  41246=>"00000000",
  41247=>"00000000",
  41248=>"00000000",
  41249=>"00000000",
  41250=>"00000000",
  41251=>"00000000",
  41252=>"00000000",
  41253=>"00000000",
  41254=>"00000000",
  41255=>"00000000",
  41256=>"00000000",
  41257=>"00000000",
  41258=>"00000000",
  41259=>"00000000",
  41260=>"00000000",
  41261=>"00000001",
  41262=>"00000000",
  41263=>"00000000",
  41264=>"00000001",
  41265=>"00000001",
  41266=>"00000000",
  41267=>"00000000",
  41268=>"00000000",
  41269=>"00000000",
  41270=>"00000000",
  41271=>"00000001",
  41272=>"00000000",
  41273=>"00000000",
  41274=>"00000000",
  41275=>"00000000",
  41276=>"11111111",
  41277=>"00000000",
  41278=>"00000000",
  41279=>"00000000",
  41280=>"00000001",
  41281=>"00000000",
  41282=>"00000000",
  41283=>"00000001",
  41284=>"00000000",
  41285=>"00000000",
  41286=>"00000000",
  41287=>"00000001",
  41288=>"00000000",
  41289=>"00000000",
  41290=>"00000000",
  41291=>"00000000",
  41292=>"00000000",
  41293=>"00000000",
  41294=>"00000000",
  41295=>"00000000",
  41296=>"00000000",
  41297=>"00000000",
  41298=>"00000000",
  41299=>"00000000",
  41300=>"00000001",
  41301=>"00000000",
  41302=>"00000000",
  41303=>"00000000",
  41304=>"00000000",
  41305=>"00000000",
  41306=>"00000000",
  41307=>"00000000",
  41308=>"00000000",
  41309=>"00000001",
  41310=>"00000000",
  41311=>"00000000",
  41312=>"00000000",
  41313=>"00000000",
  41314=>"00000000",
  41315=>"00000000",
  41316=>"00000000",
  41317=>"00000000",
  41318=>"00000000",
  41319=>"00000000",
  41320=>"00000000",
  41321=>"11111111",
  41322=>"00000000",
  41323=>"00000000",
  41324=>"00000000",
  41325=>"00000000",
  41326=>"00000000",
  41327=>"00000000",
  41328=>"00000000",
  41329=>"00000000",
  41330=>"00000000",
  41331=>"00000000",
  41332=>"00000000",
  41333=>"00000000",
  41334=>"00000000",
  41335=>"00000000",
  41336=>"00000000",
  41337=>"00000000",
  41338=>"00000000",
  41339=>"00000000",
  41340=>"00000000",
  41341=>"00000000",
  41342=>"00000000",
  41343=>"00000000",
  41344=>"00000000",
  41345=>"00000000",
  41346=>"00000000",
  41347=>"00000000",
  41348=>"00000000",
  41349=>"00000000",
  41350=>"00000000",
  41351=>"00000000",
  41352=>"00000000",
  41353=>"00000000",
  41354=>"00000000",
  41355=>"00000000",
  41356=>"00000000",
  41357=>"00000000",
  41358=>"00000000",
  41359=>"00000000",
  41360=>"00000000",
  41361=>"00000000",
  41362=>"00000000",
  41363=>"00000000",
  41364=>"00000000",
  41365=>"00000000",
  41366=>"00000001",
  41367=>"00000000",
  41368=>"00000000",
  41369=>"00000000",
  41370=>"00000000",
  41371=>"00000001",
  41372=>"00000000",
  41373=>"00000000",
  41374=>"00000000",
  41375=>"00000000",
  41376=>"00000000",
  41377=>"00000000",
  41378=>"00000000",
  41379=>"00000000",
  41380=>"00000000",
  41381=>"00000000",
  41382=>"00000000",
  41383=>"00000000",
  41384=>"00000000",
  41385=>"00000000",
  41386=>"00000000",
  41387=>"00000000",
  41388=>"00000000",
  41389=>"00000000",
  41390=>"00000000",
  41391=>"00000000",
  41392=>"00000000",
  41393=>"00000000",
  41394=>"00000000",
  41395=>"00000000",
  41396=>"00000000",
  41397=>"00000000",
  41398=>"00000000",
  41399=>"00000000",
  41400=>"00000000",
  41401=>"00000000",
  41402=>"00000000",
  41403=>"00000000",
  41404=>"00000000",
  41405=>"00000000",
  41406=>"00000000",
  41407=>"00000000",
  41408=>"00000000",
  41409=>"00000000",
  41410=>"00000000",
  41411=>"00000000",
  41412=>"00000000",
  41413=>"00000000",
  41414=>"00000000",
  41415=>"00000000",
  41416=>"00000000",
  41417=>"00000000",
  41418=>"00000000",
  41419=>"00000000",
  41420=>"00000000",
  41421=>"00000000",
  41422=>"00000000",
  41423=>"00000000",
  41424=>"00000000",
  41425=>"00000000",
  41426=>"00000000",
  41427=>"00000000",
  41428=>"00000000",
  41429=>"00000000",
  41430=>"00000000",
  41431=>"00000000",
  41432=>"00000000",
  41433=>"00000000",
  41434=>"00000000",
  41435=>"00000000",
  41436=>"00000000",
  41437=>"00000000",
  41438=>"00000000",
  41439=>"00000000",
  41440=>"00000000",
  41441=>"00000000",
  41442=>"00000000",
  41443=>"11111111",
  41444=>"11111111",
  41445=>"00000000",
  41446=>"00000000",
  41447=>"00000001",
  41448=>"00000000",
  41449=>"00000000",
  41450=>"00000000",
  41451=>"00000000",
  41452=>"00000000",
  41453=>"00000000",
  41454=>"00000000",
  41455=>"00000000",
  41456=>"00000000",
  41457=>"00000000",
  41458=>"00000000",
  41459=>"00000000",
  41460=>"00000000",
  41461=>"00000000",
  41462=>"00000000",
  41463=>"00000000",
  41464=>"00000000",
  41465=>"00000000",
  41466=>"00000000",
  41467=>"00000000",
  41468=>"00000000",
  41469=>"00000000",
  41470=>"00000000",
  41471=>"00000000",
  41472=>"00000000",
  41473=>"00000000",
  41474=>"00000000",
  41475=>"00000000",
  41476=>"00000000",
  41477=>"00000000",
  41478=>"00000000",
  41479=>"00000000",
  41480=>"00000000",
  41481=>"00000000",
  41482=>"11111111",
  41483=>"11111111",
  41484=>"00000000",
  41485=>"00000000",
  41486=>"00000000",
  41487=>"00000000",
  41488=>"00000000",
  41489=>"00000000",
  41490=>"00000000",
  41491=>"00000000",
  41492=>"00000000",
  41493=>"00000000",
  41494=>"00000000",
  41495=>"00000000",
  41496=>"00000000",
  41497=>"00000000",
  41498=>"11111111",
  41499=>"00000000",
  41500=>"11111111",
  41501=>"00000000",
  41502=>"00000000",
  41503=>"00000000",
  41504=>"00000000",
  41505=>"00000000",
  41506=>"00000000",
  41507=>"00000000",
  41508=>"00000000",
  41509=>"00000000",
  41510=>"00000000",
  41511=>"00000000",
  41512=>"00000000",
  41513=>"00000000",
  41514=>"00000000",
  41515=>"00000000",
  41516=>"00000000",
  41517=>"00000000",
  41518=>"11111111",
  41519=>"00000000",
  41520=>"00000000",
  41521=>"11111111",
  41522=>"00000000",
  41523=>"11111111",
  41524=>"00000000",
  41525=>"00000000",
  41526=>"00000000",
  41527=>"00000000",
  41528=>"00000000",
  41529=>"00000000",
  41530=>"00000000",
  41531=>"00000001",
  41532=>"00000000",
  41533=>"00000000",
  41534=>"11111111",
  41535=>"00000000",
  41536=>"00000000",
  41537=>"11111111",
  41538=>"00000000",
  41539=>"00000001",
  41540=>"00000000",
  41541=>"00000000",
  41542=>"00000000",
  41543=>"00000000",
  41544=>"00000001",
  41545=>"00000000",
  41546=>"11111111",
  41547=>"00000000",
  41548=>"00000000",
  41549=>"00000000",
  41550=>"00000000",
  41551=>"00000001",
  41552=>"00000000",
  41553=>"00000000",
  41554=>"00000000",
  41555=>"00000000",
  41556=>"00000000",
  41557=>"00000000",
  41558=>"00000000",
  41559=>"00000001",
  41560=>"00000000",
  41561=>"00000000",
  41562=>"11111111",
  41563=>"00000000",
  41564=>"00000000",
  41565=>"00000000",
  41566=>"00000000",
  41567=>"00000000",
  41568=>"00000000",
  41569=>"00000000",
  41570=>"00000000",
  41571=>"00000000",
  41572=>"00000000",
  41573=>"00000000",
  41574=>"00000001",
  41575=>"00000000",
  41576=>"00000000",
  41577=>"00000000",
  41578=>"00000000",
  41579=>"00000000",
  41580=>"00000000",
  41581=>"00000000",
  41582=>"00000000",
  41583=>"00000000",
  41584=>"00000000",
  41585=>"00000000",
  41586=>"00000000",
  41587=>"11111111",
  41588=>"00000000",
  41589=>"00000000",
  41590=>"00000000",
  41591=>"00000000",
  41592=>"00000000",
  41593=>"00000000",
  41594=>"00000000",
  41595=>"00000000",
  41596=>"00000000",
  41597=>"00000000",
  41598=>"00000000",
  41599=>"00000000",
  41600=>"00000000",
  41601=>"00000000",
  41602=>"00000000",
  41603=>"00000000",
  41604=>"00000000",
  41605=>"00000000",
  41606=>"00000000",
  41607=>"00000000",
  41608=>"00000000",
  41609=>"00000000",
  41610=>"00000000",
  41611=>"00000000",
  41612=>"00000000",
  41613=>"00000000",
  41614=>"00000000",
  41615=>"00000000",
  41616=>"00000000",
  41617=>"00000000",
  41618=>"00000000",
  41619=>"00000000",
  41620=>"00000000",
  41621=>"00000000",
  41622=>"00000000",
  41623=>"00000000",
  41624=>"00000000",
  41625=>"00000000",
  41626=>"00000000",
  41627=>"00000000",
  41628=>"00000000",
  41629=>"00000000",
  41630=>"00000000",
  41631=>"00000000",
  41632=>"00000001",
  41633=>"00000000",
  41634=>"00000000",
  41635=>"00000000",
  41636=>"00000000",
  41637=>"00000000",
  41638=>"00000000",
  41639=>"00000000",
  41640=>"00000000",
  41641=>"00000000",
  41642=>"00000000",
  41643=>"00000001",
  41644=>"00000000",
  41645=>"00000000",
  41646=>"00000000",
  41647=>"00000000",
  41648=>"00000000",
  41649=>"00000000",
  41650=>"00000000",
  41651=>"00000000",
  41652=>"00000001",
  41653=>"00000000",
  41654=>"00000000",
  41655=>"00000000",
  41656=>"00000000",
  41657=>"00000000",
  41658=>"00000001",
  41659=>"00000000",
  41660=>"00000000",
  41661=>"00000001",
  41662=>"00000000",
  41663=>"00000000",
  41664=>"00000000",
  41665=>"00000000",
  41666=>"00000000",
  41667=>"00000000",
  41668=>"00000000",
  41669=>"00000000",
  41670=>"00000000",
  41671=>"00000000",
  41672=>"00000000",
  41673=>"00000000",
  41674=>"00000000",
  41675=>"00000000",
  41676=>"00000000",
  41677=>"00000000",
  41678=>"00000000",
  41679=>"00000000",
  41680=>"00000000",
  41681=>"00000000",
  41682=>"00000000",
  41683=>"00000000",
  41684=>"00000000",
  41685=>"00000000",
  41686=>"11111111",
  41687=>"00000000",
  41688=>"00000000",
  41689=>"00000000",
  41690=>"11111111",
  41691=>"00000000",
  41692=>"00000000",
  41693=>"00000001",
  41694=>"00000000",
  41695=>"00000000",
  41696=>"00000000",
  41697=>"00000000",
  41698=>"00000000",
  41699=>"00000000",
  41700=>"00000000",
  41701=>"00000000",
  41702=>"00000000",
  41703=>"00000000",
  41704=>"00000000",
  41705=>"00000000",
  41706=>"00000000",
  41707=>"00000000",
  41708=>"00000000",
  41709=>"00000000",
  41710=>"00000000",
  41711=>"00000000",
  41712=>"00000000",
  41713=>"00000000",
  41714=>"00000000",
  41715=>"00000000",
  41716=>"00000000",
  41717=>"00000000",
  41718=>"00000000",
  41719=>"00000000",
  41720=>"00000000",
  41721=>"00000000",
  41722=>"00000000",
  41723=>"00000000",
  41724=>"00000000",
  41725=>"00000000",
  41726=>"00000000",
  41727=>"00000000",
  41728=>"00000000",
  41729=>"00000000",
  41730=>"00000000",
  41731=>"00000000",
  41732=>"00000000",
  41733=>"00000000",
  41734=>"00000000",
  41735=>"00000000",
  41736=>"00000000",
  41737=>"00000000",
  41738=>"00000000",
  41739=>"00000000",
  41740=>"00000000",
  41741=>"00000000",
  41742=>"00000000",
  41743=>"00000001",
  41744=>"00000000",
  41745=>"00000000",
  41746=>"00000000",
  41747=>"00000000",
  41748=>"00000000",
  41749=>"00000000",
  41750=>"00000000",
  41751=>"00000000",
  41752=>"00000000",
  41753=>"00000000",
  41754=>"00000000",
  41755=>"00000000",
  41756=>"00000000",
  41757=>"00000000",
  41758=>"00000000",
  41759=>"00000000",
  41760=>"00000000",
  41761=>"00000000",
  41762=>"00000001",
  41763=>"11111111",
  41764=>"00000000",
  41765=>"00000000",
  41766=>"00000000",
  41767=>"00000000",
  41768=>"00000000",
  41769=>"00000000",
  41770=>"00000000",
  41771=>"00000000",
  41772=>"00000000",
  41773=>"00000000",
  41774=>"00000000",
  41775=>"00000000",
  41776=>"00000000",
  41777=>"00000000",
  41778=>"00000000",
  41779=>"00000000",
  41780=>"00000000",
  41781=>"00000000",
  41782=>"00000000",
  41783=>"00000000",
  41784=>"11111111",
  41785=>"00000000",
  41786=>"11111111",
  41787=>"00000000",
  41788=>"00000000",
  41789=>"00000000",
  41790=>"00000001",
  41791=>"00000000",
  41792=>"00000000",
  41793=>"00000000",
  41794=>"00000000",
  41795=>"00000000",
  41796=>"00000000",
  41797=>"00000000",
  41798=>"00000000",
  41799=>"00000000",
  41800=>"00000000",
  41801=>"00000000",
  41802=>"00000000",
  41803=>"00000000",
  41804=>"00000000",
  41805=>"00000001",
  41806=>"00000000",
  41807=>"00000000",
  41808=>"00000000",
  41809=>"00000000",
  41810=>"00000000",
  41811=>"00000000",
  41812=>"00000000",
  41813=>"00000000",
  41814=>"11111111",
  41815=>"00000000",
  41816=>"00000000",
  41817=>"00000000",
  41818=>"00000000",
  41819=>"00000000",
  41820=>"00000000",
  41821=>"00000000",
  41822=>"00000000",
  41823=>"00000000",
  41824=>"00000000",
  41825=>"00000000",
  41826=>"00000000",
  41827=>"00000000",
  41828=>"00000000",
  41829=>"00000000",
  41830=>"00000001",
  41831=>"00000000",
  41832=>"00000000",
  41833=>"00000000",
  41834=>"00000000",
  41835=>"00000000",
  41836=>"00000000",
  41837=>"00000000",
  41838=>"00000000",
  41839=>"00000000",
  41840=>"00000000",
  41841=>"00000000",
  41842=>"00000000",
  41843=>"00000000",
  41844=>"00000001",
  41845=>"00000000",
  41846=>"00000000",
  41847=>"00000000",
  41848=>"00000000",
  41849=>"00000000",
  41850=>"00000000",
  41851=>"00000000",
  41852=>"00000000",
  41853=>"00000000",
  41854=>"00000000",
  41855=>"00000000",
  41856=>"00000001",
  41857=>"00000000",
  41858=>"00000001",
  41859=>"00000000",
  41860=>"00000000",
  41861=>"00000001",
  41862=>"00000000",
  41863=>"00000000",
  41864=>"00000000",
  41865=>"00000000",
  41866=>"00000000",
  41867=>"11111111",
  41868=>"00000000",
  41869=>"11111111",
  41870=>"00000000",
  41871=>"00000000",
  41872=>"00000000",
  41873=>"00000000",
  41874=>"00000000",
  41875=>"00000001",
  41876=>"00000000",
  41877=>"00000000",
  41878=>"11111111",
  41879=>"00000000",
  41880=>"00000000",
  41881=>"00000000",
  41882=>"00000000",
  41883=>"00000000",
  41884=>"00000000",
  41885=>"00000000",
  41886=>"00000000",
  41887=>"00000000",
  41888=>"00000000",
  41889=>"00000000",
  41890=>"00000000",
  41891=>"00000000",
  41892=>"11111111",
  41893=>"00000000",
  41894=>"00000000",
  41895=>"00000000",
  41896=>"00000000",
  41897=>"00000001",
  41898=>"00000001",
  41899=>"00000000",
  41900=>"00000000",
  41901=>"00000000",
  41902=>"00000000",
  41903=>"00000000",
  41904=>"11111111",
  41905=>"00000000",
  41906=>"00000000",
  41907=>"00000000",
  41908=>"00000000",
  41909=>"00000000",
  41910=>"00000000",
  41911=>"00000000",
  41912=>"00000000",
  41913=>"00000000",
  41914=>"00000000",
  41915=>"00000000",
  41916=>"00000000",
  41917=>"00000000",
  41918=>"00000000",
  41919=>"00000000",
  41920=>"00000000",
  41921=>"00000000",
  41922=>"00000000",
  41923=>"00000001",
  41924=>"00000000",
  41925=>"00000001",
  41926=>"00000000",
  41927=>"00000001",
  41928=>"00000000",
  41929=>"00000000",
  41930=>"00000000",
  41931=>"00000000",
  41932=>"00000000",
  41933=>"00000000",
  41934=>"00000000",
  41935=>"00000000",
  41936=>"11111111",
  41937=>"00000000",
  41938=>"00000000",
  41939=>"00000000",
  41940=>"11111111",
  41941=>"00000000",
  41942=>"00000000",
  41943=>"00000000",
  41944=>"00000001",
  41945=>"00000000",
  41946=>"00000000",
  41947=>"00000000",
  41948=>"00000000",
  41949=>"11111111",
  41950=>"00000000",
  41951=>"00000000",
  41952=>"00000000",
  41953=>"00000000",
  41954=>"00000000",
  41955=>"00000000",
  41956=>"00000001",
  41957=>"00000000",
  41958=>"00000000",
  41959=>"00000000",
  41960=>"00000000",
  41961=>"00000000",
  41962=>"11111111",
  41963=>"00000000",
  41964=>"00000000",
  41965=>"00000000",
  41966=>"00000000",
  41967=>"00000000",
  41968=>"00000000",
  41969=>"00000001",
  41970=>"00000000",
  41971=>"00000001",
  41972=>"00000000",
  41973=>"11111111",
  41974=>"00000000",
  41975=>"00000000",
  41976=>"00000000",
  41977=>"00000000",
  41978=>"00000000",
  41979=>"00000000",
  41980=>"00000000",
  41981=>"00000000",
  41982=>"00000000",
  41983=>"00000000",
  41984=>"11111001",
  41985=>"00000000",
  41986=>"00000000",
  41987=>"11111111",
  41988=>"00000011",
  41989=>"00000001",
  41990=>"11111010",
  41991=>"11111010",
  41992=>"11111111",
  41993=>"00000000",
  41994=>"11111101",
  41995=>"11111101",
  41996=>"00000011",
  41997=>"11111101",
  41998=>"11111110",
  41999=>"00000010",
  42000=>"00000010",
  42001=>"00000001",
  42002=>"00000001",
  42003=>"00000010",
  42004=>"00000011",
  42005=>"11111111",
  42006=>"11111111",
  42007=>"00000001",
  42008=>"11111110",
  42009=>"11111110",
  42010=>"00000011",
  42011=>"11111110",
  42012=>"00000000",
  42013=>"11111110",
  42014=>"00000001",
  42015=>"11111100",
  42016=>"00000010",
  42017=>"00000001",
  42018=>"00000000",
  42019=>"00000000",
  42020=>"11111011",
  42021=>"00000010",
  42022=>"00000010",
  42023=>"00000000",
  42024=>"00000011",
  42025=>"11111101",
  42026=>"00000010",
  42027=>"11111100",
  42028=>"11111100",
  42029=>"11110100",
  42030=>"11111011",
  42031=>"11111101",
  42032=>"11111110",
  42033=>"00000001",
  42034=>"00000010",
  42035=>"00000011",
  42036=>"11110111",
  42037=>"11111111",
  42038=>"11111010",
  42039=>"11111101",
  42040=>"00000100",
  42041=>"00000000",
  42042=>"00000000",
  42043=>"00000001",
  42044=>"11111111",
  42045=>"11111101",
  42046=>"00000010",
  42047=>"11111110",
  42048=>"11111111",
  42049=>"00000010",
  42050=>"00000100",
  42051=>"11111011",
  42052=>"11111110",
  42053=>"11111111",
  42054=>"00000010",
  42055=>"00000010",
  42056=>"00000011",
  42057=>"00000000",
  42058=>"11111101",
  42059=>"00000010",
  42060=>"00000010",
  42061=>"11111111",
  42062=>"11111010",
  42063=>"11111110",
  42064=>"11111100",
  42065=>"11111010",
  42066=>"00000000",
  42067=>"00000010",
  42068=>"00000001",
  42069=>"11111101",
  42070=>"00000010",
  42071=>"11111100",
  42072=>"11111110",
  42073=>"11111111",
  42074=>"11111110",
  42075=>"00000001",
  42076=>"11111100",
  42077=>"11111100",
  42078=>"00000001",
  42079=>"00000100",
  42080=>"00000000",
  42081=>"00000010",
  42082=>"00000010",
  42083=>"11111111",
  42084=>"11111110",
  42085=>"00000100",
  42086=>"11111101",
  42087=>"11111110",
  42088=>"11111110",
  42089=>"00000010",
  42090=>"11111011",
  42091=>"11111110",
  42092=>"00000011",
  42093=>"11111101",
  42094=>"00000001",
  42095=>"11111010",
  42096=>"00000000",
  42097=>"11111101",
  42098=>"11111101",
  42099=>"00000100",
  42100=>"11111010",
  42101=>"11111110",
  42102=>"11111110",
  42103=>"00000001",
  42104=>"00000010",
  42105=>"11111101",
  42106=>"11111110",
  42107=>"11111110",
  42108=>"00000000",
  42109=>"11111001",
  42110=>"11111111",
  42111=>"11111110",
  42112=>"00000011",
  42113=>"11111110",
  42114=>"00000000",
  42115=>"11111011",
  42116=>"11111100",
  42117=>"11111110",
  42118=>"11111011",
  42119=>"00000001",
  42120=>"00000010",
  42121=>"00000001",
  42122=>"00000010",
  42123=>"00000000",
  42124=>"11111110",
  42125=>"11111100",
  42126=>"00000010",
  42127=>"00000001",
  42128=>"11111100",
  42129=>"00000011",
  42130=>"11111100",
  42131=>"00000000",
  42132=>"11111110",
  42133=>"00000010",
  42134=>"11111110",
  42135=>"00000001",
  42136=>"11111101",
  42137=>"00000001",
  42138=>"00000011",
  42139=>"11111111",
  42140=>"11111101",
  42141=>"11111111",
  42142=>"11111010",
  42143=>"00000000",
  42144=>"11111011",
  42145=>"00000001",
  42146=>"11111011",
  42147=>"11111111",
  42148=>"11111110",
  42149=>"00000010",
  42150=>"00000010",
  42151=>"00000010",
  42152=>"00000000",
  42153=>"11111101",
  42154=>"11111010",
  42155=>"11111110",
  42156=>"11111100",
  42157=>"11111110",
  42158=>"00000000",
  42159=>"11111011",
  42160=>"00000001",
  42161=>"00000011",
  42162=>"00000001",
  42163=>"00000011",
  42164=>"00000001",
  42165=>"11111110",
  42166=>"00000010",
  42167=>"00000001",
  42168=>"00000011",
  42169=>"11111100",
  42170=>"11111110",
  42171=>"00000010",
  42172=>"11111110",
  42173=>"11111011",
  42174=>"11111011",
  42175=>"00000001",
  42176=>"11111111",
  42177=>"11111011",
  42178=>"11111111",
  42179=>"11111100",
  42180=>"11111010",
  42181=>"00000001",
  42182=>"00000010",
  42183=>"11111111",
  42184=>"00000010",
  42185=>"00000010",
  42186=>"11111010",
  42187=>"11111011",
  42188=>"00000001",
  42189=>"11111011",
  42190=>"11111010",
  42191=>"11111111",
  42192=>"11111100",
  42193=>"11111111",
  42194=>"11111010",
  42195=>"00000010",
  42196=>"11111010",
  42197=>"00000000",
  42198=>"00000000",
  42199=>"11111111",
  42200=>"11111111",
  42201=>"11111110",
  42202=>"11111101",
  42203=>"00000000",
  42204=>"00000010",
  42205=>"11111111",
  42206=>"00000000",
  42207=>"00000010",
  42208=>"00000001",
  42209=>"11111110",
  42210=>"11111100",
  42211=>"00000010",
  42212=>"11111101",
  42213=>"00000010",
  42214=>"00000000",
  42215=>"00000000",
  42216=>"11111011",
  42217=>"00000010",
  42218=>"00000011",
  42219=>"11111001",
  42220=>"11110110",
  42221=>"00000100",
  42222=>"11111101",
  42223=>"11111011",
  42224=>"00000001",
  42225=>"00000001",
  42226=>"00000100",
  42227=>"11111011",
  42228=>"11111110",
  42229=>"11111110",
  42230=>"00000000",
  42231=>"00000001",
  42232=>"00000000",
  42233=>"11111101",
  42234=>"00000000",
  42235=>"11111101",
  42236=>"00000101",
  42237=>"11111100",
  42238=>"00000010",
  42239=>"11111111",
  42240=>"00000000",
  42241=>"00000001",
  42242=>"00000000",
  42243=>"11111100",
  42244=>"11111011",
  42245=>"11111111",
  42246=>"00000011",
  42247=>"00000010",
  42248=>"11111110",
  42249=>"00000110",
  42250=>"00000001",
  42251=>"11111110",
  42252=>"00000000",
  42253=>"11111100",
  42254=>"11111101",
  42255=>"11111111",
  42256=>"00000000",
  42257=>"11111111",
  42258=>"00000010",
  42259=>"00000010",
  42260=>"00000011",
  42261=>"11111001",
  42262=>"11111100",
  42263=>"00000001",
  42264=>"00000010",
  42265=>"11111011",
  42266=>"11111100",
  42267=>"11111101",
  42268=>"00000100",
  42269=>"11111110",
  42270=>"11111110",
  42271=>"00000011",
  42272=>"00000000",
  42273=>"00000000",
  42274=>"00000010",
  42275=>"11111101",
  42276=>"00000001",
  42277=>"00000011",
  42278=>"11111110",
  42279=>"11111101",
  42280=>"11111111",
  42281=>"11111100",
  42282=>"11111110",
  42283=>"11111101",
  42284=>"11111101",
  42285=>"11111010",
  42286=>"00000001",
  42287=>"11111110",
  42288=>"11111111",
  42289=>"00000001",
  42290=>"00000010",
  42291=>"11111110",
  42292=>"00000000",
  42293=>"11111110",
  42294=>"11111111",
  42295=>"11111110",
  42296=>"00000000",
  42297=>"00000000",
  42298=>"11110111",
  42299=>"00000001",
  42300=>"11111100",
  42301=>"11111100",
  42302=>"00000000",
  42303=>"11111001",
  42304=>"11111001",
  42305=>"00000000",
  42306=>"00000000",
  42307=>"11111110",
  42308=>"11111001",
  42309=>"11111111",
  42310=>"00000100",
  42311=>"00000001",
  42312=>"00000000",
  42313=>"11111100",
  42314=>"11111110",
  42315=>"11111010",
  42316=>"11111111",
  42317=>"11111011",
  42318=>"11111011",
  42319=>"00000001",
  42320=>"11111111",
  42321=>"11111101",
  42322=>"00000001",
  42323=>"00000011",
  42324=>"00000001",
  42325=>"11111001",
  42326=>"11111100",
  42327=>"11111110",
  42328=>"00000001",
  42329=>"11111001",
  42330=>"11111111",
  42331=>"11111110",
  42332=>"11111111",
  42333=>"00000010",
  42334=>"11111101",
  42335=>"00000001",
  42336=>"11111110",
  42337=>"11111111",
  42338=>"00000001",
  42339=>"00000001",
  42340=>"11111101",
  42341=>"11111010",
  42342=>"00000010",
  42343=>"11111000",
  42344=>"11111010",
  42345=>"11111111",
  42346=>"11111001",
  42347=>"00000000",
  42348=>"00000001",
  42349=>"11111011",
  42350=>"00000000",
  42351=>"11111100",
  42352=>"11111110",
  42353=>"11111101",
  42354=>"00000001",
  42355=>"11111100",
  42356=>"11111101",
  42357=>"00000100",
  42358=>"00000000",
  42359=>"11111100",
  42360=>"11111101",
  42361=>"00000000",
  42362=>"11111111",
  42363=>"11111111",
  42364=>"11111110",
  42365=>"00000001",
  42366=>"11111100",
  42367=>"00000010",
  42368=>"00000010",
  42369=>"00000001",
  42370=>"11111111",
  42371=>"11111100",
  42372=>"00000011",
  42373=>"00000001",
  42374=>"11111101",
  42375=>"11111001",
  42376=>"11111001",
  42377=>"00000001",
  42378=>"00000010",
  42379=>"11110111",
  42380=>"11111110",
  42381=>"11111011",
  42382=>"00000000",
  42383=>"11111110",
  42384=>"11111011",
  42385=>"00000010",
  42386=>"00000000",
  42387=>"00000000",
  42388=>"11111111",
  42389=>"00000001",
  42390=>"00000000",
  42391=>"11111111",
  42392=>"11111111",
  42393=>"00000010",
  42394=>"11111100",
  42395=>"11111011",
  42396=>"11111010",
  42397=>"00000010",
  42398=>"11111010",
  42399=>"00000001",
  42400=>"11111111",
  42401=>"11111100",
  42402=>"11111110",
  42403=>"00000001",
  42404=>"11110101",
  42405=>"11111111",
  42406=>"00000010",
  42407=>"11111101",
  42408=>"11111101",
  42409=>"11111111",
  42410=>"00000011",
  42411=>"00000011",
  42412=>"11111111",
  42413=>"11111101",
  42414=>"11111110",
  42415=>"11111101",
  42416=>"00000100",
  42417=>"00000000",
  42418=>"11111110",
  42419=>"11111100",
  42420=>"00000000",
  42421=>"00000011",
  42422=>"11111110",
  42423=>"11111101",
  42424=>"00000000",
  42425=>"11111110",
  42426=>"11111110",
  42427=>"11111101",
  42428=>"11111100",
  42429=>"00000010",
  42430=>"11111101",
  42431=>"11111100",
  42432=>"00000000",
  42433=>"00000001",
  42434=>"00000000",
  42435=>"00000011",
  42436=>"11111101",
  42437=>"11111111",
  42438=>"11111000",
  42439=>"11111111",
  42440=>"11111110",
  42441=>"11111111",
  42442=>"00000000",
  42443=>"11111010",
  42444=>"11111001",
  42445=>"11111100",
  42446=>"11111101",
  42447=>"11111110",
  42448=>"11111010",
  42449=>"11111110",
  42450=>"00000001",
  42451=>"00000000",
  42452=>"11111001",
  42453=>"00000001",
  42454=>"11111111",
  42455=>"00000001",
  42456=>"11111001",
  42457=>"11111110",
  42458=>"11110111",
  42459=>"00000011",
  42460=>"11111110",
  42461=>"00000010",
  42462=>"11111100",
  42463=>"00000000",
  42464=>"00000000",
  42465=>"11111110",
  42466=>"11111100",
  42467=>"11111011",
  42468=>"11111001",
  42469=>"11111101",
  42470=>"11111010",
  42471=>"11111100",
  42472=>"11111101",
  42473=>"11111111",
  42474=>"11111100",
  42475=>"00000000",
  42476=>"00000011",
  42477=>"00000001",
  42478=>"11111111",
  42479=>"00000100",
  42480=>"11111001",
  42481=>"11111111",
  42482=>"11111101",
  42483=>"11111101",
  42484=>"00000000",
  42485=>"11111110",
  42486=>"00000010",
  42487=>"00000001",
  42488=>"11111111",
  42489=>"00000001",
  42490=>"11111111",
  42491=>"00000000",
  42492=>"11111011",
  42493=>"11111111",
  42494=>"11111111",
  42495=>"00000000",
  42496=>"11111010",
  42497=>"00000010",
  42498=>"00000011",
  42499=>"11111111",
  42500=>"00000000",
  42501=>"11111011",
  42502=>"00000001",
  42503=>"00000001",
  42504=>"11111111",
  42505=>"11111101",
  42506=>"11111010",
  42507=>"11111001",
  42508=>"00000010",
  42509=>"00000001",
  42510=>"11111111",
  42511=>"00000011",
  42512=>"11111110",
  42513=>"00000001",
  42514=>"11111100",
  42515=>"11111111",
  42516=>"00000000",
  42517=>"11111100",
  42518=>"11111110",
  42519=>"00000001",
  42520=>"11111110",
  42521=>"00000000",
  42522=>"11111101",
  42523=>"11111011",
  42524=>"11111011",
  42525=>"00000010",
  42526=>"11111001",
  42527=>"00000000",
  42528=>"00000100",
  42529=>"11111001",
  42530=>"00000001",
  42531=>"00000010",
  42532=>"11111100",
  42533=>"00000001",
  42534=>"11111100",
  42535=>"11111111",
  42536=>"00000000",
  42537=>"00000001",
  42538=>"00000000",
  42539=>"11111101",
  42540=>"11111110",
  42541=>"00000000",
  42542=>"11111110",
  42543=>"11111100",
  42544=>"00000001",
  42545=>"00000001",
  42546=>"11111011",
  42547=>"11111010",
  42548=>"00000010",
  42549=>"00000000",
  42550=>"00000000",
  42551=>"11111100",
  42552=>"00000000",
  42553=>"11111010",
  42554=>"11111010",
  42555=>"11111111",
  42556=>"11111011",
  42557=>"11111111",
  42558=>"11111010",
  42559=>"11111000",
  42560=>"11111111",
  42561=>"11111111",
  42562=>"11111111",
  42563=>"11111110",
  42564=>"11111101",
  42565=>"11111111",
  42566=>"00000100",
  42567=>"00000001",
  42568=>"00000010",
  42569=>"11111010",
  42570=>"00000010",
  42571=>"11111110",
  42572=>"11111101",
  42573=>"11111100",
  42574=>"11111111",
  42575=>"11111110",
  42576=>"11111100",
  42577=>"00000001",
  42578=>"11111010",
  42579=>"11111010",
  42580=>"11111101",
  42581=>"00000001",
  42582=>"00000010",
  42583=>"11111101",
  42584=>"11111110",
  42585=>"00000010",
  42586=>"11111011",
  42587=>"00000001",
  42588=>"11111111",
  42589=>"11111101",
  42590=>"00000000",
  42591=>"11111111",
  42592=>"00000000",
  42593=>"00000000",
  42594=>"00000110",
  42595=>"00000010",
  42596=>"00000000",
  42597=>"00000010",
  42598=>"11111011",
  42599=>"00000001",
  42600=>"11111101",
  42601=>"00000000",
  42602=>"11111100",
  42603=>"11111110",
  42604=>"00000000",
  42605=>"11111010",
  42606=>"11111110",
  42607=>"00000001",
  42608=>"00000011",
  42609=>"00000000",
  42610=>"00000010",
  42611=>"11111110",
  42612=>"11111000",
  42613=>"00000000",
  42614=>"00000010",
  42615=>"11111111",
  42616=>"11111111",
  42617=>"11111000",
  42618=>"00000011",
  42619=>"00000011",
  42620=>"11111001",
  42621=>"11111100",
  42622=>"00000010",
  42623=>"11111011",
  42624=>"11111101",
  42625=>"11111010",
  42626=>"00000000",
  42627=>"00000101",
  42628=>"00000110",
  42629=>"00000000",
  42630=>"11111111",
  42631=>"11111010",
  42632=>"00000001",
  42633=>"00000011",
  42634=>"11111110",
  42635=>"00000000",
  42636=>"11111000",
  42637=>"00000000",
  42638=>"00000100",
  42639=>"11111101",
  42640=>"11111011",
  42641=>"00000001",
  42642=>"00000001",
  42643=>"11111010",
  42644=>"11111111",
  42645=>"00000001",
  42646=>"00000010",
  42647=>"00000010",
  42648=>"00000010",
  42649=>"00000001",
  42650=>"00000001",
  42651=>"00000001",
  42652=>"00000110",
  42653=>"00000000",
  42654=>"11111100",
  42655=>"11111100",
  42656=>"11111011",
  42657=>"11111010",
  42658=>"11111111",
  42659=>"11111111",
  42660=>"00000000",
  42661=>"00000000",
  42662=>"11111001",
  42663=>"11111111",
  42664=>"11111111",
  42665=>"00000010",
  42666=>"11111100",
  42667=>"11111100",
  42668=>"11111101",
  42669=>"11111101",
  42670=>"11110110",
  42671=>"11111111",
  42672=>"00000000",
  42673=>"11111101",
  42674=>"00000000",
  42675=>"11111001",
  42676=>"00000010",
  42677=>"00000011",
  42678=>"00000001",
  42679=>"11111011",
  42680=>"11111101",
  42681=>"00000000",
  42682=>"11111100",
  42683=>"11111011",
  42684=>"00000010",
  42685=>"11111111",
  42686=>"00000000",
  42687=>"11111011",
  42688=>"11111011",
  42689=>"11111110",
  42690=>"00000000",
  42691=>"11111010",
  42692=>"11111101",
  42693=>"00000001",
  42694=>"00000000",
  42695=>"00000011",
  42696=>"00000011",
  42697=>"00000000",
  42698=>"11111111",
  42699=>"11111111",
  42700=>"00000001",
  42701=>"00000010",
  42702=>"11111111",
  42703=>"11111101",
  42704=>"11111000",
  42705=>"00000000",
  42706=>"11111111",
  42707=>"00000010",
  42708=>"00000000",
  42709=>"00000000",
  42710=>"11111011",
  42711=>"00000000",
  42712=>"11111111",
  42713=>"00000000",
  42714=>"11111101",
  42715=>"11111011",
  42716=>"11111110",
  42717=>"11111101",
  42718=>"11111100",
  42719=>"00000000",
  42720=>"00000001",
  42721=>"11111010",
  42722=>"00000010",
  42723=>"00000001",
  42724=>"11111111",
  42725=>"11111010",
  42726=>"00000000",
  42727=>"00000000",
  42728=>"11111100",
  42729=>"00000000",
  42730=>"00000001",
  42731=>"11111111",
  42732=>"00000001",
  42733=>"00000100",
  42734=>"00000000",
  42735=>"00000010",
  42736=>"00000001",
  42737=>"11111111",
  42738=>"11111101",
  42739=>"11111000",
  42740=>"00000011",
  42741=>"00000010",
  42742=>"11111111",
  42743=>"11111110",
  42744=>"00000001",
  42745=>"11111110",
  42746=>"11111011",
  42747=>"00000000",
  42748=>"11111010",
  42749=>"00000001",
  42750=>"11111011",
  42751=>"00000001",
  42752=>"00000010",
  42753=>"00000010",
  42754=>"11111111",
  42755=>"00000000",
  42756=>"11111101",
  42757=>"11111011",
  42758=>"11111111",
  42759=>"11111011",
  42760=>"11111100",
  42761=>"11111111",
  42762=>"11111110",
  42763=>"00000110",
  42764=>"11111111",
  42765=>"11111110",
  42766=>"00000011",
  42767=>"11111111",
  42768=>"00000000",
  42769=>"00000001",
  42770=>"11111101",
  42771=>"00000000",
  42772=>"00000000",
  42773=>"00000000",
  42774=>"11111111",
  42775=>"11111101",
  42776=>"00000101",
  42777=>"00000010",
  42778=>"00000001",
  42779=>"00000011",
  42780=>"11111111",
  42781=>"00000010",
  42782=>"00000011",
  42783=>"11111011",
  42784=>"00000000",
  42785=>"11111111",
  42786=>"11111101",
  42787=>"11111100",
  42788=>"11111111",
  42789=>"00000000",
  42790=>"00000010",
  42791=>"00000001",
  42792=>"11111101",
  42793=>"00000000",
  42794=>"00000001",
  42795=>"11111011",
  42796=>"00000001",
  42797=>"11111111",
  42798=>"11111110",
  42799=>"11111100",
  42800=>"00000001",
  42801=>"00000001",
  42802=>"00000000",
  42803=>"00000101",
  42804=>"11111000",
  42805=>"00000001",
  42806=>"11111100",
  42807=>"11111111",
  42808=>"00000001",
  42809=>"11111000",
  42810=>"11111000",
  42811=>"00000000",
  42812=>"00000000",
  42813=>"11111011",
  42814=>"00000000",
  42815=>"11111101",
  42816=>"00000001",
  42817=>"00000010",
  42818=>"11111110",
  42819=>"11111101",
  42820=>"11111110",
  42821=>"11111011",
  42822=>"00000010",
  42823=>"00000100",
  42824=>"00000001",
  42825=>"11111010",
  42826=>"11111011",
  42827=>"11111111",
  42828=>"11111010",
  42829=>"11111110",
  42830=>"00000001",
  42831=>"00000000",
  42832=>"00000010",
  42833=>"11111101",
  42834=>"11111111",
  42835=>"00000100",
  42836=>"11111010",
  42837=>"11111111",
  42838=>"11111011",
  42839=>"00000001",
  42840=>"00000001",
  42841=>"11111011",
  42842=>"00000001",
  42843=>"11111111",
  42844=>"11111100",
  42845=>"11111110",
  42846=>"11111101",
  42847=>"00000000",
  42848=>"11111011",
  42849=>"00000000",
  42850=>"00000011",
  42851=>"11111111",
  42852=>"00000011",
  42853=>"11111110",
  42854=>"00000000",
  42855=>"11111111",
  42856=>"11111100",
  42857=>"00000001",
  42858=>"11111011",
  42859=>"11111110",
  42860=>"00000001",
  42861=>"00000010",
  42862=>"00000011",
  42863=>"00000001",
  42864=>"00000011",
  42865=>"00000001",
  42866=>"11111110",
  42867=>"11111110",
  42868=>"00000001",
  42869=>"00000001",
  42870=>"00000010",
  42871=>"11111110",
  42872=>"00000010",
  42873=>"11111111",
  42874=>"11111110",
  42875=>"11111011",
  42876=>"00000010",
  42877=>"11111111",
  42878=>"00000001",
  42879=>"00000011",
  42880=>"11111010",
  42881=>"00000100",
  42882=>"00000000",
  42883=>"11111110",
  42884=>"11111100",
  42885=>"00000011",
  42886=>"11111111",
  42887=>"00000000",
  42888=>"11111110",
  42889=>"11111101",
  42890=>"11111010",
  42891=>"11111101",
  42892=>"00000010",
  42893=>"11111100",
  42894=>"00000000",
  42895=>"11111110",
  42896=>"11111010",
  42897=>"00000011",
  42898=>"00000010",
  42899=>"11111100",
  42900=>"00000000",
  42901=>"00000010",
  42902=>"11111011",
  42903=>"00000001",
  42904=>"11111110",
  42905=>"11111111",
  42906=>"00000000",
  42907=>"11111111",
  42908=>"00000001",
  42909=>"00000000",
  42910=>"00000001",
  42911=>"11111011",
  42912=>"00000000",
  42913=>"11111010",
  42914=>"00000010",
  42915=>"11111000",
  42916=>"11111010",
  42917=>"11111010",
  42918=>"00000011",
  42919=>"11111011",
  42920=>"11111011",
  42921=>"00000011",
  42922=>"00000001",
  42923=>"11111100",
  42924=>"11111110",
  42925=>"00000010",
  42926=>"11111110",
  42927=>"11111110",
  42928=>"00000011",
  42929=>"11111011",
  42930=>"00000001",
  42931=>"00000000",
  42932=>"00000000",
  42933=>"00000001",
  42934=>"11111101",
  42935=>"00000110",
  42936=>"11111100",
  42937=>"11111111",
  42938=>"11111110",
  42939=>"11111010",
  42940=>"11111100",
  42941=>"00000000",
  42942=>"11111011",
  42943=>"00000011",
  42944=>"00000010",
  42945=>"11111111",
  42946=>"00000000",
  42947=>"11111110",
  42948=>"00000000",
  42949=>"11111111",
  42950=>"11111111",
  42951=>"11111001",
  42952=>"00000100",
  42953=>"11111100",
  42954=>"00000000",
  42955=>"00000000",
  42956=>"11111010",
  42957=>"00000010",
  42958=>"11111110",
  42959=>"11111010",
  42960=>"11111000",
  42961=>"11111110",
  42962=>"00000101",
  42963=>"00000000",
  42964=>"11111001",
  42965=>"00000000",
  42966=>"00000011",
  42967=>"00000000",
  42968=>"11111101",
  42969=>"00000000",
  42970=>"11111110",
  42971=>"00000000",
  42972=>"11111001",
  42973=>"00000011",
  42974=>"11111101",
  42975=>"00000000",
  42976=>"11111111",
  42977=>"00000001",
  42978=>"00000000",
  42979=>"11111100",
  42980=>"11111011",
  42981=>"11111100",
  42982=>"00000001",
  42983=>"11111100",
  42984=>"11111100",
  42985=>"00000000",
  42986=>"00000001",
  42987=>"00000001",
  42988=>"00000000",
  42989=>"11111011",
  42990=>"00000100",
  42991=>"00000000",
  42992=>"11111101",
  42993=>"00000010",
  42994=>"00000010",
  42995=>"11111101",
  42996=>"11111011",
  42997=>"00000010",
  42998=>"00000000",
  42999=>"11111111",
  43000=>"11111101",
  43001=>"11110111",
  43002=>"11111111",
  43003=>"11111111",
  43004=>"00000011",
  43005=>"00000110",
  43006=>"11111111",
  43007=>"11111100",
  43008=>"11111110",
  43009=>"11111111",
  43010=>"00000000",
  43011=>"00000001",
  43012=>"11111110",
  43013=>"11111100",
  43014=>"00000001",
  43015=>"00000010",
  43016=>"11111101",
  43017=>"11111111",
  43018=>"00000000",
  43019=>"00000011",
  43020=>"11111111",
  43021=>"11111101",
  43022=>"00000010",
  43023=>"00000000",
  43024=>"00000001",
  43025=>"00000011",
  43026=>"11111110",
  43027=>"11111101",
  43028=>"11111111",
  43029=>"00000001",
  43030=>"00000000",
  43031=>"00000001",
  43032=>"00000001",
  43033=>"00000011",
  43034=>"11111111",
  43035=>"00000000",
  43036=>"11111111",
  43037=>"00000010",
  43038=>"00000010",
  43039=>"00000101",
  43040=>"11111110",
  43041=>"11111111",
  43042=>"00000000",
  43043=>"00000001",
  43044=>"00000000",
  43045=>"00000000",
  43046=>"00000000",
  43047=>"11111111",
  43048=>"00000001",
  43049=>"11111101",
  43050=>"11111111",
  43051=>"11111111",
  43052=>"11111110",
  43053=>"11111110",
  43054=>"11111110",
  43055=>"00000100",
  43056=>"00000011",
  43057=>"11111101",
  43058=>"00000010",
  43059=>"11111101",
  43060=>"00000010",
  43061=>"00000001",
  43062=>"11111101",
  43063=>"00000000",
  43064=>"11111110",
  43065=>"11111111",
  43066=>"11111101",
  43067=>"00000010",
  43068=>"11111110",
  43069=>"00000010",
  43070=>"00000010",
  43071=>"11111111",
  43072=>"11111101",
  43073=>"11111110",
  43074=>"11111111",
  43075=>"00000001",
  43076=>"00000001",
  43077=>"11111101",
  43078=>"00000001",
  43079=>"11111110",
  43080=>"11111101",
  43081=>"11111110",
  43082=>"00000010",
  43083=>"11111111",
  43084=>"11111110",
  43085=>"00000011",
  43086=>"11111111",
  43087=>"11111110",
  43088=>"11111110",
  43089=>"11111110",
  43090=>"11111110",
  43091=>"11111011",
  43092=>"00000000",
  43093=>"11111111",
  43094=>"11111111",
  43095=>"00000100",
  43096=>"00000010",
  43097=>"00000000",
  43098=>"00000010",
  43099=>"11111100",
  43100=>"11111111",
  43101=>"00000010",
  43102=>"00000000",
  43103=>"00000011",
  43104=>"11111111",
  43105=>"11111110",
  43106=>"11111110",
  43107=>"00000100",
  43108=>"11111111",
  43109=>"11111111",
  43110=>"11111110",
  43111=>"11111111",
  43112=>"11111111",
  43113=>"00000101",
  43114=>"00000001",
  43115=>"00000011",
  43116=>"00000100",
  43117=>"11111111",
  43118=>"11111101",
  43119=>"11111110",
  43120=>"11111110",
  43121=>"11111111",
  43122=>"11111101",
  43123=>"00000101",
  43124=>"00000010",
  43125=>"00000000",
  43126=>"00000010",
  43127=>"00000011",
  43128=>"11111110",
  43129=>"00000001",
  43130=>"00000011",
  43131=>"00000100",
  43132=>"11111111",
  43133=>"00000001",
  43134=>"00000000",
  43135=>"00000001",
  43136=>"11111111",
  43137=>"00000010",
  43138=>"11111111",
  43139=>"00000010",
  43140=>"11111110",
  43141=>"11111111",
  43142=>"11111111",
  43143=>"00000011",
  43144=>"00000000",
  43145=>"11111101",
  43146=>"00000001",
  43147=>"11111110",
  43148=>"11111110",
  43149=>"00000000",
  43150=>"11111111",
  43151=>"11111110",
  43152=>"00000000",
  43153=>"00000001",
  43154=>"11111111",
  43155=>"11111110",
  43156=>"11111110",
  43157=>"11111111",
  43158=>"00000001",
  43159=>"11111110",
  43160=>"11111101",
  43161=>"00000000",
  43162=>"11111101",
  43163=>"00000001",
  43164=>"11111110",
  43165=>"00000001",
  43166=>"11111111",
  43167=>"00000010",
  43168=>"00000000",
  43169=>"00000010",
  43170=>"00000000",
  43171=>"11111111",
  43172=>"11111101",
  43173=>"00000010",
  43174=>"11111110",
  43175=>"00000001",
  43176=>"11111101",
  43177=>"00000000",
  43178=>"00000010",
  43179=>"11111111",
  43180=>"11111110",
  43181=>"00000000",
  43182=>"00000001",
  43183=>"11111111",
  43184=>"00000100",
  43185=>"11111101",
  43186=>"00000000",
  43187=>"11111110",
  43188=>"00000000",
  43189=>"11111110",
  43190=>"00000001",
  43191=>"00000000",
  43192=>"00000010",
  43193=>"00000010",
  43194=>"11111110",
  43195=>"00000001",
  43196=>"11111111",
  43197=>"00000000",
  43198=>"00000000",
  43199=>"11111110",
  43200=>"11111101",
  43201=>"11111111",
  43202=>"00000000",
  43203=>"11111111",
  43204=>"11111110",
  43205=>"00000001",
  43206=>"00000110",
  43207=>"11111110",
  43208=>"11111110",
  43209=>"00000000",
  43210=>"00000000",
  43211=>"11111111",
  43212=>"11111101",
  43213=>"11111101",
  43214=>"00000010",
  43215=>"00000101",
  43216=>"11111110",
  43217=>"11111110",
  43218=>"11111110",
  43219=>"11111111",
  43220=>"11111111",
  43221=>"11111111",
  43222=>"11111101",
  43223=>"11111110",
  43224=>"11111110",
  43225=>"11111111",
  43226=>"11111110",
  43227=>"00000011",
  43228=>"00000100",
  43229=>"00000001",
  43230=>"00000001",
  43231=>"11111101",
  43232=>"11111110",
  43233=>"11111110",
  43234=>"11111110",
  43235=>"11111111",
  43236=>"00000010",
  43237=>"00000001",
  43238=>"00000001",
  43239=>"11111101",
  43240=>"00000000",
  43241=>"11111101",
  43242=>"00000001",
  43243=>"00000000",
  43244=>"11111111",
  43245=>"11111111",
  43246=>"00000000",
  43247=>"00000000",
  43248=>"11111111",
  43249=>"00000001",
  43250=>"11111100",
  43251=>"00000100",
  43252=>"11111110",
  43253=>"11111110",
  43254=>"11111110",
  43255=>"11111111",
  43256=>"00000011",
  43257=>"00000000",
  43258=>"11111101",
  43259=>"00000000",
  43260=>"11111110",
  43261=>"00000100",
  43262=>"11111111",
  43263=>"00000011",
  43264=>"11111111",
  43265=>"00000000",
  43266=>"11111100",
  43267=>"11111110",
  43268=>"00000001",
  43269=>"00000011",
  43270=>"11111101",
  43271=>"11111111",
  43272=>"11111110",
  43273=>"00000001",
  43274=>"00000010",
  43275=>"00000000",
  43276=>"11111110",
  43277=>"11111110",
  43278=>"00000011",
  43279=>"00000000",
  43280=>"00000011",
  43281=>"00000011",
  43282=>"00000000",
  43283=>"11111101",
  43284=>"11111100",
  43285=>"00000011",
  43286=>"11111111",
  43287=>"00000010",
  43288=>"11111111",
  43289=>"00000000",
  43290=>"11111110",
  43291=>"00000001",
  43292=>"00000100",
  43293=>"00000010",
  43294=>"11111110",
  43295=>"00000011",
  43296=>"11111111",
  43297=>"11111110",
  43298=>"11111101",
  43299=>"00000100",
  43300=>"11111101",
  43301=>"11111101",
  43302=>"11111110",
  43303=>"11111110",
  43304=>"11111111",
  43305=>"00000001",
  43306=>"00000101",
  43307=>"11111110",
  43308=>"11111101",
  43309=>"00000001",
  43310=>"00000001",
  43311=>"11111101",
  43312=>"00000011",
  43313=>"11111111",
  43314=>"11111111",
  43315=>"00000001",
  43316=>"11111111",
  43317=>"00000000",
  43318=>"00000010",
  43319=>"00000000",
  43320=>"11111110",
  43321=>"11111111",
  43322=>"11111110",
  43323=>"00000010",
  43324=>"11111101",
  43325=>"11111111",
  43326=>"00000001",
  43327=>"00000000",
  43328=>"00000001",
  43329=>"00000000",
  43330=>"00000001",
  43331=>"00000001",
  43332=>"11111110",
  43333=>"00000001",
  43334=>"00000101",
  43335=>"11111110",
  43336=>"11111111",
  43337=>"00000010",
  43338=>"11111111",
  43339=>"00000000",
  43340=>"11111111",
  43341=>"11111110",
  43342=>"00000010",
  43343=>"11111100",
  43344=>"00000000",
  43345=>"00000011",
  43346=>"00000010",
  43347=>"00000000",
  43348=>"11111111",
  43349=>"11111110",
  43350=>"11111110",
  43351=>"00000000",
  43352=>"00000011",
  43353=>"11111110",
  43354=>"11111111",
  43355=>"11111101",
  43356=>"11111110",
  43357=>"11111101",
  43358=>"00000001",
  43359=>"00000010",
  43360=>"00000010",
  43361=>"11111101",
  43362=>"00000010",
  43363=>"11111101",
  43364=>"00000010",
  43365=>"00000010",
  43366=>"11111110",
  43367=>"11111111",
  43368=>"11111111",
  43369=>"00000010",
  43370=>"00000011",
  43371=>"00000001",
  43372=>"00000010",
  43373=>"00000010",
  43374=>"00000001",
  43375=>"11111111",
  43376=>"00000000",
  43377=>"00000010",
  43378=>"11111101",
  43379=>"00000010",
  43380=>"00000010",
  43381=>"11111110",
  43382=>"00000000",
  43383=>"00000010",
  43384=>"00000000",
  43385=>"11111101",
  43386=>"00000001",
  43387=>"00000010",
  43388=>"11111110",
  43389=>"11111111",
  43390=>"00000100",
  43391=>"11111100",
  43392=>"11111111",
  43393=>"00000001",
  43394=>"11111101",
  43395=>"11111111",
  43396=>"11111111",
  43397=>"11111110",
  43398=>"11111111",
  43399=>"00000001",
  43400=>"11111101",
  43401=>"11111110",
  43402=>"00000000",
  43403=>"00000011",
  43404=>"11111110",
  43405=>"00000000",
  43406=>"11111111",
  43407=>"00000001",
  43408=>"11111111",
  43409=>"11111111",
  43410=>"11111111",
  43411=>"00000000",
  43412=>"00000000",
  43413=>"11111111",
  43414=>"00000011",
  43415=>"11111101",
  43416=>"11111111",
  43417=>"00000100",
  43418=>"00000010",
  43419=>"00000010",
  43420=>"11111110",
  43421=>"00000010",
  43422=>"00000010",
  43423=>"00000000",
  43424=>"11111111",
  43425=>"00000001",
  43426=>"00000001",
  43427=>"00000001",
  43428=>"11111110",
  43429=>"11111110",
  43430=>"11111110",
  43431=>"11111101",
  43432=>"00000100",
  43433=>"00000001",
  43434=>"00000010",
  43435=>"00000010",
  43436=>"00000000",
  43437=>"11111111",
  43438=>"00000000",
  43439=>"00000000",
  43440=>"00000000",
  43441=>"11111100",
  43442=>"00000011",
  43443=>"11111110",
  43444=>"11111111",
  43445=>"00000100",
  43446=>"11111110",
  43447=>"00000001",
  43448=>"00000011",
  43449=>"00000000",
  43450=>"11111110",
  43451=>"00000000",
  43452=>"11111111",
  43453=>"00000001",
  43454=>"11111111",
  43455=>"00000001",
  43456=>"11111111",
  43457=>"11111110",
  43458=>"11111111",
  43459=>"00000001",
  43460=>"00000000",
  43461=>"00000000",
  43462=>"00000010",
  43463=>"11111101",
  43464=>"00000000",
  43465=>"00000010",
  43466=>"11111110",
  43467=>"11111101",
  43468=>"00000001",
  43469=>"00000001",
  43470=>"00000100",
  43471=>"00000010",
  43472=>"00000011",
  43473=>"00000000",
  43474=>"00000011",
  43475=>"11111110",
  43476=>"11111110",
  43477=>"11111110",
  43478=>"00000110",
  43479=>"00000010",
  43480=>"00000001",
  43481=>"11111111",
  43482=>"11111111",
  43483=>"00000111",
  43484=>"00000011",
  43485=>"00000000",
  43486=>"00000001",
  43487=>"11111110",
  43488=>"00000000",
  43489=>"00000010",
  43490=>"00000011",
  43491=>"00000010",
  43492=>"00000010",
  43493=>"00000000",
  43494=>"11111110",
  43495=>"00000000",
  43496=>"11111110",
  43497=>"11111110",
  43498=>"00000011",
  43499=>"00000011",
  43500=>"00000010",
  43501=>"11111111",
  43502=>"00000010",
  43503=>"00000001",
  43504=>"00000011",
  43505=>"11111111",
  43506=>"11111101",
  43507=>"11111111",
  43508=>"00000000",
  43509=>"00000010",
  43510=>"00000010",
  43511=>"00000110",
  43512=>"11111100",
  43513=>"11111110",
  43514=>"00000001",
  43515=>"00000100",
  43516=>"00000001",
  43517=>"11111111",
  43518=>"11111110",
  43519=>"11111110",
  43520=>"11111111",
  43521=>"11111110",
  43522=>"11111110",
  43523=>"11111101",
  43524=>"00000011",
  43525=>"00000000",
  43526=>"00000010",
  43527=>"00000000",
  43528=>"11111111",
  43529=>"00000000",
  43530=>"00000001",
  43531=>"11111110",
  43532=>"00000100",
  43533=>"11111110",
  43534=>"00000011",
  43535=>"00000010",
  43536=>"00000000",
  43537=>"00000111",
  43538=>"11111101",
  43539=>"00000010",
  43540=>"00000100",
  43541=>"11111110",
  43542=>"00000010",
  43543=>"00001000",
  43544=>"00000000",
  43545=>"00000000",
  43546=>"00000100",
  43547=>"11111110",
  43548=>"11111110",
  43549=>"11111110",
  43550=>"11111111",
  43551=>"00000000",
  43552=>"11111101",
  43553=>"00000000",
  43554=>"00000001",
  43555=>"00000110",
  43556=>"00000001",
  43557=>"11111111",
  43558=>"00000010",
  43559=>"11111101",
  43560=>"11111101",
  43561=>"00000000",
  43562=>"00000000",
  43563=>"11111101",
  43564=>"00000001",
  43565=>"11111110",
  43566=>"00001000",
  43567=>"11111101",
  43568=>"11111110",
  43569=>"11111110",
  43570=>"00000010",
  43571=>"11111111",
  43572=>"11111111",
  43573=>"00000001",
  43574=>"11111111",
  43575=>"00000000",
  43576=>"00000010",
  43577=>"11111110",
  43578=>"00000010",
  43579=>"00000010",
  43580=>"11111110",
  43581=>"11111101",
  43582=>"11111110",
  43583=>"00000000",
  43584=>"00000000",
  43585=>"00000010",
  43586=>"11111111",
  43587=>"11111110",
  43588=>"11111111",
  43589=>"11111101",
  43590=>"11111111",
  43591=>"00000010",
  43592=>"00000010",
  43593=>"00000010",
  43594=>"00000000",
  43595=>"11111111",
  43596=>"00000100",
  43597=>"11111111",
  43598=>"11111110",
  43599=>"11111111",
  43600=>"00000000",
  43601=>"11111110",
  43602=>"00000001",
  43603=>"00000010",
  43604=>"11111110",
  43605=>"00000011",
  43606=>"11111111",
  43607=>"00000011",
  43608=>"00000011",
  43609=>"00000110",
  43610=>"11111111",
  43611=>"11111110",
  43612=>"11111101",
  43613=>"00000000",
  43614=>"00000001",
  43615=>"00000000",
  43616=>"00000010",
  43617=>"11111110",
  43618=>"11111101",
  43619=>"00000110",
  43620=>"11111111",
  43621=>"00000000",
  43622=>"11111111",
  43623=>"00000110",
  43624=>"11111101",
  43625=>"00000011",
  43626=>"11111101",
  43627=>"11111110",
  43628=>"11111110",
  43629=>"11111111",
  43630=>"11111111",
  43631=>"00000010",
  43632=>"11111110",
  43633=>"11111101",
  43634=>"00000001",
  43635=>"11111111",
  43636=>"00000010",
  43637=>"00000010",
  43638=>"11111101",
  43639=>"00000001",
  43640=>"00000011",
  43641=>"00000000",
  43642=>"00000110",
  43643=>"00000110",
  43644=>"11111101",
  43645=>"11111111",
  43646=>"11111110",
  43647=>"00000001",
  43648=>"00000010",
  43649=>"00000000",
  43650=>"11111111",
  43651=>"11111110",
  43652=>"11111101",
  43653=>"00000010",
  43654=>"11111101",
  43655=>"11111111",
  43656=>"00000001",
  43657=>"11111101",
  43658=>"00000000",
  43659=>"11111101",
  43660=>"11111111",
  43661=>"00000010",
  43662=>"00000010",
  43663=>"00000000",
  43664=>"00000010",
  43665=>"11111110",
  43666=>"11111110",
  43667=>"00000001",
  43668=>"11111110",
  43669=>"11111111",
  43670=>"00000001",
  43671=>"00000101",
  43672=>"00000010",
  43673=>"11111111",
  43674=>"11111111",
  43675=>"00000011",
  43676=>"00000001",
  43677=>"11111110",
  43678=>"11111111",
  43679=>"00000010",
  43680=>"00000001",
  43681=>"00000011",
  43682=>"00000010",
  43683=>"00000100",
  43684=>"00000000",
  43685=>"00000100",
  43686=>"11111110",
  43687=>"00000010",
  43688=>"11111101",
  43689=>"00000001",
  43690=>"11111111",
  43691=>"11111111",
  43692=>"00000001",
  43693=>"00000000",
  43694=>"11111111",
  43695=>"00000000",
  43696=>"00000100",
  43697=>"11111111",
  43698=>"11111111",
  43699=>"11111110",
  43700=>"00000001",
  43701=>"00000101",
  43702=>"00000110",
  43703=>"00000000",
  43704=>"00000001",
  43705=>"00000000",
  43706=>"11111111",
  43707=>"00000011",
  43708=>"00000000",
  43709=>"00000000",
  43710=>"00000000",
  43711=>"00000000",
  43712=>"11111111",
  43713=>"11111111",
  43714=>"00000000",
  43715=>"11111110",
  43716=>"11111111",
  43717=>"00000000",
  43718=>"11111111",
  43719=>"11111110",
  43720=>"11111111",
  43721=>"11111110",
  43722=>"00000010",
  43723=>"11111100",
  43724=>"00000001",
  43725=>"11111100",
  43726=>"00000001",
  43727=>"00000001",
  43728=>"00000000",
  43729=>"00000100",
  43730=>"00000001",
  43731=>"11111110",
  43732=>"00000010",
  43733=>"00000000",
  43734=>"00000001",
  43735=>"00000010",
  43736=>"11111101",
  43737=>"00000010",
  43738=>"00000000",
  43739=>"00000101",
  43740=>"00000000",
  43741=>"11111110",
  43742=>"00000000",
  43743=>"00000010",
  43744=>"00000000",
  43745=>"00000100",
  43746=>"00000010",
  43747=>"00000100",
  43748=>"00000000",
  43749=>"11111111",
  43750=>"11111111",
  43751=>"11111100",
  43752=>"00000000",
  43753=>"11111110",
  43754=>"11111111",
  43755=>"11111101",
  43756=>"11111110",
  43757=>"00000100",
  43758=>"00000001",
  43759=>"00000010",
  43760=>"00000010",
  43761=>"11111111",
  43762=>"00000001",
  43763=>"00000000",
  43764=>"11111101",
  43765=>"11111110",
  43766=>"11111110",
  43767=>"11111110",
  43768=>"11111101",
  43769=>"00000001",
  43770=>"11111111",
  43771=>"00000000",
  43772=>"00000001",
  43773=>"00000010",
  43774=>"00000000",
  43775=>"11111110",
  43776=>"00000110",
  43777=>"11111111",
  43778=>"11111101",
  43779=>"11111111",
  43780=>"00000011",
  43781=>"11111111",
  43782=>"00000000",
  43783=>"11111101",
  43784=>"00000000",
  43785=>"00000001",
  43786=>"11111111",
  43787=>"00000000",
  43788=>"11111110",
  43789=>"00000101",
  43790=>"11111110",
  43791=>"11111101",
  43792=>"11111110",
  43793=>"11111111",
  43794=>"11111111",
  43795=>"11111110",
  43796=>"00000001",
  43797=>"00000000",
  43798=>"00000000",
  43799=>"00000010",
  43800=>"11111110",
  43801=>"00000011",
  43802=>"00000011",
  43803=>"11111100",
  43804=>"00000000",
  43805=>"00000010",
  43806=>"11111110",
  43807=>"00000000",
  43808=>"11111111",
  43809=>"11111110",
  43810=>"00000010",
  43811=>"00000001",
  43812=>"00000001",
  43813=>"00000000",
  43814=>"00000101",
  43815=>"11111110",
  43816=>"00000001",
  43817=>"11111101",
  43818=>"11111100",
  43819=>"11111111",
  43820=>"11111100",
  43821=>"00000000",
  43822=>"00000000",
  43823=>"00000000",
  43824=>"00000100",
  43825=>"11111100",
  43826=>"00000010",
  43827=>"11111110",
  43828=>"00000001",
  43829=>"00000000",
  43830=>"11111110",
  43831=>"11111100",
  43832=>"11111111",
  43833=>"00000001",
  43834=>"11111110",
  43835=>"11111110",
  43836=>"00000000",
  43837=>"11111111",
  43838=>"00000000",
  43839=>"00000001",
  43840=>"00000101",
  43841=>"11111110",
  43842=>"11111111",
  43843=>"00000000",
  43844=>"00000010",
  43845=>"00000000",
  43846=>"00000001",
  43847=>"00000100",
  43848=>"00000001",
  43849=>"00000010",
  43850=>"11111110",
  43851=>"00000000",
  43852=>"11111111",
  43853=>"00000001",
  43854=>"00000011",
  43855=>"11111111",
  43856=>"00000000",
  43857=>"00000000",
  43858=>"00000001",
  43859=>"11111110",
  43860=>"11111100",
  43861=>"00000010",
  43862=>"11111111",
  43863=>"11111111",
  43864=>"00000001",
  43865=>"00000000",
  43866=>"00000001",
  43867=>"11111100",
  43868=>"00000011",
  43869=>"11111110",
  43870=>"00000001",
  43871=>"00000000",
  43872=>"00000011",
  43873=>"11111101",
  43874=>"11111101",
  43875=>"00000000",
  43876=>"00000011",
  43877=>"00000010",
  43878=>"00000000",
  43879=>"11111110",
  43880=>"00000011",
  43881=>"00000100",
  43882=>"00000000",
  43883=>"11111101",
  43884=>"11111111",
  43885=>"11111111",
  43886=>"11111111",
  43887=>"11111101",
  43888=>"11111011",
  43889=>"00000010",
  43890=>"00000000",
  43891=>"11111110",
  43892=>"00000000",
  43893=>"00000010",
  43894=>"00000011",
  43895=>"00000100",
  43896=>"11111110",
  43897=>"11111101",
  43898=>"11111100",
  43899=>"00000000",
  43900=>"11111111",
  43901=>"00000001",
  43902=>"11111101",
  43903=>"11111100",
  43904=>"00000010",
  43905=>"11111101",
  43906=>"00000001",
  43907=>"00000000",
  43908=>"11111111",
  43909=>"11111110",
  43910=>"00000001",
  43911=>"00000010",
  43912=>"11111101",
  43913=>"00000000",
  43914=>"11111101",
  43915=>"11111111",
  43916=>"00000101",
  43917=>"11111110",
  43918=>"00000000",
  43919=>"00000010",
  43920=>"11111110",
  43921=>"00000001",
  43922=>"00000100",
  43923=>"00000000",
  43924=>"00000010",
  43925=>"00000000",
  43926=>"00000001",
  43927=>"11111101",
  43928=>"00000010",
  43929=>"00000011",
  43930=>"11111111",
  43931=>"11111110",
  43932=>"11111111",
  43933=>"00000010",
  43934=>"00000010",
  43935=>"11111110",
  43936=>"00000001",
  43937=>"11111111",
  43938=>"00000011",
  43939=>"00000010",
  43940=>"00000000",
  43941=>"00000010",
  43942=>"00000000",
  43943=>"00000001",
  43944=>"00000100",
  43945=>"00000100",
  43946=>"11111110",
  43947=>"00000011",
  43948=>"11111101",
  43949=>"00000001",
  43950=>"00000000",
  43951=>"11111101",
  43952=>"00000000",
  43953=>"00000000",
  43954=>"00000001",
  43955=>"11111101",
  43956=>"11111110",
  43957=>"11111110",
  43958=>"11111111",
  43959=>"00000111",
  43960=>"11111101",
  43961=>"00000010",
  43962=>"11111110",
  43963=>"11111111",
  43964=>"00000000",
  43965=>"00000101",
  43966=>"00000010",
  43967=>"11111101",
  43968=>"00000100",
  43969=>"00000010",
  43970=>"11111100",
  43971=>"00000001",
  43972=>"11111110",
  43973=>"00000011",
  43974=>"11111111",
  43975=>"11111110",
  43976=>"11111111",
  43977=>"00000001",
  43978=>"00000011",
  43979=>"00000010",
  43980=>"11111101",
  43981=>"00000001",
  43982=>"00000010",
  43983=>"11111111",
  43984=>"11111101",
  43985=>"00000010",
  43986=>"00000100",
  43987=>"11111110",
  43988=>"11111101",
  43989=>"11111101",
  43990=>"11111101",
  43991=>"11111100",
  43992=>"00000011",
  43993=>"11111101",
  43994=>"11111111",
  43995=>"11111110",
  43996=>"00000010",
  43997=>"11111101",
  43998=>"11111111",
  43999=>"00000001",
  44000=>"00000001",
  44001=>"11111111",
  44002=>"11111111",
  44003=>"00000010",
  44004=>"11111101",
  44005=>"00000001",
  44006=>"00000000",
  44007=>"00000000",
  44008=>"00000000",
  44009=>"11111110",
  44010=>"11111111",
  44011=>"11111110",
  44012=>"00000001",
  44013=>"11111101",
  44014=>"00000111",
  44015=>"00000001",
  44016=>"00000011",
  44017=>"11111111",
  44018=>"00000100",
  44019=>"00000010",
  44020=>"00000001",
  44021=>"00000010",
  44022=>"00000001",
  44023=>"11111111",
  44024=>"11111100",
  44025=>"11111111",
  44026=>"00000000",
  44027=>"00000011",
  44028=>"11111111",
  44029=>"00000001",
  44030=>"00000010",
  44031=>"11111101",
  44032=>"00000010",
  44033=>"11111101",
  44034=>"11111100",
  44035=>"00000100",
  44036=>"00000011",
  44037=>"11111101",
  44038=>"00000000",
  44039=>"11111110",
  44040=>"11111111",
  44041=>"00000100",
  44042=>"00000001",
  44043=>"11111110",
  44044=>"11111101",
  44045=>"11111111",
  44046=>"00000100",
  44047=>"00000001",
  44048=>"11111100",
  44049=>"00000100",
  44050=>"00000000",
  44051=>"00000001",
  44052=>"00000011",
  44053=>"00000000",
  44054=>"11111101",
  44055=>"00000001",
  44056=>"00000010",
  44057=>"00000000",
  44058=>"11111111",
  44059=>"00000011",
  44060=>"11111110",
  44061=>"11111110",
  44062=>"00000011",
  44063=>"11111101",
  44064=>"11111110",
  44065=>"00000110",
  44066=>"11111101",
  44067=>"11111110",
  44068=>"11111110",
  44069=>"00000010",
  44070=>"11111110",
  44071=>"00000000",
  44072=>"00000001",
  44073=>"00000010",
  44074=>"00000010",
  44075=>"00000001",
  44076=>"11111110",
  44077=>"00000000",
  44078=>"00000001",
  44079=>"00000001",
  44080=>"11111111",
  44081=>"11111110",
  44082=>"11111101",
  44083=>"11111100",
  44084=>"00000011",
  44085=>"11111110",
  44086=>"00000010",
  44087=>"00000000",
  44088=>"00000010",
  44089=>"11111111",
  44090=>"00000001",
  44091=>"00000100",
  44092=>"00000000",
  44093=>"00000000",
  44094=>"11111101",
  44095=>"00000010",
  44096=>"00000000",
  44097=>"11111110",
  44098=>"00000010",
  44099=>"00000000",
  44100=>"00000011",
  44101=>"11111111",
  44102=>"11111110",
  44103=>"00000001",
  44104=>"11111110",
  44105=>"00000011",
  44106=>"00000000",
  44107=>"11111111",
  44108=>"00000001",
  44109=>"11111110",
  44110=>"00000011",
  44111=>"00000010",
  44112=>"00000001",
  44113=>"11111101",
  44114=>"00000011",
  44115=>"00000001",
  44116=>"11111110",
  44117=>"00000010",
  44118=>"11111100",
  44119=>"00000001",
  44120=>"11111101",
  44121=>"00000001",
  44122=>"00000000",
  44123=>"00000001",
  44124=>"00000110",
  44125=>"00000000",
  44126=>"11111110",
  44127=>"11111111",
  44128=>"00000001",
  44129=>"11111110",
  44130=>"11111101",
  44131=>"00000010",
  44132=>"00000000",
  44133=>"11111111",
  44134=>"11111111",
  44135=>"00000001",
  44136=>"11111111",
  44137=>"00000011",
  44138=>"11111110",
  44139=>"00000100",
  44140=>"11111111",
  44141=>"11111111",
  44142=>"00000010",
  44143=>"00000010",
  44144=>"11111110",
  44145=>"00000010",
  44146=>"11111111",
  44147=>"11111111",
  44148=>"00000000",
  44149=>"11111111",
  44150=>"11111101",
  44151=>"00000000",
  44152=>"00000010",
  44153=>"00000010",
  44154=>"11111110",
  44155=>"00000011",
  44156=>"11111101",
  44157=>"00000000",
  44158=>"11111111",
  44159=>"00000010",
  44160=>"00000000",
  44161=>"11111111",
  44162=>"00000000",
  44163=>"11111111",
  44164=>"00000001",
  44165=>"11111101",
  44166=>"00000010",
  44167=>"11111100",
  44168=>"11111101",
  44169=>"11111110",
  44170=>"11111110",
  44171=>"11111111",
  44172=>"00000000",
  44173=>"00000011",
  44174=>"11111101",
  44175=>"00000000",
  44176=>"00000010",
  44177=>"11111111",
  44178=>"11111111",
  44179=>"11111111",
  44180=>"00000011",
  44181=>"11111110",
  44182=>"11111101",
  44183=>"11111111",
  44184=>"00000101",
  44185=>"11111110",
  44186=>"00000000",
  44187=>"11111101",
  44188=>"00000001",
  44189=>"00000010",
  44190=>"00000100",
  44191=>"11111110",
  44192=>"11111110",
  44193=>"00000010",
  44194=>"00000001",
  44195=>"00000011",
  44196=>"00000001",
  44197=>"00000001",
  44198=>"11111101",
  44199=>"00000100",
  44200=>"00000001",
  44201=>"11111101",
  44202=>"11111110",
  44203=>"11111111",
  44204=>"11111110",
  44205=>"11111111",
  44206=>"11111110",
  44207=>"00000011",
  44208=>"00000001",
  44209=>"11111110",
  44210=>"11111110",
  44211=>"11111111",
  44212=>"00000010",
  44213=>"00000000",
  44214=>"11111101",
  44215=>"00000001",
  44216=>"00000000",
  44217=>"00000001",
  44218=>"00000000",
  44219=>"11111111",
  44220=>"11111111",
  44221=>"00000001",
  44222=>"00000001",
  44223=>"00000001",
  44224=>"11111110",
  44225=>"11111111",
  44226=>"00000000",
  44227=>"11111110",
  44228=>"00000001",
  44229=>"11111111",
  44230=>"00000011",
  44231=>"11111110",
  44232=>"00000001",
  44233=>"00000100",
  44234=>"00000001",
  44235=>"00000001",
  44236=>"11111110",
  44237=>"00000001",
  44238=>"00000000",
  44239=>"00000000",
  44240=>"00000011",
  44241=>"00000010",
  44242=>"11111111",
  44243=>"00000001",
  44244=>"11111111",
  44245=>"00000000",
  44246=>"11111110",
  44247=>"11111101",
  44248=>"11111101",
  44249=>"00000010",
  44250=>"11111110",
  44251=>"00000000",
  44252=>"00000000",
  44253=>"00000011",
  44254=>"11111110",
  44255=>"00000001",
  44256=>"11111110",
  44257=>"00000001",
  44258=>"00000010",
  44259=>"00000010",
  44260=>"11111110",
  44261=>"11111111",
  44262=>"11111111",
  44263=>"00000001",
  44264=>"11111111",
  44265=>"00000010",
  44266=>"11111111",
  44267=>"00000000",
  44268=>"11111111",
  44269=>"11111101",
  44270=>"11111110",
  44271=>"11111111",
  44272=>"00000001",
  44273=>"11111111",
  44274=>"00000100",
  44275=>"11111111",
  44276=>"00000010",
  44277=>"11111110",
  44278=>"00000000",
  44279=>"00000100",
  44280=>"00000101",
  44281=>"00000000",
  44282=>"11111111",
  44283=>"00000000",
  44284=>"00000010",
  44285=>"00000001",
  44286=>"11111101",
  44287=>"00000001",
  44288=>"11111111",
  44289=>"00000001",
  44290=>"00000010",
  44291=>"11111111",
  44292=>"00000000",
  44293=>"00000010",
  44294=>"11111110",
  44295=>"00000010",
  44296=>"00000001",
  44297=>"11111111",
  44298=>"11111111",
  44299=>"11111110",
  44300=>"00000000",
  44301=>"00000000",
  44302=>"11111111",
  44303=>"00000000",
  44304=>"11111101",
  44305=>"11111111",
  44306=>"00000100",
  44307=>"11111100",
  44308=>"00000000",
  44309=>"11111101",
  44310=>"00000011",
  44311=>"00000000",
  44312=>"00000010",
  44313=>"11111111",
  44314=>"11111101",
  44315=>"11111111",
  44316=>"11111101",
  44317=>"11111110",
  44318=>"11111101",
  44319=>"11111111",
  44320=>"11111111",
  44321=>"00000010",
  44322=>"00000001",
  44323=>"00000000",
  44324=>"11111111",
  44325=>"00000011",
  44326=>"00000001",
  44327=>"11111100",
  44328=>"11111111",
  44329=>"00000011",
  44330=>"11111101",
  44331=>"00000011",
  44332=>"11111111",
  44333=>"00000000",
  44334=>"11111111",
  44335=>"11111111",
  44336=>"00000010",
  44337=>"11111110",
  44338=>"00000010",
  44339=>"11111111",
  44340=>"11111110",
  44341=>"11111111",
  44342=>"00000100",
  44343=>"11111110",
  44344=>"11111110",
  44345=>"11111101",
  44346=>"11111111",
  44347=>"11111100",
  44348=>"11111111",
  44349=>"00000000",
  44350=>"00000000",
  44351=>"11111111",
  44352=>"11111110",
  44353=>"11111101",
  44354=>"00000100",
  44355=>"11111111",
  44356=>"00000011",
  44357=>"11111110",
  44358=>"11111110",
  44359=>"11111111",
  44360=>"11111110",
  44361=>"00000000",
  44362=>"11111110",
  44363=>"00000000",
  44364=>"00000100",
  44365=>"00000001",
  44366=>"00000000",
  44367=>"00000001",
  44368=>"00000001",
  44369=>"00000010",
  44370=>"11111110",
  44371=>"11111101",
  44372=>"11111110",
  44373=>"11111110",
  44374=>"11111111",
  44375=>"11111110",
  44376=>"00000000",
  44377=>"11111111",
  44378=>"11111111",
  44379=>"00000000",
  44380=>"00000011",
  44381=>"00000011",
  44382=>"00000001",
  44383=>"00000010",
  44384=>"11111100",
  44385=>"00000001",
  44386=>"00000000",
  44387=>"11111101",
  44388=>"11111101",
  44389=>"11111101",
  44390=>"11111110",
  44391=>"00000000",
  44392=>"00000001",
  44393=>"00000001",
  44394=>"00000010",
  44395=>"00000000",
  44396=>"11111111",
  44397=>"11111101",
  44398=>"11111111",
  44399=>"11111101",
  44400=>"00000001",
  44401=>"00000001",
  44402=>"11111110",
  44403=>"00000011",
  44404=>"00000001",
  44405=>"11111101",
  44406=>"11111110",
  44407=>"00000011",
  44408=>"00000010",
  44409=>"00000000",
  44410=>"11111110",
  44411=>"00000001",
  44412=>"11111111",
  44413=>"11111101",
  44414=>"00000000",
  44415=>"11111111",
  44416=>"00000010",
  44417=>"00000001",
  44418=>"00000000",
  44419=>"00000010",
  44420=>"11111101",
  44421=>"00000101",
  44422=>"11111101",
  44423=>"00000001",
  44424=>"00000001",
  44425=>"11111101",
  44426=>"11111110",
  44427=>"00000010",
  44428=>"11111101",
  44429=>"00000000",
  44430=>"00000010",
  44431=>"00000010",
  44432=>"11111110",
  44433=>"11111101",
  44434=>"00000001",
  44435=>"00000010",
  44436=>"11111110",
  44437=>"00000011",
  44438=>"00000100",
  44439=>"00000100",
  44440=>"00000000",
  44441=>"11111110",
  44442=>"00000000",
  44443=>"00000011",
  44444=>"11111111",
  44445=>"00000011",
  44446=>"11111111",
  44447=>"11111110",
  44448=>"00000101",
  44449=>"11111110",
  44450=>"11111101",
  44451=>"00000001",
  44452=>"00000011",
  44453=>"11111110",
  44454=>"11111111",
  44455=>"00000000",
  44456=>"11111111",
  44457=>"00000001",
  44458=>"11111111",
  44459=>"11111110",
  44460=>"11111110",
  44461=>"11111111",
  44462=>"11111110",
  44463=>"11111111",
  44464=>"11111111",
  44465=>"00000001",
  44466=>"11111110",
  44467=>"00000001",
  44468=>"00000100",
  44469=>"00000011",
  44470=>"11111111",
  44471=>"11111101",
  44472=>"11111111",
  44473=>"00000010",
  44474=>"11111110",
  44475=>"00000000",
  44476=>"00000010",
  44477=>"00000010",
  44478=>"00000000",
  44479=>"00000010",
  44480=>"00000000",
  44481=>"00000001",
  44482=>"00000001",
  44483=>"00000000",
  44484=>"00000010",
  44485=>"11111111",
  44486=>"11111101",
  44487=>"11111110",
  44488=>"00000011",
  44489=>"00000000",
  44490=>"00000000",
  44491=>"11111111",
  44492=>"00000001",
  44493=>"00000001",
  44494=>"00000000",
  44495=>"11111101",
  44496=>"11111110",
  44497=>"00000001",
  44498=>"00000000",
  44499=>"00000101",
  44500=>"00000001",
  44501=>"00000011",
  44502=>"11111110",
  44503=>"00000010",
  44504=>"00000010",
  44505=>"00000001",
  44506=>"11111111",
  44507=>"00000000",
  44508=>"00000011",
  44509=>"00000011",
  44510=>"11111111",
  44511=>"00000011",
  44512=>"00000001",
  44513=>"11111111",
  44514=>"11111110",
  44515=>"00000001",
  44516=>"00000000",
  44517=>"11111111",
  44518=>"00000010",
  44519=>"00000000",
  44520=>"00000101",
  44521=>"11111110",
  44522=>"00000000",
  44523=>"00000000",
  44524=>"00000001",
  44525=>"11111101",
  44526=>"11111111",
  44527=>"11111100",
  44528=>"00000010",
  44529=>"11111101",
  44530=>"00000011",
  44531=>"00000000",
  44532=>"00000010",
  44533=>"11111110",
  44534=>"11111111",
  44535=>"00000010",
  44536=>"00000000",
  44537=>"00000001",
  44538=>"00000000",
  44539=>"11111111",
  44540=>"00000010",
  44541=>"00000011",
  44542=>"11111101",
  44543=>"11111111",
  44544=>"11111110",
  44545=>"11111110",
  44546=>"00000111",
  44547=>"00000010",
  44548=>"00000000",
  44549=>"00000000",
  44550=>"00000000",
  44551=>"11111100",
  44552=>"00000010",
  44553=>"00000010",
  44554=>"00000000",
  44555=>"00000000",
  44556=>"11111100",
  44557=>"11111101",
  44558=>"11111111",
  44559=>"00000010",
  44560=>"11111110",
  44561=>"00000010",
  44562=>"00000000",
  44563=>"00000100",
  44564=>"00000000",
  44565=>"00000001",
  44566=>"00000011",
  44567=>"11111110",
  44568=>"11111110",
  44569=>"11111111",
  44570=>"00000001",
  44571=>"00000011",
  44572=>"11111111",
  44573=>"00000100",
  44574=>"11111110",
  44575=>"11111111",
  44576=>"00000011",
  44577=>"11111110",
  44578=>"11111110",
  44579=>"11111110",
  44580=>"00000001",
  44581=>"00000000",
  44582=>"11111111",
  44583=>"00000010",
  44584=>"11111111",
  44585=>"00000100",
  44586=>"11111101",
  44587=>"00000000",
  44588=>"00000010",
  44589=>"00000000",
  44590=>"11111110",
  44591=>"00000011",
  44592=>"11111111",
  44593=>"11111111",
  44594=>"00000011",
  44595=>"00000100",
  44596=>"11111110",
  44597=>"00000001",
  44598=>"11111110",
  44599=>"11111111",
  44600=>"11111101",
  44601=>"00000010",
  44602=>"11111111",
  44603=>"00000001",
  44604=>"00000000",
  44605=>"11111111",
  44606=>"00000010",
  44607=>"11111110",
  44608=>"00000001",
  44609=>"11111101",
  44610=>"11111111",
  44611=>"00000000",
  44612=>"00000000",
  44613=>"00000000",
  44614=>"11111101",
  44615=>"00000010",
  44616=>"00000000",
  44617=>"11111111",
  44618=>"11111111",
  44619=>"11111110",
  44620=>"11111101",
  44621=>"11111111",
  44622=>"11111111",
  44623=>"11111111",
  44624=>"00000010",
  44625=>"11111101",
  44626=>"11111110",
  44627=>"00000011",
  44628=>"00000011",
  44629=>"00000010",
  44630=>"11111110",
  44631=>"00000011",
  44632=>"11111110",
  44633=>"00000001",
  44634=>"11111111",
  44635=>"00000000",
  44636=>"11111101",
  44637=>"11111101",
  44638=>"00000010",
  44639=>"00000000",
  44640=>"11111111",
  44641=>"11111110",
  44642=>"11111101",
  44643=>"00000001",
  44644=>"00000100",
  44645=>"11111110",
  44646=>"11111111",
  44647=>"11111110",
  44648=>"00000000",
  44649=>"00000010",
  44650=>"00000001",
  44651=>"00000001",
  44652=>"00000110",
  44653=>"00000011",
  44654=>"00000100",
  44655=>"00000001",
  44656=>"11111110",
  44657=>"11111111",
  44658=>"00000001",
  44659=>"11111101",
  44660=>"00000010",
  44661=>"11111110",
  44662=>"11111101",
  44663=>"00000001",
  44664=>"00000001",
  44665=>"11111110",
  44666=>"00000000",
  44667=>"00000001",
  44668=>"11111110",
  44669=>"11111111",
  44670=>"11111111",
  44671=>"11111111",
  44672=>"00000000",
  44673=>"00000000",
  44674=>"00000001",
  44675=>"11111110",
  44676=>"00000101",
  44677=>"11111111",
  44678=>"00000100",
  44679=>"00000000",
  44680=>"00000001",
  44681=>"11111110",
  44682=>"11111110",
  44683=>"00000101",
  44684=>"00000000",
  44685=>"11111110",
  44686=>"00000001",
  44687=>"00000000",
  44688=>"11111111",
  44689=>"11111111",
  44690=>"00000001",
  44691=>"11111110",
  44692=>"00000010",
  44693=>"00000001",
  44694=>"00000011",
  44695=>"00000010",
  44696=>"00000111",
  44697=>"11111110",
  44698=>"00000011",
  44699=>"11111110",
  44700=>"00000100",
  44701=>"11111111",
  44702=>"00000000",
  44703=>"00000001",
  44704=>"00000011",
  44705=>"11111110",
  44706=>"00000011",
  44707=>"00000001",
  44708=>"11111111",
  44709=>"00000000",
  44710=>"11111111",
  44711=>"11111110",
  44712=>"00000011",
  44713=>"00000001",
  44714=>"00000101",
  44715=>"11111101",
  44716=>"00000001",
  44717=>"00000001",
  44718=>"00000010",
  44719=>"11111100",
  44720=>"11111110",
  44721=>"11111111",
  44722=>"11111110",
  44723=>"00000000",
  44724=>"11111111",
  44725=>"11111110",
  44726=>"00000100",
  44727=>"11111101",
  44728=>"00000001",
  44729=>"00000010",
  44730=>"11111110",
  44731=>"11111111",
  44732=>"11111101",
  44733=>"00000000",
  44734=>"00000001",
  44735=>"00000000",
  44736=>"00000001",
  44737=>"00000000",
  44738=>"11111100",
  44739=>"11111110",
  44740=>"00000011",
  44741=>"11111110",
  44742=>"11111110",
  44743=>"00000000",
  44744=>"00000001",
  44745=>"11111101",
  44746=>"00000001",
  44747=>"11111111",
  44748=>"00000100",
  44749=>"00000001",
  44750=>"11111111",
  44751=>"00000011",
  44752=>"11111110",
  44753=>"00000000",
  44754=>"00000001",
  44755=>"11111110",
  44756=>"00000000",
  44757=>"00000000",
  44758=>"11111111",
  44759=>"11111110",
  44760=>"11111111",
  44761=>"11111111",
  44762=>"00000001",
  44763=>"00000001",
  44764=>"00000110",
  44765=>"00000000",
  44766=>"11111110",
  44767=>"00000000",
  44768=>"00000101",
  44769=>"11111101",
  44770=>"00000010",
  44771=>"00000011",
  44772=>"00000000",
  44773=>"00000011",
  44774=>"00000000",
  44775=>"00000101",
  44776=>"11111101",
  44777=>"11111111",
  44778=>"11111110",
  44779=>"00000001",
  44780=>"11111101",
  44781=>"11111111",
  44782=>"00000000",
  44783=>"11111110",
  44784=>"11111110",
  44785=>"11111101",
  44786=>"11111111",
  44787=>"00000000",
  44788=>"00000000",
  44789=>"00000010",
  44790=>"00000011",
  44791=>"11111110",
  44792=>"11111100",
  44793=>"00000000",
  44794=>"00000010",
  44795=>"00000100",
  44796=>"00000011",
  44797=>"00000011",
  44798=>"00000001",
  44799=>"00000010",
  44800=>"00000100",
  44801=>"11111110",
  44802=>"00000011",
  44803=>"11111110",
  44804=>"11111101",
  44805=>"11111111",
  44806=>"11111111",
  44807=>"11111110",
  44808=>"00000001",
  44809=>"00000001",
  44810=>"00000010",
  44811=>"00000100",
  44812=>"00000000",
  44813=>"11111111",
  44814=>"00000011",
  44815=>"11111110",
  44816=>"11111111",
  44817=>"11111111",
  44818=>"00000010",
  44819=>"11111110",
  44820=>"00000011",
  44821=>"00000000",
  44822=>"11111111",
  44823=>"00000010",
  44824=>"11111100",
  44825=>"11111101",
  44826=>"00000010",
  44827=>"11111100",
  44828=>"11111110",
  44829=>"11111110",
  44830=>"11111101",
  44831=>"11111101",
  44832=>"00000000",
  44833=>"00000011",
  44834=>"11111111",
  44835=>"00000010",
  44836=>"11111111",
  44837=>"00000111",
  44838=>"00000101",
  44839=>"00000001",
  44840=>"11111101",
  44841=>"00000001",
  44842=>"00000001",
  44843=>"00000001",
  44844=>"11111110",
  44845=>"00000001",
  44846=>"00000001",
  44847=>"00000010",
  44848=>"00000001",
  44849=>"11111110",
  44850=>"00000010",
  44851=>"00000000",
  44852=>"00000010",
  44853=>"11111101",
  44854=>"00000000",
  44855=>"00000011",
  44856=>"11111110",
  44857=>"00000000",
  44858=>"11111110",
  44859=>"00000000",
  44860=>"00000010",
  44861=>"11111101",
  44862=>"00000001",
  44863=>"11111111",
  44864=>"00000001",
  44865=>"00000001",
  44866=>"11111110",
  44867=>"11111101",
  44868=>"11111111",
  44869=>"11111111",
  44870=>"00000011",
  44871=>"00000101",
  44872=>"11111111",
  44873=>"00000001",
  44874=>"11111111",
  44875=>"11111111",
  44876=>"11111111",
  44877=>"00000000",
  44878=>"11111100",
  44879=>"11111101",
  44880=>"11111101",
  44881=>"00000010",
  44882=>"00000011",
  44883=>"00000011",
  44884=>"11111110",
  44885=>"11111110",
  44886=>"00000010",
  44887=>"11111111",
  44888=>"00000110",
  44889=>"00000010",
  44890=>"00000100",
  44891=>"11111111",
  44892=>"00000100",
  44893=>"00000000",
  44894=>"11111101",
  44895=>"00000011",
  44896=>"11111110",
  44897=>"11111111",
  44898=>"00000001",
  44899=>"00000011",
  44900=>"00000001",
  44901=>"00000000",
  44902=>"00000001",
  44903=>"00000010",
  44904=>"11111111",
  44905=>"00000001",
  44906=>"00000010",
  44907=>"00000000",
  44908=>"00000000",
  44909=>"00000010",
  44910=>"00000001",
  44911=>"00000001",
  44912=>"00000011",
  44913=>"00000000",
  44914=>"00000000",
  44915=>"11111110",
  44916=>"00000010",
  44917=>"11111111",
  44918=>"00000010",
  44919=>"00000001",
  44920=>"11111101",
  44921=>"00000001",
  44922=>"00000000",
  44923=>"11111110",
  44924=>"00000001",
  44925=>"11111111",
  44926=>"00000010",
  44927=>"00000011",
  44928=>"00000001",
  44929=>"00000001",
  44930=>"00000001",
  44931=>"11111110",
  44932=>"11111110",
  44933=>"11111110",
  44934=>"00000001",
  44935=>"00000010",
  44936=>"11111110",
  44937=>"00000000",
  44938=>"11111110",
  44939=>"00000010",
  44940=>"00000010",
  44941=>"00000000",
  44942=>"11111110",
  44943=>"00000000",
  44944=>"11111110",
  44945=>"00000010",
  44946=>"00000000",
  44947=>"11111110",
  44948=>"11111101",
  44949=>"11111110",
  44950=>"00000001",
  44951=>"11111111",
  44952=>"00000000",
  44953=>"00000011",
  44954=>"00000000",
  44955=>"11111111",
  44956=>"11111110",
  44957=>"11111111",
  44958=>"11111111",
  44959=>"00000100",
  44960=>"00000011",
  44961=>"00000000",
  44962=>"11111100",
  44963=>"11111101",
  44964=>"00000001",
  44965=>"00000010",
  44966=>"11111111",
  44967=>"00000010",
  44968=>"00000000",
  44969=>"00000011",
  44970=>"00000011",
  44971=>"11111110",
  44972=>"11111111",
  44973=>"11111110",
  44974=>"00000010",
  44975=>"00000001",
  44976=>"00000110",
  44977=>"00000000",
  44978=>"00000000",
  44979=>"11111101",
  44980=>"00000011",
  44981=>"11111110",
  44982=>"11111111",
  44983=>"00000001",
  44984=>"11111110",
  44985=>"00000011",
  44986=>"00000011",
  44987=>"11111110",
  44988=>"11111111",
  44989=>"11111111",
  44990=>"11111110",
  44991=>"11111110",
  44992=>"11111110",
  44993=>"11111110",
  44994=>"11111111",
  44995=>"11111110",
  44996=>"00000011",
  44997=>"00000001",
  44998=>"11111101",
  44999=>"00000000",
  45000=>"00000000",
  45001=>"00000001",
  45002=>"00000000",
  45003=>"00000011",
  45004=>"00000010",
  45005=>"11111110",
  45006=>"11111110",
  45007=>"00000010",
  45008=>"00000011",
  45009=>"00000011",
  45010=>"00000001",
  45011=>"00000000",
  45012=>"00000010",
  45013=>"11111111",
  45014=>"11111100",
  45015=>"00000011",
  45016=>"11111111",
  45017=>"00000011",
  45018=>"11111110",
  45019=>"00000010",
  45020=>"11111111",
  45021=>"00000001",
  45022=>"00000010",
  45023=>"00000011",
  45024=>"11111111",
  45025=>"11111110",
  45026=>"00000001",
  45027=>"00000000",
  45028=>"00000010",
  45029=>"00000001",
  45030=>"00000010",
  45031=>"11111110",
  45032=>"00000000",
  45033=>"11111111",
  45034=>"11111110",
  45035=>"11111110",
  45036=>"00000001",
  45037=>"11111111",
  45038=>"11111100",
  45039=>"11111110",
  45040=>"11111101",
  45041=>"00000011",
  45042=>"00000100",
  45043=>"11111101",
  45044=>"00000000",
  45045=>"00000100",
  45046=>"11111100",
  45047=>"00000001",
  45048=>"00000000",
  45049=>"11111111",
  45050=>"11111111",
  45051=>"00000110",
  45052=>"00000010",
  45053=>"00000000",
  45054=>"00000000",
  45055=>"11111110",
  45056=>"11111111",
  45057=>"11111110",
  45058=>"00000001",
  45059=>"11111101",
  45060=>"11111101",
  45061=>"11111101",
  45062=>"00000000",
  45063=>"00000000",
  45064=>"11111111",
  45065=>"11111111",
  45066=>"00000011",
  45067=>"11111101",
  45068=>"00000100",
  45069=>"00000100",
  45070=>"11111110",
  45071=>"00000010",
  45072=>"00000111",
  45073=>"11111111",
  45074=>"00000010",
  45075=>"11111110",
  45076=>"11111110",
  45077=>"00000011",
  45078=>"11111111",
  45079=>"00000100",
  45080=>"11111101",
  45081=>"11111110",
  45082=>"00000001",
  45083=>"00000010",
  45084=>"00000010",
  45085=>"00000000",
  45086=>"00000001",
  45087=>"00000010",
  45088=>"00000001",
  45089=>"11111111",
  45090=>"11111110",
  45091=>"11111100",
  45092=>"00000000",
  45093=>"11111111",
  45094=>"00000001",
  45095=>"11111101",
  45096=>"11111111",
  45097=>"11111110",
  45098=>"11111101",
  45099=>"00000001",
  45100=>"00000001",
  45101=>"00000001",
  45102=>"00000010",
  45103=>"00000001",
  45104=>"00000010",
  45105=>"00000001",
  45106=>"00000001",
  45107=>"00000011",
  45108=>"00000010",
  45109=>"00000011",
  45110=>"00000001",
  45111=>"00000011",
  45112=>"11111110",
  45113=>"00000000",
  45114=>"00000010",
  45115=>"00000011",
  45116=>"11111101",
  45117=>"00000010",
  45118=>"00000010",
  45119=>"11111101",
  45120=>"11111101",
  45121=>"00000110",
  45122=>"11111110",
  45123=>"00000000",
  45124=>"00000001",
  45125=>"00000010",
  45126=>"00000010",
  45127=>"00000000",
  45128=>"11111111",
  45129=>"11111101",
  45130=>"11111111",
  45131=>"11111101",
  45132=>"00000010",
  45133=>"11111110",
  45134=>"00000001",
  45135=>"11111110",
  45136=>"11111110",
  45137=>"00000000",
  45138=>"11111101",
  45139=>"00000001",
  45140=>"11111111",
  45141=>"11111111",
  45142=>"00000010",
  45143=>"00000001",
  45144=>"00000010",
  45145=>"00000001",
  45146=>"00000000",
  45147=>"00000100",
  45148=>"00000000",
  45149=>"00000000",
  45150=>"00000011",
  45151=>"00000000",
  45152=>"00000000",
  45153=>"11111110",
  45154=>"11111111",
  45155=>"11111101",
  45156=>"00000010",
  45157=>"00000000",
  45158=>"00000000",
  45159=>"11111111",
  45160=>"00000010",
  45161=>"00000011",
  45162=>"00000000",
  45163=>"11111111",
  45164=>"11111101",
  45165=>"11111111",
  45166=>"00000010",
  45167=>"00000001",
  45168=>"00000011",
  45169=>"00000010",
  45170=>"11111111",
  45171=>"00000000",
  45172=>"11111101",
  45173=>"11111101",
  45174=>"11111101",
  45175=>"00000100",
  45176=>"00000010",
  45177=>"00000001",
  45178=>"00000000",
  45179=>"11111111",
  45180=>"00000000",
  45181=>"00000000",
  45182=>"00000100",
  45183=>"11111100",
  45184=>"00000010",
  45185=>"11111111",
  45186=>"11111101",
  45187=>"00000001",
  45188=>"00000001",
  45189=>"00000000",
  45190=>"11111101",
  45191=>"11111111",
  45192=>"00000000",
  45193=>"00000101",
  45194=>"00000010",
  45195=>"00000000",
  45196=>"11111101",
  45197=>"00000000",
  45198=>"11111101",
  45199=>"11111100",
  45200=>"11111111",
  45201=>"11111101",
  45202=>"00000001",
  45203=>"00000001",
  45204=>"11111110",
  45205=>"00000100",
  45206=>"11111110",
  45207=>"11111101",
  45208=>"00000011",
  45209=>"00000101",
  45210=>"11111111",
  45211=>"11111110",
  45212=>"00000000",
  45213=>"11111110",
  45214=>"11111111",
  45215=>"11111101",
  45216=>"00000001",
  45217=>"11111111",
  45218=>"00000100",
  45219=>"00000000",
  45220=>"00000011",
  45221=>"00000100",
  45222=>"11111101",
  45223=>"11111111",
  45224=>"00000001",
  45225=>"11111100",
  45226=>"11111101",
  45227=>"00000001",
  45228=>"00000000",
  45229=>"11111111",
  45230=>"00000001",
  45231=>"11111110",
  45232=>"00000000",
  45233=>"11111110",
  45234=>"00000001",
  45235=>"11111101",
  45236=>"11111101",
  45237=>"00000001",
  45238=>"11111110",
  45239=>"00000010",
  45240=>"00000010",
  45241=>"11111111",
  45242=>"11111101",
  45243=>"11111101",
  45244=>"00000010",
  45245=>"00000000",
  45246=>"11111111",
  45247=>"00000000",
  45248=>"00000010",
  45249=>"00000011",
  45250=>"11111111",
  45251=>"00000000",
  45252=>"00000010",
  45253=>"11111111",
  45254=>"11111110",
  45255=>"11111111",
  45256=>"11111111",
  45257=>"11111101",
  45258=>"11111110",
  45259=>"00000001",
  45260=>"00000001",
  45261=>"00000011",
  45262=>"11111110",
  45263=>"11111111",
  45264=>"11111111",
  45265=>"11111111",
  45266=>"00000000",
  45267=>"00000100",
  45268=>"00000001",
  45269=>"11111111",
  45270=>"11111111",
  45271=>"11111101",
  45272=>"11111101",
  45273=>"00000001",
  45274=>"00000000",
  45275=>"00000010",
  45276=>"11111111",
  45277=>"00000010",
  45278=>"11111110",
  45279=>"11111110",
  45280=>"00000010",
  45281=>"00000001",
  45282=>"00000011",
  45283=>"00000001",
  45284=>"00000001",
  45285=>"11111101",
  45286=>"00000101",
  45287=>"11111110",
  45288=>"00000001",
  45289=>"00000011",
  45290=>"11111101",
  45291=>"00000000",
  45292=>"00000010",
  45293=>"11111101",
  45294=>"00000011",
  45295=>"11111111",
  45296=>"00000010",
  45297=>"00000001",
  45298=>"11111100",
  45299=>"11111111",
  45300=>"11111101",
  45301=>"00000000",
  45302=>"00000001",
  45303=>"11111101",
  45304=>"00000001",
  45305=>"11111111",
  45306=>"11111100",
  45307=>"11111110",
  45308=>"11111101",
  45309=>"11111111",
  45310=>"11111101",
  45311=>"00000010",
  45312=>"00000010",
  45313=>"11111100",
  45314=>"00000010",
  45315=>"00000001",
  45316=>"00000000",
  45317=>"11111111",
  45318=>"00000010",
  45319=>"11111101",
  45320=>"11111111",
  45321=>"11111111",
  45322=>"11111111",
  45323=>"11111110",
  45324=>"11111110",
  45325=>"11111111",
  45326=>"00000000",
  45327=>"11111101",
  45328=>"00000011",
  45329=>"00000000",
  45330=>"00000010",
  45331=>"00000001",
  45332=>"11111110",
  45333=>"00000000",
  45334=>"00000000",
  45335=>"11111101",
  45336=>"00000101",
  45337=>"11111110",
  45338=>"00000000",
  45339=>"11111110",
  45340=>"00000000",
  45341=>"00000000",
  45342=>"00000100",
  45343=>"00000100",
  45344=>"00000011",
  45345=>"00000001",
  45346=>"11111111",
  45347=>"11111110",
  45348=>"00000001",
  45349=>"11111101",
  45350=>"00000011",
  45351=>"11111100",
  45352=>"00000000",
  45353=>"00000010",
  45354=>"11111111",
  45355=>"00000001",
  45356=>"11111111",
  45357=>"00000011",
  45358=>"00000010",
  45359=>"11111101",
  45360=>"00000001",
  45361=>"00000000",
  45362=>"11111101",
  45363=>"00000011",
  45364=>"11111101",
  45365=>"11111101",
  45366=>"11111110",
  45367=>"00000010",
  45368=>"11111111",
  45369=>"11111110",
  45370=>"00000010",
  45371=>"11111101",
  45372=>"00000010",
  45373=>"00000010",
  45374=>"00000000",
  45375=>"00000001",
  45376=>"11111111",
  45377=>"00000001",
  45378=>"00000001",
  45379=>"11111110",
  45380=>"11111110",
  45381=>"11111111",
  45382=>"11111110",
  45383=>"00000001",
  45384=>"11111110",
  45385=>"00000001",
  45386=>"11111110",
  45387=>"00000001",
  45388=>"11111111",
  45389=>"11111110",
  45390=>"00000001",
  45391=>"11111101",
  45392=>"00000010",
  45393=>"00000010",
  45394=>"11111101",
  45395=>"00000101",
  45396=>"11111101",
  45397=>"11111110",
  45398=>"00000101",
  45399=>"11111111",
  45400=>"00000000",
  45401=>"00000001",
  45402=>"11111111",
  45403=>"11111110",
  45404=>"00000001",
  45405=>"11111101",
  45406=>"00000001",
  45407=>"11111100",
  45408=>"00000101",
  45409=>"00000000",
  45410=>"11111110",
  45411=>"11111100",
  45412=>"11111110",
  45413=>"11111111",
  45414=>"00000010",
  45415=>"00000000",
  45416=>"11111101",
  45417=>"00000001",
  45418=>"00000011",
  45419=>"00000010",
  45420=>"11111100",
  45421=>"00000000",
  45422=>"00000010",
  45423=>"00000010",
  45424=>"00000001",
  45425=>"00000010",
  45426=>"00000001",
  45427=>"00000001",
  45428=>"11111101",
  45429=>"00000011",
  45430=>"11111111",
  45431=>"00000001",
  45432=>"11111111",
  45433=>"00000000",
  45434=>"00000011",
  45435=>"11111101",
  45436=>"00000001",
  45437=>"00000001",
  45438=>"11111101",
  45439=>"11111111",
  45440=>"00000100",
  45441=>"11111100",
  45442=>"00000001",
  45443=>"00000010",
  45444=>"00000010",
  45445=>"11111110",
  45446=>"11111101",
  45447=>"00000001",
  45448=>"00000010",
  45449=>"00000000",
  45450=>"00000000",
  45451=>"11111101",
  45452=>"00000010",
  45453=>"11111110",
  45454=>"11111101",
  45455=>"11111111",
  45456=>"11111111",
  45457=>"00000100",
  45458=>"11111111",
  45459=>"11111111",
  45460=>"11111111",
  45461=>"11111110",
  45462=>"11111110",
  45463=>"00000010",
  45464=>"00000001",
  45465=>"11111101",
  45466=>"00000001",
  45467=>"00000000",
  45468=>"11111101",
  45469=>"11111101",
  45470=>"11111110",
  45471=>"00000101",
  45472=>"11111111",
  45473=>"00000001",
  45474=>"00000000",
  45475=>"11111100",
  45476=>"00000000",
  45477=>"00000010",
  45478=>"00000011",
  45479=>"00000000",
  45480=>"11111100",
  45481=>"00000011",
  45482=>"00000001",
  45483=>"00000001",
  45484=>"00000010",
  45485=>"00000010",
  45486=>"11111111",
  45487=>"00000011",
  45488=>"00000010",
  45489=>"00000000",
  45490=>"11111111",
  45491=>"11111101",
  45492=>"00000001",
  45493=>"00000010",
  45494=>"11111110",
  45495=>"00000010",
  45496=>"00000101",
  45497=>"11111110",
  45498=>"11111111",
  45499=>"00000001",
  45500=>"11111110",
  45501=>"11111101",
  45502=>"00000000",
  45503=>"00000000",
  45504=>"11111101",
  45505=>"11111101",
  45506=>"00000000",
  45507=>"00000100",
  45508=>"11111100",
  45509=>"11111110",
  45510=>"00000000",
  45511=>"11111100",
  45512=>"00000100",
  45513=>"00000001",
  45514=>"00000101",
  45515=>"00000001",
  45516=>"11111110",
  45517=>"00000000",
  45518=>"00000000",
  45519=>"11111100",
  45520=>"00000010",
  45521=>"11111110",
  45522=>"11111101",
  45523=>"00000001",
  45524=>"00000000",
  45525=>"11111111",
  45526=>"00000000",
  45527=>"11111111",
  45528=>"00000000",
  45529=>"00000001",
  45530=>"11111101",
  45531=>"00000010",
  45532=>"11111111",
  45533=>"00000001",
  45534=>"11111110",
  45535=>"11111111",
  45536=>"00000010",
  45537=>"00000010",
  45538=>"11111111",
  45539=>"00000010",
  45540=>"11111110",
  45541=>"00000011",
  45542=>"00000000",
  45543=>"11111101",
  45544=>"11111110",
  45545=>"00000010",
  45546=>"00000001",
  45547=>"00000011",
  45548=>"11111111",
  45549=>"11111110",
  45550=>"00000000",
  45551=>"11111011",
  45552=>"11111111",
  45553=>"00000001",
  45554=>"00000010",
  45555=>"00000001",
  45556=>"00000000",
  45557=>"00000000",
  45558=>"11111100",
  45559=>"00000010",
  45560=>"00000001",
  45561=>"11111111",
  45562=>"00000001",
  45563=>"00000001",
  45564=>"00000101",
  45565=>"00000011",
  45566=>"11111111",
  45567=>"00000100",
  45568=>"00000001",
  45569=>"00000000",
  45570=>"11111110",
  45571=>"11111110",
  45572=>"00000000",
  45573=>"11111110",
  45574=>"11111110",
  45575=>"00000011",
  45576=>"00000001",
  45577=>"00000011",
  45578=>"11111111",
  45579=>"00000010",
  45580=>"11111110",
  45581=>"11111110",
  45582=>"11111100",
  45583=>"00000001",
  45584=>"11111110",
  45585=>"00000010",
  45586=>"11111111",
  45587=>"11111101",
  45588=>"11111110",
  45589=>"00000001",
  45590=>"11111111",
  45591=>"00000001",
  45592=>"00000010",
  45593=>"00000110",
  45594=>"00000001",
  45595=>"00000010",
  45596=>"00000010",
  45597=>"00000001",
  45598=>"11111111",
  45599=>"00000001",
  45600=>"11111110",
  45601=>"00000000",
  45602=>"00000010",
  45603=>"00000010",
  45604=>"00000000",
  45605=>"11111101",
  45606=>"00000001",
  45607=>"11111110",
  45608=>"00000010",
  45609=>"11111101",
  45610=>"11111101",
  45611=>"11111101",
  45612=>"11111110",
  45613=>"11111110",
  45614=>"00000001",
  45615=>"11111101",
  45616=>"11111101",
  45617=>"00000001",
  45618=>"00000010",
  45619=>"00000000",
  45620=>"11111100",
  45621=>"00000100",
  45622=>"00000000",
  45623=>"00000010",
  45624=>"00000011",
  45625=>"11111101",
  45626=>"00000001",
  45627=>"00000001",
  45628=>"00000010",
  45629=>"00000001",
  45630=>"00000000",
  45631=>"11111101",
  45632=>"00000000",
  45633=>"00000000",
  45634=>"11111110",
  45635=>"00000010",
  45636=>"11111110",
  45637=>"00000000",
  45638=>"11111110",
  45639=>"00000010",
  45640=>"00000000",
  45641=>"00000000",
  45642=>"00000000",
  45643=>"00000010",
  45644=>"00000001",
  45645=>"11111111",
  45646=>"11111111",
  45647=>"11111110",
  45648=>"00000001",
  45649=>"00000011",
  45650=>"00000010",
  45651=>"00000001",
  45652=>"00000011",
  45653=>"11111110",
  45654=>"00000001",
  45655=>"00000001",
  45656=>"11111110",
  45657=>"11111111",
  45658=>"00000001",
  45659=>"11111101",
  45660=>"11111100",
  45661=>"11111110",
  45662=>"11111110",
  45663=>"00000000",
  45664=>"00000000",
  45665=>"11111111",
  45666=>"11111111",
  45667=>"00000001",
  45668=>"11111101",
  45669=>"00000011",
  45670=>"11111111",
  45671=>"00000100",
  45672=>"11111111",
  45673=>"00000101",
  45674=>"00000001",
  45675=>"11111111",
  45676=>"11111111",
  45677=>"11111110",
  45678=>"11111101",
  45679=>"11111101",
  45680=>"00000110",
  45681=>"00000100",
  45682=>"00000001",
  45683=>"00000001",
  45684=>"11111111",
  45685=>"00000000",
  45686=>"00000001",
  45687=>"11111110",
  45688=>"00000100",
  45689=>"00000000",
  45690=>"00000001",
  45691=>"11111101",
  45692=>"00000011",
  45693=>"00000010",
  45694=>"00000000",
  45695=>"00000000",
  45696=>"11111110",
  45697=>"11111110",
  45698=>"11111101",
  45699=>"11111101",
  45700=>"11111110",
  45701=>"00000010",
  45702=>"11111101",
  45703=>"00000000",
  45704=>"11111111",
  45705=>"00000101",
  45706=>"11111111",
  45707=>"00000000",
  45708=>"00000010",
  45709=>"00000010",
  45710=>"00000110",
  45711=>"00000110",
  45712=>"00000000",
  45713=>"00000000",
  45714=>"00000101",
  45715=>"00000001",
  45716=>"00000001",
  45717=>"00000000",
  45718=>"11111110",
  45719=>"11111111",
  45720=>"11111110",
  45721=>"00000010",
  45722=>"00000011",
  45723=>"11111110",
  45724=>"00000000",
  45725=>"11111101",
  45726=>"00000010",
  45727=>"11111101",
  45728=>"00000000",
  45729=>"11111110",
  45730=>"11111111",
  45731=>"11111110",
  45732=>"00000000",
  45733=>"00000000",
  45734=>"00000001",
  45735=>"11111100",
  45736=>"11111111",
  45737=>"11111101",
  45738=>"00000011",
  45739=>"11111101",
  45740=>"00000011",
  45741=>"00000011",
  45742=>"11111101",
  45743=>"00000000",
  45744=>"00000001",
  45745=>"00000001",
  45746=>"00000000",
  45747=>"00000001",
  45748=>"11111111",
  45749=>"00000000",
  45750=>"11111101",
  45751=>"00000001",
  45752=>"00000000",
  45753=>"00000011",
  45754=>"00000011",
  45755=>"11111111",
  45756=>"11111111",
  45757=>"11111111",
  45758=>"00000000",
  45759=>"11111101",
  45760=>"00000000",
  45761=>"00000001",
  45762=>"00000000",
  45763=>"11111110",
  45764=>"11111111",
  45765=>"11111101",
  45766=>"11111101",
  45767=>"00000010",
  45768=>"00000011",
  45769=>"00000010",
  45770=>"00000011",
  45771=>"11111111",
  45772=>"00000000",
  45773=>"00000111",
  45774=>"00000010",
  45775=>"00000011",
  45776=>"00000010",
  45777=>"11111111",
  45778=>"00000000",
  45779=>"11111110",
  45780=>"11111101",
  45781=>"00000000",
  45782=>"00000011",
  45783=>"00000001",
  45784=>"11111101",
  45785=>"00000101",
  45786=>"11111110",
  45787=>"00000001",
  45788=>"11111101",
  45789=>"00000000",
  45790=>"00000010",
  45791=>"00000001",
  45792=>"11111111",
  45793=>"11111111",
  45794=>"00000110",
  45795=>"00000100",
  45796=>"00000000",
  45797=>"11111100",
  45798=>"00000001",
  45799=>"11111110",
  45800=>"11111100",
  45801=>"00000001",
  45802=>"00000000",
  45803=>"00000001",
  45804=>"00000010",
  45805=>"00000000",
  45806=>"00000001",
  45807=>"11111111",
  45808=>"00000001",
  45809=>"00000000",
  45810=>"00000000",
  45811=>"00000010",
  45812=>"11111011",
  45813=>"00000001",
  45814=>"00000001",
  45815=>"11111110",
  45816=>"00000000",
  45817=>"00000100",
  45818=>"11111110",
  45819=>"00000000",
  45820=>"11111111",
  45821=>"00000010",
  45822=>"11111111",
  45823=>"00000001",
  45824=>"00000000",
  45825=>"00000001",
  45826=>"00000011",
  45827=>"00000011",
  45828=>"11111111",
  45829=>"00000000",
  45830=>"11111110",
  45831=>"00000000",
  45832=>"11111111",
  45833=>"11111111",
  45834=>"11111110",
  45835=>"00000011",
  45836=>"11111111",
  45837=>"00000001",
  45838=>"11111111",
  45839=>"00000101",
  45840=>"11111100",
  45841=>"11111111",
  45842=>"00000011",
  45843=>"11111101",
  45844=>"11111101",
  45845=>"00000001",
  45846=>"11111110",
  45847=>"11111111",
  45848=>"00000000",
  45849=>"11111110",
  45850=>"11111110",
  45851=>"11111111",
  45852=>"11111111",
  45853=>"11111100",
  45854=>"11111111",
  45855=>"00000010",
  45856=>"11111111",
  45857=>"11111110",
  45858=>"00000010",
  45859=>"11111110",
  45860=>"00000010",
  45861=>"00000010",
  45862=>"00000001",
  45863=>"11111110",
  45864=>"11111110",
  45865=>"00000001",
  45866=>"00000010",
  45867=>"00000001",
  45868=>"00000010",
  45869=>"00000010",
  45870=>"00000000",
  45871=>"00000000",
  45872=>"11111101",
  45873=>"11111111",
  45874=>"00000010",
  45875=>"11111101",
  45876=>"11111101",
  45877=>"11111101",
  45878=>"00000000",
  45879=>"00000000",
  45880=>"00000011",
  45881=>"11111111",
  45882=>"11111101",
  45883=>"00000011",
  45884=>"11111111",
  45885=>"00000000",
  45886=>"11111111",
  45887=>"00000010",
  45888=>"00000001",
  45889=>"00000010",
  45890=>"11111101",
  45891=>"00000001",
  45892=>"00000010",
  45893=>"00000001",
  45894=>"11111101",
  45895=>"11111110",
  45896=>"00000010",
  45897=>"11111111",
  45898=>"11111111",
  45899=>"11111110",
  45900=>"11111110",
  45901=>"00000010",
  45902=>"00000010",
  45903=>"11111110",
  45904=>"11111110",
  45905=>"00000011",
  45906=>"11111110",
  45907=>"11111111",
  45908=>"11111110",
  45909=>"11111101",
  45910=>"00000001",
  45911=>"11111101",
  45912=>"11111111",
  45913=>"00000010",
  45914=>"11111111",
  45915=>"00000010",
  45916=>"11111111",
  45917=>"11111111",
  45918=>"11111111",
  45919=>"11111111",
  45920=>"11111111",
  45921=>"00000010",
  45922=>"11111110",
  45923=>"11111111",
  45924=>"11111110",
  45925=>"11111111",
  45926=>"00000000",
  45927=>"00000011",
  45928=>"00000010",
  45929=>"00000010",
  45930=>"11111111",
  45931=>"11111110",
  45932=>"00000001",
  45933=>"11111100",
  45934=>"11111110",
  45935=>"00000011",
  45936=>"11111010",
  45937=>"00000000",
  45938=>"11111111",
  45939=>"11111110",
  45940=>"00000001",
  45941=>"11111110",
  45942=>"00000001",
  45943=>"00000010",
  45944=>"11111100",
  45945=>"00000001",
  45946=>"00000000",
  45947=>"00000000",
  45948=>"00000101",
  45949=>"11111101",
  45950=>"00000110",
  45951=>"11111111",
  45952=>"00000001",
  45953=>"11111100",
  45954=>"00000010",
  45955=>"11111101",
  45956=>"00000001",
  45957=>"00000001",
  45958=>"11111100",
  45959=>"00000000",
  45960=>"00000000",
  45961=>"11111110",
  45962=>"00000000",
  45963=>"11111111",
  45964=>"00000001",
  45965=>"00000010",
  45966=>"00000000",
  45967=>"11111111",
  45968=>"00000001",
  45969=>"00000000",
  45970=>"11111011",
  45971=>"11111111",
  45972=>"00000001",
  45973=>"00000000",
  45974=>"11111110",
  45975=>"00000010",
  45976=>"00000000",
  45977=>"00000001",
  45978=>"11111110",
  45979=>"00000101",
  45980=>"00000100",
  45981=>"11111111",
  45982=>"11111110",
  45983=>"00000000",
  45984=>"11111111",
  45985=>"11111101",
  45986=>"00000000",
  45987=>"11111110",
  45988=>"00000010",
  45989=>"00000000",
  45990=>"00000100",
  45991=>"11111110",
  45992=>"00000001",
  45993=>"11111101",
  45994=>"00000000",
  45995=>"11111110",
  45996=>"11111100",
  45997=>"00000001",
  45998=>"00000001",
  45999=>"00000000",
  46000=>"00000000",
  46001=>"00000000",
  46002=>"00000010",
  46003=>"11111111",
  46004=>"11111111",
  46005=>"11111100",
  46006=>"11111111",
  46007=>"11111110",
  46008=>"00000010",
  46009=>"00000001",
  46010=>"11111101",
  46011=>"00000001",
  46012=>"11111110",
  46013=>"11111110",
  46014=>"11111111",
  46015=>"00000001",
  46016=>"00000001",
  46017=>"00000001",
  46018=>"00000011",
  46019=>"11111110",
  46020=>"00000000",
  46021=>"11111111",
  46022=>"11111111",
  46023=>"11111111",
  46024=>"00000000",
  46025=>"11111110",
  46026=>"11111111",
  46027=>"00000010",
  46028=>"11111101",
  46029=>"11111101",
  46030=>"00000001",
  46031=>"00000000",
  46032=>"00000001",
  46033=>"11111110",
  46034=>"11111100",
  46035=>"11111111",
  46036=>"00000000",
  46037=>"00000001",
  46038=>"00000000",
  46039=>"11111101",
  46040=>"11111110",
  46041=>"00000010",
  46042=>"00000011",
  46043=>"11111110",
  46044=>"11111101",
  46045=>"11111110",
  46046=>"00000010",
  46047=>"11111111",
  46048=>"11111110",
  46049=>"00000001",
  46050=>"00000001",
  46051=>"00000010",
  46052=>"11111110",
  46053=>"11111110",
  46054=>"00000110",
  46055=>"00000011",
  46056=>"11111111",
  46057=>"11111111",
  46058=>"00000001",
  46059=>"11111110",
  46060=>"00000000",
  46061=>"11111101",
  46062=>"00001000",
  46063=>"00000000",
  46064=>"11111110",
  46065=>"00000100",
  46066=>"00000001",
  46067=>"00000011",
  46068=>"11111111",
  46069=>"11111111",
  46070=>"11111101",
  46071=>"11111111",
  46072=>"11111110",
  46073=>"11111110",
  46074=>"00000110",
  46075=>"00000001",
  46076=>"00000010",
  46077=>"00000101",
  46078=>"11111101",
  46079=>"00000000",
  46080=>"00000000",
  46081=>"00000010",
  46082=>"11111111",
  46083=>"00000011",
  46084=>"00000101",
  46085=>"11111101",
  46086=>"00000011",
  46087=>"00000011",
  46088=>"00000001",
  46089=>"00000000",
  46090=>"11111111",
  46091=>"11111101",
  46092=>"00000001",
  46093=>"11111111",
  46094=>"00000000",
  46095=>"11111110",
  46096=>"11111101",
  46097=>"11111110",
  46098=>"11111111",
  46099=>"00000000",
  46100=>"00000110",
  46101=>"00000001",
  46102=>"11111110",
  46103=>"11111111",
  46104=>"00000010",
  46105=>"00000011",
  46106=>"00000100",
  46107=>"11111110",
  46108=>"00000001",
  46109=>"11111101",
  46110=>"00000001",
  46111=>"00000001",
  46112=>"00000011",
  46113=>"11111111",
  46114=>"11111110",
  46115=>"00000000",
  46116=>"11111110",
  46117=>"11111101",
  46118=>"00000000",
  46119=>"00000010",
  46120=>"00000001",
  46121=>"00000000",
  46122=>"00000000",
  46123=>"00000010",
  46124=>"00000010",
  46125=>"11111110",
  46126=>"11111101",
  46127=>"11111101",
  46128=>"00000001",
  46129=>"11111111",
  46130=>"00000010",
  46131=>"00000010",
  46132=>"00000011",
  46133=>"00000010",
  46134=>"11111110",
  46135=>"00000001",
  46136=>"00000001",
  46137=>"11111100",
  46138=>"00000011",
  46139=>"11111111",
  46140=>"11111101",
  46141=>"00000001",
  46142=>"00000101",
  46143=>"00000010",
  46144=>"00000101",
  46145=>"11111101",
  46146=>"11111101",
  46147=>"11111101",
  46148=>"11111111",
  46149=>"00000000",
  46150=>"00000010",
  46151=>"11111101",
  46152=>"11111101",
  46153=>"00000000",
  46154=>"00000001",
  46155=>"00000010",
  46156=>"00000001",
  46157=>"00000111",
  46158=>"00000011",
  46159=>"00000000",
  46160=>"00000001",
  46161=>"00000000",
  46162=>"11111101",
  46163=>"11111110",
  46164=>"11111110",
  46165=>"11111101",
  46166=>"11111110",
  46167=>"00000010",
  46168=>"11111101",
  46169=>"11111101",
  46170=>"11111110",
  46171=>"11111101",
  46172=>"00000011",
  46173=>"00000001",
  46174=>"11111110",
  46175=>"00000001",
  46176=>"11111110",
  46177=>"11111110",
  46178=>"00000100",
  46179=>"00000010",
  46180=>"00000010",
  46181=>"00000011",
  46182=>"00000000",
  46183=>"00000001",
  46184=>"11111111",
  46185=>"00000100",
  46186=>"00000001",
  46187=>"11111111",
  46188=>"11111111",
  46189=>"00000000",
  46190=>"00000001",
  46191=>"00000010",
  46192=>"00000011",
  46193=>"00000100",
  46194=>"11111111",
  46195=>"11111111",
  46196=>"00000000",
  46197=>"11111110",
  46198=>"11111101",
  46199=>"11111111",
  46200=>"11111111",
  46201=>"11111110",
  46202=>"00000100",
  46203=>"11111111",
  46204=>"00000001",
  46205=>"00000100",
  46206=>"11111110",
  46207=>"00000010",
  46208=>"00000001",
  46209=>"00000101",
  46210=>"00000001",
  46211=>"00000000",
  46212=>"00000010",
  46213=>"00000000",
  46214=>"11111110",
  46215=>"11111111",
  46216=>"11111110",
  46217=>"00000001",
  46218=>"00000000",
  46219=>"00000101",
  46220=>"11111110",
  46221=>"11111111",
  46222=>"00000001",
  46223=>"11111101",
  46224=>"11111110",
  46225=>"00000010",
  46226=>"11111111",
  46227=>"00000010",
  46228=>"11111101",
  46229=>"11111101",
  46230=>"00000011",
  46231=>"11111111",
  46232=>"00000000",
  46233=>"00000000",
  46234=>"00000000",
  46235=>"11111110",
  46236=>"00000000",
  46237=>"00000011",
  46238=>"11111111",
  46239=>"11111110",
  46240=>"00000011",
  46241=>"00000100",
  46242=>"00000001",
  46243=>"00000000",
  46244=>"00000000",
  46245=>"11111100",
  46246=>"00000010",
  46247=>"00000000",
  46248=>"00000001",
  46249=>"00000000",
  46250=>"11111111",
  46251=>"11111111",
  46252=>"00000010",
  46253=>"00000011",
  46254=>"00000000",
  46255=>"11111110",
  46256=>"00000010",
  46257=>"00000000",
  46258=>"00000010",
  46259=>"00000100",
  46260=>"00000100",
  46261=>"00000000",
  46262=>"11111111",
  46263=>"00000010",
  46264=>"11111100",
  46265=>"11111111",
  46266=>"00000010",
  46267=>"11111111",
  46268=>"00000010",
  46269=>"11111110",
  46270=>"00000010",
  46271=>"00000001",
  46272=>"11111101",
  46273=>"00000000",
  46274=>"11111111",
  46275=>"00000010",
  46276=>"00000000",
  46277=>"11111111",
  46278=>"11111101",
  46279=>"00000000",
  46280=>"00000000",
  46281=>"00000001",
  46282=>"00000001",
  46283=>"11111111",
  46284=>"00000000",
  46285=>"00000010",
  46286=>"00000000",
  46287=>"11111110",
  46288=>"00000001",
  46289=>"11111110",
  46290=>"11111111",
  46291=>"00000000",
  46292=>"00000001",
  46293=>"11111111",
  46294=>"11111100",
  46295=>"00000001",
  46296=>"00000001",
  46297=>"00000100",
  46298=>"11111101",
  46299=>"11111111",
  46300=>"11111101",
  46301=>"00000010",
  46302=>"11111101",
  46303=>"11111110",
  46304=>"11111110",
  46305=>"11111111",
  46306=>"00000100",
  46307=>"00000001",
  46308=>"00000001",
  46309=>"11111111",
  46310=>"11111100",
  46311=>"11111100",
  46312=>"11111101",
  46313=>"00000000",
  46314=>"00000000",
  46315=>"00000001",
  46316=>"00000010",
  46317=>"11111100",
  46318=>"00000011",
  46319=>"11111111",
  46320=>"11111111",
  46321=>"11111111",
  46322=>"00000000",
  46323=>"00000100",
  46324=>"00000001",
  46325=>"00000000",
  46326=>"00000000",
  46327=>"11111110",
  46328=>"11111111",
  46329=>"00000001",
  46330=>"00000011",
  46331=>"00000001",
  46332=>"11111111",
  46333=>"00000010",
  46334=>"00000010",
  46335=>"00000001",
  46336=>"11111111",
  46337=>"00000011",
  46338=>"11111110",
  46339=>"00000011",
  46340=>"11111111",
  46341=>"00000000",
  46342=>"00000010",
  46343=>"11111101",
  46344=>"00000001",
  46345=>"11111101",
  46346=>"00000010",
  46347=>"11111101",
  46348=>"11111111",
  46349=>"00000010",
  46350=>"11111110",
  46351=>"00000000",
  46352=>"11111110",
  46353=>"00000011",
  46354=>"00000001",
  46355=>"00000001",
  46356=>"11111111",
  46357=>"11111101",
  46358=>"11111110",
  46359=>"00000101",
  46360=>"00000100",
  46361=>"00000011",
  46362=>"00000001",
  46363=>"11111111",
  46364=>"00000011",
  46365=>"00000001",
  46366=>"00000001",
  46367=>"11111101",
  46368=>"00000001",
  46369=>"11111110",
  46370=>"00000100",
  46371=>"00000101",
  46372=>"00000000",
  46373=>"00000001",
  46374=>"11111101",
  46375=>"11111101",
  46376=>"11111110",
  46377=>"00000101",
  46378=>"11111110",
  46379=>"00000000",
  46380=>"00000010",
  46381=>"11111111",
  46382=>"00000100",
  46383=>"00000001",
  46384=>"11111110",
  46385=>"11111111",
  46386=>"00000100",
  46387=>"00000010",
  46388=>"00000000",
  46389=>"00000011",
  46390=>"00000000",
  46391=>"11111111",
  46392=>"00000000",
  46393=>"11111101",
  46394=>"00000001",
  46395=>"00000000",
  46396=>"00000011",
  46397=>"00000000",
  46398=>"00000010",
  46399=>"00000001",
  46400=>"00000000",
  46401=>"00000000",
  46402=>"11111111",
  46403=>"11111110",
  46404=>"11111111",
  46405=>"00000000",
  46406=>"11111110",
  46407=>"11111111",
  46408=>"11111111",
  46409=>"11111111",
  46410=>"00000100",
  46411=>"11111111",
  46412=>"00000100",
  46413=>"00000010",
  46414=>"00000000",
  46415=>"11111100",
  46416=>"11111101",
  46417=>"00000011",
  46418=>"00000001",
  46419=>"00000000",
  46420=>"00000001",
  46421=>"11111110",
  46422=>"11111110",
  46423=>"00000000",
  46424=>"00000010",
  46425=>"00000010",
  46426=>"11111101",
  46427=>"11111111",
  46428=>"11111101",
  46429=>"00000100",
  46430=>"00000010",
  46431=>"11111111",
  46432=>"11111111",
  46433=>"11111111",
  46434=>"00000011",
  46435=>"00000011",
  46436=>"00000100",
  46437=>"11111101",
  46438=>"11111100",
  46439=>"00000000",
  46440=>"00000011",
  46441=>"00000100",
  46442=>"00000000",
  46443=>"11111111",
  46444=>"00000000",
  46445=>"00000110",
  46446=>"11111111",
  46447=>"00000001",
  46448=>"00000011",
  46449=>"11111101",
  46450=>"00000001",
  46451=>"00000001",
  46452=>"11111111",
  46453=>"00000001",
  46454=>"11111110",
  46455=>"00000010",
  46456=>"00000000",
  46457=>"00000000",
  46458=>"11111110",
  46459=>"00000000",
  46460=>"11111110",
  46461=>"11111110",
  46462=>"11111110",
  46463=>"00000010",
  46464=>"00000001",
  46465=>"00000001",
  46466=>"11111110",
  46467=>"00000001",
  46468=>"00000010",
  46469=>"00000000",
  46470=>"00000101",
  46471=>"00000001",
  46472=>"00000000",
  46473=>"00000010",
  46474=>"00000100",
  46475=>"00000101",
  46476=>"11111111",
  46477=>"11111111",
  46478=>"00000010",
  46479=>"11111101",
  46480=>"11111111",
  46481=>"00000000",
  46482=>"00000010",
  46483=>"00000010",
  46484=>"11111110",
  46485=>"00000100",
  46486=>"11111111",
  46487=>"00000010",
  46488=>"11111110",
  46489=>"00000001",
  46490=>"00000000",
  46491=>"00000001",
  46492=>"11111100",
  46493=>"00000000",
  46494=>"11111110",
  46495=>"00000010",
  46496=>"11111110",
  46497=>"11111111",
  46498=>"11111110",
  46499=>"00000000",
  46500=>"00000010",
  46501=>"11111101",
  46502=>"00000010",
  46503=>"11111110",
  46504=>"11111111",
  46505=>"00000000",
  46506=>"11111100",
  46507=>"00000001",
  46508=>"11111110",
  46509=>"00000100",
  46510=>"00000011",
  46511=>"00000000",
  46512=>"11111110",
  46513=>"00000101",
  46514=>"00000010",
  46515=>"11111111",
  46516=>"00000001",
  46517=>"00000010",
  46518=>"11111101",
  46519=>"00000010",
  46520=>"11111111",
  46521=>"00000000",
  46522=>"11111111",
  46523=>"11111110",
  46524=>"11111110",
  46525=>"11111111",
  46526=>"00000011",
  46527=>"00000000",
  46528=>"00000011",
  46529=>"11111101",
  46530=>"00000100",
  46531=>"00000000",
  46532=>"11111101",
  46533=>"00000010",
  46534=>"00000011",
  46535=>"00000001",
  46536=>"00000000",
  46537=>"00000001",
  46538=>"11111110",
  46539=>"00000010",
  46540=>"11111111",
  46541=>"11111110",
  46542=>"00000101",
  46543=>"00000001",
  46544=>"00000011",
  46545=>"00000101",
  46546=>"00000010",
  46547=>"00000001",
  46548=>"11111111",
  46549=>"11111101",
  46550=>"00000011",
  46551=>"00000010",
  46552=>"00000000",
  46553=>"00000100",
  46554=>"00000010",
  46555=>"11111111",
  46556=>"11111111",
  46557=>"00000001",
  46558=>"11111111",
  46559=>"11111101",
  46560=>"00000000",
  46561=>"11111111",
  46562=>"00000001",
  46563=>"00000001",
  46564=>"11111110",
  46565=>"11111111",
  46566=>"11111110",
  46567=>"00000001",
  46568=>"00000010",
  46569=>"00000000",
  46570=>"11111110",
  46571=>"00000010",
  46572=>"11111111",
  46573=>"00000001",
  46574=>"00000010",
  46575=>"00000000",
  46576=>"11111111",
  46577=>"00000100",
  46578=>"11111101",
  46579=>"00000010",
  46580=>"00000010",
  46581=>"00000010",
  46582=>"11111101",
  46583=>"00000010",
  46584=>"00000000",
  46585=>"11111101",
  46586=>"11111101",
  46587=>"00000010",
  46588=>"00000001",
  46589=>"11111111",
  46590=>"11111111",
  46591=>"11111110",
  46592=>"00000000",
  46593=>"00000001",
  46594=>"00000001",
  46595=>"00000010",
  46596=>"00000110",
  46597=>"00000101",
  46598=>"11111111",
  46599=>"00000010",
  46600=>"00000010",
  46601=>"00000010",
  46602=>"00000011",
  46603=>"00000100",
  46604=>"11111100",
  46605=>"00000001",
  46606=>"00000001",
  46607=>"11111110",
  46608=>"00000000",
  46609=>"00000001",
  46610=>"11111101",
  46611=>"11111110",
  46612=>"00000001",
  46613=>"00000001",
  46614=>"11111111",
  46615=>"00000010",
  46616=>"00000001",
  46617=>"00000001",
  46618=>"00000010",
  46619=>"11111110",
  46620=>"00000010",
  46621=>"00000011",
  46622=>"00000000",
  46623=>"11111101",
  46624=>"11111111",
  46625=>"11111111",
  46626=>"00000010",
  46627=>"00000100",
  46628=>"11111101",
  46629=>"00000000",
  46630=>"11111101",
  46631=>"00000000",
  46632=>"11111101",
  46633=>"11111101",
  46634=>"11111111",
  46635=>"11111110",
  46636=>"00000010",
  46637=>"00000010",
  46638=>"00000010",
  46639=>"00000000",
  46640=>"11111111",
  46641=>"00000100",
  46642=>"00000001",
  46643=>"00000010",
  46644=>"00000010",
  46645=>"11111111",
  46646=>"00000010",
  46647=>"11111101",
  46648=>"00000010",
  46649=>"00000001",
  46650=>"11111111",
  46651=>"00000010",
  46652=>"00000001",
  46653=>"00000001",
  46654=>"00000101",
  46655=>"11111111",
  46656=>"00000001",
  46657=>"00000011",
  46658=>"00000011",
  46659=>"11111101",
  46660=>"11111110",
  46661=>"00000100",
  46662=>"11111110",
  46663=>"11111111",
  46664=>"11111101",
  46665=>"00000010",
  46666=>"11111111",
  46667=>"00000100",
  46668=>"00000001",
  46669=>"11111101",
  46670=>"11111110",
  46671=>"11111111",
  46672=>"00000011",
  46673=>"00000000",
  46674=>"11111101",
  46675=>"00000000",
  46676=>"11111110",
  46677=>"00000010",
  46678=>"00000000",
  46679=>"00000011",
  46680=>"00000001",
  46681=>"00000010",
  46682=>"00000000",
  46683=>"11111111",
  46684=>"11111111",
  46685=>"00000001",
  46686=>"11111111",
  46687=>"11111111",
  46688=>"00000001",
  46689=>"11111110",
  46690=>"00000000",
  46691=>"00000000",
  46692=>"11111110",
  46693=>"11111100",
  46694=>"00000010",
  46695=>"11111101",
  46696=>"00000100",
  46697=>"11111110",
  46698=>"11111110",
  46699=>"00000010",
  46700=>"11111111",
  46701=>"11111111",
  46702=>"11111101",
  46703=>"00000000",
  46704=>"00000001",
  46705=>"11111110",
  46706=>"00000011",
  46707=>"11111111",
  46708=>"11111110",
  46709=>"11111111",
  46710=>"11111110",
  46711=>"00000001",
  46712=>"11111111",
  46713=>"00000001",
  46714=>"00000100",
  46715=>"00000001",
  46716=>"11111111",
  46717=>"11111110",
  46718=>"11111110",
  46719=>"00000011",
  46720=>"00000000",
  46721=>"00000001",
  46722=>"11111111",
  46723=>"00000011",
  46724=>"00000010",
  46725=>"11111110",
  46726=>"00000000",
  46727=>"00000100",
  46728=>"00000001",
  46729=>"11111101",
  46730=>"00000001",
  46731=>"00000011",
  46732=>"00000010",
  46733=>"00000001",
  46734=>"11111101",
  46735=>"11111101",
  46736=>"00000001",
  46737=>"11111101",
  46738=>"11111111",
  46739=>"00000001",
  46740=>"00000001",
  46741=>"00000001",
  46742=>"11111110",
  46743=>"00000001",
  46744=>"11111111",
  46745=>"11111101",
  46746=>"11111110",
  46747=>"00000011",
  46748=>"11111110",
  46749=>"11111111",
  46750=>"00000000",
  46751=>"00000011",
  46752=>"11111111",
  46753=>"11111101",
  46754=>"00000011",
  46755=>"11111101",
  46756=>"11111111",
  46757=>"00000011",
  46758=>"00000101",
  46759=>"00000010",
  46760=>"00000101",
  46761=>"11111111",
  46762=>"00000010",
  46763=>"00000000",
  46764=>"11111101",
  46765=>"11111101",
  46766=>"00000001",
  46767=>"00000010",
  46768=>"11111101",
  46769=>"11111111",
  46770=>"00000000",
  46771=>"00000000",
  46772=>"00000101",
  46773=>"00000101",
  46774=>"11111101",
  46775=>"00000000",
  46776=>"00000011",
  46777=>"11111111",
  46778=>"11111111",
  46779=>"00000001",
  46780=>"00000001",
  46781=>"00000001",
  46782=>"11111111",
  46783=>"11111101",
  46784=>"00000011",
  46785=>"11111100",
  46786=>"11111101",
  46787=>"11111110",
  46788=>"00000001",
  46789=>"00000011",
  46790=>"11111110",
  46791=>"00000001",
  46792=>"11111111",
  46793=>"00000001",
  46794=>"00000010",
  46795=>"00000000",
  46796=>"00000010",
  46797=>"11111110",
  46798=>"11111101",
  46799=>"00000001",
  46800=>"11111111",
  46801=>"00000000",
  46802=>"11111110",
  46803=>"11111110",
  46804=>"11111111",
  46805=>"11111111",
  46806=>"00000010",
  46807=>"11111110",
  46808=>"00000001",
  46809=>"00000010",
  46810=>"00000010",
  46811=>"00000001",
  46812=>"00000001",
  46813=>"11111110",
  46814=>"00000000",
  46815=>"00000001",
  46816=>"11111110",
  46817=>"00000000",
  46818=>"00000011",
  46819=>"00000010",
  46820=>"00000000",
  46821=>"11111101",
  46822=>"00000010",
  46823=>"00000000",
  46824=>"00000010",
  46825=>"11111101",
  46826=>"11111100",
  46827=>"00000001",
  46828=>"11111110",
  46829=>"11111101",
  46830=>"11111111",
  46831=>"00000001",
  46832=>"00000010",
  46833=>"00000010",
  46834=>"00000001",
  46835=>"11111101",
  46836=>"11111101",
  46837=>"11111101",
  46838=>"00000000",
  46839=>"00000001",
  46840=>"11111111",
  46841=>"11111111",
  46842=>"11111110",
  46843=>"11111110",
  46844=>"00000010",
  46845=>"00000011",
  46846=>"00000100",
  46847=>"00000001",
  46848=>"11111100",
  46849=>"00000001",
  46850=>"00000100",
  46851=>"00000001",
  46852=>"00000110",
  46853=>"11111111",
  46854=>"00000010",
  46855=>"00000010",
  46856=>"00000010",
  46857=>"00000001",
  46858=>"11111111",
  46859=>"00000000",
  46860=>"00000010",
  46861=>"00000110",
  46862=>"11111101",
  46863=>"11111111",
  46864=>"00000010",
  46865=>"00000010",
  46866=>"00000001",
  46867=>"11111100",
  46868=>"11111110",
  46869=>"11111101",
  46870=>"00000010",
  46871=>"00000000",
  46872=>"11111111",
  46873=>"11111101",
  46874=>"00000010",
  46875=>"11111110",
  46876=>"00000011",
  46877=>"00000010",
  46878=>"11111110",
  46879=>"00000000",
  46880=>"00000010",
  46881=>"00000010",
  46882=>"11111110",
  46883=>"00000001",
  46884=>"11111111",
  46885=>"00000010",
  46886=>"11111111",
  46887=>"00000011",
  46888=>"11111110",
  46889=>"00000100",
  46890=>"11111111",
  46891=>"11111101",
  46892=>"00000001",
  46893=>"00000001",
  46894=>"00000000",
  46895=>"00000000",
  46896=>"11111101",
  46897=>"00000100",
  46898=>"00000010",
  46899=>"00000000",
  46900=>"11111110",
  46901=>"00000000",
  46902=>"00000011",
  46903=>"00000011",
  46904=>"11111111",
  46905=>"00000010",
  46906=>"00000011",
  46907=>"11111111",
  46908=>"00000100",
  46909=>"11111101",
  46910=>"00000010",
  46911=>"11111110",
  46912=>"00000111",
  46913=>"00000010",
  46914=>"00000001",
  46915=>"11111110",
  46916=>"00000001",
  46917=>"11111111",
  46918=>"11111110",
  46919=>"11111101",
  46920=>"11111100",
  46921=>"00000001",
  46922=>"11111110",
  46923=>"00000010",
  46924=>"00000011",
  46925=>"00000000",
  46926=>"00000010",
  46927=>"11111101",
  46928=>"11111111",
  46929=>"11111110",
  46930=>"00000000",
  46931=>"00000000",
  46932=>"00000000",
  46933=>"11111111",
  46934=>"11111111",
  46935=>"11111101",
  46936=>"11111110",
  46937=>"11111110",
  46938=>"00000000",
  46939=>"00000001",
  46940=>"11111110",
  46941=>"11111111",
  46942=>"00000101",
  46943=>"00000000",
  46944=>"00000000",
  46945=>"00000001",
  46946=>"00000001",
  46947=>"11111110",
  46948=>"11111110",
  46949=>"00000001",
  46950=>"11111110",
  46951=>"11111111",
  46952=>"11111110",
  46953=>"11111110",
  46954=>"11111110",
  46955=>"11111110",
  46956=>"00000001",
  46957=>"00000001",
  46958=>"11111101",
  46959=>"11111101",
  46960=>"00000000",
  46961=>"00000011",
  46962=>"00000001",
  46963=>"11111110",
  46964=>"00000000",
  46965=>"00000011",
  46966=>"00000011",
  46967=>"00000011",
  46968=>"11111110",
  46969=>"11111110",
  46970=>"00000001",
  46971=>"00000000",
  46972=>"00000010",
  46973=>"00000000",
  46974=>"00000000",
  46975=>"00000010",
  46976=>"11111111",
  46977=>"11111110",
  46978=>"11111100",
  46979=>"00000000",
  46980=>"11111110",
  46981=>"11111101",
  46982=>"00000000",
  46983=>"11111111",
  46984=>"11111111",
  46985=>"00000110",
  46986=>"00000000",
  46987=>"00000011",
  46988=>"00000000",
  46989=>"00000010",
  46990=>"11111101",
  46991=>"11111110",
  46992=>"00000010",
  46993=>"00000100",
  46994=>"00000011",
  46995=>"00000000",
  46996=>"00000001",
  46997=>"11111111",
  46998=>"11111111",
  46999=>"00000010",
  47000=>"11111111",
  47001=>"00000100",
  47002=>"11111101",
  47003=>"11111101",
  47004=>"00000000",
  47005=>"00000011",
  47006=>"11111101",
  47007=>"00000001",
  47008=>"11111100",
  47009=>"11111110",
  47010=>"11111101",
  47011=>"11111110",
  47012=>"11111110",
  47013=>"00000100",
  47014=>"11111110",
  47015=>"00000000",
  47016=>"00000011",
  47017=>"00000011",
  47018=>"11111110",
  47019=>"11111111",
  47020=>"00000001",
  47021=>"11111111",
  47022=>"00000011",
  47023=>"11111111",
  47024=>"11111110",
  47025=>"00000001",
  47026=>"00000001",
  47027=>"00000100",
  47028=>"00000011",
  47029=>"00000010",
  47030=>"00000001",
  47031=>"00000000",
  47032=>"00000100",
  47033=>"00000001",
  47034=>"11111111",
  47035=>"00000011",
  47036=>"00000010",
  47037=>"11111111",
  47038=>"00000000",
  47039=>"00000010",
  47040=>"11111111",
  47041=>"00000001",
  47042=>"00000011",
  47043=>"00000010",
  47044=>"00000010",
  47045=>"11111111",
  47046=>"11111110",
  47047=>"00000001",
  47048=>"00000011",
  47049=>"11111111",
  47050=>"11111101",
  47051=>"00000001",
  47052=>"00000011",
  47053=>"00000011",
  47054=>"11111101",
  47055=>"11111110",
  47056=>"00000000",
  47057=>"00000100",
  47058=>"11111100",
  47059=>"11111111",
  47060=>"00000010",
  47061=>"00000000",
  47062=>"00000001",
  47063=>"11111110",
  47064=>"00000001",
  47065=>"11111110",
  47066=>"11111110",
  47067=>"11111110",
  47068=>"00000010",
  47069=>"00000010",
  47070=>"00000001",
  47071=>"11111110",
  47072=>"00000000",
  47073=>"00000001",
  47074=>"00000001",
  47075=>"11111110",
  47076=>"00000010",
  47077=>"11111101",
  47078=>"00000001",
  47079=>"00000110",
  47080=>"00000000",
  47081=>"00000010",
  47082=>"11111111",
  47083=>"00000001",
  47084=>"00000010",
  47085=>"11111111",
  47086=>"00000100",
  47087=>"00000000",
  47088=>"11111111",
  47089=>"00000001",
  47090=>"00000101",
  47091=>"00000011",
  47092=>"00000001",
  47093=>"00000010",
  47094=>"11111101",
  47095=>"11111101",
  47096=>"00000100",
  47097=>"00000001",
  47098=>"11111110",
  47099=>"00000001",
  47100=>"11111110",
  47101=>"11111110",
  47102=>"00000100",
  47103=>"00000000",
  47104=>"00000011",
  47105=>"00000010",
  47106=>"00000010",
  47107=>"00000001",
  47108=>"00000010",
  47109=>"00000000",
  47110=>"00000000",
  47111=>"11111111",
  47112=>"00000000",
  47113=>"11111101",
  47114=>"00000011",
  47115=>"11111110",
  47116=>"11111111",
  47117=>"00000000",
  47118=>"00000001",
  47119=>"00000000",
  47120=>"11111111",
  47121=>"00000010",
  47122=>"00000001",
  47123=>"00000011",
  47124=>"11111111",
  47125=>"00000011",
  47126=>"11111101",
  47127=>"11111110",
  47128=>"11111111",
  47129=>"11111111",
  47130=>"00000010",
  47131=>"11111111",
  47132=>"00000001",
  47133=>"00000001",
  47134=>"00000001",
  47135=>"00000000",
  47136=>"11111111",
  47137=>"00000000",
  47138=>"11111111",
  47139=>"11111110",
  47140=>"11111110",
  47141=>"11111111",
  47142=>"00000001",
  47143=>"11111111",
  47144=>"11111101",
  47145=>"11111111",
  47146=>"00000011",
  47147=>"00000000",
  47148=>"11111101",
  47149=>"11111111",
  47150=>"11111110",
  47151=>"11111111",
  47152=>"11111110",
  47153=>"00000001",
  47154=>"00000001",
  47155=>"00000010",
  47156=>"00000000",
  47157=>"00000001",
  47158=>"00000001",
  47159=>"00000001",
  47160=>"11111100",
  47161=>"00000000",
  47162=>"11111110",
  47163=>"00000010",
  47164=>"11111111",
  47165=>"11111111",
  47166=>"00000000",
  47167=>"00000001",
  47168=>"00000010",
  47169=>"00000010",
  47170=>"11111101",
  47171=>"11111101",
  47172=>"00000010",
  47173=>"00000010",
  47174=>"00000001",
  47175=>"11111101",
  47176=>"11111111",
  47177=>"11111110",
  47178=>"11111111",
  47179=>"11111110",
  47180=>"00000001",
  47181=>"00000001",
  47182=>"00000001",
  47183=>"00000001",
  47184=>"00000000",
  47185=>"11111111",
  47186=>"11111110",
  47187=>"00000100",
  47188=>"00000010",
  47189=>"11111101",
  47190=>"00000101",
  47191=>"11111101",
  47192=>"00000001",
  47193=>"11111111",
  47194=>"00000001",
  47195=>"00000000",
  47196=>"00000000",
  47197=>"11111110",
  47198=>"00000011",
  47199=>"11111111",
  47200=>"00000110",
  47201=>"11111101",
  47202=>"11111110",
  47203=>"00000010",
  47204=>"00000010",
  47205=>"00000010",
  47206=>"00000010",
  47207=>"11111101",
  47208=>"11111110",
  47209=>"11111111",
  47210=>"11111111",
  47211=>"00000010",
  47212=>"11111101",
  47213=>"11111110",
  47214=>"00000000",
  47215=>"00000000",
  47216=>"00000001",
  47217=>"00000011",
  47218=>"00000000",
  47219=>"00000000",
  47220=>"11111101",
  47221=>"11111111",
  47222=>"00000000",
  47223=>"00000001",
  47224=>"00000010",
  47225=>"11111111",
  47226=>"00000011",
  47227=>"00000011",
  47228=>"11111111",
  47229=>"00000010",
  47230=>"11111111",
  47231=>"11111111",
  47232=>"11111110",
  47233=>"11111111",
  47234=>"11111111",
  47235=>"00000010",
  47236=>"11111111",
  47237=>"11111110",
  47238=>"11111110",
  47239=>"11111111",
  47240=>"00000010",
  47241=>"00000001",
  47242=>"11111111",
  47243=>"00000011",
  47244=>"00000100",
  47245=>"11111101",
  47246=>"11111111",
  47247=>"00000001",
  47248=>"11111110",
  47249=>"00000010",
  47250=>"00000000",
  47251=>"11111101",
  47252=>"11111111",
  47253=>"11111110",
  47254=>"00000101",
  47255=>"00000100",
  47256=>"11111111",
  47257=>"00000010",
  47258=>"00000001",
  47259=>"00000010",
  47260=>"00000010",
  47261=>"11111101",
  47262=>"00000000",
  47263=>"00000100",
  47264=>"00000000",
  47265=>"00000010",
  47266=>"00000001",
  47267=>"11111111",
  47268=>"11111110",
  47269=>"00000010",
  47270=>"00000001",
  47271=>"00000010",
  47272=>"00000001",
  47273=>"11111101",
  47274=>"00000001",
  47275=>"11111111",
  47276=>"11111110",
  47277=>"11111110",
  47278=>"11111111",
  47279=>"11111111",
  47280=>"11111110",
  47281=>"00000000",
  47282=>"00000010",
  47283=>"11111111",
  47284=>"00000000",
  47285=>"00000000",
  47286=>"00000000",
  47287=>"11111101",
  47288=>"11111110",
  47289=>"11111111",
  47290=>"11111101",
  47291=>"00000000",
  47292=>"11111111",
  47293=>"00000000",
  47294=>"11111111",
  47295=>"11111101",
  47296=>"11111111",
  47297=>"11111110",
  47298=>"11111101",
  47299=>"00000010",
  47300=>"00000100",
  47301=>"00000001",
  47302=>"00000000",
  47303=>"00000000",
  47304=>"00000011",
  47305=>"11111110",
  47306=>"11111101",
  47307=>"11111110",
  47308=>"00000010",
  47309=>"11111110",
  47310=>"00000001",
  47311=>"00000000",
  47312=>"00000001",
  47313=>"11111101",
  47314=>"11111101",
  47315=>"11111111",
  47316=>"00000001",
  47317=>"11111111",
  47318=>"11111110",
  47319=>"11111110",
  47320=>"00000001",
  47321=>"11111111",
  47322=>"00000000",
  47323=>"00000011",
  47324=>"00000100",
  47325=>"00000000",
  47326=>"00000010",
  47327=>"00000000",
  47328=>"00000010",
  47329=>"11111101",
  47330=>"00000100",
  47331=>"00000010",
  47332=>"00000011",
  47333=>"00000000",
  47334=>"00000000",
  47335=>"00000011",
  47336=>"00000010",
  47337=>"11111110",
  47338=>"11111110",
  47339=>"11111111",
  47340=>"00000000",
  47341=>"00000011",
  47342=>"00000011",
  47343=>"11111110",
  47344=>"00000010",
  47345=>"00000010",
  47346=>"00000001",
  47347=>"00000000",
  47348=>"11111111",
  47349=>"00000001",
  47350=>"00000001",
  47351=>"00000010",
  47352=>"11111110",
  47353=>"11111110",
  47354=>"00000010",
  47355=>"11111111",
  47356=>"00000010",
  47357=>"00000010",
  47358=>"11111111",
  47359=>"00000001",
  47360=>"00000100",
  47361=>"00000000",
  47362=>"00000000",
  47363=>"00000010",
  47364=>"11111110",
  47365=>"00000001",
  47366=>"00000011",
  47367=>"00000011",
  47368=>"00000011",
  47369=>"11111111",
  47370=>"11111110",
  47371=>"11111111",
  47372=>"00000011",
  47373=>"00000011",
  47374=>"11111111",
  47375=>"00000000",
  47376=>"00000001",
  47377=>"00000010",
  47378=>"11111111",
  47379=>"11111101",
  47380=>"00000001",
  47381=>"11111110",
  47382=>"00000011",
  47383=>"11111101",
  47384=>"11111111",
  47385=>"00000001",
  47386=>"00000000",
  47387=>"11111111",
  47388=>"00000001",
  47389=>"00000011",
  47390=>"11111110",
  47391=>"00000000",
  47392=>"11111111",
  47393=>"00000000",
  47394=>"00000000",
  47395=>"00000000",
  47396=>"00000000",
  47397=>"00000010",
  47398=>"11111111",
  47399=>"00000010",
  47400=>"11111111",
  47401=>"00000000",
  47402=>"00000100",
  47403=>"11111110",
  47404=>"00000010",
  47405=>"11111111",
  47406=>"00000010",
  47407=>"11111111",
  47408=>"00000000",
  47409=>"00000000",
  47410=>"00000000",
  47411=>"11111101",
  47412=>"11111111",
  47413=>"11111111",
  47414=>"11111111",
  47415=>"00000100",
  47416=>"11111110",
  47417=>"00000011",
  47418=>"11111110",
  47419=>"00000000",
  47420=>"11111111",
  47421=>"11111110",
  47422=>"11111111",
  47423=>"00000010",
  47424=>"00000001",
  47425=>"00000010",
  47426=>"11111110",
  47427=>"00000001",
  47428=>"11111111",
  47429=>"00000001",
  47430=>"11111111",
  47431=>"00000001",
  47432=>"11111110",
  47433=>"00000000",
  47434=>"11111101",
  47435=>"00000001",
  47436=>"00000001",
  47437=>"11111101",
  47438=>"11111101",
  47439=>"11111111",
  47440=>"11111111",
  47441=>"11111111",
  47442=>"11111101",
  47443=>"00000001",
  47444=>"00000001",
  47445=>"00000001",
  47446=>"00000000",
  47447=>"00000001",
  47448=>"00000001",
  47449=>"00000001",
  47450=>"00000001",
  47451=>"11111111",
  47452=>"00000110",
  47453=>"11111101",
  47454=>"11111101",
  47455=>"00000001",
  47456=>"11111110",
  47457=>"11111111",
  47458=>"11111110",
  47459=>"00000000",
  47460=>"11111110",
  47461=>"00000010",
  47462=>"11111110",
  47463=>"11111111",
  47464=>"11111110",
  47465=>"11111111",
  47466=>"11111101",
  47467=>"11111101",
  47468=>"11111111",
  47469=>"11111110",
  47470=>"11111101",
  47471=>"00000001",
  47472=>"00000000",
  47473=>"11111111",
  47474=>"11111111",
  47475=>"11111110",
  47476=>"00000010",
  47477=>"11111101",
  47478=>"11111110",
  47479=>"00000001",
  47480=>"00000001",
  47481=>"00000010",
  47482=>"11111101",
  47483=>"00000001",
  47484=>"00000011",
  47485=>"11111110",
  47486=>"11111111",
  47487=>"00000011",
  47488=>"00000010",
  47489=>"00000000",
  47490=>"11111111",
  47491=>"00000001",
  47492=>"11111111",
  47493=>"00000000",
  47494=>"11111110",
  47495=>"00000000",
  47496=>"00000011",
  47497=>"11111101",
  47498=>"00000000",
  47499=>"11111101",
  47500=>"11111111",
  47501=>"00000010",
  47502=>"00000001",
  47503=>"00000001",
  47504=>"11111110",
  47505=>"11111110",
  47506=>"11111110",
  47507=>"00000011",
  47508=>"11111110",
  47509=>"11111110",
  47510=>"00000011",
  47511=>"00000010",
  47512=>"11111101",
  47513=>"00000000",
  47514=>"00000010",
  47515=>"11111101",
  47516=>"00000010",
  47517=>"11111101",
  47518=>"11111101",
  47519=>"00000001",
  47520=>"00000001",
  47521=>"00000000",
  47522=>"11111111",
  47523=>"00000100",
  47524=>"11111101",
  47525=>"00000001",
  47526=>"00000000",
  47527=>"00000001",
  47528=>"00000010",
  47529=>"11111111",
  47530=>"11111110",
  47531=>"00000100",
  47532=>"11111110",
  47533=>"00000001",
  47534=>"00000010",
  47535=>"11111111",
  47536=>"11111101",
  47537=>"00000010",
  47538=>"11111110",
  47539=>"11111111",
  47540=>"11111101",
  47541=>"00000001",
  47542=>"11111111",
  47543=>"11111110",
  47544=>"00000001",
  47545=>"00000100",
  47546=>"00000000",
  47547=>"00000001",
  47548=>"00000011",
  47549=>"11111111",
  47550=>"11111111",
  47551=>"00000000",
  47552=>"00000011",
  47553=>"00000001",
  47554=>"11111111",
  47555=>"00000010",
  47556=>"00000000",
  47557=>"11111101",
  47558=>"00000001",
  47559=>"11111100",
  47560=>"00000000",
  47561=>"00000010",
  47562=>"11111101",
  47563=>"11111111",
  47564=>"00000001",
  47565=>"00000001",
  47566=>"00000000",
  47567=>"00000000",
  47568=>"00000001",
  47569=>"00000010",
  47570=>"11111101",
  47571=>"00000001",
  47572=>"00000011",
  47573=>"11111111",
  47574=>"11111110",
  47575=>"11111111",
  47576=>"11111110",
  47577=>"00000001",
  47578=>"11111110",
  47579=>"11111110",
  47580=>"11111100",
  47581=>"11111110",
  47582=>"00000011",
  47583=>"00000010",
  47584=>"11111101",
  47585=>"11111111",
  47586=>"00000010",
  47587=>"00000000",
  47588=>"00000000",
  47589=>"00000001",
  47590=>"11111111",
  47591=>"00000010",
  47592=>"00000010",
  47593=>"00000000",
  47594=>"11111111",
  47595=>"00000001",
  47596=>"11111110",
  47597=>"00000100",
  47598=>"11111110",
  47599=>"11111101",
  47600=>"00000010",
  47601=>"11111110",
  47602=>"00000010",
  47603=>"00000000",
  47604=>"11111111",
  47605=>"11111110",
  47606=>"00000100",
  47607=>"00000001",
  47608=>"00000010",
  47609=>"11111101",
  47610=>"00000100",
  47611=>"00000011",
  47612=>"11111111",
  47613=>"00000000",
  47614=>"00000011",
  47615=>"00000000",
  47616=>"00000010",
  47617=>"00000001",
  47618=>"11111101",
  47619=>"11111110",
  47620=>"11111110",
  47621=>"11111111",
  47622=>"11111110",
  47623=>"00000010",
  47624=>"11111101",
  47625=>"11111111",
  47626=>"11111111",
  47627=>"11111111",
  47628=>"11111110",
  47629=>"00000000",
  47630=>"00000000",
  47631=>"11111101",
  47632=>"11111111",
  47633=>"11111110",
  47634=>"00000010",
  47635=>"00000001",
  47636=>"11111111",
  47637=>"00000000",
  47638=>"00000000",
  47639=>"11111101",
  47640=>"00000010",
  47641=>"11111101",
  47642=>"00000010",
  47643=>"11111110",
  47644=>"00000010",
  47645=>"11111111",
  47646=>"00000010",
  47647=>"00000010",
  47648=>"00000001",
  47649=>"00000011",
  47650=>"00000011",
  47651=>"11111111",
  47652=>"00000000",
  47653=>"11111110",
  47654=>"00000000",
  47655=>"11111111",
  47656=>"00000000",
  47657=>"00000010",
  47658=>"00000001",
  47659=>"00000100",
  47660=>"11111110",
  47661=>"11111110",
  47662=>"11111110",
  47663=>"00000000",
  47664=>"11111111",
  47665=>"00000011",
  47666=>"11111111",
  47667=>"00000010",
  47668=>"11111111",
  47669=>"00000001",
  47670=>"11111101",
  47671=>"11111110",
  47672=>"00000010",
  47673=>"00000011",
  47674=>"11111111",
  47675=>"00000001",
  47676=>"00000000",
  47677=>"11111110",
  47678=>"00000000",
  47679=>"00000010",
  47680=>"11111110",
  47681=>"11111110",
  47682=>"00000000",
  47683=>"00000001",
  47684=>"00000000",
  47685=>"00000001",
  47686=>"00000101",
  47687=>"11111110",
  47688=>"00000000",
  47689=>"00000001",
  47690=>"00000011",
  47691=>"00000010",
  47692=>"00000011",
  47693=>"00000010",
  47694=>"00000011",
  47695=>"00000000",
  47696=>"00000001",
  47697=>"11111110",
  47698=>"11111111",
  47699=>"11111101",
  47700=>"00000011",
  47701=>"11111111",
  47702=>"11111110",
  47703=>"00000001",
  47704=>"11111110",
  47705=>"00000011",
  47706=>"00000001",
  47707=>"00000001",
  47708=>"00000001",
  47709=>"11111110",
  47710=>"11111111",
  47711=>"00000010",
  47712=>"00000001",
  47713=>"00000001",
  47714=>"00000000",
  47715=>"11111110",
  47716=>"11111111",
  47717=>"00000000",
  47718=>"11111110",
  47719=>"00000001",
  47720=>"11111110",
  47721=>"11111110",
  47722=>"11111101",
  47723=>"11111101",
  47724=>"11111110",
  47725=>"11111101",
  47726=>"00000010",
  47727=>"00000000",
  47728=>"11111110",
  47729=>"00000011",
  47730=>"00000000",
  47731=>"11111111",
  47732=>"11111111",
  47733=>"11111110",
  47734=>"11111111",
  47735=>"00000000",
  47736=>"00000001",
  47737=>"00000001",
  47738=>"11111110",
  47739=>"11111110",
  47740=>"00000010",
  47741=>"00000011",
  47742=>"11111111",
  47743=>"00000000",
  47744=>"00000000",
  47745=>"00000011",
  47746=>"00000000",
  47747=>"00000001",
  47748=>"00000010",
  47749=>"00000010",
  47750=>"11111110",
  47751=>"00000000",
  47752=>"00000001",
  47753=>"11111111",
  47754=>"00000001",
  47755=>"00000001",
  47756=>"11111111",
  47757=>"11111111",
  47758=>"11111111",
  47759=>"00000001",
  47760=>"11111110",
  47761=>"11111111",
  47762=>"00000101",
  47763=>"00000000",
  47764=>"11111110",
  47765=>"11111101",
  47766=>"11111110",
  47767=>"00000100",
  47768=>"11111100",
  47769=>"00000001",
  47770=>"11111111",
  47771=>"00000010",
  47772=>"11111111",
  47773=>"00000100",
  47774=>"11111111",
  47775=>"00000001",
  47776=>"00000010",
  47777=>"11111101",
  47778=>"11111110",
  47779=>"11111111",
  47780=>"00000001",
  47781=>"00000001",
  47782=>"00000010",
  47783=>"11111111",
  47784=>"11111101",
  47785=>"00000011",
  47786=>"11111110",
  47787=>"00000000",
  47788=>"00000100",
  47789=>"00000001",
  47790=>"11111111",
  47791=>"11111110",
  47792=>"11111101",
  47793=>"11111110",
  47794=>"00000001",
  47795=>"11111111",
  47796=>"00000000",
  47797=>"00000010",
  47798=>"11111110",
  47799=>"11111111",
  47800=>"11111111",
  47801=>"00000001",
  47802=>"11111111",
  47803=>"00000001",
  47804=>"00000001",
  47805=>"00000011",
  47806=>"00000011",
  47807=>"00000000",
  47808=>"00000010",
  47809=>"00000010",
  47810=>"00000001",
  47811=>"00000000",
  47812=>"00000000",
  47813=>"00000001",
  47814=>"11111101",
  47815=>"11111111",
  47816=>"11111110",
  47817=>"11111110",
  47818=>"00000001",
  47819=>"11111110",
  47820=>"11111101",
  47821=>"11111110",
  47822=>"11111111",
  47823=>"11111101",
  47824=>"00000000",
  47825=>"11111110",
  47826=>"00000000",
  47827=>"00000001",
  47828=>"11111111",
  47829=>"00000011",
  47830=>"11111111",
  47831=>"00000000",
  47832=>"11111111",
  47833=>"00000010",
  47834=>"11111111",
  47835=>"11111101",
  47836=>"00000000",
  47837=>"00000001",
  47838=>"00000001",
  47839=>"11111111",
  47840=>"00000000",
  47841=>"11111111",
  47842=>"11111101",
  47843=>"00000011",
  47844=>"00000011",
  47845=>"11111110",
  47846=>"11111110",
  47847=>"11111110",
  47848=>"11111111",
  47849=>"11111110",
  47850=>"11111111",
  47851=>"11111111",
  47852=>"00000001",
  47853=>"00000001",
  47854=>"00000010",
  47855=>"00000010",
  47856=>"00000100",
  47857=>"00000010",
  47858=>"00000010",
  47859=>"11111110",
  47860=>"11111111",
  47861=>"11111110",
  47862=>"00000001",
  47863=>"00000010",
  47864=>"00000001",
  47865=>"00000100",
  47866=>"11111110",
  47867=>"11111111",
  47868=>"00000000",
  47869=>"11111111",
  47870=>"00000011",
  47871=>"11111110",
  47872=>"00000011",
  47873=>"00000101",
  47874=>"00000011",
  47875=>"00000011",
  47876=>"11111110",
  47877=>"11111111",
  47878=>"11111110",
  47879=>"00000000",
  47880=>"11111111",
  47881=>"00000000",
  47882=>"00000010",
  47883=>"00000001",
  47884=>"11111110",
  47885=>"11111111",
  47886=>"00000010",
  47887=>"11111111",
  47888=>"11111110",
  47889=>"00000001",
  47890=>"00000000",
  47891=>"00000001",
  47892=>"00000000",
  47893=>"11111110",
  47894=>"00000001",
  47895=>"11111111",
  47896=>"11111101",
  47897=>"00000001",
  47898=>"00000011",
  47899=>"00000010",
  47900=>"11111111",
  47901=>"00000000",
  47902=>"00000001",
  47903=>"11111110",
  47904=>"00000000",
  47905=>"00000011",
  47906=>"11111111",
  47907=>"00000000",
  47908=>"11111101",
  47909=>"00000010",
  47910=>"11111101",
  47911=>"11111111",
  47912=>"11111101",
  47913=>"11111101",
  47914=>"11111111",
  47915=>"00000000",
  47916=>"00000000",
  47917=>"00000001",
  47918=>"11111111",
  47919=>"00000010",
  47920=>"11111110",
  47921=>"00000000",
  47922=>"11111111",
  47923=>"00000100",
  47924=>"00000010",
  47925=>"00000000",
  47926=>"11111110",
  47927=>"00000010",
  47928=>"00000011",
  47929=>"00000010",
  47930=>"00000000",
  47931=>"11111111",
  47932=>"00000000",
  47933=>"00000000",
  47934=>"00000001",
  47935=>"11111110",
  47936=>"11111111",
  47937=>"00000011",
  47938=>"00000010",
  47939=>"11111111",
  47940=>"11111111",
  47941=>"11111101",
  47942=>"00000001",
  47943=>"11111111",
  47944=>"11111101",
  47945=>"11111110",
  47946=>"11111110",
  47947=>"11111111",
  47948=>"00000011",
  47949=>"11111110",
  47950=>"11111110",
  47951=>"11111110",
  47952=>"00000000",
  47953=>"00000010",
  47954=>"11111101",
  47955=>"00000000",
  47956=>"11111101",
  47957=>"11111110",
  47958=>"11111111",
  47959=>"11111101",
  47960=>"11111101",
  47961=>"00000011",
  47962=>"11111111",
  47963=>"00000000",
  47964=>"00000000",
  47965=>"11111101",
  47966=>"00000100",
  47967=>"00000011",
  47968=>"00000010",
  47969=>"00000001",
  47970=>"11111111",
  47971=>"11111111",
  47972=>"00000001",
  47973=>"11111110",
  47974=>"00000100",
  47975=>"00000001",
  47976=>"11111111",
  47977=>"11111101",
  47978=>"11111111",
  47979=>"11111110",
  47980=>"11111110",
  47981=>"00000000",
  47982=>"00000001",
  47983=>"00000100",
  47984=>"00000000",
  47985=>"00000001",
  47986=>"11111111",
  47987=>"00000010",
  47988=>"00000010",
  47989=>"00000001",
  47990=>"11111111",
  47991=>"11111101",
  47992=>"00000001",
  47993=>"00000001",
  47994=>"00000001",
  47995=>"11111110",
  47996=>"00000001",
  47997=>"00000001",
  47998=>"11111101",
  47999=>"00000010",
  48000=>"00000000",
  48001=>"11111111",
  48002=>"11111110",
  48003=>"11111111",
  48004=>"00000011",
  48005=>"11111110",
  48006=>"11111101",
  48007=>"11111110",
  48008=>"11111111",
  48009=>"11111111",
  48010=>"11111111",
  48011=>"00000000",
  48012=>"11111101",
  48013=>"00000010",
  48014=>"00000000",
  48015=>"00000000",
  48016=>"00000001",
  48017=>"00000001",
  48018=>"11111100",
  48019=>"00000000",
  48020=>"11111111",
  48021=>"00000000",
  48022=>"00000000",
  48023=>"11111110",
  48024=>"11111110",
  48025=>"11111110",
  48026=>"11111111",
  48027=>"11111101",
  48028=>"11111100",
  48029=>"11111110",
  48030=>"11111101",
  48031=>"00000000",
  48032=>"00000010",
  48033=>"11111110",
  48034=>"00000010",
  48035=>"00000000",
  48036=>"00000000",
  48037=>"00000001",
  48038=>"11111111",
  48039=>"00000001",
  48040=>"11111111",
  48041=>"11111100",
  48042=>"11111111",
  48043=>"11111111",
  48044=>"00000010",
  48045=>"00000010",
  48046=>"00000010",
  48047=>"00000000",
  48048=>"00000011",
  48049=>"11111100",
  48050=>"11111101",
  48051=>"00000000",
  48052=>"11111111",
  48053=>"11111111",
  48054=>"00000000",
  48055=>"00000010",
  48056=>"00000010",
  48057=>"00000001",
  48058=>"11111101",
  48059=>"00000010",
  48060=>"00000010",
  48061=>"11111101",
  48062=>"00000000",
  48063=>"00000000",
  48064=>"11111111",
  48065=>"11111101",
  48066=>"11111110",
  48067=>"00000001",
  48068=>"00000011",
  48069=>"00000011",
  48070=>"00000000",
  48071=>"11111111",
  48072=>"00000010",
  48073=>"11111101",
  48074=>"00000001",
  48075=>"00000001",
  48076=>"00000011",
  48077=>"00000010",
  48078=>"11111111",
  48079=>"00000001",
  48080=>"00000001",
  48081=>"11111110",
  48082=>"00000000",
  48083=>"11111110",
  48084=>"00000010",
  48085=>"00000000",
  48086=>"11111110",
  48087=>"00000010",
  48088=>"11111110",
  48089=>"11111101",
  48090=>"00000000",
  48091=>"11111111",
  48092=>"11111101",
  48093=>"11111101",
  48094=>"00000010",
  48095=>"11111111",
  48096=>"11111111",
  48097=>"11111110",
  48098=>"11111110",
  48099=>"11111110",
  48100=>"00000001",
  48101=>"00000001",
  48102=>"11111111",
  48103=>"00000001",
  48104=>"00000001",
  48105=>"00000100",
  48106=>"11111111",
  48107=>"00000100",
  48108=>"00000001",
  48109=>"00000001",
  48110=>"00000001",
  48111=>"11111111",
  48112=>"11111101",
  48113=>"00000001",
  48114=>"11111111",
  48115=>"00000010",
  48116=>"00000000",
  48117=>"11111110",
  48118=>"00000011",
  48119=>"00000001",
  48120=>"11111111",
  48121=>"11111111",
  48122=>"00000100",
  48123=>"00000000",
  48124=>"11111110",
  48125=>"00000001",
  48126=>"00000100",
  48127=>"00000000",
  48128=>"00000010",
  48129=>"11111101",
  48130=>"11111111",
  48131=>"00000010",
  48132=>"00000010",
  48133=>"00000101",
  48134=>"00000000",
  48135=>"00000000",
  48136=>"00000010",
  48137=>"00000010",
  48138=>"11111111",
  48139=>"11111111",
  48140=>"00000000",
  48141=>"00000001",
  48142=>"11111111",
  48143=>"00000000",
  48144=>"00000000",
  48145=>"11111100",
  48146=>"00000001",
  48147=>"00000000",
  48148=>"00000000",
  48149=>"11111110",
  48150=>"00000010",
  48151=>"11111101",
  48152=>"00000010",
  48153=>"00000010",
  48154=>"00000010",
  48155=>"00000010",
  48156=>"00000001",
  48157=>"00000000",
  48158=>"11111111",
  48159=>"11111111",
  48160=>"00000011",
  48161=>"00000010",
  48162=>"00000000",
  48163=>"11111111",
  48164=>"00000001",
  48165=>"11111101",
  48166=>"11111101",
  48167=>"00000000",
  48168=>"11111101",
  48169=>"11111111",
  48170=>"00000110",
  48171=>"00000001",
  48172=>"11111111",
  48173=>"11111111",
  48174=>"11111111",
  48175=>"11111101",
  48176=>"11111111",
  48177=>"11111110",
  48178=>"11111111",
  48179=>"00000010",
  48180=>"11111111",
  48181=>"11111101",
  48182=>"00000100",
  48183=>"00000011",
  48184=>"00001000",
  48185=>"11111111",
  48186=>"00000100",
  48187=>"00000001",
  48188=>"11111110",
  48189=>"11111111",
  48190=>"11111101",
  48191=>"00000011",
  48192=>"11111111",
  48193=>"00000001",
  48194=>"11111101",
  48195=>"11111111",
  48196=>"00000010",
  48197=>"00000000",
  48198=>"11111111",
  48199=>"00000011",
  48200=>"00000001",
  48201=>"11111111",
  48202=>"00000010",
  48203=>"11111101",
  48204=>"00000010",
  48205=>"11111101",
  48206=>"11111110",
  48207=>"11111111",
  48208=>"11111110",
  48209=>"11111111",
  48210=>"11111110",
  48211=>"00000001",
  48212=>"00000001",
  48213=>"11111110",
  48214=>"11111110",
  48215=>"11111111",
  48216=>"00000001",
  48217=>"11111110",
  48218=>"11111111",
  48219=>"00000001",
  48220=>"00000001",
  48221=>"00000001",
  48222=>"00000000",
  48223=>"11111101",
  48224=>"11111111",
  48225=>"00000011",
  48226=>"00000000",
  48227=>"11111111",
  48228=>"11111110",
  48229=>"11111110",
  48230=>"00000000",
  48231=>"00000010",
  48232=>"11111111",
  48233=>"00000101",
  48234=>"00000010",
  48235=>"11111111",
  48236=>"11111011",
  48237=>"00000001",
  48238=>"00000000",
  48239=>"11111101",
  48240=>"11111110",
  48241=>"00000111",
  48242=>"00000001",
  48243=>"00000110",
  48244=>"11111110",
  48245=>"00000101",
  48246=>"00000000",
  48247=>"00000010",
  48248=>"11111111",
  48249=>"00000001",
  48250=>"00000011",
  48251=>"11111110",
  48252=>"11111101",
  48253=>"00000000",
  48254=>"11111111",
  48255=>"11111111",
  48256=>"11111110",
  48257=>"00000101",
  48258=>"00000110",
  48259=>"00000001",
  48260=>"00000011",
  48261=>"11111111",
  48262=>"11111111",
  48263=>"00000010",
  48264=>"11111110",
  48265=>"11111110",
  48266=>"00000000",
  48267=>"11111110",
  48268=>"11111101",
  48269=>"11111111",
  48270=>"11111101",
  48271=>"00000000",
  48272=>"11111111",
  48273=>"00000010",
  48274=>"11111111",
  48275=>"00000001",
  48276=>"00000001",
  48277=>"00000001",
  48278=>"00000000",
  48279=>"11111101",
  48280=>"11111111",
  48281=>"11111110",
  48282=>"11111111",
  48283=>"00000101",
  48284=>"00000010",
  48285=>"00000100",
  48286=>"11111110",
  48287=>"00000000",
  48288=>"00000000",
  48289=>"11111101",
  48290=>"00000010",
  48291=>"00000001",
  48292=>"11111110",
  48293=>"11111110",
  48294=>"00000000",
  48295=>"00000100",
  48296=>"00000000",
  48297=>"11111111",
  48298=>"00000000",
  48299=>"00000000",
  48300=>"00000011",
  48301=>"11111101",
  48302=>"11111111",
  48303=>"11111111",
  48304=>"00000011",
  48305=>"00000010",
  48306=>"00000011",
  48307=>"00000000",
  48308=>"00000010",
  48309=>"00000000",
  48310=>"00000101",
  48311=>"11111100",
  48312=>"00000001",
  48313=>"11111111",
  48314=>"00000000",
  48315=>"00000100",
  48316=>"11111101",
  48317=>"00000010",
  48318=>"11111101",
  48319=>"00000000",
  48320=>"11111101",
  48321=>"00000010",
  48322=>"11111101",
  48323=>"00000000",
  48324=>"11111110",
  48325=>"00000110",
  48326=>"00000011",
  48327=>"11111111",
  48328=>"11111111",
  48329=>"11111111",
  48330=>"11111110",
  48331=>"00000000",
  48332=>"00000000",
  48333=>"11111111",
  48334=>"00000010",
  48335=>"11111111",
  48336=>"11111101",
  48337=>"00000010",
  48338=>"11111111",
  48339=>"00000000",
  48340=>"11111111",
  48341=>"11111101",
  48342=>"00000001",
  48343=>"11111111",
  48344=>"11111111",
  48345=>"00000001",
  48346=>"11111101",
  48347=>"00000000",
  48348=>"11111110",
  48349=>"11111101",
  48350=>"11111111",
  48351=>"11111111",
  48352=>"11111110",
  48353=>"00000000",
  48354=>"00000001",
  48355=>"11111110",
  48356=>"00000001",
  48357=>"00000001",
  48358=>"00000001",
  48359=>"11111111",
  48360=>"11111111",
  48361=>"00000010",
  48362=>"00000010",
  48363=>"00000010",
  48364=>"00000000",
  48365=>"00000001",
  48366=>"11111111",
  48367=>"00000000",
  48368=>"11111111",
  48369=>"00000001",
  48370=>"11111110",
  48371=>"00000010",
  48372=>"11111110",
  48373=>"00000001",
  48374=>"11111110",
  48375=>"00000000",
  48376=>"11111110",
  48377=>"00000000",
  48378=>"11111101",
  48379=>"00000000",
  48380=>"00000100",
  48381=>"00000000",
  48382=>"11111101",
  48383=>"11111111",
  48384=>"11111111",
  48385=>"00000010",
  48386=>"00000000",
  48387=>"00000011",
  48388=>"00000000",
  48389=>"00000000",
  48390=>"00000110",
  48391=>"00000011",
  48392=>"11111111",
  48393=>"00000011",
  48394=>"00000011",
  48395=>"00000001",
  48396=>"11111110",
  48397=>"11111110",
  48398=>"11111111",
  48399=>"00000001",
  48400=>"11111101",
  48401=>"11111110",
  48402=>"00000000",
  48403=>"11111101",
  48404=>"11111110",
  48405=>"00000001",
  48406=>"00000001",
  48407=>"00000001",
  48408=>"11111110",
  48409=>"00000001",
  48410=>"11111101",
  48411=>"00000001",
  48412=>"00000100",
  48413=>"11111101",
  48414=>"11111110",
  48415=>"00000000",
  48416=>"00000001",
  48417=>"00000100",
  48418=>"00000001",
  48419=>"11111111",
  48420=>"00000001",
  48421=>"11111110",
  48422=>"11111110",
  48423=>"00000010",
  48424=>"11111111",
  48425=>"00000011",
  48426=>"00000001",
  48427=>"00000010",
  48428=>"11111110",
  48429=>"00000011",
  48430=>"11111111",
  48431=>"00000001",
  48432=>"11111110",
  48433=>"11111100",
  48434=>"00000010",
  48435=>"11111111",
  48436=>"00000110",
  48437=>"11111101",
  48438=>"00000010",
  48439=>"11111110",
  48440=>"00000110",
  48441=>"00000001",
  48442=>"00000010",
  48443=>"11111111",
  48444=>"00000001",
  48445=>"11111110",
  48446=>"11111110",
  48447=>"00000010",
  48448=>"11111110",
  48449=>"00000001",
  48450=>"11111110",
  48451=>"11111111",
  48452=>"11111111",
  48453=>"00000001",
  48454=>"11111110",
  48455=>"00000001",
  48456=>"11111110",
  48457=>"11111101",
  48458=>"11111101",
  48459=>"00000000",
  48460=>"11111101",
  48461=>"00000000",
  48462=>"00000010",
  48463=>"11111110",
  48464=>"00000010",
  48465=>"11111110",
  48466=>"00000011",
  48467=>"11111111",
  48468=>"11111110",
  48469=>"00000000",
  48470=>"00000000",
  48471=>"11111101",
  48472=>"00000000",
  48473=>"00000000",
  48474=>"00000001",
  48475=>"11111110",
  48476=>"00000000",
  48477=>"00000010",
  48478=>"11111101",
  48479=>"00000000",
  48480=>"00000000",
  48481=>"11111110",
  48482=>"11111100",
  48483=>"11111101",
  48484=>"00000001",
  48485=>"00000000",
  48486=>"00000000",
  48487=>"00000001",
  48488=>"00000010",
  48489=>"11111101",
  48490=>"00000000",
  48491=>"00000000",
  48492=>"00000001",
  48493=>"11111101",
  48494=>"11111101",
  48495=>"11111110",
  48496=>"00000000",
  48497=>"00000001",
  48498=>"00000010",
  48499=>"00000010",
  48500=>"11111110",
  48501=>"11111110",
  48502=>"00000001",
  48503=>"00000010",
  48504=>"00000010",
  48505=>"11111111",
  48506=>"11111101",
  48507=>"11111110",
  48508=>"11111101",
  48509=>"11111101",
  48510=>"00000010",
  48511=>"00000010",
  48512=>"11111111",
  48513=>"00000001",
  48514=>"00000000",
  48515=>"11111101",
  48516=>"11111111",
  48517=>"11111111",
  48518=>"11111101",
  48519=>"00000011",
  48520=>"00000000",
  48521=>"11111111",
  48522=>"00000001",
  48523=>"11111110",
  48524=>"00000001",
  48525=>"00000010",
  48526=>"00000001",
  48527=>"11111101",
  48528=>"00000000",
  48529=>"11111100",
  48530=>"00000000",
  48531=>"00000000",
  48532=>"11111101",
  48533=>"00000000",
  48534=>"00000010",
  48535=>"11111101",
  48536=>"00000010",
  48537=>"00000000",
  48538=>"11111110",
  48539=>"11111110",
  48540=>"00000011",
  48541=>"00000001",
  48542=>"00000001",
  48543=>"11111110",
  48544=>"00000010",
  48545=>"00000000",
  48546=>"11111111",
  48547=>"11111101",
  48548=>"11111101",
  48549=>"11111111",
  48550=>"11111101",
  48551=>"00000000",
  48552=>"00000010",
  48553=>"00000000",
  48554=>"11111111",
  48555=>"00000010",
  48556=>"00000000",
  48557=>"11111110",
  48558=>"00000000",
  48559=>"00000001",
  48560=>"11111100",
  48561=>"00000010",
  48562=>"00000001",
  48563=>"11111111",
  48564=>"11111101",
  48565=>"11111101",
  48566=>"11111110",
  48567=>"11111100",
  48568=>"00000000",
  48569=>"00000000",
  48570=>"11111101",
  48571=>"11111111",
  48572=>"00000001",
  48573=>"00000000",
  48574=>"00000000",
  48575=>"11111111",
  48576=>"11111110",
  48577=>"00000101",
  48578=>"11111111",
  48579=>"11111101",
  48580=>"11111110",
  48581=>"00000001",
  48582=>"00000001",
  48583=>"11111111",
  48584=>"11111110",
  48585=>"11111111",
  48586=>"00000010",
  48587=>"00000000",
  48588=>"00000000",
  48589=>"11111111",
  48590=>"00000000",
  48591=>"00000011",
  48592=>"00000011",
  48593=>"11111110",
  48594=>"11111100",
  48595=>"11111100",
  48596=>"11111101",
  48597=>"00000000",
  48598=>"11111101",
  48599=>"00000010",
  48600=>"11111110",
  48601=>"11111101",
  48602=>"11111111",
  48603=>"00000001",
  48604=>"00000001",
  48605=>"00000001",
  48606=>"11111110",
  48607=>"11111101",
  48608=>"00000001",
  48609=>"00000000",
  48610=>"11111110",
  48611=>"00000001",
  48612=>"11111110",
  48613=>"11111101",
  48614=>"00000010",
  48615=>"00000000",
  48616=>"00000001",
  48617=>"11111111",
  48618=>"00000000",
  48619=>"11111101",
  48620=>"00000001",
  48621=>"00000101",
  48622=>"00000010",
  48623=>"00000101",
  48624=>"11111101",
  48625=>"00000010",
  48626=>"00000000",
  48627=>"00000000",
  48628=>"11111111",
  48629=>"00000100",
  48630=>"11111101",
  48631=>"11111110",
  48632=>"00000000",
  48633=>"11111111",
  48634=>"11111101",
  48635=>"00000000",
  48636=>"11111110",
  48637=>"11111101",
  48638=>"00000100",
  48639=>"00000001",
  48640=>"00000001",
  48641=>"00000010",
  48642=>"00000000",
  48643=>"00000110",
  48644=>"11111110",
  48645=>"11111111",
  48646=>"11111111",
  48647=>"00000001",
  48648=>"00000010",
  48649=>"00000001",
  48650=>"00000001",
  48651=>"00000001",
  48652=>"00000011",
  48653=>"11111111",
  48654=>"11111101",
  48655=>"00000000",
  48656=>"00000000",
  48657=>"00000001",
  48658=>"00000011",
  48659=>"00000000",
  48660=>"11111111",
  48661=>"11111110",
  48662=>"00000010",
  48663=>"11111111",
  48664=>"11111111",
  48665=>"00000001",
  48666=>"00000001",
  48667=>"00000001",
  48668=>"11111101",
  48669=>"00000001",
  48670=>"00000000",
  48671=>"00000000",
  48672=>"11111111",
  48673=>"11111101",
  48674=>"00000010",
  48675=>"00000000",
  48676=>"00000001",
  48677=>"11111111",
  48678=>"11111101",
  48679=>"11111110",
  48680=>"11111110",
  48681=>"11111100",
  48682=>"00000000",
  48683=>"00000010",
  48684=>"00000000",
  48685=>"00000010",
  48686=>"00000001",
  48687=>"00000100",
  48688=>"11111111",
  48689=>"00000001",
  48690=>"11111111",
  48691=>"00000011",
  48692=>"00000010",
  48693=>"11111110",
  48694=>"00000100",
  48695=>"00000000",
  48696=>"11111111",
  48697=>"00000010",
  48698=>"00000010",
  48699=>"11111110",
  48700=>"11111111",
  48701=>"11111111",
  48702=>"11111101",
  48703=>"00000010",
  48704=>"11111110",
  48705=>"00000001",
  48706=>"11111111",
  48707=>"00000001",
  48708=>"11111110",
  48709=>"00000000",
  48710=>"00000111",
  48711=>"11111111",
  48712=>"00000001",
  48713=>"00000000",
  48714=>"11111110",
  48715=>"11111100",
  48716=>"11111110",
  48717=>"00000010",
  48718=>"11111101",
  48719=>"00000000",
  48720=>"00000001",
  48721=>"11111111",
  48722=>"11111111",
  48723=>"11111111",
  48724=>"00000010",
  48725=>"00000001",
  48726=>"00000010",
  48727=>"00000110",
  48728=>"11111110",
  48729=>"00000000",
  48730=>"11111110",
  48731=>"00000000",
  48732=>"00000001",
  48733=>"11111111",
  48734=>"11111111",
  48735=>"11111110",
  48736=>"11111101",
  48737=>"00000001",
  48738=>"11111101",
  48739=>"11111111",
  48740=>"00000010",
  48741=>"11111101",
  48742=>"00000010",
  48743=>"11111101",
  48744=>"00000001",
  48745=>"11111101",
  48746=>"11111110",
  48747=>"00000010",
  48748=>"11111101",
  48749=>"11111110",
  48750=>"00000001",
  48751=>"00000000",
  48752=>"00000001",
  48753=>"11111100",
  48754=>"11111110",
  48755=>"00000000",
  48756=>"11111111",
  48757=>"00000001",
  48758=>"00000000",
  48759=>"00000010",
  48760=>"11111111",
  48761=>"00000010",
  48762=>"11111111",
  48763=>"00000001",
  48764=>"00000011",
  48765=>"00000010",
  48766=>"00000000",
  48767=>"11111110",
  48768=>"00000001",
  48769=>"00000101",
  48770=>"11111111",
  48771=>"00000010",
  48772=>"11111100",
  48773=>"11111110",
  48774=>"00000011",
  48775=>"00000010",
  48776=>"00000001",
  48777=>"11111100",
  48778=>"00000001",
  48779=>"00000000",
  48780=>"11111111",
  48781=>"00000000",
  48782=>"11111110",
  48783=>"00000001",
  48784=>"11111111",
  48785=>"11111111",
  48786=>"11111111",
  48787=>"00000011",
  48788=>"11111110",
  48789=>"00000001",
  48790=>"00000000",
  48791=>"00000001",
  48792=>"11111111",
  48793=>"11111101",
  48794=>"11111100",
  48795=>"00000000",
  48796=>"00001000",
  48797=>"00000001",
  48798=>"00000000",
  48799=>"11111111",
  48800=>"00000001",
  48801=>"11111101",
  48802=>"11111111",
  48803=>"00000000",
  48804=>"11111111",
  48805=>"00000000",
  48806=>"00000000",
  48807=>"00000001",
  48808=>"00000011",
  48809=>"00000001",
  48810=>"11111110",
  48811=>"00000001",
  48812=>"00000001",
  48813=>"00000000",
  48814=>"00000010",
  48815=>"11111111",
  48816=>"11111100",
  48817=>"11111101",
  48818=>"11111101",
  48819=>"11111111",
  48820=>"00000100",
  48821=>"00000001",
  48822=>"00000100",
  48823=>"00000001",
  48824=>"00000100",
  48825=>"00000010",
  48826=>"00000010",
  48827=>"00000100",
  48828=>"00000000",
  48829=>"11111110",
  48830=>"11111101",
  48831=>"11111111",
  48832=>"00000000",
  48833=>"00000010",
  48834=>"11111110",
  48835=>"00000100",
  48836=>"11111101",
  48837=>"00000001",
  48838=>"00000001",
  48839=>"00000000",
  48840=>"00000010",
  48841=>"11111101",
  48842=>"00000000",
  48843=>"00000010",
  48844=>"00000000",
  48845=>"11111111",
  48846=>"00000010",
  48847=>"00000001",
  48848=>"00000000",
  48849=>"00000100",
  48850=>"00000010",
  48851=>"11111110",
  48852=>"00000011",
  48853=>"00000010",
  48854=>"00000010",
  48855=>"00000000",
  48856=>"00000000",
  48857=>"11111111",
  48858=>"11111110",
  48859=>"11111110",
  48860=>"11111100",
  48861=>"00000000",
  48862=>"00000000",
  48863=>"00000010",
  48864=>"11111110",
  48865=>"00000011",
  48866=>"11111110",
  48867=>"11111110",
  48868=>"11111110",
  48869=>"11111101",
  48870=>"00000010",
  48871=>"11111110",
  48872=>"11111101",
  48873=>"00000000",
  48874=>"00000010",
  48875=>"00000010",
  48876=>"00000001",
  48877=>"00000111",
  48878=>"11111111",
  48879=>"11111101",
  48880=>"00000000",
  48881=>"11111110",
  48882=>"00000001",
  48883=>"11111101",
  48884=>"11111110",
  48885=>"11111110",
  48886=>"00000000",
  48887=>"00000000",
  48888=>"11111101",
  48889=>"00000010",
  48890=>"00000001",
  48891=>"11111101",
  48892=>"11111111",
  48893=>"00000001",
  48894=>"00000000",
  48895=>"11111111",
  48896=>"00000000",
  48897=>"11111101",
  48898=>"00000010",
  48899=>"00000010",
  48900=>"11111110",
  48901=>"00000000",
  48902=>"00000011",
  48903=>"11111110",
  48904=>"00000000",
  48905=>"00000001",
  48906=>"00000001",
  48907=>"11111110",
  48908=>"11111111",
  48909=>"11111100",
  48910=>"11111111",
  48911=>"00000010",
  48912=>"11111111",
  48913=>"11111101",
  48914=>"11111101",
  48915=>"00000000",
  48916=>"00000000",
  48917=>"11111111",
  48918=>"11111101",
  48919=>"00000000",
  48920=>"11111111",
  48921=>"11111100",
  48922=>"00000000",
  48923=>"00000000",
  48924=>"00000001",
  48925=>"11111110",
  48926=>"00000011",
  48927=>"00000100",
  48928=>"00000001",
  48929=>"00000011",
  48930=>"00000000",
  48931=>"11111111",
  48932=>"00000011",
  48933=>"00000000",
  48934=>"00000010",
  48935=>"00000001",
  48936=>"11111111",
  48937=>"00000000",
  48938=>"00000101",
  48939=>"00000010",
  48940=>"00000000",
  48941=>"11111111",
  48942=>"00000001",
  48943=>"11111101",
  48944=>"11111111",
  48945=>"00001000",
  48946=>"00000011",
  48947=>"00000011",
  48948=>"00000000",
  48949=>"00000000",
  48950=>"00000001",
  48951=>"00000001",
  48952=>"00000001",
  48953=>"11111110",
  48954=>"00000000",
  48955=>"11111111",
  48956=>"00000001",
  48957=>"11111110",
  48958=>"11111110",
  48959=>"11111110",
  48960=>"00000000",
  48961=>"00000001",
  48962=>"00000000",
  48963=>"00000000",
  48964=>"11111111",
  48965=>"00000000",
  48966=>"11111110",
  48967=>"00000000",
  48968=>"00000010",
  48969=>"11111110",
  48970=>"11111111",
  48971=>"00000000",
  48972=>"00000001",
  48973=>"11111111",
  48974=>"00000011",
  48975=>"00000001",
  48976=>"11111110",
  48977=>"00000000",
  48978=>"00000100",
  48979=>"00000010",
  48980=>"11111110",
  48981=>"00000000",
  48982=>"00000000",
  48983=>"00000101",
  48984=>"11111111",
  48985=>"00000010",
  48986=>"11111101",
  48987=>"11111101",
  48988=>"11111101",
  48989=>"00000001",
  48990=>"00000000",
  48991=>"00000011",
  48992=>"11111111",
  48993=>"00000001",
  48994=>"11111110",
  48995=>"00000000",
  48996=>"11111111",
  48997=>"00000001",
  48998=>"11111110",
  48999=>"11111111",
  49000=>"00000010",
  49001=>"00000001",
  49002=>"00000001",
  49003=>"11111111",
  49004=>"11111111",
  49005=>"00000000",
  49006=>"11111111",
  49007=>"00000010",
  49008=>"11111111",
  49009=>"11111101",
  49010=>"11111111",
  49011=>"11111110",
  49012=>"00000001",
  49013=>"00000011",
  49014=>"00000000",
  49015=>"11111110",
  49016=>"00000000",
  49017=>"00000001",
  49018=>"11111111",
  49019=>"00000010",
  49020=>"11111101",
  49021=>"00000001",
  49022=>"00000001",
  49023=>"00000010",
  49024=>"00000000",
  49025=>"11111101",
  49026=>"11111110",
  49027=>"00000001",
  49028=>"00000001",
  49029=>"00000000",
  49030=>"00000011",
  49031=>"00000001",
  49032=>"11111111",
  49033=>"00000100",
  49034=>"11111110",
  49035=>"00000001",
  49036=>"00000000",
  49037=>"11111111",
  49038=>"11111110",
  49039=>"00000010",
  49040=>"00000010",
  49041=>"00000001",
  49042=>"11111101",
  49043=>"00000001",
  49044=>"00000001",
  49045=>"11111111",
  49046=>"00000100",
  49047=>"11111111",
  49048=>"11111110",
  49049=>"11111111",
  49050=>"11111101",
  49051=>"11111110",
  49052=>"00000001",
  49053=>"00000010",
  49054=>"00000101",
  49055=>"00000000",
  49056=>"00000000",
  49057=>"11111111",
  49058=>"11111101",
  49059=>"00000000",
  49060=>"00000010",
  49061=>"00000010",
  49062=>"11111110",
  49063=>"00000001",
  49064=>"11111111",
  49065=>"00000000",
  49066=>"11111111",
  49067=>"00000001",
  49068=>"00000010",
  49069=>"11111111",
  49070=>"11111110",
  49071=>"00000001",
  49072=>"11111110",
  49073=>"00000011",
  49074=>"11111110",
  49075=>"00000110",
  49076=>"11111101",
  49077=>"11111110",
  49078=>"00000011",
  49079=>"11111101",
  49080=>"00000000",
  49081=>"00000101",
  49082=>"00000000",
  49083=>"00000000",
  49084=>"00000010",
  49085=>"00000000",
  49086=>"00000010",
  49087=>"00000001",
  49088=>"00000010",
  49089=>"11111111",
  49090=>"11111110",
  49091=>"00000001",
  49092=>"00000010",
  49093=>"00000001",
  49094=>"11111110",
  49095=>"00000010",
  49096=>"00000011",
  49097=>"00000001",
  49098=>"00000000",
  49099=>"00000001",
  49100=>"00000101",
  49101=>"00000010",
  49102=>"00000000",
  49103=>"11111101",
  49104=>"00000000",
  49105=>"00000001",
  49106=>"00000101",
  49107=>"00000000",
  49108=>"00000010",
  49109=>"00000001",
  49110=>"00000101",
  49111=>"11111110",
  49112=>"00000011",
  49113=>"11111111",
  49114=>"00000001",
  49115=>"11111110",
  49116=>"00000011",
  49117=>"00000000",
  49118=>"00000011",
  49119=>"00000001",
  49120=>"00000010",
  49121=>"00000100",
  49122=>"00000000",
  49123=>"11111111",
  49124=>"11111110",
  49125=>"00000110",
  49126=>"11111110",
  49127=>"00000010",
  49128=>"11111110",
  49129=>"00000010",
  49130=>"00000000",
  49131=>"11111110",
  49132=>"00000010",
  49133=>"11111101",
  49134=>"11111110",
  49135=>"11111110",
  49136=>"00000010",
  49137=>"11111110",
  49138=>"00000011",
  49139=>"00000001",
  49140=>"00000110",
  49141=>"11111111",
  49142=>"00000011",
  49143=>"11111111",
  49144=>"00000010",
  49145=>"00000000",
  49146=>"00000001",
  49147=>"00000001",
  49148=>"11111100",
  49149=>"00000000",
  49150=>"00000000",
  49151=>"00000010",
  49152=>"00000000",
  49153=>"11111101",
  49154=>"11111110",
  49155=>"00000001",
  49156=>"00000110",
  49157=>"00000010",
  49158=>"11111111",
  49159=>"11111110",
  49160=>"00000000",
  49161=>"11111110",
  49162=>"00000000",
  49163=>"00000000",
  49164=>"11111100",
  49165=>"00000010",
  49166=>"11111111",
  49167=>"00000011",
  49168=>"11111101",
  49169=>"11111111",
  49170=>"00000000",
  49171=>"11111110",
  49172=>"11111100",
  49173=>"00000000",
  49174=>"00000010",
  49175=>"00000001",
  49176=>"11111101",
  49177=>"00000010",
  49178=>"00000011",
  49179=>"11111110",
  49180=>"11111111",
  49181=>"11111110",
  49182=>"00000101",
  49183=>"00000100",
  49184=>"11111110",
  49185=>"11111111",
  49186=>"11111111",
  49187=>"11111111",
  49188=>"00000101",
  49189=>"00000100",
  49190=>"11111111",
  49191=>"11111111",
  49192=>"11111100",
  49193=>"11111101",
  49194=>"00000100",
  49195=>"11111101",
  49196=>"00000101",
  49197=>"11111111",
  49198=>"11111110",
  49199=>"11111111",
  49200=>"00000011",
  49201=>"00000010",
  49202=>"11111101",
  49203=>"00000011",
  49204=>"11111111",
  49205=>"11111111",
  49206=>"00000001",
  49207=>"00000000",
  49208=>"00000011",
  49209=>"11111111",
  49210=>"00000001",
  49211=>"11111101",
  49212=>"00000000",
  49213=>"00000000",
  49214=>"11111100",
  49215=>"00000101",
  49216=>"00000010",
  49217=>"11111110",
  49218=>"11111101",
  49219=>"00000010",
  49220=>"11111111",
  49221=>"00000000",
  49222=>"11111101",
  49223=>"00000010",
  49224=>"11111111",
  49225=>"11111110",
  49226=>"00000010",
  49227=>"00000001",
  49228=>"00000001",
  49229=>"00000000",
  49230=>"00000000",
  49231=>"00000000",
  49232=>"11111111",
  49233=>"00000010",
  49234=>"00000000",
  49235=>"00000010",
  49236=>"00000001",
  49237=>"11111110",
  49238=>"11111111",
  49239=>"00000010",
  49240=>"00000000",
  49241=>"11111101",
  49242=>"00000011",
  49243=>"11111011",
  49244=>"00000011",
  49245=>"00000011",
  49246=>"00000010",
  49247=>"00000000",
  49248=>"11111110",
  49249=>"00000100",
  49250=>"00000010",
  49251=>"00000100",
  49252=>"00000000",
  49253=>"00000100",
  49254=>"11111111",
  49255=>"00000010",
  49256=>"00000010",
  49257=>"11111011",
  49258=>"11111111",
  49259=>"00000000",
  49260=>"00000100",
  49261=>"00000100",
  49262=>"11111110",
  49263=>"00000000",
  49264=>"00000010",
  49265=>"11111110",
  49266=>"00000000",
  49267=>"00000100",
  49268=>"00000000",
  49269=>"00000011",
  49270=>"00000000",
  49271=>"11111100",
  49272=>"11111100",
  49273=>"00000000",
  49274=>"11111111",
  49275=>"00000010",
  49276=>"11111110",
  49277=>"11111100",
  49278=>"11111111",
  49279=>"00000100",
  49280=>"00000001",
  49281=>"00000011",
  49282=>"00000001",
  49283=>"11111111",
  49284=>"00000010",
  49285=>"11111110",
  49286=>"11111110",
  49287=>"00000100",
  49288=>"11111111",
  49289=>"11111111",
  49290=>"00000000",
  49291=>"00000001",
  49292=>"00000001",
  49293=>"00000000",
  49294=>"00000100",
  49295=>"11111110",
  49296=>"00000110",
  49297=>"00000001",
  49298=>"11111110",
  49299=>"11111111",
  49300=>"11111101",
  49301=>"00000001",
  49302=>"00000010",
  49303=>"11111110",
  49304=>"11111111",
  49305=>"00000001",
  49306=>"11111101",
  49307=>"00000000",
  49308=>"00000001",
  49309=>"00000000",
  49310=>"00000000",
  49311=>"00000000",
  49312=>"00000010",
  49313=>"11111110",
  49314=>"00000001",
  49315=>"00000001",
  49316=>"00000000",
  49317=>"00000011",
  49318=>"11111111",
  49319=>"00000000",
  49320=>"11111110",
  49321=>"00000010",
  49322=>"11111101",
  49323=>"00000010",
  49324=>"11111110",
  49325=>"00000010",
  49326=>"11111101",
  49327=>"11111110",
  49328=>"11111111",
  49329=>"11111101",
  49330=>"00000001",
  49331=>"11111111",
  49332=>"00000100",
  49333=>"11111110",
  49334=>"00000010",
  49335=>"11111100",
  49336=>"11111011",
  49337=>"00000010",
  49338=>"00000010",
  49339=>"00000100",
  49340=>"00000000",
  49341=>"11111110",
  49342=>"00000000",
  49343=>"11111110",
  49344=>"11111111",
  49345=>"11111111",
  49346=>"00000000",
  49347=>"11111110",
  49348=>"11111111",
  49349=>"00000101",
  49350=>"00000011",
  49351=>"00000000",
  49352=>"00000010",
  49353=>"00000101",
  49354=>"00000000",
  49355=>"00000010",
  49356=>"00000011",
  49357=>"00000000",
  49358=>"11111101",
  49359=>"11111100",
  49360=>"00000010",
  49361=>"00000011",
  49362=>"00000000",
  49363=>"00000000",
  49364=>"11111110",
  49365=>"11111101",
  49366=>"00000011",
  49367=>"11111110",
  49368=>"11111100",
  49369=>"11111111",
  49370=>"00000010",
  49371=>"00000011",
  49372=>"00000001",
  49373=>"11111110",
  49374=>"00000001",
  49375=>"11111100",
  49376=>"00000000",
  49377=>"11111110",
  49378=>"11111110",
  49379=>"00000001",
  49380=>"11111110",
  49381=>"11111101",
  49382=>"00000000",
  49383=>"00000010",
  49384=>"00000100",
  49385=>"00000010",
  49386=>"00000010",
  49387=>"00000010",
  49388=>"11111111",
  49389=>"00000011",
  49390=>"11111100",
  49391=>"11111110",
  49392=>"11111110",
  49393=>"11111110",
  49394=>"00000011",
  49395=>"00000001",
  49396=>"00000000",
  49397=>"00000000",
  49398=>"00000001",
  49399=>"00000001",
  49400=>"00000011",
  49401=>"00000000",
  49402=>"11111101",
  49403=>"00000000",
  49404=>"00000101",
  49405=>"00000100",
  49406=>"00000001",
  49407=>"11111111",
  49408=>"11111111",
  49409=>"00000001",
  49410=>"11111101",
  49411=>"11111101",
  49412=>"00000001",
  49413=>"00000000",
  49414=>"00000100",
  49415=>"00000101",
  49416=>"00000000",
  49417=>"11111110",
  49418=>"00000011",
  49419=>"00000010",
  49420=>"11111110",
  49421=>"00000000",
  49422=>"11111101",
  49423=>"00000000",
  49424=>"11111110",
  49425=>"00000010",
  49426=>"11111101",
  49427=>"00000010",
  49428=>"11111111",
  49429=>"00000001",
  49430=>"00000001",
  49431=>"11111111",
  49432=>"11111101",
  49433=>"00000011",
  49434=>"00000011",
  49435=>"11111111",
  49436=>"00000100",
  49437=>"00000000",
  49438=>"00000010",
  49439=>"00000001",
  49440=>"11111101",
  49441=>"00000001",
  49442=>"11111100",
  49443=>"00000010",
  49444=>"11111110",
  49445=>"00000100",
  49446=>"00000001",
  49447=>"00000100",
  49448=>"00000000",
  49449=>"11111111",
  49450=>"00000010",
  49451=>"11111111",
  49452=>"11111101",
  49453=>"11111110",
  49454=>"00000001",
  49455=>"11111111",
  49456=>"00000011",
  49457=>"11111111",
  49458=>"11111101",
  49459=>"11111110",
  49460=>"00000000",
  49461=>"00000100",
  49462=>"00000000",
  49463=>"00000001",
  49464=>"00000011",
  49465=>"11111101",
  49466=>"11111101",
  49467=>"00000010",
  49468=>"00000001",
  49469=>"00000000",
  49470=>"00000100",
  49471=>"00000001",
  49472=>"00000000",
  49473=>"00000010",
  49474=>"00000100",
  49475=>"11111101",
  49476=>"00000000",
  49477=>"00000001",
  49478=>"11111110",
  49479=>"00000000",
  49480=>"00000001",
  49481=>"00000100",
  49482=>"00000001",
  49483=>"00000010",
  49484=>"00000010",
  49485=>"11111111",
  49486=>"11111111",
  49487=>"00000011",
  49488=>"11111100",
  49489=>"11111111",
  49490=>"00000001",
  49491=>"11111110",
  49492=>"00000001",
  49493=>"00000000",
  49494=>"11111110",
  49495=>"00000000",
  49496=>"00000101",
  49497=>"11111110",
  49498=>"11111101",
  49499=>"00000001",
  49500=>"00000100",
  49501=>"00000001",
  49502=>"11111111",
  49503=>"00000000",
  49504=>"00000001",
  49505=>"11111110",
  49506=>"00000001",
  49507=>"11111111",
  49508=>"00000001",
  49509=>"00000000",
  49510=>"11111101",
  49511=>"00000000",
  49512=>"00000010",
  49513=>"11111101",
  49514=>"11111111",
  49515=>"11111111",
  49516=>"00000011",
  49517=>"00000001",
  49518=>"11111111",
  49519=>"11111111",
  49520=>"11111111",
  49521=>"00000000",
  49522=>"00000101",
  49523=>"00000010",
  49524=>"11111101",
  49525=>"11111110",
  49526=>"00000010",
  49527=>"00000011",
  49528=>"11111111",
  49529=>"00000101",
  49530=>"11111111",
  49531=>"00000000",
  49532=>"00000000",
  49533=>"00000010",
  49534=>"11111110",
  49535=>"00000110",
  49536=>"00000011",
  49537=>"00000010",
  49538=>"00000001",
  49539=>"00000000",
  49540=>"11111110",
  49541=>"11111101",
  49542=>"00000000",
  49543=>"00000010",
  49544=>"11111110",
  49545=>"00000000",
  49546=>"11111111",
  49547=>"00000000",
  49548=>"11111101",
  49549=>"00000001",
  49550=>"11111111",
  49551=>"11111111",
  49552=>"11111110",
  49553=>"11111101",
  49554=>"00000010",
  49555=>"11111100",
  49556=>"00000000",
  49557=>"00000100",
  49558=>"11111100",
  49559=>"00000101",
  49560=>"00000100",
  49561=>"00000001",
  49562=>"00000000",
  49563=>"00000000",
  49564=>"11111101",
  49565=>"11111111",
  49566=>"00000001",
  49567=>"00000100",
  49568=>"11111110",
  49569=>"11111110",
  49570=>"11111111",
  49571=>"11111111",
  49572=>"00000000",
  49573=>"11111101",
  49574=>"11111101",
  49575=>"00000001",
  49576=>"11111111",
  49577=>"11111111",
  49578=>"11111111",
  49579=>"00000001",
  49580=>"11111111",
  49581=>"00000010",
  49582=>"00000100",
  49583=>"11111110",
  49584=>"00000011",
  49585=>"11111111",
  49586=>"11111111",
  49587=>"00000000",
  49588=>"00000000",
  49589=>"11111110",
  49590=>"11111111",
  49591=>"00000000",
  49592=>"00000010",
  49593=>"00000010",
  49594=>"11111111",
  49595=>"00000010",
  49596=>"00000000",
  49597=>"00000000",
  49598=>"00000010",
  49599=>"00000000",
  49600=>"11111101",
  49601=>"11111110",
  49602=>"00000010",
  49603=>"00000000",
  49604=>"11111111",
  49605=>"11111111",
  49606=>"11111110",
  49607=>"00000011",
  49608=>"11111111",
  49609=>"00000001",
  49610=>"11111110",
  49611=>"00000001",
  49612=>"00000010",
  49613=>"11111101",
  49614=>"00000010",
  49615=>"00000000",
  49616=>"00000001",
  49617=>"11111110",
  49618=>"00000011",
  49619=>"11111111",
  49620=>"00000000",
  49621=>"11111110",
  49622=>"11111101",
  49623=>"11111110",
  49624=>"11111101",
  49625=>"11111101",
  49626=>"11111110",
  49627=>"00000010",
  49628=>"00000010",
  49629=>"00000010",
  49630=>"11111111",
  49631=>"00000011",
  49632=>"11111101",
  49633=>"11111101",
  49634=>"11111111",
  49635=>"00000000",
  49636=>"11111111",
  49637=>"00000001",
  49638=>"00000000",
  49639=>"00000010",
  49640=>"00000010",
  49641=>"00000001",
  49642=>"00000001",
  49643=>"00000001",
  49644=>"00000010",
  49645=>"00000010",
  49646=>"11111111",
  49647=>"00000000",
  49648=>"00000001",
  49649=>"11111101",
  49650=>"11111110",
  49651=>"11111110",
  49652=>"00000000",
  49653=>"11111110",
  49654=>"11111111",
  49655=>"00000001",
  49656=>"11111111",
  49657=>"11111111",
  49658=>"11111101",
  49659=>"11111110",
  49660=>"11111111",
  49661=>"11111110",
  49662=>"11111111",
  49663=>"00000000",
  49664=>"11111111",
  49665=>"00000001",
  49666=>"11111110",
  49667=>"00000010",
  49668=>"11111110",
  49669=>"00000001",
  49670=>"11111110",
  49671=>"00000100",
  49672=>"11111110",
  49673=>"11111101",
  49674=>"00000001",
  49675=>"11111110",
  49676=>"00000010",
  49677=>"11111101",
  49678=>"00000100",
  49679=>"11111101",
  49680=>"00000000",
  49681=>"11111100",
  49682=>"00000001",
  49683=>"00000011",
  49684=>"11111110",
  49685=>"00000001",
  49686=>"11111110",
  49687=>"00000001",
  49688=>"00000000",
  49689=>"00000000",
  49690=>"11111110",
  49691=>"00000010",
  49692=>"00000001",
  49693=>"00000010",
  49694=>"00000001",
  49695=>"00000001",
  49696=>"11111101",
  49697=>"00000001",
  49698=>"11111111",
  49699=>"00000001",
  49700=>"11111111",
  49701=>"00000110",
  49702=>"11111111",
  49703=>"00000100",
  49704=>"11111101",
  49705=>"00000100",
  49706=>"00000001",
  49707=>"00000001",
  49708=>"11111100",
  49709=>"00000000",
  49710=>"00000001",
  49711=>"11111110",
  49712=>"00000101",
  49713=>"11111110",
  49714=>"11111101",
  49715=>"11111110",
  49716=>"11111101",
  49717=>"11111111",
  49718=>"11111101",
  49719=>"00000001",
  49720=>"00000001",
  49721=>"11111110",
  49722=>"00000001",
  49723=>"00000010",
  49724=>"00000001",
  49725=>"11111101",
  49726=>"11111111",
  49727=>"00000010",
  49728=>"11111100",
  49729=>"00000010",
  49730=>"11111110",
  49731=>"11111111",
  49732=>"00000010",
  49733=>"11111111",
  49734=>"11111101",
  49735=>"00000001",
  49736=>"11111111",
  49737=>"00000010",
  49738=>"00000000",
  49739=>"11111110",
  49740=>"00000000",
  49741=>"11111111",
  49742=>"00000011",
  49743=>"11111111",
  49744=>"00000000",
  49745=>"00000000",
  49746=>"00000000",
  49747=>"00000100",
  49748=>"11111110",
  49749=>"11111111",
  49750=>"00000010",
  49751=>"00000010",
  49752=>"00000010",
  49753=>"11111101",
  49754=>"11111110",
  49755=>"00000001",
  49756=>"11111111",
  49757=>"00000000",
  49758=>"11111110",
  49759=>"00000000",
  49760=>"00000000",
  49761=>"00000000",
  49762=>"11111101",
  49763=>"00000100",
  49764=>"11111100",
  49765=>"11111100",
  49766=>"00000000",
  49767=>"00000001",
  49768=>"11111101",
  49769=>"00000011",
  49770=>"11111110",
  49771=>"00000001",
  49772=>"11111110",
  49773=>"00000010",
  49774=>"11111110",
  49775=>"00000110",
  49776=>"00000000",
  49777=>"00000001",
  49778=>"00000100",
  49779=>"00000000",
  49780=>"11111110",
  49781=>"00000001",
  49782=>"11111111",
  49783=>"00000101",
  49784=>"00000001",
  49785=>"00000010",
  49786=>"11111111",
  49787=>"11111111",
  49788=>"11111111",
  49789=>"00000010",
  49790=>"00000110",
  49791=>"11111101",
  49792=>"00000001",
  49793=>"11111110",
  49794=>"11111111",
  49795=>"00000011",
  49796=>"11111100",
  49797=>"11111101",
  49798=>"11111110",
  49799=>"11111111",
  49800=>"11111101",
  49801=>"11111110",
  49802=>"11111101",
  49803=>"11111111",
  49804=>"11111110",
  49805=>"11111101",
  49806=>"11111111",
  49807=>"11111111",
  49808=>"00000000",
  49809=>"11111101",
  49810=>"11111110",
  49811=>"00000001",
  49812=>"00000100",
  49813=>"00000001",
  49814=>"11111111",
  49815=>"00000011",
  49816=>"00000000",
  49817=>"00001000",
  49818=>"00000001",
  49819=>"00000010",
  49820=>"00000110",
  49821=>"00000001",
  49822=>"11111101",
  49823=>"00000000",
  49824=>"00000010",
  49825=>"00000001",
  49826=>"00000011",
  49827=>"11111101",
  49828=>"00000001",
  49829=>"11111101",
  49830=>"00000000",
  49831=>"00000101",
  49832=>"11111110",
  49833=>"11111111",
  49834=>"11111110",
  49835=>"11111111",
  49836=>"11111111",
  49837=>"00000000",
  49838=>"11111101",
  49839=>"11111101",
  49840=>"00000001",
  49841=>"11111101",
  49842=>"00000010",
  49843=>"00000001",
  49844=>"00000010",
  49845=>"11111101",
  49846=>"11111110",
  49847=>"00000010",
  49848=>"11111110",
  49849=>"11111101",
  49850=>"11111111",
  49851=>"00000001",
  49852=>"00000000",
  49853=>"11111110",
  49854=>"11111110",
  49855=>"00000001",
  49856=>"11111101",
  49857=>"11111101",
  49858=>"00000101",
  49859=>"00000010",
  49860=>"11111110",
  49861=>"11111101",
  49862=>"00000000",
  49863=>"00000000",
  49864=>"00000000",
  49865=>"00000001",
  49866=>"11111101",
  49867=>"11111100",
  49868=>"11111111",
  49869=>"11111110",
  49870=>"11111100",
  49871=>"11111101",
  49872=>"11111111",
  49873=>"00000000",
  49874=>"00000010",
  49875=>"11111111",
  49876=>"00000100",
  49877=>"00000110",
  49878=>"00000010",
  49879=>"11111110",
  49880=>"00000011",
  49881=>"11111110",
  49882=>"11111110",
  49883=>"00000110",
  49884=>"11111110",
  49885=>"11111111",
  49886=>"00000000",
  49887=>"00000100",
  49888=>"11111111",
  49889=>"00000000",
  49890=>"11111101",
  49891=>"00000000",
  49892=>"00000000",
  49893=>"00000011",
  49894=>"11111110",
  49895=>"00000011",
  49896=>"00000000",
  49897=>"00000000",
  49898=>"00000100",
  49899=>"00000010",
  49900=>"00000010",
  49901=>"11111101",
  49902=>"00000101",
  49903=>"00000001",
  49904=>"00000010",
  49905=>"00000001",
  49906=>"00000000",
  49907=>"00000001",
  49908=>"00000001",
  49909=>"11111101",
  49910=>"00000011",
  49911=>"00000000",
  49912=>"11111111",
  49913=>"11111111",
  49914=>"00000000",
  49915=>"00000011",
  49916=>"11111111",
  49917=>"11111101",
  49918=>"11111110",
  49919=>"00000001",
  49920=>"00000000",
  49921=>"00000010",
  49922=>"00000000",
  49923=>"00000100",
  49924=>"11111111",
  49925=>"00000100",
  49926=>"00000100",
  49927=>"11111101",
  49928=>"11111110",
  49929=>"00000011",
  49930=>"00000010",
  49931=>"11111011",
  49932=>"00000011",
  49933=>"00000001",
  49934=>"00000000",
  49935=>"00000001",
  49936=>"00000000",
  49937=>"00000011",
  49938=>"11111111",
  49939=>"11111100",
  49940=>"11111100",
  49941=>"11111110",
  49942=>"00000001",
  49943=>"00000000",
  49944=>"11111101",
  49945=>"11111110",
  49946=>"00000001",
  49947=>"00000001",
  49948=>"11111110",
  49949=>"00000010",
  49950=>"11111111",
  49951=>"00000001",
  49952=>"00000101",
  49953=>"11111101",
  49954=>"11111111",
  49955=>"11111110",
  49956=>"00000101",
  49957=>"11111101",
  49958=>"11111101",
  49959=>"11111110",
  49960=>"00000011",
  49961=>"11111100",
  49962=>"11111111",
  49963=>"00000010",
  49964=>"00000001",
  49965=>"00000000",
  49966=>"00000000",
  49967=>"11111110",
  49968=>"11111111",
  49969=>"00000100",
  49970=>"11111111",
  49971=>"00000010",
  49972=>"11111110",
  49973=>"11111100",
  49974=>"11111110",
  49975=>"00000000",
  49976=>"11111100",
  49977=>"00000001",
  49978=>"11111111",
  49979=>"11111111",
  49980=>"00000000",
  49981=>"00000010",
  49982=>"00000001",
  49983=>"11111110",
  49984=>"00000101",
  49985=>"11111110",
  49986=>"11111111",
  49987=>"00000110",
  49988=>"11111111",
  49989=>"00000001",
  49990=>"11111101",
  49991=>"11111110",
  49992=>"00000001",
  49993=>"00000001",
  49994=>"11111110",
  49995=>"00000000",
  49996=>"11111111",
  49997=>"00000010",
  49998=>"00000110",
  49999=>"00000001",
  50000=>"00000000",
  50001=>"11111101",
  50002=>"11111111",
  50003=>"00000100",
  50004=>"11111110",
  50005=>"00000001",
  50006=>"00000001",
  50007=>"11111110",
  50008=>"11111110",
  50009=>"00000011",
  50010=>"00000011",
  50011=>"00000000",
  50012=>"00000010",
  50013=>"00000001",
  50014=>"11111110",
  50015=>"00000010",
  50016=>"00000001",
  50017=>"00000000",
  50018=>"11111111",
  50019=>"11111110",
  50020=>"11111101",
  50021=>"00000010",
  50022=>"11111111",
  50023=>"00000110",
  50024=>"00000000",
  50025=>"00000010",
  50026=>"00000000",
  50027=>"00000010",
  50028=>"00000001",
  50029=>"11111101",
  50030=>"00000001",
  50031=>"11111110",
  50032=>"11111110",
  50033=>"00000000",
  50034=>"11111111",
  50035=>"00000000",
  50036=>"00000010",
  50037=>"00001000",
  50038=>"00000010",
  50039=>"11111101",
  50040=>"00000010",
  50041=>"00000001",
  50042=>"00000100",
  50043=>"00000010",
  50044=>"11111101",
  50045=>"00000010",
  50046=>"11111111",
  50047=>"00000100",
  50048=>"11111111",
  50049=>"11111100",
  50050=>"11111101",
  50051=>"00000000",
  50052=>"11111110",
  50053=>"00000000",
  50054=>"00000000",
  50055=>"00000000",
  50056=>"00000001",
  50057=>"00000100",
  50058=>"00000001",
  50059=>"11111110",
  50060=>"11111110",
  50061=>"00000001",
  50062=>"11111110",
  50063=>"00000000",
  50064=>"00000001",
  50065=>"00000010",
  50066=>"11111111",
  50067=>"00000001",
  50068=>"00000010",
  50069=>"11111110",
  50070=>"00000001",
  50071=>"00000000",
  50072=>"00000101",
  50073=>"00000010",
  50074=>"11111111",
  50075=>"00000011",
  50076=>"11111111",
  50077=>"00000011",
  50078=>"00000011",
  50079=>"11111101",
  50080=>"11111101",
  50081=>"00000001",
  50082=>"00000000",
  50083=>"11111110",
  50084=>"11111111",
  50085=>"11111110",
  50086=>"00000000",
  50087=>"00000001",
  50088=>"11111100",
  50089=>"11111110",
  50090=>"00000010",
  50091=>"11111101",
  50092=>"00000001",
  50093=>"00000001",
  50094=>"00000011",
  50095=>"00000001",
  50096=>"11111110",
  50097=>"00000011",
  50098=>"00000000",
  50099=>"00000010",
  50100=>"11111101",
  50101=>"11111101",
  50102=>"11111110",
  50103=>"00000110",
  50104=>"00000001",
  50105=>"00000011",
  50106=>"00000010",
  50107=>"11111110",
  50108=>"00000000",
  50109=>"00000001",
  50110=>"11111110",
  50111=>"11111111",
  50112=>"11111101",
  50113=>"00000011",
  50114=>"00000010",
  50115=>"00000000",
  50116=>"11111101",
  50117=>"11111111",
  50118=>"11111111",
  50119=>"11111110",
  50120=>"00000001",
  50121=>"11111110",
  50122=>"11111111",
  50123=>"00000000",
  50124=>"00000000",
  50125=>"00000011",
  50126=>"11111100",
  50127=>"00000001",
  50128=>"00000100",
  50129=>"11111111",
  50130=>"11111111",
  50131=>"11111101",
  50132=>"11111111",
  50133=>"00000011",
  50134=>"00000101",
  50135=>"00000100",
  50136=>"11111111",
  50137=>"00000011",
  50138=>"11111110",
  50139=>"00000111",
  50140=>"11111110",
  50141=>"00000000",
  50142=>"00000000",
  50143=>"11111111",
  50144=>"00000000",
  50145=>"00000000",
  50146=>"00000010",
  50147=>"00000000",
  50148=>"00000010",
  50149=>"11111110",
  50150=>"00000001",
  50151=>"11111111",
  50152=>"00000000",
  50153=>"11111110",
  50154=>"00000110",
  50155=>"00000110",
  50156=>"11111101",
  50157=>"11111100",
  50158=>"11111110",
  50159=>"00000001",
  50160=>"11111111",
  50161=>"00000000",
  50162=>"00000011",
  50163=>"00000001",
  50164=>"11111101",
  50165=>"00000010",
  50166=>"00000011",
  50167=>"00000000",
  50168=>"00000000",
  50169=>"00000011",
  50170=>"00000011",
  50171=>"00000010",
  50172=>"00000001",
  50173=>"11111100",
  50174=>"00000001",
  50175=>"11111100",
  50176=>"00000001",
  50177=>"00000010",
  50178=>"00000000",
  50179=>"11111111",
  50180=>"11111101",
  50181=>"00000000",
  50182=>"00000100",
  50183=>"00000000",
  50184=>"11111111",
  50185=>"00000100",
  50186=>"11111111",
  50187=>"00000010",
  50188=>"00000101",
  50189=>"00000100",
  50190=>"00000000",
  50191=>"00000001",
  50192=>"11111111",
  50193=>"11111111",
  50194=>"00000001",
  50195=>"00000100",
  50196=>"11111110",
  50197=>"00000000",
  50198=>"00000000",
  50199=>"00000110",
  50200=>"00000000",
  50201=>"11111111",
  50202=>"11111111",
  50203=>"11111100",
  50204=>"00000000",
  50205=>"00000000",
  50206=>"11111101",
  50207=>"11111110",
  50208=>"11111111",
  50209=>"00000010",
  50210=>"00000010",
  50211=>"00000000",
  50212=>"11111101",
  50213=>"00000000",
  50214=>"00000101",
  50215=>"00000011",
  50216=>"00000100",
  50217=>"11111111",
  50218=>"11111110",
  50219=>"00000000",
  50220=>"11111110",
  50221=>"00000010",
  50222=>"00000101",
  50223=>"00000000",
  50224=>"11111110",
  50225=>"00000110",
  50226=>"11111111",
  50227=>"00000011",
  50228=>"00000001",
  50229=>"11111110",
  50230=>"00000001",
  50231=>"11111101",
  50232=>"11111111",
  50233=>"11111101",
  50234=>"11111110",
  50235=>"00000010",
  50236=>"00000101",
  50237=>"11111110",
  50238=>"11111111",
  50239=>"11111101",
  50240=>"00000001",
  50241=>"00000101",
  50242=>"00000001",
  50243=>"00000011",
  50244=>"00000001",
  50245=>"11111111",
  50246=>"11111111",
  50247=>"11111101",
  50248=>"00000010",
  50249=>"00000100",
  50250=>"00000001",
  50251=>"00000100",
  50252=>"00000000",
  50253=>"00000000",
  50254=>"11111110",
  50255=>"00000011",
  50256=>"11111111",
  50257=>"00000011",
  50258=>"00000000",
  50259=>"11111100",
  50260=>"00000101",
  50261=>"00000000",
  50262=>"11111101",
  50263=>"11111101",
  50264=>"00000000",
  50265=>"11111101",
  50266=>"11111101",
  50267=>"11111101",
  50268=>"11111110",
  50269=>"11111110",
  50270=>"11111110",
  50271=>"11111011",
  50272=>"11111110",
  50273=>"00000010",
  50274=>"00000001",
  50275=>"00000001",
  50276=>"11111110",
  50277=>"00000001",
  50278=>"00000010",
  50279=>"00000100",
  50280=>"11111111",
  50281=>"00000000",
  50282=>"00000001",
  50283=>"00000100",
  50284=>"11111101",
  50285=>"11111101",
  50286=>"00000010",
  50287=>"00000001",
  50288=>"00000011",
  50289=>"00000000",
  50290=>"00000010",
  50291=>"11111111",
  50292=>"00000010",
  50293=>"00000011",
  50294=>"00000010",
  50295=>"00000001",
  50296=>"00000101",
  50297=>"00000001",
  50298=>"00000000",
  50299=>"11111101",
  50300=>"00000101",
  50301=>"00000010",
  50302=>"11111110",
  50303=>"11111101",
  50304=>"00000010",
  50305=>"11111101",
  50306=>"00000001",
  50307=>"11111100",
  50308=>"00000000",
  50309=>"00000000",
  50310=>"00000011",
  50311=>"00000011",
  50312=>"00000000",
  50313=>"00000011",
  50314=>"00000000",
  50315=>"00000000",
  50316=>"00000001",
  50317=>"00000001",
  50318=>"00000001",
  50319=>"00000000",
  50320=>"11111101",
  50321=>"11111100",
  50322=>"11111101",
  50323=>"11111101",
  50324=>"00000001",
  50325=>"00000100",
  50326=>"11111111",
  50327=>"00000100",
  50328=>"11111111",
  50329=>"11111111",
  50330=>"11111101",
  50331=>"11111110",
  50332=>"11111110",
  50333=>"11111111",
  50334=>"11111110",
  50335=>"00000010",
  50336=>"00000000",
  50337=>"11111101",
  50338=>"00000011",
  50339=>"11111100",
  50340=>"00000010",
  50341=>"00000100",
  50342=>"00000100",
  50343=>"00000001",
  50344=>"00000000",
  50345=>"00000011",
  50346=>"00000000",
  50347=>"11111111",
  50348=>"11111110",
  50349=>"11111110",
  50350=>"00000010",
  50351=>"11111111",
  50352=>"11111110",
  50353=>"00000101",
  50354=>"11111110",
  50355=>"11111100",
  50356=>"00000000",
  50357=>"00000010",
  50358=>"00000001",
  50359=>"11111101",
  50360=>"00000000",
  50361=>"00000011",
  50362=>"00000000",
  50363=>"11111101",
  50364=>"00000000",
  50365=>"00000001",
  50366=>"11111101",
  50367=>"00000001",
  50368=>"00000010",
  50369=>"00000011",
  50370=>"00000011",
  50371=>"11111111",
  50372=>"00000011",
  50373=>"00000010",
  50374=>"00000000",
  50375=>"11111111",
  50376=>"00000001",
  50377=>"11111101",
  50378=>"00000001",
  50379=>"00000011",
  50380=>"00000001",
  50381=>"00000000",
  50382=>"11111111",
  50383=>"00000000",
  50384=>"11111111",
  50385=>"00000000",
  50386=>"00000010",
  50387=>"11111110",
  50388=>"00000010",
  50389=>"00000010",
  50390=>"11111100",
  50391=>"11111110",
  50392=>"00000100",
  50393=>"11111111",
  50394=>"00000110",
  50395=>"11111101",
  50396=>"00000010",
  50397=>"00000010",
  50398=>"00000010",
  50399=>"00000000",
  50400=>"00000100",
  50401=>"00000010",
  50402=>"11111101",
  50403=>"00000011",
  50404=>"00000000",
  50405=>"00000010",
  50406=>"11111111",
  50407=>"11111110",
  50408=>"11111111",
  50409=>"00000110",
  50410=>"11111100",
  50411=>"00000011",
  50412=>"11111111",
  50413=>"11111110",
  50414=>"00000001",
  50415=>"00000011",
  50416=>"00000010",
  50417=>"11111111",
  50418=>"11111100",
  50419=>"00000000",
  50420=>"11111111",
  50421=>"11111110",
  50422=>"11111101",
  50423=>"00000011",
  50424=>"11111111",
  50425=>"00000011",
  50426=>"00000100",
  50427=>"00000001",
  50428=>"00000010",
  50429=>"00000001",
  50430=>"00000000",
  50431=>"00000010",
  50432=>"11111111",
  50433=>"11111110",
  50434=>"11111111",
  50435=>"00000010",
  50436=>"11111110",
  50437=>"00000001",
  50438=>"11111101",
  50439=>"11111111",
  50440=>"00000000",
  50441=>"11111100",
  50442=>"11111110",
  50443=>"00000010",
  50444=>"11111111",
  50445=>"00000010",
  50446=>"00000100",
  50447=>"11111101",
  50448=>"11111110",
  50449=>"00000010",
  50450=>"00000011",
  50451=>"00000011",
  50452=>"11111111",
  50453=>"11111110",
  50454=>"00000000",
  50455=>"00000001",
  50456=>"00000001",
  50457=>"00000000",
  50458=>"11111111",
  50459=>"00000010",
  50460=>"11111110",
  50461=>"00000010",
  50462=>"00000000",
  50463=>"00000000",
  50464=>"00000011",
  50465=>"11111101",
  50466=>"00000001",
  50467=>"11111101",
  50468=>"00000011",
  50469=>"00000111",
  50470=>"00000000",
  50471=>"00000001",
  50472=>"00000001",
  50473=>"00000000",
  50474=>"11111111",
  50475=>"11111101",
  50476=>"00000010",
  50477=>"11111111",
  50478=>"00000011",
  50479=>"11111101",
  50480=>"11111101",
  50481=>"00000000",
  50482=>"00000001",
  50483=>"11111110",
  50484=>"00000000",
  50485=>"11111101",
  50486=>"11111101",
  50487=>"11111111",
  50488=>"00000010",
  50489=>"00000010",
  50490=>"11111111",
  50491=>"11111111",
  50492=>"11111110",
  50493=>"00000010",
  50494=>"00000001",
  50495=>"00000011",
  50496=>"11111110",
  50497=>"00000000",
  50498=>"00000010",
  50499=>"00000100",
  50500=>"11111111",
  50501=>"11111111",
  50502=>"11111110",
  50503=>"11111101",
  50504=>"00000100",
  50505=>"00000001",
  50506=>"11111110",
  50507=>"00000001",
  50508=>"11111100",
  50509=>"00000010",
  50510=>"00000000",
  50511=>"00000000",
  50512=>"11111110",
  50513=>"11111111",
  50514=>"00000000",
  50515=>"00000100",
  50516=>"00000000",
  50517=>"00000000",
  50518=>"11111110",
  50519=>"00000000",
  50520=>"11111110",
  50521=>"11111111",
  50522=>"11111111",
  50523=>"11111101",
  50524=>"11111110",
  50525=>"11111110",
  50526=>"00000000",
  50527=>"11111110",
  50528=>"00000011",
  50529=>"11111111",
  50530=>"11111110",
  50531=>"11111110",
  50532=>"11111111",
  50533=>"00000000",
  50534=>"11111111",
  50535=>"00000000",
  50536=>"11111111",
  50537=>"00000000",
  50538=>"00000011",
  50539=>"11111110",
  50540=>"00000011",
  50541=>"11111111",
  50542=>"00000010",
  50543=>"00000010",
  50544=>"00000010",
  50545=>"11111110",
  50546=>"11111111",
  50547=>"11111110",
  50548=>"00000100",
  50549=>"00000011",
  50550=>"00000011",
  50551=>"11111101",
  50552=>"11111101",
  50553=>"11111100",
  50554=>"11111110",
  50555=>"11111111",
  50556=>"11111110",
  50557=>"11111111",
  50558=>"00000010",
  50559=>"11111110",
  50560=>"11111111",
  50561=>"11111110",
  50562=>"11111111",
  50563=>"00000010",
  50564=>"00000001",
  50565=>"00000000",
  50566=>"11111110",
  50567=>"11111110",
  50568=>"11111101",
  50569=>"11111110",
  50570=>"11111111",
  50571=>"00000000",
  50572=>"00000010",
  50573=>"11111110",
  50574=>"11111111",
  50575=>"11111101",
  50576=>"00000000",
  50577=>"00000011",
  50578=>"00000001",
  50579=>"11111110",
  50580=>"00000000",
  50581=>"11111110",
  50582=>"11111110",
  50583=>"00000000",
  50584=>"11111110",
  50585=>"11111111",
  50586=>"11111101",
  50587=>"00000000",
  50588=>"00000010",
  50589=>"00000000",
  50590=>"00000010",
  50591=>"11111101",
  50592=>"11111101",
  50593=>"11111111",
  50594=>"11111101",
  50595=>"00000011",
  50596=>"00000000",
  50597=>"11111110",
  50598=>"11111101",
  50599=>"00000011",
  50600=>"11111111",
  50601=>"11111111",
  50602=>"11111111",
  50603=>"11111100",
  50604=>"00000001",
  50605=>"00000000",
  50606=>"11111110",
  50607=>"11111101",
  50608=>"11111110",
  50609=>"00000010",
  50610=>"11111110",
  50611=>"00000100",
  50612=>"11111110",
  50613=>"00000000",
  50614=>"00000000",
  50615=>"11111110",
  50616=>"11111100",
  50617=>"11111110",
  50618=>"00000011",
  50619=>"00000010",
  50620=>"11111111",
  50621=>"00000011",
  50622=>"11111111",
  50623=>"11111110",
  50624=>"00000011",
  50625=>"11111111",
  50626=>"11111100",
  50627=>"00000011",
  50628=>"00000001",
  50629=>"00000001",
  50630=>"11111111",
  50631=>"11111100",
  50632=>"00000101",
  50633=>"00000010",
  50634=>"11111110",
  50635=>"00000001",
  50636=>"11111110",
  50637=>"11111111",
  50638=>"11111111",
  50639=>"00000001",
  50640=>"11111111",
  50641=>"00000010",
  50642=>"00000001",
  50643=>"11111111",
  50644=>"11111111",
  50645=>"00000101",
  50646=>"00000000",
  50647=>"11111110",
  50648=>"00000000",
  50649=>"11111111",
  50650=>"11111110",
  50651=>"00000001",
  50652=>"11111111",
  50653=>"11111111",
  50654=>"11111100",
  50655=>"11111110",
  50656=>"00000000",
  50657=>"11111111",
  50658=>"00000001",
  50659=>"00000000",
  50660=>"00000000",
  50661=>"00000000",
  50662=>"11111111",
  50663=>"11111111",
  50664=>"11111101",
  50665=>"00000010",
  50666=>"00000000",
  50667=>"11111111",
  50668=>"00000100",
  50669=>"11111111",
  50670=>"11111110",
  50671=>"11111101",
  50672=>"11111101",
  50673=>"00000000",
  50674=>"00000011",
  50675=>"11111111",
  50676=>"00000010",
  50677=>"11111110",
  50678=>"00000001",
  50679=>"11111101",
  50680=>"00000010",
  50681=>"00000010",
  50682=>"00000010",
  50683=>"11111100",
  50684=>"11111100",
  50685=>"00000010",
  50686=>"11111111",
  50687=>"00000011",
  50688=>"11111111",
  50689=>"11111111",
  50690=>"11111101",
  50691=>"00000001",
  50692=>"00000000",
  50693=>"00000001",
  50694=>"11111100",
  50695=>"00000011",
  50696=>"11111111",
  50697=>"00000001",
  50698=>"11111111",
  50699=>"11111110",
  50700=>"11111110",
  50701=>"00000000",
  50702=>"11111111",
  50703=>"11111101",
  50704=>"11111100",
  50705=>"11111101",
  50706=>"00000001",
  50707=>"00000011",
  50708=>"11111110",
  50709=>"11111111",
  50710=>"00000011",
  50711=>"11111101",
  50712=>"11111101",
  50713=>"11111111",
  50714=>"11111110",
  50715=>"11111111",
  50716=>"00000001",
  50717=>"11111110",
  50718=>"00000010",
  50719=>"00000001",
  50720=>"00000001",
  50721=>"11111110",
  50722=>"00000010",
  50723=>"11111110",
  50724=>"00000011",
  50725=>"00000010",
  50726=>"00000101",
  50727=>"11111101",
  50728=>"00000010",
  50729=>"11111101",
  50730=>"00000000",
  50731=>"00000011",
  50732=>"11111111",
  50733=>"00000111",
  50734=>"11111111",
  50735=>"11111111",
  50736=>"11111100",
  50737=>"00000101",
  50738=>"11111110",
  50739=>"11111111",
  50740=>"11111110",
  50741=>"00000010",
  50742=>"00000000",
  50743=>"11111111",
  50744=>"00000001",
  50745=>"00000000",
  50746=>"11111111",
  50747=>"11111111",
  50748=>"00000010",
  50749=>"11111111",
  50750=>"11111110",
  50751=>"11111111",
  50752=>"00000001",
  50753=>"00000010",
  50754=>"00000001",
  50755=>"00000001",
  50756=>"00000011",
  50757=>"00000000",
  50758=>"00000011",
  50759=>"11111111",
  50760=>"00000000",
  50761=>"11111110",
  50762=>"11111111",
  50763=>"00000010",
  50764=>"11111101",
  50765=>"00000001",
  50766=>"11111111",
  50767=>"11111110",
  50768=>"00000001",
  50769=>"00000000",
  50770=>"00000010",
  50771=>"11111110",
  50772=>"11111110",
  50773=>"11111101",
  50774=>"11111111",
  50775=>"00000010",
  50776=>"11111111",
  50777=>"00000001",
  50778=>"11111110",
  50779=>"11111101",
  50780=>"11111101",
  50781=>"11111111",
  50782=>"00000011",
  50783=>"00000100",
  50784=>"11111110",
  50785=>"11111111",
  50786=>"00000000",
  50787=>"00000001",
  50788=>"00000000",
  50789=>"00000100",
  50790=>"00000000",
  50791=>"11111100",
  50792=>"11111100",
  50793=>"00000100",
  50794=>"00000011",
  50795=>"11111110",
  50796=>"00000010",
  50797=>"11111111",
  50798=>"11111111",
  50799=>"11111110",
  50800=>"00000100",
  50801=>"11111101",
  50802=>"11111111",
  50803=>"11111110",
  50804=>"11111110",
  50805=>"00000001",
  50806=>"11111101",
  50807=>"00000000",
  50808=>"11111110",
  50809=>"11111111",
  50810=>"00000010",
  50811=>"11111111",
  50812=>"00000010",
  50813=>"11111111",
  50814=>"11111101",
  50815=>"00000011",
  50816=>"00000000",
  50817=>"11111110",
  50818=>"00000101",
  50819=>"11111101",
  50820=>"11111101",
  50821=>"11111110",
  50822=>"11111110",
  50823=>"11111101",
  50824=>"11111110",
  50825=>"11111111",
  50826=>"11111111",
  50827=>"00000001",
  50828=>"11111111",
  50829=>"00000010",
  50830=>"00000000",
  50831=>"00000000",
  50832=>"00000010",
  50833=>"11111111",
  50834=>"11111110",
  50835=>"00000011",
  50836=>"11111100",
  50837=>"00000000",
  50838=>"00000001",
  50839=>"11111110",
  50840=>"00000010",
  50841=>"11111110",
  50842=>"00000011",
  50843=>"00000001",
  50844=>"00000011",
  50845=>"00000100",
  50846=>"00000000",
  50847=>"00000000",
  50848=>"11111110",
  50849=>"00000000",
  50850=>"00000010",
  50851=>"11111111",
  50852=>"00000011",
  50853=>"00000001",
  50854=>"11111110",
  50855=>"00000100",
  50856=>"00000010",
  50857=>"11111111",
  50858=>"00000001",
  50859=>"11111110",
  50860=>"11111110",
  50861=>"00000001",
  50862=>"00000000",
  50863=>"11111111",
  50864=>"11111111",
  50865=>"11111101",
  50866=>"11111110",
  50867=>"11111111",
  50868=>"00000000",
  50869=>"00000000",
  50870=>"00000001",
  50871=>"00000001",
  50872=>"11111101",
  50873=>"00000000",
  50874=>"11111111",
  50875=>"11111101",
  50876=>"11111110",
  50877=>"00000101",
  50878=>"00000001",
  50879=>"11111110",
  50880=>"11111110",
  50881=>"00000001",
  50882=>"00000010",
  50883=>"11111110",
  50884=>"11111111",
  50885=>"00000011",
  50886=>"00000101",
  50887=>"11111101",
  50888=>"11111100",
  50889=>"00000001",
  50890=>"00000000",
  50891=>"00000000",
  50892=>"11111110",
  50893=>"11111110",
  50894=>"00000011",
  50895=>"00000001",
  50896=>"00000000",
  50897=>"00000000",
  50898=>"11111101",
  50899=>"11111110",
  50900=>"00000000",
  50901=>"00000001",
  50902=>"00000010",
  50903=>"00000000",
  50904=>"11111110",
  50905=>"00000101",
  50906=>"00000010",
  50907=>"11111111",
  50908=>"00000010",
  50909=>"11111111",
  50910=>"00000001",
  50911=>"11111101",
  50912=>"00000000",
  50913=>"11111110",
  50914=>"11111100",
  50915=>"00000001",
  50916=>"00000010",
  50917=>"11111101",
  50918=>"00000101",
  50919=>"11111101",
  50920=>"00000001",
  50921=>"00000001",
  50922=>"00000000",
  50923=>"11111110",
  50924=>"00000001",
  50925=>"11111101",
  50926=>"00000010",
  50927=>"11111101",
  50928=>"11111101",
  50929=>"11111101",
  50930=>"00000000",
  50931=>"00000001",
  50932=>"00000001",
  50933=>"11111111",
  50934=>"11111110",
  50935=>"00000100",
  50936=>"11111111",
  50937=>"00000000",
  50938=>"00000000",
  50939=>"00000011",
  50940=>"11111110",
  50941=>"11111110",
  50942=>"00000011",
  50943=>"00000011",
  50944=>"11111110",
  50945=>"00000010",
  50946=>"11111111",
  50947=>"11111110",
  50948=>"11111101",
  50949=>"11111111",
  50950=>"00000000",
  50951=>"00000010",
  50952=>"00000001",
  50953=>"00000010",
  50954=>"11111100",
  50955=>"11111111",
  50956=>"11111100",
  50957=>"00000010",
  50958=>"00000001",
  50959=>"11111111",
  50960=>"00000110",
  50961=>"11111111",
  50962=>"00000011",
  50963=>"00000011",
  50964=>"11111110",
  50965=>"00000011",
  50966=>"00000000",
  50967=>"11111111",
  50968=>"00000101",
  50969=>"00000101",
  50970=>"11111110",
  50971=>"00000100",
  50972=>"11111101",
  50973=>"11111101",
  50974=>"11111111",
  50975=>"00000000",
  50976=>"11111110",
  50977=>"11111101",
  50978=>"00000010",
  50979=>"11111110",
  50980=>"11111111",
  50981=>"11111110",
  50982=>"11111101",
  50983=>"11111111",
  50984=>"00000101",
  50985=>"11111100",
  50986=>"00000010",
  50987=>"11111101",
  50988=>"00000111",
  50989=>"00000010",
  50990=>"11111110",
  50991=>"00000011",
  50992=>"00000010",
  50993=>"00000010",
  50994=>"00000000",
  50995=>"11111101",
  50996=>"00000010",
  50997=>"11111110",
  50998=>"00000000",
  50999=>"00000000",
  51000=>"11111110",
  51001=>"00000010",
  51002=>"11111110",
  51003=>"11111110",
  51004=>"11111101",
  51005=>"00000010",
  51006=>"00000010",
  51007=>"00000000",
  51008=>"00000001",
  51009=>"00000001",
  51010=>"00000000",
  51011=>"11111101",
  51012=>"00000001",
  51013=>"00000000",
  51014=>"00000001",
  51015=>"00000001",
  51016=>"00000001",
  51017=>"00000000",
  51018=>"00000000",
  51019=>"00000000",
  51020=>"11111110",
  51021=>"00000001",
  51022=>"11111111",
  51023=>"00000001",
  51024=>"00000100",
  51025=>"11111101",
  51026=>"00000100",
  51027=>"00000001",
  51028=>"00000000",
  51029=>"00000000",
  51030=>"00000011",
  51031=>"00000010",
  51032=>"11111101",
  51033=>"11111110",
  51034=>"11111101",
  51035=>"11111111",
  51036=>"00000001",
  51037=>"11111111",
  51038=>"00000000",
  51039=>"00000000",
  51040=>"00000001",
  51041=>"00000010",
  51042=>"00000011",
  51043=>"00000000",
  51044=>"11111111",
  51045=>"11111110",
  51046=>"11111101",
  51047=>"00000010",
  51048=>"00000000",
  51049=>"00000010",
  51050=>"00000000",
  51051=>"00000010",
  51052=>"00000001",
  51053=>"00000011",
  51054=>"00000100",
  51055=>"11111110",
  51056=>"11111101",
  51057=>"00000001",
  51058=>"00000001",
  51059=>"00000001",
  51060=>"00000001",
  51061=>"00000000",
  51062=>"11111111",
  51063=>"11111101",
  51064=>"00000001",
  51065=>"00000000",
  51066=>"11111111",
  51067=>"00000000",
  51068=>"00000000",
  51069=>"00000010",
  51070=>"11111100",
  51071=>"11111111",
  51072=>"00000010",
  51073=>"00000011",
  51074=>"00000011",
  51075=>"00000000",
  51076=>"11111101",
  51077=>"00000100",
  51078=>"11111111",
  51079=>"00000000",
  51080=>"00000001",
  51081=>"00000001",
  51082=>"11111111",
  51083=>"11111111",
  51084=>"00000000",
  51085=>"00000011",
  51086=>"11111110",
  51087=>"00000100",
  51088=>"00000000",
  51089=>"11111110",
  51090=>"11111111",
  51091=>"11111111",
  51092=>"00000001",
  51093=>"00000100",
  51094=>"11111111",
  51095=>"11111111",
  51096=>"11111110",
  51097=>"00000001",
  51098=>"00000101",
  51099=>"00000101",
  51100=>"00000001",
  51101=>"00000010",
  51102=>"00000000",
  51103=>"00000001",
  51104=>"00000001",
  51105=>"11111111",
  51106=>"00000100",
  51107=>"00000010",
  51108=>"11111110",
  51109=>"11111110",
  51110=>"00000010",
  51111=>"00000010",
  51112=>"11111101",
  51113=>"00000011",
  51114=>"11111101",
  51115=>"00000001",
  51116=>"00000011",
  51117=>"11111111",
  51118=>"00000001",
  51119=>"11111110",
  51120=>"00000000",
  51121=>"11111110",
  51122=>"11111110",
  51123=>"00000000",
  51124=>"00000011",
  51125=>"00000100",
  51126=>"11111110",
  51127=>"11111111",
  51128=>"00000010",
  51129=>"11111100",
  51130=>"11111110",
  51131=>"11111111",
  51132=>"00000010",
  51133=>"00000000",
  51134=>"00000100",
  51135=>"00000000",
  51136=>"11111110",
  51137=>"00000011",
  51138=>"00000000",
  51139=>"11111110",
  51140=>"11111110",
  51141=>"11111101",
  51142=>"11111111",
  51143=>"11111111",
  51144=>"00000100",
  51145=>"11111111",
  51146=>"11111101",
  51147=>"00000001",
  51148=>"00000001",
  51149=>"00000010",
  51150=>"00000101",
  51151=>"00000000",
  51152=>"00000011",
  51153=>"11111111",
  51154=>"11111100",
  51155=>"00000010",
  51156=>"11111111",
  51157=>"11111110",
  51158=>"11111110",
  51159=>"00000011",
  51160=>"11111111",
  51161=>"11111111",
  51162=>"11111110",
  51163=>"11111110",
  51164=>"11111101",
  51165=>"11111110",
  51166=>"00000001",
  51167=>"11111111",
  51168=>"11111110",
  51169=>"11111111",
  51170=>"00000010",
  51171=>"11111111",
  51172=>"11111111",
  51173=>"00000100",
  51174=>"11111111",
  51175=>"11111110",
  51176=>"11111101",
  51177=>"00000000",
  51178=>"11111101",
  51179=>"11111100",
  51180=>"11111111",
  51181=>"00000101",
  51182=>"00000001",
  51183=>"11111110",
  51184=>"11111110",
  51185=>"00000011",
  51186=>"11111110",
  51187=>"00000001",
  51188=>"11111101",
  51189=>"11111110",
  51190=>"00000000",
  51191=>"00000000",
  51192=>"00000011",
  51193=>"00000000",
  51194=>"11111111",
  51195=>"11111110",
  51196=>"00000101",
  51197=>"11111101",
  51198=>"11111111",
  51199=>"00000011",
  51200=>"00000001",
  51201=>"11111110",
  51202=>"11111100",
  51203=>"11111110",
  51204=>"00000011",
  51205=>"11111111",
  51206=>"00000000",
  51207=>"11111111",
  51208=>"11111100",
  51209=>"00000000",
  51210=>"11111110",
  51211=>"11111111",
  51212=>"11111101",
  51213=>"00000100",
  51214=>"00000010",
  51215=>"00000100",
  51216=>"11111111",
  51217=>"00000001",
  51218=>"11111101",
  51219=>"00000001",
  51220=>"11111111",
  51221=>"00000001",
  51222=>"11111110",
  51223=>"11111101",
  51224=>"11111110",
  51225=>"00000001",
  51226=>"11111111",
  51227=>"11111101",
  51228=>"11111101",
  51229=>"00000011",
  51230=>"00000010",
  51231=>"00000010",
  51232=>"00000010",
  51233=>"11111101",
  51234=>"00000100",
  51235=>"00000100",
  51236=>"00000010",
  51237=>"00000000",
  51238=>"11111101",
  51239=>"00000010",
  51240=>"00000101",
  51241=>"11111110",
  51242=>"11111100",
  51243=>"11111111",
  51244=>"00000011",
  51245=>"00000010",
  51246=>"00000011",
  51247=>"00000001",
  51248=>"00000000",
  51249=>"11111111",
  51250=>"11111101",
  51251=>"00000101",
  51252=>"00000001",
  51253=>"11111111",
  51254=>"11111111",
  51255=>"00000011",
  51256=>"00000010",
  51257=>"00000000",
  51258=>"11111110",
  51259=>"00000100",
  51260=>"00000000",
  51261=>"00000011",
  51262=>"00000001",
  51263=>"11111111",
  51264=>"00000010",
  51265=>"00000010",
  51266=>"11111101",
  51267=>"00000010",
  51268=>"11111111",
  51269=>"11111110",
  51270=>"00000010",
  51271=>"11111110",
  51272=>"11111111",
  51273=>"11111111",
  51274=>"00000010",
  51275=>"00000000",
  51276=>"11111110",
  51277=>"11111111",
  51278=>"00000011",
  51279=>"00000011",
  51280=>"00000000",
  51281=>"11111110",
  51282=>"00000110",
  51283=>"11111111",
  51284=>"00000001",
  51285=>"11111110",
  51286=>"11111111",
  51287=>"00000000",
  51288=>"00000010",
  51289=>"00000001",
  51290=>"00000000",
  51291=>"00000010",
  51292=>"11111111",
  51293=>"11111110",
  51294=>"11111110",
  51295=>"00000000",
  51296=>"11111101",
  51297=>"00000000",
  51298=>"00000111",
  51299=>"11111110",
  51300=>"00000000",
  51301=>"11111110",
  51302=>"11111111",
  51303=>"11111101",
  51304=>"00000010",
  51305=>"00000100",
  51306=>"00000001",
  51307=>"00000010",
  51308=>"00000001",
  51309=>"11111111",
  51310=>"00000110",
  51311=>"00000011",
  51312=>"00000010",
  51313=>"00000010",
  51314=>"11111111",
  51315=>"11111100",
  51316=>"00000001",
  51317=>"00000101",
  51318=>"00000000",
  51319=>"11111110",
  51320=>"00000000",
  51321=>"11111101",
  51322=>"11111101",
  51323=>"00000000",
  51324=>"11111111",
  51325=>"11111110",
  51326=>"00000100",
  51327=>"00000001",
  51328=>"00000001",
  51329=>"00000001",
  51330=>"00000000",
  51331=>"00000000",
  51332=>"00000010",
  51333=>"11111110",
  51334=>"11111111",
  51335=>"11111111",
  51336=>"11111101",
  51337=>"00000001",
  51338=>"11111111",
  51339=>"11111110",
  51340=>"11111101",
  51341=>"11111101",
  51342=>"00000000",
  51343=>"00000101",
  51344=>"00000000",
  51345=>"00000011",
  51346=>"00000010",
  51347=>"11111110",
  51348=>"00000000",
  51349=>"11111110",
  51350=>"00000001",
  51351=>"00000110",
  51352=>"11111111",
  51353=>"00000010",
  51354=>"11111111",
  51355=>"00000010",
  51356=>"11111110",
  51357=>"11111111",
  51358=>"11111110",
  51359=>"00000011",
  51360=>"11111111",
  51361=>"11111101",
  51362=>"11111111",
  51363=>"11111111",
  51364=>"11111110",
  51365=>"00000010",
  51366=>"00000011",
  51367=>"11111111",
  51368=>"00000001",
  51369=>"11111111",
  51370=>"00000001",
  51371=>"00000010",
  51372=>"11111110",
  51373=>"00000010",
  51374=>"11111111",
  51375=>"11111101",
  51376=>"00000000",
  51377=>"11111110",
  51378=>"00000000",
  51379=>"11111110",
  51380=>"00000000",
  51381=>"11111110",
  51382=>"11111100",
  51383=>"00000000",
  51384=>"11111101",
  51385=>"00000010",
  51386=>"11111110",
  51387=>"11111111",
  51388=>"11111110",
  51389=>"00000000",
  51390=>"11111111",
  51391=>"00000001",
  51392=>"00000000",
  51393=>"00000000",
  51394=>"11111101",
  51395=>"00000001",
  51396=>"11111101",
  51397=>"11111110",
  51398=>"00000001",
  51399=>"00000010",
  51400=>"00000000",
  51401=>"11111110",
  51402=>"11111110",
  51403=>"00000011",
  51404=>"11111100",
  51405=>"11111111",
  51406=>"00000010",
  51407=>"00000010",
  51408=>"00000000",
  51409=>"11111110",
  51410=>"00000010",
  51411=>"11111111",
  51412=>"00000000",
  51413=>"11111100",
  51414=>"11111111",
  51415=>"00000000",
  51416=>"00000011",
  51417=>"00000011",
  51418=>"00000010",
  51419=>"00000001",
  51420=>"00000000",
  51421=>"11111110",
  51422=>"00000000",
  51423=>"00000100",
  51424=>"11111111",
  51425=>"00000001",
  51426=>"00000000",
  51427=>"00000001",
  51428=>"00000001",
  51429=>"11111110",
  51430=>"11111110",
  51431=>"11111111",
  51432=>"00000000",
  51433=>"11111111",
  51434=>"00000010",
  51435=>"00000001",
  51436=>"00000011",
  51437=>"00000000",
  51438=>"11111110",
  51439=>"00000000",
  51440=>"00000011",
  51441=>"11111100",
  51442=>"00000010",
  51443=>"11111110",
  51444=>"11111110",
  51445=>"00000000",
  51446=>"00000011",
  51447=>"00000010",
  51448=>"11111101",
  51449=>"00000000",
  51450=>"00000001",
  51451=>"00000000",
  51452=>"00000001",
  51453=>"11111111",
  51454=>"11111110",
  51455=>"00000000",
  51456=>"11111110",
  51457=>"00000100",
  51458=>"11111110",
  51459=>"11111101",
  51460=>"11111111",
  51461=>"00000000",
  51462=>"11111101",
  51463=>"00000011",
  51464=>"11111101",
  51465=>"00000001",
  51466=>"11111110",
  51467=>"11111101",
  51468=>"11111111",
  51469=>"00000011",
  51470=>"11111111",
  51471=>"11111101",
  51472=>"00000101",
  51473=>"11111111",
  51474=>"11111110",
  51475=>"00000011",
  51476=>"00000111",
  51477=>"11111111",
  51478=>"00000000",
  51479=>"00000011",
  51480=>"00000101",
  51481=>"00000001",
  51482=>"00000000",
  51483=>"00000010",
  51484=>"00000001",
  51485=>"00000010",
  51486=>"00000000",
  51487=>"11111100",
  51488=>"00000010",
  51489=>"00000011",
  51490=>"11111110",
  51491=>"11111100",
  51492=>"11111111",
  51493=>"11111111",
  51494=>"00000001",
  51495=>"00000011",
  51496=>"11111100",
  51497=>"11111101",
  51498=>"11111111",
  51499=>"11111111",
  51500=>"00000001",
  51501=>"11111110",
  51502=>"00000000",
  51503=>"00000000",
  51504=>"00000000",
  51505=>"00000011",
  51506=>"11111110",
  51507=>"11111110",
  51508=>"11111100",
  51509=>"00000011",
  51510=>"11111111",
  51511=>"00000100",
  51512=>"11111111",
  51513=>"00000011",
  51514=>"00000010",
  51515=>"11111110",
  51516=>"00000010",
  51517=>"11111111",
  51518=>"11111111",
  51519=>"00000001",
  51520=>"00000010",
  51521=>"11111111",
  51522=>"00000001",
  51523=>"11111110",
  51524=>"00000010",
  51525=>"00000000",
  51526=>"00000000",
  51527=>"00000011",
  51528=>"11111111",
  51529=>"11111110",
  51530=>"00000000",
  51531=>"11111110",
  51532=>"11111111",
  51533=>"00000011",
  51534=>"00000000",
  51535=>"00000111",
  51536=>"00000000",
  51537=>"00000001",
  51538=>"11111101",
  51539=>"00000011",
  51540=>"00000010",
  51541=>"00000100",
  51542=>"00000010",
  51543=>"11111101",
  51544=>"00000000",
  51545=>"11111110",
  51546=>"00000010",
  51547=>"11111111",
  51548=>"00000001",
  51549=>"00000001",
  51550=>"00000100",
  51551=>"11111111",
  51552=>"11111110",
  51553=>"00000010",
  51554=>"00000001",
  51555=>"11111111",
  51556=>"00000011",
  51557=>"11111111",
  51558=>"11111110",
  51559=>"00000000",
  51560=>"00000001",
  51561=>"00000001",
  51562=>"00000001",
  51563=>"00000100",
  51564=>"00000000",
  51565=>"11111110",
  51566=>"00000010",
  51567=>"11111110",
  51568=>"00000011",
  51569=>"00000101",
  51570=>"00000000",
  51571=>"00000010",
  51572=>"11111111",
  51573=>"00000010",
  51574=>"00000010",
  51575=>"11111101",
  51576=>"00000101",
  51577=>"11111110",
  51578=>"00000001",
  51579=>"11111111",
  51580=>"00000101",
  51581=>"11111110",
  51582=>"11111101",
  51583=>"11111110",
  51584=>"00000011",
  51585=>"00000010",
  51586=>"00000001",
  51587=>"00000000",
  51588=>"11111101",
  51589=>"00000010",
  51590=>"00000011",
  51591=>"00000001",
  51592=>"00000001",
  51593=>"11111110",
  51594=>"11111110",
  51595=>"11111110",
  51596=>"00000000",
  51597=>"11111110",
  51598=>"11111111",
  51599=>"00000011",
  51600=>"11111110",
  51601=>"00000001",
  51602=>"11111111",
  51603=>"00000011",
  51604=>"00000000",
  51605=>"11111110",
  51606=>"00000000",
  51607=>"11111111",
  51608=>"00000000",
  51609=>"11111101",
  51610=>"00000100",
  51611=>"11111110",
  51612=>"11111111",
  51613=>"00000011",
  51614=>"11111111",
  51615=>"11111100",
  51616=>"00000000",
  51617=>"11111101",
  51618=>"00000001",
  51619=>"00000000",
  51620=>"11111110",
  51621=>"00000001",
  51622=>"11111101",
  51623=>"00000010",
  51624=>"11111011",
  51625=>"11111111",
  51626=>"00000000",
  51627=>"00000011",
  51628=>"00000000",
  51629=>"00000001",
  51630=>"11111111",
  51631=>"00000010",
  51632=>"00000011",
  51633=>"00000000",
  51634=>"11111111",
  51635=>"11111110",
  51636=>"00000101",
  51637=>"11111110",
  51638=>"00000010",
  51639=>"00000100",
  51640=>"11111110",
  51641=>"11111111",
  51642=>"11111101",
  51643=>"00000001",
  51644=>"11111101",
  51645=>"11111111",
  51646=>"00000000",
  51647=>"00000000",
  51648=>"00000000",
  51649=>"11111111",
  51650=>"11111100",
  51651=>"00000000",
  51652=>"00000011",
  51653=>"11111110",
  51654=>"11111110",
  51655=>"00000101",
  51656=>"00000100",
  51657=>"00000010",
  51658=>"00000000",
  51659=>"11111110",
  51660=>"00000011",
  51661=>"00000100",
  51662=>"00000011",
  51663=>"11111111",
  51664=>"00000000",
  51665=>"11111110",
  51666=>"00000001",
  51667=>"11111111",
  51668=>"11111111",
  51669=>"00000001",
  51670=>"11111111",
  51671=>"00000001",
  51672=>"00000001",
  51673=>"00000000",
  51674=>"00000000",
  51675=>"11111111",
  51676=>"00000110",
  51677=>"00000010",
  51678=>"11111100",
  51679=>"00000100",
  51680=>"00000001",
  51681=>"11111100",
  51682=>"11111110",
  51683=>"11111101",
  51684=>"11111110",
  51685=>"00000000",
  51686=>"11111110",
  51687=>"00000001",
  51688=>"00000010",
  51689=>"00000100",
  51690=>"00000011",
  51691=>"11111101",
  51692=>"00000001",
  51693=>"00000010",
  51694=>"00000001",
  51695=>"11111101",
  51696=>"11111110",
  51697=>"11111111",
  51698=>"00000010",
  51699=>"00000000",
  51700=>"00000011",
  51701=>"00000011",
  51702=>"00000000",
  51703=>"11111111",
  51704=>"00000000",
  51705=>"00000001",
  51706=>"00000010",
  51707=>"11111111",
  51708=>"00000010",
  51709=>"00000000",
  51710=>"11111100",
  51711=>"00000001",
  51712=>"00000010",
  51713=>"11111110",
  51714=>"11111100",
  51715=>"00000010",
  51716=>"00000000",
  51717=>"11111101",
  51718=>"00000001",
  51719=>"11111011",
  51720=>"00000001",
  51721=>"00000000",
  51722=>"11111101",
  51723=>"00000001",
  51724=>"11111111",
  51725=>"00000001",
  51726=>"00000110",
  51727=>"00000011",
  51728=>"11111101",
  51729=>"11111111",
  51730=>"00000000",
  51731=>"00000011",
  51732=>"00000011",
  51733=>"00000100",
  51734=>"00000000",
  51735=>"00000011",
  51736=>"00000000",
  51737=>"00000010",
  51738=>"11111111",
  51739=>"11111110",
  51740=>"00000010",
  51741=>"00000000",
  51742=>"11111101",
  51743=>"00000100",
  51744=>"00000001",
  51745=>"11111110",
  51746=>"00000001",
  51747=>"11111110",
  51748=>"00000000",
  51749=>"11111110",
  51750=>"00000000",
  51751=>"11111110",
  51752=>"00000011",
  51753=>"11111110",
  51754=>"00000100",
  51755=>"11111111",
  51756=>"00000000",
  51757=>"00000011",
  51758=>"00000000",
  51759=>"11111111",
  51760=>"00000011",
  51761=>"11111101",
  51762=>"11111111",
  51763=>"11111110",
  51764=>"00000101",
  51765=>"11111110",
  51766=>"11111100",
  51767=>"00000000",
  51768=>"11111111",
  51769=>"11111110",
  51770=>"00000001",
  51771=>"00000000",
  51772=>"00000011",
  51773=>"00000100",
  51774=>"00000010",
  51775=>"00000000",
  51776=>"00000010",
  51777=>"00000000",
  51778=>"00000011",
  51779=>"00000001",
  51780=>"00000011",
  51781=>"11111110",
  51782=>"00000000",
  51783=>"00000000",
  51784=>"00000010",
  51785=>"00000000",
  51786=>"00000001",
  51787=>"11111100",
  51788=>"00000000",
  51789=>"00000000",
  51790=>"00000001",
  51791=>"00000010",
  51792=>"00000001",
  51793=>"00000100",
  51794=>"00000010",
  51795=>"00000001",
  51796=>"11111110",
  51797=>"00000011",
  51798=>"11111101",
  51799=>"11111111",
  51800=>"00000000",
  51801=>"11111100",
  51802=>"00000001",
  51803=>"11111100",
  51804=>"00000010",
  51805=>"11111111",
  51806=>"00000001",
  51807=>"00000101",
  51808=>"00000011",
  51809=>"11111111",
  51810=>"11111101",
  51811=>"00000000",
  51812=>"00000000",
  51813=>"00000100",
  51814=>"00000000",
  51815=>"00000101",
  51816=>"11111110",
  51817=>"00000000",
  51818=>"00000000",
  51819=>"00000000",
  51820=>"11111110",
  51821=>"00000100",
  51822=>"00000001",
  51823=>"11111101",
  51824=>"11111110",
  51825=>"11111101",
  51826=>"00000101",
  51827=>"00000010",
  51828=>"00000010",
  51829=>"11111101",
  51830=>"00000100",
  51831=>"00000000",
  51832=>"11111110",
  51833=>"00000000",
  51834=>"11111101",
  51835=>"11111100",
  51836=>"11111110",
  51837=>"00000010",
  51838=>"00000110",
  51839=>"11111101",
  51840=>"11111110",
  51841=>"11111110",
  51842=>"00000011",
  51843=>"00000100",
  51844=>"00000110",
  51845=>"11111101",
  51846=>"11111110",
  51847=>"11111101",
  51848=>"00000001",
  51849=>"00000010",
  51850=>"00000001",
  51851=>"00000000",
  51852=>"00000000",
  51853=>"00000010",
  51854=>"11111101",
  51855=>"00000101",
  51856=>"11111101",
  51857=>"00000000",
  51858=>"11111111",
  51859=>"00000011",
  51860=>"11111110",
  51861=>"00000001",
  51862=>"11111101",
  51863=>"11111110",
  51864=>"11111111",
  51865=>"11111111",
  51866=>"11111111",
  51867=>"11111101",
  51868=>"11111110",
  51869=>"00000001",
  51870=>"11111111",
  51871=>"11111110",
  51872=>"00000000",
  51873=>"00000011",
  51874=>"11111101",
  51875=>"00000000",
  51876=>"11111101",
  51877=>"11111110",
  51878=>"00000001",
  51879=>"00000101",
  51880=>"11111100",
  51881=>"11111101",
  51882=>"11111101",
  51883=>"00000010",
  51884=>"11111101",
  51885=>"00000000",
  51886=>"00000001",
  51887=>"11111101",
  51888=>"00000100",
  51889=>"11111100",
  51890=>"11111101",
  51891=>"00000011",
  51892=>"00000000",
  51893=>"11111101",
  51894=>"11111110",
  51895=>"11111111",
  51896=>"00000001",
  51897=>"00000001",
  51898=>"00000001",
  51899=>"00000001",
  51900=>"11111100",
  51901=>"00001000",
  51902=>"11111101",
  51903=>"00000010",
  51904=>"00000011",
  51905=>"11111111",
  51906=>"11111110",
  51907=>"00000011",
  51908=>"00000000",
  51909=>"00000100",
  51910=>"00000011",
  51911=>"00000001",
  51912=>"00000101",
  51913=>"00000110",
  51914=>"11111110",
  51915=>"11111101",
  51916=>"11111111",
  51917=>"00000001",
  51918=>"11111111",
  51919=>"11111100",
  51920=>"00000010",
  51921=>"11111110",
  51922=>"00000100",
  51923=>"00000000",
  51924=>"11111111",
  51925=>"11111110",
  51926=>"00000010",
  51927=>"11111100",
  51928=>"00000100",
  51929=>"00000001",
  51930=>"00000010",
  51931=>"11111101",
  51932=>"00000010",
  51933=>"00000010",
  51934=>"00000001",
  51935=>"11111111",
  51936=>"00000100",
  51937=>"00000011",
  51938=>"11111111",
  51939=>"00000000",
  51940=>"00000000",
  51941=>"11111111",
  51942=>"11111110",
  51943=>"00000010",
  51944=>"11111110",
  51945=>"11111110",
  51946=>"00000001",
  51947=>"00000001",
  51948=>"00000010",
  51949=>"00000010",
  51950=>"00000100",
  51951=>"11111111",
  51952=>"00000100",
  51953=>"00000001",
  51954=>"00000010",
  51955=>"11111111",
  51956=>"00000000",
  51957=>"00000011",
  51958=>"00000000",
  51959=>"11111100",
  51960=>"11111111",
  51961=>"11111110",
  51962=>"11111110",
  51963=>"00000010",
  51964=>"11111110",
  51965=>"00000011",
  51966=>"00000000",
  51967=>"11111101",
  51968=>"00000001",
  51969=>"00000001",
  51970=>"00000000",
  51971=>"11111111",
  51972=>"11111110",
  51973=>"00000001",
  51974=>"00000011",
  51975=>"00000001",
  51976=>"00000010",
  51977=>"00000010",
  51978=>"11111101",
  51979=>"00000111",
  51980=>"11111110",
  51981=>"11111100",
  51982=>"11111101",
  51983=>"11111110",
  51984=>"00000101",
  51985=>"00000010",
  51986=>"00000001",
  51987=>"00000010",
  51988=>"00000001",
  51989=>"11111111",
  51990=>"00001000",
  51991=>"00000011",
  51992=>"11111110",
  51993=>"11111100",
  51994=>"00000000",
  51995=>"00000000",
  51996=>"11111101",
  51997=>"00000010",
  51998=>"00000000",
  51999=>"00000100",
  52000=>"00000010",
  52001=>"11111101",
  52002=>"11111111",
  52003=>"00000011",
  52004=>"00000000",
  52005=>"11111101",
  52006=>"11111110",
  52007=>"00000010",
  52008=>"00000100",
  52009=>"00000010",
  52010=>"11111111",
  52011=>"11111110",
  52012=>"11111111",
  52013=>"11111110",
  52014=>"00000000",
  52015=>"00000000",
  52016=>"11111111",
  52017=>"11111101",
  52018=>"11111100",
  52019=>"00000101",
  52020=>"11111111",
  52021=>"11111101",
  52022=>"00000010",
  52023=>"00000011",
  52024=>"11111110",
  52025=>"11111111",
  52026=>"11111110",
  52027=>"00000001",
  52028=>"11111101",
  52029=>"00000001",
  52030=>"11111101",
  52031=>"00000101",
  52032=>"00000001",
  52033=>"00000010",
  52034=>"00000010",
  52035=>"11111101",
  52036=>"11111101",
  52037=>"11111110",
  52038=>"00000010",
  52039=>"00000011",
  52040=>"11111111",
  52041=>"00000011",
  52042=>"11111101",
  52043=>"11111100",
  52044=>"11111110",
  52045=>"00000001",
  52046=>"11111110",
  52047=>"11111111",
  52048=>"00000011",
  52049=>"00000000",
  52050=>"11111111",
  52051=>"00000011",
  52052=>"00000011",
  52053=>"11111101",
  52054=>"00000001",
  52055=>"00000111",
  52056=>"00000000",
  52057=>"00000000",
  52058=>"00000001",
  52059=>"00000001",
  52060=>"11111110",
  52061=>"00000011",
  52062=>"00000001",
  52063=>"00000011",
  52064=>"11111101",
  52065=>"11111110",
  52066=>"00000100",
  52067=>"11111110",
  52068=>"11111110",
  52069=>"00000010",
  52070=>"11111101",
  52071=>"11111100",
  52072=>"00000000",
  52073=>"11111111",
  52074=>"11111110",
  52075=>"00000000",
  52076=>"00000010",
  52077=>"11111111",
  52078=>"11111111",
  52079=>"00000011",
  52080=>"00000100",
  52081=>"00000000",
  52082=>"00000001",
  52083=>"00000001",
  52084=>"00000000",
  52085=>"11111101",
  52086=>"00000000",
  52087=>"11111110",
  52088=>"00000101",
  52089=>"00000001",
  52090=>"00000010",
  52091=>"11111110",
  52092=>"11111111",
  52093=>"11111111",
  52094=>"00000011",
  52095=>"00000011",
  52096=>"00000001",
  52097=>"00000110",
  52098=>"11111101",
  52099=>"11111111",
  52100=>"11111111",
  52101=>"11111110",
  52102=>"11111111",
  52103=>"00000001",
  52104=>"00000001",
  52105=>"11111110",
  52106=>"00000000",
  52107=>"00000011",
  52108=>"00000001",
  52109=>"00000001",
  52110=>"11111110",
  52111=>"00000011",
  52112=>"11111101",
  52113=>"00000101",
  52114=>"00000001",
  52115=>"00000001",
  52116=>"11111111",
  52117=>"00000010",
  52118=>"00000001",
  52119=>"11111100",
  52120=>"00000001",
  52121=>"11111110",
  52122=>"00000000",
  52123=>"11111110",
  52124=>"00000010",
  52125=>"11111100",
  52126=>"11111100",
  52127=>"00000000",
  52128=>"00001000",
  52129=>"11111110",
  52130=>"00000011",
  52131=>"00000000",
  52132=>"11111111",
  52133=>"00000001",
  52134=>"11111110",
  52135=>"00000001",
  52136=>"11111110",
  52137=>"00000001",
  52138=>"11111111",
  52139=>"00000011",
  52140=>"00000000",
  52141=>"00000000",
  52142=>"00000001",
  52143=>"00000000",
  52144=>"11111111",
  52145=>"11111110",
  52146=>"11111100",
  52147=>"11111111",
  52148=>"00000100",
  52149=>"00000101",
  52150=>"00000000",
  52151=>"00000001",
  52152=>"11111101",
  52153=>"00000000",
  52154=>"11111110",
  52155=>"00000010",
  52156=>"00000001",
  52157=>"11111111",
  52158=>"11111111",
  52159=>"00000001",
  52160=>"00000010",
  52161=>"00000010",
  52162=>"11111111",
  52163=>"00000000",
  52164=>"00000010",
  52165=>"00000000",
  52166=>"11111111",
  52167=>"11111101",
  52168=>"00000011",
  52169=>"00000010",
  52170=>"11111100",
  52171=>"11111101",
  52172=>"11111110",
  52173=>"00000010",
  52174=>"00000000",
  52175=>"00000010",
  52176=>"00000010",
  52177=>"11111111",
  52178=>"00000011",
  52179=>"00000001",
  52180=>"11111111",
  52181=>"11111100",
  52182=>"11111111",
  52183=>"11111111",
  52184=>"00000001",
  52185=>"00000000",
  52186=>"00000001",
  52187=>"11111111",
  52188=>"00000011",
  52189=>"00000011",
  52190=>"11111111",
  52191=>"11111110",
  52192=>"00000000",
  52193=>"11111110",
  52194=>"00000010",
  52195=>"00000000",
  52196=>"00000010",
  52197=>"11111110",
  52198=>"11111111",
  52199=>"11111111",
  52200=>"00000011",
  52201=>"00000010",
  52202=>"11111111",
  52203=>"00000000",
  52204=>"11111110",
  52205=>"00000100",
  52206=>"11111111",
  52207=>"00000100",
  52208=>"00000000",
  52209=>"11111110",
  52210=>"00000000",
  52211=>"00000011",
  52212=>"11111111",
  52213=>"11111101",
  52214=>"11111111",
  52215=>"00000110",
  52216=>"00000001",
  52217=>"00000011",
  52218=>"11111101",
  52219=>"00000000",
  52220=>"00000010",
  52221=>"11111110",
  52222=>"00000011",
  52223=>"11111111",
  52224=>"00000000",
  52225=>"00000001",
  52226=>"00000100",
  52227=>"00000000",
  52228=>"00000000",
  52229=>"11111111",
  52230=>"00000010",
  52231=>"00000001",
  52232=>"00000001",
  52233=>"11111110",
  52234=>"00000010",
  52235=>"11111101",
  52236=>"11111101",
  52237=>"00000000",
  52238=>"11111101",
  52239=>"00000011",
  52240=>"00000001",
  52241=>"00000000",
  52242=>"00000001",
  52243=>"11111101",
  52244=>"00000000",
  52245=>"11111101",
  52246=>"11111110",
  52247=>"00000001",
  52248=>"11111110",
  52249=>"11111111",
  52250=>"11111101",
  52251=>"00000010",
  52252=>"00000101",
  52253=>"00000010",
  52254=>"11111110",
  52255=>"11111110",
  52256=>"11111111",
  52257=>"11111101",
  52258=>"00000110",
  52259=>"11111110",
  52260=>"00000000",
  52261=>"00000000",
  52262=>"00000100",
  52263=>"11111111",
  52264=>"00000011",
  52265=>"00000011",
  52266=>"11111111",
  52267=>"11111101",
  52268=>"11111111",
  52269=>"00000000",
  52270=>"00000001",
  52271=>"11111110",
  52272=>"11111110",
  52273=>"11111111",
  52274=>"11111111",
  52275=>"11111101",
  52276=>"11111111",
  52277=>"11111110",
  52278=>"00000000",
  52279=>"11111111",
  52280=>"00000001",
  52281=>"00000011",
  52282=>"11111111",
  52283=>"00000000",
  52284=>"00000000",
  52285=>"00000000",
  52286=>"11111101",
  52287=>"11111101",
  52288=>"00000001",
  52289=>"00000001",
  52290=>"11111110",
  52291=>"11111110",
  52292=>"00000001",
  52293=>"11111110",
  52294=>"11111111",
  52295=>"11111111",
  52296=>"11111110",
  52297=>"11111110",
  52298=>"00000000",
  52299=>"00000000",
  52300=>"00000000",
  52301=>"11111110",
  52302=>"00000001",
  52303=>"00000010",
  52304=>"00000001",
  52305=>"00000011",
  52306=>"00000100",
  52307=>"11111101",
  52308=>"11111110",
  52309=>"00000001",
  52310=>"00000001",
  52311=>"11111101",
  52312=>"11111111",
  52313=>"11111100",
  52314=>"00000001",
  52315=>"00000001",
  52316=>"00000000",
  52317=>"00000001",
  52318=>"11111101",
  52319=>"11111110",
  52320=>"00000000",
  52321=>"11111111",
  52322=>"11111111",
  52323=>"11111101",
  52324=>"00000001",
  52325=>"11111110",
  52326=>"00000010",
  52327=>"00000001",
  52328=>"11111111",
  52329=>"11111110",
  52330=>"11111111",
  52331=>"00000100",
  52332=>"11111111",
  52333=>"11111110",
  52334=>"00000010",
  52335=>"11111111",
  52336=>"11111110",
  52337=>"00000001",
  52338=>"00000000",
  52339=>"11111111",
  52340=>"11111111",
  52341=>"11111100",
  52342=>"00000101",
  52343=>"00000000",
  52344=>"11111011",
  52345=>"11111111",
  52346=>"00000000",
  52347=>"00000000",
  52348=>"00000101",
  52349=>"00000001",
  52350=>"11111100",
  52351=>"00000010",
  52352=>"11111111",
  52353=>"00000000",
  52354=>"00000001",
  52355=>"00000001",
  52356=>"00000010",
  52357=>"00000000",
  52358=>"00000000",
  52359=>"11111101",
  52360=>"00000000",
  52361=>"00000011",
  52362=>"11111110",
  52363=>"11111111",
  52364=>"11111101",
  52365=>"11111101",
  52366=>"00000100",
  52367=>"11111101",
  52368=>"00000001",
  52369=>"11111101",
  52370=>"00000001",
  52371=>"11111111",
  52372=>"11111110",
  52373=>"11111100",
  52374=>"00000011",
  52375=>"11111110",
  52376=>"11111110",
  52377=>"00000010",
  52378=>"00000110",
  52379=>"11111111",
  52380=>"11111111",
  52381=>"00000010",
  52382=>"00000010",
  52383=>"11111110",
  52384=>"00000000",
  52385=>"00000000",
  52386=>"11111101",
  52387=>"11111111",
  52388=>"11111101",
  52389=>"00000001",
  52390=>"00000000",
  52391=>"00000010",
  52392=>"11111111",
  52393=>"00000011",
  52394=>"00000000",
  52395=>"11111111",
  52396=>"00000011",
  52397=>"11111110",
  52398=>"00000000",
  52399=>"00000011",
  52400=>"11111111",
  52401=>"11111101",
  52402=>"11111101",
  52403=>"00000001",
  52404=>"11111110",
  52405=>"11111110",
  52406=>"11111101",
  52407=>"00000001",
  52408=>"00000100",
  52409=>"00000011",
  52410=>"00000000",
  52411=>"00000001",
  52412=>"00000011",
  52413=>"00000010",
  52414=>"11111111",
  52415=>"11111111",
  52416=>"00000001",
  52417=>"11111110",
  52418=>"00000010",
  52419=>"00000000",
  52420=>"00000010",
  52421=>"00000000",
  52422=>"11111111",
  52423=>"11111110",
  52424=>"11111101",
  52425=>"00000011",
  52426=>"00000001",
  52427=>"11111111",
  52428=>"11111101",
  52429=>"11111111",
  52430=>"11111110",
  52431=>"00000000",
  52432=>"00000000",
  52433=>"11111111",
  52434=>"00000000",
  52435=>"00000100",
  52436=>"11111110",
  52437=>"00000000",
  52438=>"00000011",
  52439=>"00000010",
  52440=>"00000000",
  52441=>"00000000",
  52442=>"00000001",
  52443=>"11111111",
  52444=>"00000000",
  52445=>"00000100",
  52446=>"00000110",
  52447=>"11111101",
  52448=>"11111111",
  52449=>"00000011",
  52450=>"00000001",
  52451=>"11111101",
  52452=>"11111111",
  52453=>"11111101",
  52454=>"11111111",
  52455=>"00000010",
  52456=>"11111101",
  52457=>"11111101",
  52458=>"11111110",
  52459=>"11111110",
  52460=>"00000000",
  52461=>"11111110",
  52462=>"00000001",
  52463=>"11111110",
  52464=>"00000000",
  52465=>"00000100",
  52466=>"00000010",
  52467=>"00000000",
  52468=>"00000010",
  52469=>"11111111",
  52470=>"11111111",
  52471=>"11111111",
  52472=>"11111111",
  52473=>"11111101",
  52474=>"00000101",
  52475=>"00000001",
  52476=>"11111101",
  52477=>"00000001",
  52478=>"00000100",
  52479=>"11111101",
  52480=>"11111111",
  52481=>"00000001",
  52482=>"00000010",
  52483=>"00000010",
  52484=>"00000001",
  52485=>"00000001",
  52486=>"00000010",
  52487=>"00000000",
  52488=>"00000011",
  52489=>"00000001",
  52490=>"00000011",
  52491=>"00000000",
  52492=>"11111110",
  52493=>"00000001",
  52494=>"00000000",
  52495=>"00000010",
  52496=>"00000101",
  52497=>"11111111",
  52498=>"11111110",
  52499=>"00000100",
  52500=>"00000010",
  52501=>"00000000",
  52502=>"11111101",
  52503=>"11111110",
  52504=>"11111111",
  52505=>"00000000",
  52506=>"00000010",
  52507=>"00000000",
  52508=>"11111110",
  52509=>"00000010",
  52510=>"00000010",
  52511=>"00000100",
  52512=>"11111110",
  52513=>"11111110",
  52514=>"00000011",
  52515=>"00000011",
  52516=>"11111101",
  52517=>"00000000",
  52518=>"11111111",
  52519=>"11111101",
  52520=>"00000000",
  52521=>"11111111",
  52522=>"00000001",
  52523=>"00000001",
  52524=>"00000010",
  52525=>"11111110",
  52526=>"11111111",
  52527=>"00000110",
  52528=>"00000000",
  52529=>"00000000",
  52530=>"11111111",
  52531=>"11111111",
  52532=>"11111101",
  52533=>"11111111",
  52534=>"00000001",
  52535=>"00000000",
  52536=>"11111110",
  52537=>"00000010",
  52538=>"11111110",
  52539=>"00000011",
  52540=>"11111111",
  52541=>"11111101",
  52542=>"00000000",
  52543=>"00000000",
  52544=>"11111111",
  52545=>"00000100",
  52546=>"00000000",
  52547=>"00000000",
  52548=>"11111110",
  52549=>"00000010",
  52550=>"00000110",
  52551=>"00000000",
  52552=>"11111110",
  52553=>"11111101",
  52554=>"00000000",
  52555=>"00000010",
  52556=>"11111110",
  52557=>"00000010",
  52558=>"00000000",
  52559=>"00000000",
  52560=>"00000010",
  52561=>"11111110",
  52562=>"11111111",
  52563=>"00000000",
  52564=>"00000001",
  52565=>"11111101",
  52566=>"11111110",
  52567=>"00000100",
  52568=>"00000001",
  52569=>"00000001",
  52570=>"00000000",
  52571=>"11111110",
  52572=>"00000000",
  52573=>"11111110",
  52574=>"00000010",
  52575=>"00000111",
  52576=>"11111111",
  52577=>"11111110",
  52578=>"11111111",
  52579=>"00000001",
  52580=>"11111110",
  52581=>"11111101",
  52582=>"00000001",
  52583=>"11111111",
  52584=>"11111110",
  52585=>"11111101",
  52586=>"11111110",
  52587=>"00000010",
  52588=>"11111100",
  52589=>"00000010",
  52590=>"11111110",
  52591=>"00000000",
  52592=>"11111110",
  52593=>"00000001",
  52594=>"11111110",
  52595=>"00000001",
  52596=>"00000010",
  52597=>"11111110",
  52598=>"00000011",
  52599=>"00000001",
  52600=>"00000010",
  52601=>"11111111",
  52602=>"00000001",
  52603=>"11111111",
  52604=>"00000000",
  52605=>"00000010",
  52606=>"00000000",
  52607=>"11111101",
  52608=>"00000101",
  52609=>"00000100",
  52610=>"00000011",
  52611=>"11111110",
  52612=>"00000100",
  52613=>"11111101",
  52614=>"11111111",
  52615=>"11111110",
  52616=>"11111111",
  52617=>"00000010",
  52618=>"00000100",
  52619=>"11111110",
  52620=>"00000001",
  52621=>"11111101",
  52622=>"00000010",
  52623=>"00000000",
  52624=>"00000001",
  52625=>"11111110",
  52626=>"00000001",
  52627=>"00000001",
  52628=>"11111111",
  52629=>"11111110",
  52630=>"11111111",
  52631=>"11111111",
  52632=>"00000000",
  52633=>"11111111",
  52634=>"11111100",
  52635=>"11111110",
  52636=>"00000010",
  52637=>"00000001",
  52638=>"11111111",
  52639=>"00001000",
  52640=>"11111111",
  52641=>"11111111",
  52642=>"00000101",
  52643=>"11111110",
  52644=>"11111111",
  52645=>"11111110",
  52646=>"00000000",
  52647=>"00000010",
  52648=>"00000001",
  52649=>"11111111",
  52650=>"00000010",
  52651=>"11111110",
  52652=>"11111110",
  52653=>"00000010",
  52654=>"00000001",
  52655=>"11111101",
  52656=>"00000000",
  52657=>"11111110",
  52658=>"00000001",
  52659=>"11111111",
  52660=>"00000000",
  52661=>"11111101",
  52662=>"00000011",
  52663=>"11111111",
  52664=>"11111110",
  52665=>"00000011",
  52666=>"00000000",
  52667=>"00000010",
  52668=>"00000000",
  52669=>"00001001",
  52670=>"00000011",
  52671=>"00000100",
  52672=>"11111110",
  52673=>"00000000",
  52674=>"11111110",
  52675=>"00000011",
  52676=>"11111101",
  52677=>"00000001",
  52678=>"11111111",
  52679=>"11111110",
  52680=>"11111100",
  52681=>"11111111",
  52682=>"11111111",
  52683=>"11111111",
  52684=>"11111101",
  52685=>"11111111",
  52686=>"11111111",
  52687=>"00000001",
  52688=>"00000001",
  52689=>"11111110",
  52690=>"11111101",
  52691=>"00000001",
  52692=>"11111110",
  52693=>"11111110",
  52694=>"00000001",
  52695=>"11111110",
  52696=>"11111101",
  52697=>"11111101",
  52698=>"11111111",
  52699=>"00000000",
  52700=>"11111101",
  52701=>"11111101",
  52702=>"11111111",
  52703=>"11111110",
  52704=>"00000001",
  52705=>"00000001",
  52706=>"00000001",
  52707=>"00000010",
  52708=>"00000000",
  52709=>"11111101",
  52710=>"00000010",
  52711=>"00000010",
  52712=>"11111101",
  52713=>"11111111",
  52714=>"11111101",
  52715=>"11111110",
  52716=>"00000100",
  52717=>"11111110",
  52718=>"11111101",
  52719=>"00000010",
  52720=>"00000000",
  52721=>"11111110",
  52722=>"00000011",
  52723=>"00000011",
  52724=>"00000001",
  52725=>"00000000",
  52726=>"11111101",
  52727=>"11111111",
  52728=>"00000001",
  52729=>"00000011",
  52730=>"11111101",
  52731=>"00000001",
  52732=>"11111111",
  52733=>"00000010",
  52734=>"00000001",
  52735=>"00000010",
  52736=>"11111111",
  52737=>"00000001",
  52738=>"11111110",
  52739=>"00000010",
  52740=>"00000001",
  52741=>"11111111",
  52742=>"00000001",
  52743=>"11111110",
  52744=>"00000011",
  52745=>"00000010",
  52746=>"11111111",
  52747=>"00000001",
  52748=>"11111110",
  52749=>"11111111",
  52750=>"11111101",
  52751=>"00000011",
  52752=>"00000001",
  52753=>"11111111",
  52754=>"00000001",
  52755=>"11111101",
  52756=>"11111111",
  52757=>"00000010",
  52758=>"00000001",
  52759=>"11111110",
  52760=>"11111111",
  52761=>"00000111",
  52762=>"00000010",
  52763=>"11111110",
  52764=>"11111111",
  52765=>"00000001",
  52766=>"00000001",
  52767=>"00000001",
  52768=>"11111111",
  52769=>"11111110",
  52770=>"00000001",
  52771=>"11111101",
  52772=>"00000001",
  52773=>"11111111",
  52774=>"11111110",
  52775=>"00000000",
  52776=>"11111110",
  52777=>"11111111",
  52778=>"11111101",
  52779=>"11111111",
  52780=>"00000010",
  52781=>"11111110",
  52782=>"11111111",
  52783=>"00000000",
  52784=>"11111110",
  52785=>"11111101",
  52786=>"00000010",
  52787=>"00000001",
  52788=>"00000010",
  52789=>"00000001",
  52790=>"11111110",
  52791=>"11111111",
  52792=>"00000000",
  52793=>"00000010",
  52794=>"11111111",
  52795=>"00000001",
  52796=>"00000100",
  52797=>"11111101",
  52798=>"00000000",
  52799=>"11111111",
  52800=>"00000000",
  52801=>"00000000",
  52802=>"00000001",
  52803=>"00000000",
  52804=>"00000000",
  52805=>"00000010",
  52806=>"00000000",
  52807=>"00000001",
  52808=>"00000000",
  52809=>"00000000",
  52810=>"11111110",
  52811=>"11111111",
  52812=>"00000010",
  52813=>"00000000",
  52814=>"11111101",
  52815=>"11111101",
  52816=>"00000001",
  52817=>"11111101",
  52818=>"00000011",
  52819=>"00000000",
  52820=>"00000001",
  52821=>"00000010",
  52822=>"00000100",
  52823=>"11111110",
  52824=>"00000010",
  52825=>"11111111",
  52826=>"11111110",
  52827=>"00000011",
  52828=>"00000110",
  52829=>"00000001",
  52830=>"11111101",
  52831=>"11111110",
  52832=>"00000001",
  52833=>"00000010",
  52834=>"11111111",
  52835=>"11111111",
  52836=>"00000001",
  52837=>"00000101",
  52838=>"00000000",
  52839=>"11111100",
  52840=>"00000011",
  52841=>"00000001",
  52842=>"00000000",
  52843=>"00000000",
  52844=>"11111101",
  52845=>"00000000",
  52846=>"11111111",
  52847=>"00000010",
  52848=>"00000001",
  52849=>"00000000",
  52850=>"11111111",
  52851=>"11111111",
  52852=>"11111111",
  52853=>"11111111",
  52854=>"00000010",
  52855=>"11111101",
  52856=>"11111101",
  52857=>"11111101",
  52858=>"11111110",
  52859=>"00000000",
  52860=>"00000001",
  52861=>"11111101",
  52862=>"11111101",
  52863=>"00000001",
  52864=>"00000010",
  52865=>"00000000",
  52866=>"11111110",
  52867=>"11111110",
  52868=>"00000000",
  52869=>"11111111",
  52870=>"11111111",
  52871=>"11111110",
  52872=>"11111110",
  52873=>"00000011",
  52874=>"00000000",
  52875=>"11111111",
  52876=>"00000000",
  52877=>"11111110",
  52878=>"11111110",
  52879=>"11111111",
  52880=>"00000000",
  52881=>"00000010",
  52882=>"11111111",
  52883=>"00000010",
  52884=>"11111101",
  52885=>"11111110",
  52886=>"00000000",
  52887=>"11111101",
  52888=>"00000000",
  52889=>"11111110",
  52890=>"00000011",
  52891=>"11111110",
  52892=>"11111110",
  52893=>"11111110",
  52894=>"00000001",
  52895=>"11111101",
  52896=>"00000001",
  52897=>"11111111",
  52898=>"11111111",
  52899=>"11111110",
  52900=>"00000000",
  52901=>"00000000",
  52902=>"11111111",
  52903=>"00000000",
  52904=>"11111111",
  52905=>"11111101",
  52906=>"11111111",
  52907=>"00000001",
  52908=>"11111110",
  52909=>"00000000",
  52910=>"00000010",
  52911=>"00000001",
  52912=>"11111101",
  52913=>"00000001",
  52914=>"00000010",
  52915=>"11111110",
  52916=>"00000000",
  52917=>"11111101",
  52918=>"11111111",
  52919=>"11111111",
  52920=>"11111111",
  52921=>"11111111",
  52922=>"11111110",
  52923=>"00000001",
  52924=>"11111111",
  52925=>"11111101",
  52926=>"00000001",
  52927=>"11111110",
  52928=>"11111110",
  52929=>"11111110",
  52930=>"00000010",
  52931=>"00000001",
  52932=>"00000001",
  52933=>"00000011",
  52934=>"00000011",
  52935=>"11111101",
  52936=>"11111100",
  52937=>"00000010",
  52938=>"00000010",
  52939=>"11111110",
  52940=>"11111111",
  52941=>"00000011",
  52942=>"11111110",
  52943=>"00000000",
  52944=>"11111110",
  52945=>"00000001",
  52946=>"00000001",
  52947=>"00000001",
  52948=>"00000001",
  52949=>"11111110",
  52950=>"00000010",
  52951=>"11111110",
  52952=>"00000000",
  52953=>"11111110",
  52954=>"00000001",
  52955=>"11111101",
  52956=>"11111110",
  52957=>"00000000",
  52958=>"11111110",
  52959=>"00000000",
  52960=>"00000010",
  52961=>"00000001",
  52962=>"00000001",
  52963=>"00000000",
  52964=>"00000001",
  52965=>"11111110",
  52966=>"00000000",
  52967=>"00000000",
  52968=>"11111101",
  52969=>"00000000",
  52970=>"11111100",
  52971=>"00000000",
  52972=>"11111110",
  52973=>"11111101",
  52974=>"11111111",
  52975=>"00000000",
  52976=>"00000010",
  52977=>"00000001",
  52978=>"11111110",
  52979=>"00000001",
  52980=>"00000001",
  52981=>"00000100",
  52982=>"00000001",
  52983=>"00000000",
  52984=>"11111101",
  52985=>"00000000",
  52986=>"11111110",
  52987=>"11111111",
  52988=>"11111111",
  52989=>"00000001",
  52990=>"11111110",
  52991=>"00000010",
  52992=>"11111110",
  52993=>"11111111",
  52994=>"11111111",
  52995=>"00000101",
  52996=>"00000000",
  52997=>"11111101",
  52998=>"00000000",
  52999=>"00000001",
  53000=>"00000000",
  53001=>"00000001",
  53002=>"11111111",
  53003=>"00000011",
  53004=>"00000010",
  53005=>"00000000",
  53006=>"11111110",
  53007=>"00000010",
  53008=>"00000001",
  53009=>"11111110",
  53010=>"11111110",
  53011=>"00000000",
  53012=>"11111110",
  53013=>"11111101",
  53014=>"11111111",
  53015=>"11111110",
  53016=>"00000010",
  53017=>"00000011",
  53018=>"00000000",
  53019=>"00000001",
  53020=>"11111101",
  53021=>"00000101",
  53022=>"00000001",
  53023=>"11111110",
  53024=>"11111110",
  53025=>"11111111",
  53026=>"11111111",
  53027=>"00000001",
  53028=>"11111111",
  53029=>"00000010",
  53030=>"00000000",
  53031=>"11111101",
  53032=>"00000001",
  53033=>"00000000",
  53034=>"11111101",
  53035=>"11111111",
  53036=>"11111111",
  53037=>"11111110",
  53038=>"11111101",
  53039=>"11111110",
  53040=>"00000001",
  53041=>"11111111",
  53042=>"00000100",
  53043=>"11111111",
  53044=>"00000000",
  53045=>"11111101",
  53046=>"00000010",
  53047=>"11111101",
  53048=>"00000100",
  53049=>"00000001",
  53050=>"11111101",
  53051=>"00000010",
  53052=>"00000000",
  53053=>"00000100",
  53054=>"11111110",
  53055=>"00000011",
  53056=>"11111110",
  53057=>"11111111",
  53058=>"00000001",
  53059=>"00000010",
  53060=>"11111111",
  53061=>"11111111",
  53062=>"00000010",
  53063=>"11111101",
  53064=>"11111101",
  53065=>"11111101",
  53066=>"00000001",
  53067=>"00000011",
  53068=>"11111111",
  53069=>"00000001",
  53070=>"00000001",
  53071=>"00000001",
  53072=>"00000000",
  53073=>"00000000",
  53074=>"11111110",
  53075=>"11111111",
  53076=>"00000000",
  53077=>"11111110",
  53078=>"00000010",
  53079=>"11111101",
  53080=>"11111100",
  53081=>"00000010",
  53082=>"11111100",
  53083=>"00000100",
  53084=>"00000010",
  53085=>"11111111",
  53086=>"00000000",
  53087=>"11111101",
  53088=>"00000010",
  53089=>"00000001",
  53090=>"00000010",
  53091=>"11111111",
  53092=>"00000001",
  53093=>"00000001",
  53094=>"00000001",
  53095=>"00000001",
  53096=>"00000011",
  53097=>"11111110",
  53098=>"11111111",
  53099=>"11111111",
  53100=>"11111110",
  53101=>"00000000",
  53102=>"00000100",
  53103=>"11111110",
  53104=>"00000001",
  53105=>"11111100",
  53106=>"00000010",
  53107=>"11111100",
  53108=>"11111111",
  53109=>"00000001",
  53110=>"11111110",
  53111=>"11111111",
  53112=>"00000000",
  53113=>"11111111",
  53114=>"11111101",
  53115=>"00000000",
  53116=>"00000100",
  53117=>"00000001",
  53118=>"00000010",
  53119=>"11111111",
  53120=>"11111110",
  53121=>"11111111",
  53122=>"11111101",
  53123=>"00000001",
  53124=>"11111111",
  53125=>"00000010",
  53126=>"00000011",
  53127=>"11111111",
  53128=>"11111101",
  53129=>"11111110",
  53130=>"11111111",
  53131=>"11111111",
  53132=>"11111110",
  53133=>"11111101",
  53134=>"00000100",
  53135=>"00000010",
  53136=>"11111110",
  53137=>"00000000",
  53138=>"00000110",
  53139=>"00000000",
  53140=>"11111111",
  53141=>"11111110",
  53142=>"00000010",
  53143=>"00000011",
  53144=>"11111111",
  53145=>"11111101",
  53146=>"11111111",
  53147=>"11111111",
  53148=>"00000000",
  53149=>"00000011",
  53150=>"00000011",
  53151=>"00000010",
  53152=>"11111110",
  53153=>"00000010",
  53154=>"00000001",
  53155=>"00000000",
  53156=>"00000010",
  53157=>"11111111",
  53158=>"00000000",
  53159=>"00000010",
  53160=>"00000001",
  53161=>"11111110",
  53162=>"11111110",
  53163=>"00000010",
  53164=>"11111111",
  53165=>"00000110",
  53166=>"00000010",
  53167=>"00000000",
  53168=>"11111111",
  53169=>"00000001",
  53170=>"00000001",
  53171=>"00000010",
  53172=>"11111100",
  53173=>"11111111",
  53174=>"00000010",
  53175=>"11111111",
  53176=>"11111110",
  53177=>"11111110",
  53178=>"00000010",
  53179=>"00000010",
  53180=>"11111110",
  53181=>"00000000",
  53182=>"00000001",
  53183=>"00000001",
  53184=>"00000001",
  53185=>"00000000",
  53186=>"11111110",
  53187=>"00000000",
  53188=>"11111110",
  53189=>"11111110",
  53190=>"11111111",
  53191=>"00000001",
  53192=>"11111110",
  53193=>"00000000",
  53194=>"00000000",
  53195=>"00000000",
  53196=>"00000001",
  53197=>"11111111",
  53198=>"11111111",
  53199=>"11111110",
  53200=>"11111111",
  53201=>"00000000",
  53202=>"11111101",
  53203=>"00000000",
  53204=>"00000001",
  53205=>"11111100",
  53206=>"11111101",
  53207=>"00000010",
  53208=>"11111110",
  53209=>"00000001",
  53210=>"00000001",
  53211=>"11111111",
  53212=>"00000000",
  53213=>"11111111",
  53214=>"00000001",
  53215=>"11111111",
  53216=>"11111101",
  53217=>"11111101",
  53218=>"00000001",
  53219=>"00000000",
  53220=>"11111110",
  53221=>"11111100",
  53222=>"00000101",
  53223=>"00000001",
  53224=>"00000001",
  53225=>"00000000",
  53226=>"11111111",
  53227=>"11111101",
  53228=>"11111110",
  53229=>"00000011",
  53230=>"00000000",
  53231=>"00000100",
  53232=>"11111111",
  53233=>"00000011",
  53234=>"11111101",
  53235=>"11111101",
  53236=>"00000001",
  53237=>"11111111",
  53238=>"00000010",
  53239=>"00000001",
  53240=>"11111110",
  53241=>"00000000",
  53242=>"11111111",
  53243=>"00000000",
  53244=>"11111101",
  53245=>"11111111",
  53246=>"00000001",
  53247=>"11111111",
  53248=>"11111111",
  53249=>"00000000",
  53250=>"00000001",
  53251=>"00000001",
  53252=>"00000000",
  53253=>"11111111",
  53254=>"11111111",
  53255=>"11111111",
  53256=>"11111101",
  53257=>"00000010",
  53258=>"00000000",
  53259=>"11111111",
  53260=>"00000001",
  53261=>"11111101",
  53262=>"00000110",
  53263=>"00000010",
  53264=>"00000010",
  53265=>"11111101",
  53266=>"00000010",
  53267=>"11111111",
  53268=>"00000000",
  53269=>"00000001",
  53270=>"11111111",
  53271=>"11111111",
  53272=>"11111111",
  53273=>"00000001",
  53274=>"00000000",
  53275=>"00000001",
  53276=>"11111101",
  53277=>"11111111",
  53278=>"00000100",
  53279=>"00000000",
  53280=>"00000000",
  53281=>"00000000",
  53282=>"11111111",
  53283=>"11111111",
  53284=>"11111110",
  53285=>"11111111",
  53286=>"11111110",
  53287=>"11111110",
  53288=>"11111101",
  53289=>"00000010",
  53290=>"11111111",
  53291=>"00000100",
  53292=>"00000101",
  53293=>"00000001",
  53294=>"00000001",
  53295=>"00000001",
  53296=>"00000011",
  53297=>"00000000",
  53298=>"11111100",
  53299=>"11111110",
  53300=>"00000000",
  53301=>"11111111",
  53302=>"00000001",
  53303=>"00000010",
  53304=>"00000000",
  53305=>"00000011",
  53306=>"00000000",
  53307=>"00000010",
  53308=>"00000100",
  53309=>"00000001",
  53310=>"00000001",
  53311=>"00000001",
  53312=>"11111110",
  53313=>"00000010",
  53314=>"00000000",
  53315=>"11111110",
  53316=>"00000000",
  53317=>"00000011",
  53318=>"11111110",
  53319=>"00000001",
  53320=>"00000001",
  53321=>"00000010",
  53322=>"00000000",
  53323=>"00000000",
  53324=>"00000000",
  53325=>"00000011",
  53326=>"11111111",
  53327=>"11111110",
  53328=>"00000000",
  53329=>"11111110",
  53330=>"11111110",
  53331=>"00000110",
  53332=>"00000010",
  53333=>"11111110",
  53334=>"00000100",
  53335=>"11111110",
  53336=>"00000011",
  53337=>"00000001",
  53338=>"11111111",
  53339=>"00000010",
  53340=>"00000011",
  53341=>"11111111",
  53342=>"00000010",
  53343=>"00000111",
  53344=>"11111110",
  53345=>"11111110",
  53346=>"11111011",
  53347=>"00000000",
  53348=>"11111111",
  53349=>"11111110",
  53350=>"11111111",
  53351=>"00000010",
  53352=>"00000010",
  53353=>"00000000",
  53354=>"00000000",
  53355=>"00000010",
  53356=>"00000000",
  53357=>"00000001",
  53358=>"11111101",
  53359=>"11111101",
  53360=>"11111110",
  53361=>"00000001",
  53362=>"00000101",
  53363=>"00000011",
  53364=>"00000001",
  53365=>"00000001",
  53366=>"00000011",
  53367=>"00000000",
  53368=>"11111101",
  53369=>"00000000",
  53370=>"00000000",
  53371=>"11111100",
  53372=>"00000010",
  53373=>"11111101",
  53374=>"00000010",
  53375=>"11111100",
  53376=>"11111101",
  53377=>"00000011",
  53378=>"00000000",
  53379=>"00000001",
  53380=>"11111111",
  53381=>"00000101",
  53382=>"00000000",
  53383=>"00000100",
  53384=>"00000000",
  53385=>"00000011",
  53386=>"11111111",
  53387=>"00000100",
  53388=>"00000001",
  53389=>"00000011",
  53390=>"11111110",
  53391=>"00000001",
  53392=>"11111111",
  53393=>"00000011",
  53394=>"00000000",
  53395=>"00000101",
  53396=>"00000010",
  53397=>"00000000",
  53398=>"00000010",
  53399=>"00000100",
  53400=>"11111110",
  53401=>"00000001",
  53402=>"00000011",
  53403=>"00000001",
  53404=>"00000010",
  53405=>"00000100",
  53406=>"00000011",
  53407=>"11111111",
  53408=>"00000011",
  53409=>"00000010",
  53410=>"00000010",
  53411=>"11111110",
  53412=>"00000000",
  53413=>"00000101",
  53414=>"11111101",
  53415=>"11111100",
  53416=>"00000101",
  53417=>"00000001",
  53418=>"11111110",
  53419=>"11111111",
  53420=>"00000001",
  53421=>"11111101",
  53422=>"11111101",
  53423=>"00000010",
  53424=>"11111111",
  53425=>"00000010",
  53426=>"00000100",
  53427=>"00000011",
  53428=>"11111101",
  53429=>"11111110",
  53430=>"00000010",
  53431=>"00000001",
  53432=>"11111110",
  53433=>"00000001",
  53434=>"00000000",
  53435=>"11111110",
  53436=>"00000010",
  53437=>"11111111",
  53438=>"00000000",
  53439=>"11111110",
  53440=>"00000010",
  53441=>"11111110",
  53442=>"00000100",
  53443=>"11111111",
  53444=>"11111110",
  53445=>"00000010",
  53446=>"00000000",
  53447=>"00000100",
  53448=>"00000011",
  53449=>"00000000",
  53450=>"00000000",
  53451=>"11111110",
  53452=>"00000100",
  53453=>"00000010",
  53454=>"11111111",
  53455=>"00000101",
  53456=>"11111111",
  53457=>"11111110",
  53458=>"00000010",
  53459=>"00000010",
  53460=>"00000001",
  53461=>"00000011",
  53462=>"00000001",
  53463=>"00000001",
  53464=>"00000000",
  53465=>"00000000",
  53466=>"11111110",
  53467=>"11111101",
  53468=>"00000010",
  53469=>"00000010",
  53470=>"00000000",
  53471=>"00000100",
  53472=>"00000001",
  53473=>"00000000",
  53474=>"11111111",
  53475=>"11111110",
  53476=>"00000000",
  53477=>"00000100",
  53478=>"11111100",
  53479=>"11111110",
  53480=>"00000001",
  53481=>"11111111",
  53482=>"00000000",
  53483=>"00000000",
  53484=>"11111111",
  53485=>"00000011",
  53486=>"11111111",
  53487=>"00000001",
  53488=>"00000111",
  53489=>"11111110",
  53490=>"00000001",
  53491=>"00000000",
  53492=>"00000001",
  53493=>"00000101",
  53494=>"00000001",
  53495=>"11111101",
  53496=>"00000000",
  53497=>"00000010",
  53498=>"11111111",
  53499=>"00000000",
  53500=>"11111110",
  53501=>"00000010",
  53502=>"11111101",
  53503=>"00000001",
  53504=>"00000000",
  53505=>"00000000",
  53506=>"11111111",
  53507=>"00000011",
  53508=>"11111111",
  53509=>"00000001",
  53510=>"11111110",
  53511=>"11111101",
  53512=>"11111101",
  53513=>"11111110",
  53514=>"11111111",
  53515=>"00000010",
  53516=>"11111111",
  53517=>"00000011",
  53518=>"11111110",
  53519=>"00000000",
  53520=>"11111110",
  53521=>"00000010",
  53522=>"00000010",
  53523=>"11111101",
  53524=>"00000100",
  53525=>"00000000",
  53526=>"11111111",
  53527=>"00000001",
  53528=>"11111110",
  53529=>"00000001",
  53530=>"00000001",
  53531=>"00000000",
  53532=>"00000010",
  53533=>"11111101",
  53534=>"11111101",
  53535=>"11111110",
  53536=>"00000001",
  53537=>"00000010",
  53538=>"00000100",
  53539=>"00000010",
  53540=>"00000010",
  53541=>"11111101",
  53542=>"00000001",
  53543=>"00000001",
  53544=>"00000000",
  53545=>"00000001",
  53546=>"00000010",
  53547=>"00000010",
  53548=>"11111111",
  53549=>"11111101",
  53550=>"11111110",
  53551=>"00000001",
  53552=>"00000010",
  53553=>"11111101",
  53554=>"00000010",
  53555=>"00000001",
  53556=>"00000000",
  53557=>"00000011",
  53558=>"00000011",
  53559=>"11111111",
  53560=>"00000000",
  53561=>"00000010",
  53562=>"11111111",
  53563=>"11111101",
  53564=>"00000100",
  53565=>"11111111",
  53566=>"11111110",
  53567=>"00000000",
  53568=>"00000010",
  53569=>"11111110",
  53570=>"11111111",
  53571=>"00000000",
  53572=>"11111111",
  53573=>"11111111",
  53574=>"00000010",
  53575=>"00000010",
  53576=>"00000000",
  53577=>"00000001",
  53578=>"00000100",
  53579=>"11111101",
  53580=>"00000011",
  53581=>"11111101",
  53582=>"00000000",
  53583=>"00000000",
  53584=>"11111101",
  53585=>"11111101",
  53586=>"11111110",
  53587=>"11111111",
  53588=>"11111111",
  53589=>"11111101",
  53590=>"00000010",
  53591=>"00000001",
  53592=>"00000010",
  53593=>"11111110",
  53594=>"11111101",
  53595=>"00000001",
  53596=>"11111111",
  53597=>"11111110",
  53598=>"11111101",
  53599=>"11111110",
  53600=>"00000001",
  53601=>"11111111",
  53602=>"00000001",
  53603=>"00000101",
  53604=>"00000001",
  53605=>"00000001",
  53606=>"00000100",
  53607=>"11111110",
  53608=>"11111101",
  53609=>"00000010",
  53610=>"11111111",
  53611=>"00000010",
  53612=>"00000001",
  53613=>"00000011",
  53614=>"00000000",
  53615=>"00000001",
  53616=>"11111110",
  53617=>"00000011",
  53618=>"11111111",
  53619=>"11111111",
  53620=>"00000011",
  53621=>"00000001",
  53622=>"11111111",
  53623=>"00000000",
  53624=>"00000000",
  53625=>"00000000",
  53626=>"11111111",
  53627=>"00000011",
  53628=>"00000000",
  53629=>"11111110",
  53630=>"11111101",
  53631=>"11111110",
  53632=>"00000000",
  53633=>"11111111",
  53634=>"11111110",
  53635=>"11111111",
  53636=>"11111101",
  53637=>"11111101",
  53638=>"00000001",
  53639=>"11111101",
  53640=>"00000010",
  53641=>"00000011",
  53642=>"11111101",
  53643=>"00000000",
  53644=>"00000001",
  53645=>"00000001",
  53646=>"11111110",
  53647=>"00000011",
  53648=>"11111111",
  53649=>"00000000",
  53650=>"11111111",
  53651=>"11111100",
  53652=>"00000001",
  53653=>"00000010",
  53654=>"00000001",
  53655=>"11111101",
  53656=>"00000100",
  53657=>"11111100",
  53658=>"00000011",
  53659=>"00000001",
  53660=>"00000000",
  53661=>"00000011",
  53662=>"00000010",
  53663=>"11111100",
  53664=>"00000000",
  53665=>"11111110",
  53666=>"11111111",
  53667=>"00000011",
  53668=>"11111111",
  53669=>"00000000",
  53670=>"00000011",
  53671=>"11111100",
  53672=>"11111111",
  53673=>"11111101",
  53674=>"11111111",
  53675=>"00000101",
  53676=>"00000000",
  53677=>"00000001",
  53678=>"00000001",
  53679=>"00000010",
  53680=>"11111110",
  53681=>"11111101",
  53682=>"00000011",
  53683=>"00000010",
  53684=>"00000011",
  53685=>"00000000",
  53686=>"00000101",
  53687=>"00000001",
  53688=>"00000000",
  53689=>"00000001",
  53690=>"11111110",
  53691=>"11111110",
  53692=>"00000001",
  53693=>"11111101",
  53694=>"11111101",
  53695=>"11111110",
  53696=>"11111111",
  53697=>"00000000",
  53698=>"11111101",
  53699=>"11111111",
  53700=>"00000111",
  53701=>"11111101",
  53702=>"00000010",
  53703=>"00000000",
  53704=>"11111101",
  53705=>"00000011",
  53706=>"11111100",
  53707=>"00000001",
  53708=>"00000001",
  53709=>"00000010",
  53710=>"00000000",
  53711=>"00000010",
  53712=>"00000010",
  53713=>"11111111",
  53714=>"00000001",
  53715=>"00000101",
  53716=>"00000010",
  53717=>"00000001",
  53718=>"11111111",
  53719=>"00000000",
  53720=>"11111111",
  53721=>"00000000",
  53722=>"00000000",
  53723=>"11111101",
  53724=>"00000010",
  53725=>"00000010",
  53726=>"11111111",
  53727=>"11111110",
  53728=>"00000111",
  53729=>"00000011",
  53730=>"00000000",
  53731=>"00000011",
  53732=>"00000001",
  53733=>"11111111",
  53734=>"11111101",
  53735=>"00000001",
  53736=>"11111100",
  53737=>"11111101",
  53738=>"00000000",
  53739=>"00000001",
  53740=>"11111100",
  53741=>"11111011",
  53742=>"00000001",
  53743=>"00000011",
  53744=>"00000000",
  53745=>"11111111",
  53746=>"00000001",
  53747=>"11111110",
  53748=>"00000011",
  53749=>"11111110",
  53750=>"00000011",
  53751=>"00000000",
  53752=>"00000010",
  53753=>"11111111",
  53754=>"00000000",
  53755=>"00000001",
  53756=>"11111101",
  53757=>"11111100",
  53758=>"11111110",
  53759=>"11111101",
  53760=>"00000001",
  53761=>"00000100",
  53762=>"00000010",
  53763=>"11111110",
  53764=>"00000011",
  53765=>"11111110",
  53766=>"11111100",
  53767=>"00000100",
  53768=>"11111110",
  53769=>"00000000",
  53770=>"00000001",
  53771=>"11111111",
  53772=>"00000000",
  53773=>"11111110",
  53774=>"11111101",
  53775=>"00000001",
  53776=>"00000000",
  53777=>"00000001",
  53778=>"00000000",
  53779=>"11111111",
  53780=>"00000011",
  53781=>"11111111",
  53782=>"00000011",
  53783=>"00000010",
  53784=>"00000001",
  53785=>"00000000",
  53786=>"11111101",
  53787=>"00000010",
  53788=>"00000000",
  53789=>"00000000",
  53790=>"11111101",
  53791=>"11111101",
  53792=>"11111111",
  53793=>"00000011",
  53794=>"00000000",
  53795=>"11111110",
  53796=>"11111101",
  53797=>"11111111",
  53798=>"11111111",
  53799=>"11111111",
  53800=>"11111110",
  53801=>"00000010",
  53802=>"00000001",
  53803=>"00000010",
  53804=>"00000000",
  53805=>"00000001",
  53806=>"00000001",
  53807=>"00000001",
  53808=>"00000000",
  53809=>"00000010",
  53810=>"11111110",
  53811=>"11111111",
  53812=>"11111110",
  53813=>"11111111",
  53814=>"00000010",
  53815=>"00000010",
  53816=>"00000000",
  53817=>"00000010",
  53818=>"00000011",
  53819=>"11111101",
  53820=>"00000000",
  53821=>"00000011",
  53822=>"00000000",
  53823=>"00000010",
  53824=>"00000010",
  53825=>"00000011",
  53826=>"11111110",
  53827=>"00000010",
  53828=>"11111111",
  53829=>"11111111",
  53830=>"11111100",
  53831=>"11111111",
  53832=>"11111111",
  53833=>"11111111",
  53834=>"00000100",
  53835=>"00000001",
  53836=>"00000100",
  53837=>"00000000",
  53838=>"11111111",
  53839=>"11111111",
  53840=>"00000001",
  53841=>"00000011",
  53842=>"00000000",
  53843=>"00000010",
  53844=>"00000011",
  53845=>"00000000",
  53846=>"00000001",
  53847=>"00000000",
  53848=>"00000001",
  53849=>"00000000",
  53850=>"00000001",
  53851=>"00000001",
  53852=>"11111110",
  53853=>"00000011",
  53854=>"00000000",
  53855=>"11111101",
  53856=>"00000001",
  53857=>"00000001",
  53858=>"11111100",
  53859=>"00000010",
  53860=>"11111110",
  53861=>"11111110",
  53862=>"11111110",
  53863=>"00000000",
  53864=>"00000010",
  53865=>"11111101",
  53866=>"11111111",
  53867=>"00000000",
  53868=>"00000010",
  53869=>"00000001",
  53870=>"00000101",
  53871=>"11111110",
  53872=>"00000000",
  53873=>"11111111",
  53874=>"00000011",
  53875=>"11111111",
  53876=>"11111110",
  53877=>"00000000",
  53878=>"00000001",
  53879=>"00000001",
  53880=>"11111110",
  53881=>"11111110",
  53882=>"11111110",
  53883=>"11111111",
  53884=>"00000100",
  53885=>"00000010",
  53886=>"00000011",
  53887=>"00000000",
  53888=>"11111111",
  53889=>"00000011",
  53890=>"00000001",
  53891=>"11111111",
  53892=>"11111101",
  53893=>"00000000",
  53894=>"11111101",
  53895=>"00000010",
  53896=>"00000011",
  53897=>"11111110",
  53898=>"00000000",
  53899=>"11111111",
  53900=>"11111110",
  53901=>"11111111",
  53902=>"11111111",
  53903=>"00000000",
  53904=>"00000100",
  53905=>"11111111",
  53906=>"00000010",
  53907=>"11111101",
  53908=>"00000011",
  53909=>"00000000",
  53910=>"11111111",
  53911=>"11111100",
  53912=>"11111110",
  53913=>"00000000",
  53914=>"11111111",
  53915=>"00000000",
  53916=>"11111110",
  53917=>"11111111",
  53918=>"11111100",
  53919=>"00000001",
  53920=>"11111110",
  53921=>"11111111",
  53922=>"11111110",
  53923=>"11111111",
  53924=>"00000010",
  53925=>"11111111",
  53926=>"11111111",
  53927=>"00000000",
  53928=>"00000011",
  53929=>"00000001",
  53930=>"00000010",
  53931=>"00000011",
  53932=>"11111110",
  53933=>"11111111",
  53934=>"00000000",
  53935=>"11111101",
  53936=>"11111111",
  53937=>"11111110",
  53938=>"11111101",
  53939=>"00000001",
  53940=>"11111111",
  53941=>"00000000",
  53942=>"00000000",
  53943=>"00000011",
  53944=>"11111110",
  53945=>"11111101",
  53946=>"00000000",
  53947=>"00000000",
  53948=>"00000010",
  53949=>"11111111",
  53950=>"00000010",
  53951=>"00000001",
  53952=>"00000001",
  53953=>"11111111",
  53954=>"00000011",
  53955=>"00000000",
  53956=>"00000010",
  53957=>"11111111",
  53958=>"11111110",
  53959=>"00000100",
  53960=>"00000011",
  53961=>"11111110",
  53962=>"00000010",
  53963=>"00001010",
  53964=>"11111110",
  53965=>"11111101",
  53966=>"11111101",
  53967=>"00000100",
  53968=>"11111111",
  53969=>"11111100",
  53970=>"00000001",
  53971=>"00000011",
  53972=>"00000000",
  53973=>"00000000",
  53974=>"00000010",
  53975=>"00000000",
  53976=>"11111101",
  53977=>"11111101",
  53978=>"11111110",
  53979=>"11111111",
  53980=>"00000010",
  53981=>"00000000",
  53982=>"11111100",
  53983=>"11111110",
  53984=>"00000010",
  53985=>"00000010",
  53986=>"11111100",
  53987=>"00000001",
  53988=>"11111111",
  53989=>"00000000",
  53990=>"00000011",
  53991=>"11111100",
  53992=>"00000000",
  53993=>"11111111",
  53994=>"11111101",
  53995=>"00000011",
  53996=>"11111111",
  53997=>"11111110",
  53998=>"00000001",
  53999=>"00000010",
  54000=>"11111110",
  54001=>"11111111",
  54002=>"00000010",
  54003=>"00000001",
  54004=>"11111110",
  54005=>"11111111",
  54006=>"11111110",
  54007=>"00000000",
  54008=>"00000010",
  54009=>"11111110",
  54010=>"00000011",
  54011=>"11111110",
  54012=>"00000010",
  54013=>"00000001",
  54014=>"00000010",
  54015=>"00000100",
  54016=>"00000010",
  54017=>"00000100",
  54018=>"00000000",
  54019=>"11111101",
  54020=>"11111111",
  54021=>"11111100",
  54022=>"11111101",
  54023=>"00000011",
  54024=>"11111111",
  54025=>"11111110",
  54026=>"00000001",
  54027=>"00000000",
  54028=>"11111110",
  54029=>"11111111",
  54030=>"00000000",
  54031=>"11111111",
  54032=>"00000010",
  54033=>"11111110",
  54034=>"11111101",
  54035=>"11111101",
  54036=>"00000010",
  54037=>"11111111",
  54038=>"00000000",
  54039=>"00000000",
  54040=>"11111111",
  54041=>"00000001",
  54042=>"11111100",
  54043=>"00000010",
  54044=>"00000001",
  54045=>"00000011",
  54046=>"11111110",
  54047=>"11111110",
  54048=>"00000001",
  54049=>"11111111",
  54050=>"11111110",
  54051=>"00000100",
  54052=>"00000000",
  54053=>"11111111",
  54054=>"00000010",
  54055=>"00000101",
  54056=>"00000001",
  54057=>"11111110",
  54058=>"11111111",
  54059=>"00000011",
  54060=>"00000010",
  54061=>"00000010",
  54062=>"11111111",
  54063=>"00000001",
  54064=>"11111101",
  54065=>"00000000",
  54066=>"00000010",
  54067=>"00000100",
  54068=>"00000001",
  54069=>"00000000",
  54070=>"00000010",
  54071=>"11111111",
  54072=>"00000010",
  54073=>"00000000",
  54074=>"00000010",
  54075=>"11111110",
  54076=>"11111111",
  54077=>"00000000",
  54078=>"11111110",
  54079=>"00000001",
  54080=>"11111110",
  54081=>"00000011",
  54082=>"11111101",
  54083=>"00000001",
  54084=>"11111110",
  54085=>"00000001",
  54086=>"00000011",
  54087=>"00000011",
  54088=>"11111111",
  54089=>"11111101",
  54090=>"00000010",
  54091=>"00000101",
  54092=>"11111111",
  54093=>"11111100",
  54094=>"00000000",
  54095=>"11111110",
  54096=>"00000000",
  54097=>"11111110",
  54098=>"11111110",
  54099=>"00000110",
  54100=>"00000000",
  54101=>"00000001",
  54102=>"11111111",
  54103=>"11111111",
  54104=>"11111110",
  54105=>"00000010",
  54106=>"11111110",
  54107=>"00000010",
  54108=>"00000000",
  54109=>"00000000",
  54110=>"11111110",
  54111=>"00000011",
  54112=>"00000000",
  54113=>"11111110",
  54114=>"00000100",
  54115=>"00000101",
  54116=>"11111101",
  54117=>"00000001",
  54118=>"11111110",
  54119=>"11111111",
  54120=>"00000001",
  54121=>"11111101",
  54122=>"11111111",
  54123=>"00000000",
  54124=>"11111100",
  54125=>"00000010",
  54126=>"11111100",
  54127=>"00000001",
  54128=>"11111100",
  54129=>"11111110",
  54130=>"11111111",
  54131=>"00000001",
  54132=>"11111110",
  54133=>"00000001",
  54134=>"11111101",
  54135=>"00000001",
  54136=>"00000000",
  54137=>"11111111",
  54138=>"00000000",
  54139=>"11111101",
  54140=>"11111111",
  54141=>"00000000",
  54142=>"11111101",
  54143=>"00000011",
  54144=>"00000010",
  54145=>"00000111",
  54146=>"11111110",
  54147=>"00000111",
  54148=>"11111111",
  54149=>"00000100",
  54150=>"11111111",
  54151=>"00000100",
  54152=>"00000100",
  54153=>"11111111",
  54154=>"00000010",
  54155=>"00000010",
  54156=>"11111111",
  54157=>"00000010",
  54158=>"00000000",
  54159=>"11111111",
  54160=>"00000010",
  54161=>"00000001",
  54162=>"11111100",
  54163=>"11111110",
  54164=>"11111111",
  54165=>"11111110",
  54166=>"00000001",
  54167=>"00000011",
  54168=>"00000001",
  54169=>"11111110",
  54170=>"00000011",
  54171=>"11111101",
  54172=>"00000001",
  54173=>"00000010",
  54174=>"11111101",
  54175=>"00000100",
  54176=>"00000100",
  54177=>"00000000",
  54178=>"11111111",
  54179=>"11111110",
  54180=>"11111111",
  54181=>"11111101",
  54182=>"11111111",
  54183=>"11111111",
  54184=>"00000001",
  54185=>"00000001",
  54186=>"11111111",
  54187=>"11111101",
  54188=>"00000011",
  54189=>"11111111",
  54190=>"00000000",
  54191=>"00000010",
  54192=>"11111100",
  54193=>"00000100",
  54194=>"00000001",
  54195=>"11111111",
  54196=>"11111101",
  54197=>"11111111",
  54198=>"11111111",
  54199=>"00000010",
  54200=>"00000010",
  54201=>"11111101",
  54202=>"00000110",
  54203=>"00000010",
  54204=>"00000011",
  54205=>"11111101",
  54206=>"00000011",
  54207=>"00000001",
  54208=>"00000001",
  54209=>"11111111",
  54210=>"11111101",
  54211=>"00000100",
  54212=>"00000000",
  54213=>"11111111",
  54214=>"11111101",
  54215=>"11111111",
  54216=>"11111110",
  54217=>"11111111",
  54218=>"11111111",
  54219=>"00000001",
  54220=>"00000010",
  54221=>"00000011",
  54222=>"00000000",
  54223=>"00000010",
  54224=>"00000011",
  54225=>"11111101",
  54226=>"11111110",
  54227=>"00000010",
  54228=>"00000001",
  54229=>"00000000",
  54230=>"00000000",
  54231=>"11111111",
  54232=>"00000000",
  54233=>"00000001",
  54234=>"00000001",
  54235=>"00000000",
  54236=>"00000001",
  54237=>"00000101",
  54238=>"00000001",
  54239=>"11111111",
  54240=>"00000010",
  54241=>"00000000",
  54242=>"11111110",
  54243=>"11111110",
  54244=>"00000001",
  54245=>"11111111",
  54246=>"11111110",
  54247=>"00000011",
  54248=>"00000010",
  54249=>"00000001",
  54250=>"00000011",
  54251=>"00000000",
  54252=>"00000001",
  54253=>"00000001",
  54254=>"11111110",
  54255=>"11111110",
  54256=>"11111101",
  54257=>"00000000",
  54258=>"11111111",
  54259=>"00000001",
  54260=>"11111110",
  54261=>"00000010",
  54262=>"11111110",
  54263=>"00000001",
  54264=>"00000000",
  54265=>"00000000",
  54266=>"11111100",
  54267=>"11111101",
  54268=>"00000000",
  54269=>"11111110",
  54270=>"00000001",
  54271=>"00000010",
  54272=>"00000010",
  54273=>"00000001",
  54274=>"00000001",
  54275=>"11111111",
  54276=>"11111100",
  54277=>"11111110",
  54278=>"11111111",
  54279=>"00000001",
  54280=>"00000001",
  54281=>"00000011",
  54282=>"00000000",
  54283=>"11111111",
  54284=>"00000101",
  54285=>"00000001",
  54286=>"00000001",
  54287=>"00000100",
  54288=>"11111110",
  54289=>"00000000",
  54290=>"00000001",
  54291=>"00000000",
  54292=>"00000001",
  54293=>"00000010",
  54294=>"00000000",
  54295=>"00000010",
  54296=>"11111110",
  54297=>"11111110",
  54298=>"00000000",
  54299=>"00000000",
  54300=>"00000100",
  54301=>"00000000",
  54302=>"11111111",
  54303=>"11111111",
  54304=>"11111101",
  54305=>"11111101",
  54306=>"00000100",
  54307=>"11111111",
  54308=>"00000000",
  54309=>"11111101",
  54310=>"11111110",
  54311=>"11111110",
  54312=>"00000101",
  54313=>"00000010",
  54314=>"11111111",
  54315=>"00000000",
  54316=>"00000000",
  54317=>"00000000",
  54318=>"00000001",
  54319=>"11111110",
  54320=>"11111111",
  54321=>"11111111",
  54322=>"00000000",
  54323=>"11111111",
  54324=>"11111101",
  54325=>"00000100",
  54326=>"00000001",
  54327=>"11111111",
  54328=>"11111101",
  54329=>"00000100",
  54330=>"11111101",
  54331=>"00000001",
  54332=>"11111111",
  54333=>"00000001",
  54334=>"11111111",
  54335=>"11111111",
  54336=>"11111101",
  54337=>"00000011",
  54338=>"00000110",
  54339=>"00000001",
  54340=>"11111111",
  54341=>"11111100",
  54342=>"00000010",
  54343=>"11111111",
  54344=>"00000001",
  54345=>"00000000",
  54346=>"11111101",
  54347=>"11111110",
  54348=>"00000010",
  54349=>"00000000",
  54350=>"11111111",
  54351=>"11111101",
  54352=>"00000010",
  54353=>"11111100",
  54354=>"11111110",
  54355=>"00000000",
  54356=>"00000100",
  54357=>"11111110",
  54358=>"00000000",
  54359=>"11111110",
  54360=>"00000001",
  54361=>"00000010",
  54362=>"11111101",
  54363=>"00000100",
  54364=>"11111101",
  54365=>"11111111",
  54366=>"11111110",
  54367=>"11111100",
  54368=>"00000100",
  54369=>"00000011",
  54370=>"00000000",
  54371=>"11111101",
  54372=>"00000010",
  54373=>"11111111",
  54374=>"00000000",
  54375=>"00000010",
  54376=>"00000011",
  54377=>"11111111",
  54378=>"11111111",
  54379=>"00000000",
  54380=>"11111110",
  54381=>"11111110",
  54382=>"00000000",
  54383=>"11111101",
  54384=>"11111111",
  54385=>"00000001",
  54386=>"00000010",
  54387=>"11111111",
  54388=>"00000011",
  54389=>"11111101",
  54390=>"00000001",
  54391=>"00000010",
  54392=>"00000010",
  54393=>"00000010",
  54394=>"11111110",
  54395=>"00000001",
  54396=>"00000001",
  54397=>"00000000",
  54398=>"00000100",
  54399=>"11111100",
  54400=>"00000011",
  54401=>"11111110",
  54402=>"11111110",
  54403=>"11111110",
  54404=>"00000001",
  54405=>"00000100",
  54406=>"00000011",
  54407=>"11111111",
  54408=>"11111110",
  54409=>"00000101",
  54410=>"11111101",
  54411=>"11111111",
  54412=>"11111111",
  54413=>"00000011",
  54414=>"00000001",
  54415=>"00000011",
  54416=>"00000001",
  54417=>"11111111",
  54418=>"11111111",
  54419=>"00000010",
  54420=>"00000001",
  54421=>"00000100",
  54422=>"11111110",
  54423=>"11111101",
  54424=>"11111111",
  54425=>"00000010",
  54426=>"00000101",
  54427=>"00000010",
  54428=>"00000000",
  54429=>"00000001",
  54430=>"00000010",
  54431=>"00000001",
  54432=>"00000000",
  54433=>"11111101",
  54434=>"11111100",
  54435=>"11111111",
  54436=>"00000010",
  54437=>"11111010",
  54438=>"11111110",
  54439=>"00000000",
  54440=>"00000001",
  54441=>"00000001",
  54442=>"00000010",
  54443=>"11111110",
  54444=>"00000001",
  54445=>"11111111",
  54446=>"11111110",
  54447=>"00000001",
  54448=>"00000001",
  54449=>"00000000",
  54450=>"11111111",
  54451=>"00000000",
  54452=>"11111101",
  54453=>"00000001",
  54454=>"11111111",
  54455=>"00000100",
  54456=>"00000110",
  54457=>"11111111",
  54458=>"00000010",
  54459=>"11111100",
  54460=>"00000010",
  54461=>"00000001",
  54462=>"00000010",
  54463=>"00000001",
  54464=>"00000011",
  54465=>"11111101",
  54466=>"11111101",
  54467=>"00000001",
  54468=>"11111111",
  54469=>"11111111",
  54470=>"00000000",
  54471=>"00000110",
  54472=>"00000100",
  54473=>"00000000",
  54474=>"11111110",
  54475=>"00000001",
  54476=>"00000100",
  54477=>"11111110",
  54478=>"00000001",
  54479=>"00000000",
  54480=>"00000000",
  54481=>"00000000",
  54482=>"11111101",
  54483=>"00000100",
  54484=>"00000001",
  54485=>"00000011",
  54486=>"00000011",
  54487=>"11111111",
  54488=>"11111100",
  54489=>"00000010",
  54490=>"00000000",
  54491=>"00000011",
  54492=>"00000000",
  54493=>"11111111",
  54494=>"00000001",
  54495=>"11111110",
  54496=>"00000001",
  54497=>"00000011",
  54498=>"11111110",
  54499=>"00000011",
  54500=>"11111101",
  54501=>"11111101",
  54502=>"00000001",
  54503=>"11111110",
  54504=>"00000001",
  54505=>"00000011",
  54506=>"00000000",
  54507=>"11111111",
  54508=>"11111110",
  54509=>"11111111",
  54510=>"11111101",
  54511=>"00000010",
  54512=>"00000001",
  54513=>"11111011",
  54514=>"00000000",
  54515=>"11111111",
  54516=>"00000100",
  54517=>"00000101",
  54518=>"00000100",
  54519=>"00000100",
  54520=>"00000000",
  54521=>"11111111",
  54522=>"00000100",
  54523=>"11111111",
  54524=>"11111110",
  54525=>"00000001",
  54526=>"00000101",
  54527=>"11111110",
  54528=>"11111111",
  54529=>"00000100",
  54530=>"00000100",
  54531=>"11111110",
  54532=>"00000010",
  54533=>"11111111",
  54534=>"00000000",
  54535=>"11111111",
  54536=>"11111110",
  54537=>"11111011",
  54538=>"11111110",
  54539=>"11111111",
  54540=>"00000001",
  54541=>"11111100",
  54542=>"11111110",
  54543=>"11111111",
  54544=>"11111101",
  54545=>"00000010",
  54546=>"00000001",
  54547=>"00000100",
  54548=>"00000000",
  54549=>"11111111",
  54550=>"00000010",
  54551=>"11111111",
  54552=>"00000000",
  54553=>"00000001",
  54554=>"00000001",
  54555=>"11111111",
  54556=>"11111101",
  54557=>"00000000",
  54558=>"11111111",
  54559=>"00000000",
  54560=>"11111111",
  54561=>"11111110",
  54562=>"00000000",
  54563=>"11111011",
  54564=>"00000011",
  54565=>"11111111",
  54566=>"00000000",
  54567=>"00000010",
  54568=>"11111110",
  54569=>"00000000",
  54570=>"11111111",
  54571=>"00000010",
  54572=>"00000010",
  54573=>"00000000",
  54574=>"11111100",
  54575=>"00000010",
  54576=>"11111111",
  54577=>"00000011",
  54578=>"00000010",
  54579=>"00000000",
  54580=>"11111101",
  54581=>"00000000",
  54582=>"00000001",
  54583=>"00000001",
  54584=>"11111111",
  54585=>"11111110",
  54586=>"11111110",
  54587=>"00000001",
  54588=>"00000001",
  54589=>"00000001",
  54590=>"00000010",
  54591=>"00000000",
  54592=>"00000010",
  54593=>"00000011",
  54594=>"00000000",
  54595=>"00000001",
  54596=>"00000001",
  54597=>"11111110",
  54598=>"00000100",
  54599=>"11111101",
  54600=>"00000101",
  54601=>"11111101",
  54602=>"00000001",
  54603=>"00000001",
  54604=>"00000000",
  54605=>"11111101",
  54606=>"00000000",
  54607=>"00000000",
  54608=>"00000001",
  54609=>"11111111",
  54610=>"11111111",
  54611=>"00000110",
  54612=>"11111101",
  54613=>"11111111",
  54614=>"00000000",
  54615=>"00000011",
  54616=>"11111111",
  54617=>"00000011",
  54618=>"11111101",
  54619=>"00000101",
  54620=>"00000000",
  54621=>"11111110",
  54622=>"00000010",
  54623=>"00000001",
  54624=>"00000010",
  54625=>"00000001",
  54626=>"11111110",
  54627=>"00000010",
  54628=>"00000000",
  54629=>"11111101",
  54630=>"00000101",
  54631=>"11111111",
  54632=>"11111101",
  54633=>"00000000",
  54634=>"11111111",
  54635=>"00000010",
  54636=>"00000001",
  54637=>"00000001",
  54638=>"00000101",
  54639=>"00000001",
  54640=>"11111110",
  54641=>"00000001",
  54642=>"11111111",
  54643=>"11111110",
  54644=>"00000100",
  54645=>"11111100",
  54646=>"00000110",
  54647=>"11111110",
  54648=>"11111110",
  54649=>"11111110",
  54650=>"11111100",
  54651=>"00000001",
  54652=>"00000001",
  54653=>"00000010",
  54654=>"00000000",
  54655=>"11111110",
  54656=>"11111100",
  54657=>"00000001",
  54658=>"00000100",
  54659=>"00000010",
  54660=>"00000001",
  54661=>"00000011",
  54662=>"11111111",
  54663=>"00000010",
  54664=>"11111111",
  54665=>"00000001",
  54666=>"11111111",
  54667=>"00000010",
  54668=>"00000000",
  54669=>"00000001",
  54670=>"11111110",
  54671=>"00000001",
  54672=>"11111111",
  54673=>"00000010",
  54674=>"11111100",
  54675=>"00000001",
  54676=>"00000110",
  54677=>"11111101",
  54678=>"11111101",
  54679=>"11111110",
  54680=>"11111111",
  54681=>"11111110",
  54682=>"11111100",
  54683=>"00000001",
  54684=>"11111101",
  54685=>"11111111",
  54686=>"00000010",
  54687=>"11111101",
  54688=>"11111101",
  54689=>"00000010",
  54690=>"11111110",
  54691=>"00000000",
  54692=>"00000000",
  54693=>"00000010",
  54694=>"00000100",
  54695=>"00000001",
  54696=>"00000000",
  54697=>"00000010",
  54698=>"00000010",
  54699=>"11111101",
  54700=>"11111110",
  54701=>"11111100",
  54702=>"00000001",
  54703=>"11111111",
  54704=>"00000010",
  54705=>"11111100",
  54706=>"11111110",
  54707=>"00000011",
  54708=>"11111101",
  54709=>"11111100",
  54710=>"00000100",
  54711=>"11111110",
  54712=>"11111110",
  54713=>"11111100",
  54714=>"11111101",
  54715=>"00000000",
  54716=>"00000000",
  54717=>"11111110",
  54718=>"00000100",
  54719=>"00000000",
  54720=>"00000011",
  54721=>"11111101",
  54722=>"00000010",
  54723=>"00000001",
  54724=>"00000001",
  54725=>"11111111",
  54726=>"11111111",
  54727=>"11111111",
  54728=>"00000010",
  54729=>"11111101",
  54730=>"11111111",
  54731=>"00000001",
  54732=>"11111100",
  54733=>"11111111",
  54734=>"11111110",
  54735=>"11111100",
  54736=>"00000000",
  54737=>"00000001",
  54738=>"00000011",
  54739=>"00000001",
  54740=>"00000001",
  54741=>"00000011",
  54742=>"11111110",
  54743=>"11111111",
  54744=>"00000010",
  54745=>"11111101",
  54746=>"00000010",
  54747=>"11111101",
  54748=>"11111101",
  54749=>"00000001",
  54750=>"00000100",
  54751=>"11111100",
  54752=>"00000001",
  54753=>"11111111",
  54754=>"00000010",
  54755=>"00000000",
  54756=>"00000000",
  54757=>"11111101",
  54758=>"00000001",
  54759=>"11111111",
  54760=>"11111111",
  54761=>"11111111",
  54762=>"11111111",
  54763=>"00000000",
  54764=>"00000100",
  54765=>"11111111",
  54766=>"11111111",
  54767=>"00000000",
  54768=>"11111101",
  54769=>"11111101",
  54770=>"00000010",
  54771=>"00000010",
  54772=>"11111101",
  54773=>"00000001",
  54774=>"00000001",
  54775=>"11111100",
  54776=>"00000000",
  54777=>"11111101",
  54778=>"11111110",
  54779=>"11111101",
  54780=>"11111110",
  54781=>"11111111",
  54782=>"11111110",
  54783=>"00000010",
  54784=>"00000000",
  54785=>"00000010",
  54786=>"00000010",
  54787=>"00000010",
  54788=>"11111100",
  54789=>"11111111",
  54790=>"11111110",
  54791=>"11111100",
  54792=>"00000010",
  54793=>"11111111",
  54794=>"00000010",
  54795=>"00000000",
  54796=>"00000011",
  54797=>"11111110",
  54798=>"00000000",
  54799=>"00000101",
  54800=>"00000000",
  54801=>"00000000",
  54802=>"00000011",
  54803=>"00000101",
  54804=>"11111110",
  54805=>"11111101",
  54806=>"11111110",
  54807=>"11111110",
  54808=>"11111111",
  54809=>"11111110",
  54810=>"11111111",
  54811=>"00000001",
  54812=>"00000000",
  54813=>"11111111",
  54814=>"00000000",
  54815=>"00000010",
  54816=>"00000010",
  54817=>"00000010",
  54818=>"00000100",
  54819=>"11111110",
  54820=>"00000000",
  54821=>"11111111",
  54822=>"00000000",
  54823=>"11111101",
  54824=>"00000000",
  54825=>"11111110",
  54826=>"00000000",
  54827=>"00000000",
  54828=>"00000001",
  54829=>"00000000",
  54830=>"11111111",
  54831=>"11111111",
  54832=>"00000010",
  54833=>"00000000",
  54834=>"00000000",
  54835=>"11111110",
  54836=>"11111111",
  54837=>"11111110",
  54838=>"00000000",
  54839=>"11111101",
  54840=>"00000010",
  54841=>"00000001",
  54842=>"00000000",
  54843=>"11111111",
  54844=>"11111110",
  54845=>"00000010",
  54846=>"00000000",
  54847=>"11111111",
  54848=>"00000100",
  54849=>"11111111",
  54850=>"00000001",
  54851=>"11111110",
  54852=>"00000010",
  54853=>"11111111",
  54854=>"00000000",
  54855=>"00000000",
  54856=>"00000000",
  54857=>"11111110",
  54858=>"11111101",
  54859=>"11111111",
  54860=>"11111110",
  54861=>"00000000",
  54862=>"00000011",
  54863=>"00000000",
  54864=>"11111110",
  54865=>"00000000",
  54866=>"00000001",
  54867=>"11111101",
  54868=>"11111101",
  54869=>"11111101",
  54870=>"11111100",
  54871=>"00000010",
  54872=>"00000011",
  54873=>"00000001",
  54874=>"11111111",
  54875=>"00000010",
  54876=>"00000010",
  54877=>"11111101",
  54878=>"11111110",
  54879=>"00000010",
  54880=>"11111111",
  54881=>"00000101",
  54882=>"00000110",
  54883=>"11111100",
  54884=>"11111110",
  54885=>"00000101",
  54886=>"00000001",
  54887=>"00000001",
  54888=>"11111100",
  54889=>"11111111",
  54890=>"11111111",
  54891=>"00000000",
  54892=>"11111111",
  54893=>"11111110",
  54894=>"11111100",
  54895=>"00000001",
  54896=>"00000001",
  54897=>"00000010",
  54898=>"00000001",
  54899=>"00000001",
  54900=>"11111110",
  54901=>"00000010",
  54902=>"00000001",
  54903=>"00000001",
  54904=>"00000001",
  54905=>"11111110",
  54906=>"00000100",
  54907=>"11111100",
  54908=>"11111111",
  54909=>"11111110",
  54910=>"00000000",
  54911=>"00000010",
  54912=>"11111110",
  54913=>"11111111",
  54914=>"00000110",
  54915=>"11111111",
  54916=>"11111100",
  54917=>"00000011",
  54918=>"11111110",
  54919=>"11111110",
  54920=>"00000000",
  54921=>"00000010",
  54922=>"00000010",
  54923=>"00000001",
  54924=>"00000010",
  54925=>"00000011",
  54926=>"00000100",
  54927=>"00000011",
  54928=>"00000010",
  54929=>"00001000",
  54930=>"11111111",
  54931=>"00000010",
  54932=>"00000001",
  54933=>"11111101",
  54934=>"00000101",
  54935=>"11111101",
  54936=>"11111111",
  54937=>"00000011",
  54938=>"11111110",
  54939=>"00000000",
  54940=>"11111011",
  54941=>"11111110",
  54942=>"00000000",
  54943=>"11111101",
  54944=>"11111111",
  54945=>"11111111",
  54946=>"00000000",
  54947=>"11111111",
  54948=>"00000011",
  54949=>"11111100",
  54950=>"00000001",
  54951=>"11111101",
  54952=>"00000000",
  54953=>"00000001",
  54954=>"11111110",
  54955=>"00000011",
  54956=>"11111111",
  54957=>"00000010",
  54958=>"11111110",
  54959=>"00000000",
  54960=>"11111111",
  54961=>"00000001",
  54962=>"11111110",
  54963=>"11111111",
  54964=>"11111111",
  54965=>"00000001",
  54966=>"00000001",
  54967=>"00000001",
  54968=>"00000001",
  54969=>"11111111",
  54970=>"11111111",
  54971=>"00000001",
  54972=>"00000000",
  54973=>"11111111",
  54974=>"00000000",
  54975=>"00000010",
  54976=>"00000000",
  54977=>"00000011",
  54978=>"11111110",
  54979=>"11111111",
  54980=>"00000011",
  54981=>"11111011",
  54982=>"11111111",
  54983=>"00000000",
  54984=>"00000000",
  54985=>"11111111",
  54986=>"11111101",
  54987=>"11111100",
  54988=>"11111111",
  54989=>"11111110",
  54990=>"11111110",
  54991=>"11111110",
  54992=>"00000001",
  54993=>"11111111",
  54994=>"00000000",
  54995=>"11111101",
  54996=>"11111101",
  54997=>"11111110",
  54998=>"00000001",
  54999=>"00000011",
  55000=>"00000011",
  55001=>"00000101",
  55002=>"00000000",
  55003=>"11111101",
  55004=>"11111110",
  55005=>"00000001",
  55006=>"00000011",
  55007=>"00000010",
  55008=>"00000000",
  55009=>"11111110",
  55010=>"11111110",
  55011=>"11111110",
  55012=>"11111110",
  55013=>"00000010",
  55014=>"00000010",
  55015=>"00000001",
  55016=>"00000000",
  55017=>"00000010",
  55018=>"00000001",
  55019=>"11111110",
  55020=>"00000010",
  55021=>"11111110",
  55022=>"11111111",
  55023=>"00000001",
  55024=>"11111111",
  55025=>"00000101",
  55026=>"00000001",
  55027=>"00000001",
  55028=>"11111111",
  55029=>"00000010",
  55030=>"00000010",
  55031=>"00000011",
  55032=>"00000010",
  55033=>"11111110",
  55034=>"00000100",
  55035=>"00000001",
  55036=>"00000001",
  55037=>"00000010",
  55038=>"00000000",
  55039=>"00000000",
  55040=>"11111101",
  55041=>"11111110",
  55042=>"00000001",
  55043=>"11111110",
  55044=>"00000010",
  55045=>"11111110",
  55046=>"11111110",
  55047=>"00000001",
  55048=>"11111101",
  55049=>"11111101",
  55050=>"00000001",
  55051=>"11111111",
  55052=>"11111111",
  55053=>"00000001",
  55054=>"00000000",
  55055=>"00000001",
  55056=>"00000000",
  55057=>"11111111",
  55058=>"11111110",
  55059=>"00000011",
  55060=>"11111111",
  55061=>"00000010",
  55062=>"00000010",
  55063=>"11111111",
  55064=>"00000011",
  55065=>"00000100",
  55066=>"11111101",
  55067=>"00000001",
  55068=>"00000010",
  55069=>"00000100",
  55070=>"11111101",
  55071=>"00000010",
  55072=>"00000010",
  55073=>"00000001",
  55074=>"11111110",
  55075=>"00000010",
  55076=>"11111110",
  55077=>"00000001",
  55078=>"11111111",
  55079=>"11111111",
  55080=>"00000011",
  55081=>"00000100",
  55082=>"11111111",
  55083=>"00000011",
  55084=>"00000011",
  55085=>"11111111",
  55086=>"00000000",
  55087=>"00000001",
  55088=>"11111111",
  55089=>"00000010",
  55090=>"00000001",
  55091=>"11111110",
  55092=>"00000001",
  55093=>"11111110",
  55094=>"00000001",
  55095=>"00000011",
  55096=>"00000001",
  55097=>"00000001",
  55098=>"11111111",
  55099=>"11111100",
  55100=>"00000001",
  55101=>"00000010",
  55102=>"00000011",
  55103=>"00000001",
  55104=>"11111101",
  55105=>"11111100",
  55106=>"00000100",
  55107=>"00000000",
  55108=>"00000000",
  55109=>"00000011",
  55110=>"00000100",
  55111=>"11111111",
  55112=>"00000011",
  55113=>"11111111",
  55114=>"00000001",
  55115=>"00000100",
  55116=>"00000001",
  55117=>"11111100",
  55118=>"11111101",
  55119=>"00000100",
  55120=>"11111011",
  55121=>"00000010",
  55122=>"00000010",
  55123=>"00000000",
  55124=>"11111110",
  55125=>"00000001",
  55126=>"11111111",
  55127=>"11111111",
  55128=>"11111111",
  55129=>"00000001",
  55130=>"00000001",
  55131=>"11111110",
  55132=>"11111110",
  55133=>"11111110",
  55134=>"11111111",
  55135=>"00000001",
  55136=>"11111111",
  55137=>"11111111",
  55138=>"11111110",
  55139=>"11111101",
  55140=>"11111110",
  55141=>"11111100",
  55142=>"00000000",
  55143=>"11111101",
  55144=>"11111111",
  55145=>"00000010",
  55146=>"00000001",
  55147=>"11111111",
  55148=>"00000101",
  55149=>"00000001",
  55150=>"00000000",
  55151=>"00000010",
  55152=>"00000110",
  55153=>"00000010",
  55154=>"00000001",
  55155=>"00000100",
  55156=>"00000001",
  55157=>"11111101",
  55158=>"11111101",
  55159=>"00000010",
  55160=>"00000100",
  55161=>"00000000",
  55162=>"11111101",
  55163=>"11111110",
  55164=>"00000000",
  55165=>"00000001",
  55166=>"00000010",
  55167=>"11111100",
  55168=>"00000010",
  55169=>"11111110",
  55170=>"00000010",
  55171=>"11111100",
  55172=>"11111111",
  55173=>"00000010",
  55174=>"11111110",
  55175=>"00000010",
  55176=>"11111111",
  55177=>"00000010",
  55178=>"11111110",
  55179=>"00000000",
  55180=>"11111101",
  55181=>"00000100",
  55182=>"00000000",
  55183=>"00000011",
  55184=>"00000001",
  55185=>"11111101",
  55186=>"00000000",
  55187=>"11111110",
  55188=>"11111111",
  55189=>"11111100",
  55190=>"11111110",
  55191=>"11111101",
  55192=>"11111111",
  55193=>"11111110",
  55194=>"11111111",
  55195=>"00000010",
  55196=>"00000110",
  55197=>"00000000",
  55198=>"00000000",
  55199=>"00000001",
  55200=>"00000001",
  55201=>"00000001",
  55202=>"00000101",
  55203=>"00000100",
  55204=>"11111111",
  55205=>"00000001",
  55206=>"00000010",
  55207=>"11111110",
  55208=>"00000010",
  55209=>"00000010",
  55210=>"11111111",
  55211=>"00000010",
  55212=>"00000110",
  55213=>"11111110",
  55214=>"00000100",
  55215=>"00000001",
  55216=>"11111101",
  55217=>"11111111",
  55218=>"00000010",
  55219=>"00000000",
  55220=>"00000010",
  55221=>"11111011",
  55222=>"00000010",
  55223=>"11111110",
  55224=>"11111110",
  55225=>"11111110",
  55226=>"00000010",
  55227=>"11111101",
  55228=>"00000010",
  55229=>"11111110",
  55230=>"00000011",
  55231=>"00000001",
  55232=>"11111100",
  55233=>"00000010",
  55234=>"00000000",
  55235=>"00000000",
  55236=>"00000001",
  55237=>"11111111",
  55238=>"00000001",
  55239=>"00000000",
  55240=>"11111101",
  55241=>"11111110",
  55242=>"00000000",
  55243=>"11111101",
  55244=>"11111111",
  55245=>"11111111",
  55246=>"00000001",
  55247=>"00000010",
  55248=>"00000010",
  55249=>"00000000",
  55250=>"11111101",
  55251=>"00000001",
  55252=>"00000001",
  55253=>"11111101",
  55254=>"00000001",
  55255=>"00000111",
  55256=>"11111111",
  55257=>"00000000",
  55258=>"11111110",
  55259=>"11111101",
  55260=>"11111101",
  55261=>"11111100",
  55262=>"00000001",
  55263=>"11111110",
  55264=>"00000001",
  55265=>"11111110",
  55266=>"00000101",
  55267=>"00000000",
  55268=>"11111111",
  55269=>"00000010",
  55270=>"11111110",
  55271=>"00000010",
  55272=>"11111101",
  55273=>"00000000",
  55274=>"00000000",
  55275=>"11111111",
  55276=>"00000010",
  55277=>"11111111",
  55278=>"11111100",
  55279=>"00000001",
  55280=>"11111101",
  55281=>"00000001",
  55282=>"11111111",
  55283=>"00000010",
  55284=>"11111110",
  55285=>"00000000",
  55286=>"00000001",
  55287=>"00000001",
  55288=>"11111101",
  55289=>"00000010",
  55290=>"00000100",
  55291=>"11111110",
  55292=>"11111010",
  55293=>"00000001",
  55294=>"11111111",
  55295=>"00000010",
  55296=>"00000011",
  55297=>"00000001",
  55298=>"00000001",
  55299=>"11111111",
  55300=>"11111110",
  55301=>"00000000",
  55302=>"11111110",
  55303=>"11111110",
  55304=>"11111110",
  55305=>"00000001",
  55306=>"00000001",
  55307=>"11111110",
  55308=>"11111101",
  55309=>"11111111",
  55310=>"00000010",
  55311=>"11111110",
  55312=>"00000011",
  55313=>"00000001",
  55314=>"11111101",
  55315=>"11111111",
  55316=>"00000010",
  55317=>"00000010",
  55318=>"00000100",
  55319=>"11111101",
  55320=>"00000001",
  55321=>"00000010",
  55322=>"11111111",
  55323=>"00000011",
  55324=>"00000010",
  55325=>"11111101",
  55326=>"00000001",
  55327=>"00000001",
  55328=>"00000011",
  55329=>"11111110",
  55330=>"11111100",
  55331=>"00000011",
  55332=>"00000001",
  55333=>"11111110",
  55334=>"11111101",
  55335=>"00000100",
  55336=>"00000100",
  55337=>"00000100",
  55338=>"11111100",
  55339=>"00000001",
  55340=>"00000000",
  55341=>"11111101",
  55342=>"11111110",
  55343=>"11111111",
  55344=>"00000000",
  55345=>"11111110",
  55346=>"00000001",
  55347=>"11111111",
  55348=>"11111101",
  55349=>"00000001",
  55350=>"00000001",
  55351=>"00000010",
  55352=>"00000001",
  55353=>"11111101",
  55354=>"00000000",
  55355=>"11111110",
  55356=>"11111110",
  55357=>"00000000",
  55358=>"11111110",
  55359=>"00000011",
  55360=>"00000011",
  55361=>"11111110",
  55362=>"00000101",
  55363=>"11111111",
  55364=>"11111110",
  55365=>"11111101",
  55366=>"00000000",
  55367=>"00000010",
  55368=>"00000011",
  55369=>"00000001",
  55370=>"00000011",
  55371=>"00000000",
  55372=>"00000001",
  55373=>"11111101",
  55374=>"00000011",
  55375=>"00000101",
  55376=>"11111111",
  55377=>"00000001",
  55378=>"11111110",
  55379=>"11111111",
  55380=>"00000000",
  55381=>"11111110",
  55382=>"11111111",
  55383=>"11111111",
  55384=>"11111111",
  55385=>"00000101",
  55386=>"00000000",
  55387=>"00000000",
  55388=>"11111110",
  55389=>"00000001",
  55390=>"00000000",
  55391=>"11111100",
  55392=>"00000010",
  55393=>"00000000",
  55394=>"00000000",
  55395=>"11111101",
  55396=>"00000000",
  55397=>"00000100",
  55398=>"11111110",
  55399=>"11111111",
  55400=>"11111111",
  55401=>"11111100",
  55402=>"00000001",
  55403=>"00000010",
  55404=>"11111100",
  55405=>"00000011",
  55406=>"00000001",
  55407=>"00000000",
  55408=>"00000001",
  55409=>"11111101",
  55410=>"00000010",
  55411=>"11111101",
  55412=>"11111111",
  55413=>"11111101",
  55414=>"00000001",
  55415=>"00000010",
  55416=>"11111100",
  55417=>"11111110",
  55418=>"11111110",
  55419=>"11111111",
  55420=>"11111101",
  55421=>"11111110",
  55422=>"00000011",
  55423=>"00000101",
  55424=>"00000010",
  55425=>"11111101",
  55426=>"11111110",
  55427=>"11111110",
  55428=>"11111101",
  55429=>"11111111",
  55430=>"00000000",
  55431=>"11111110",
  55432=>"11111111",
  55433=>"11111111",
  55434=>"11111100",
  55435=>"11111111",
  55436=>"11111111",
  55437=>"00000010",
  55438=>"00000011",
  55439=>"11111110",
  55440=>"11111101",
  55441=>"00000000",
  55442=>"11111111",
  55443=>"11111111",
  55444=>"00000101",
  55445=>"00000001",
  55446=>"11111100",
  55447=>"11111101",
  55448=>"11111100",
  55449=>"11111110",
  55450=>"11111111",
  55451=>"11111111",
  55452=>"00000000",
  55453=>"11111101",
  55454=>"11111110",
  55455=>"00000010",
  55456=>"11111111",
  55457=>"11111110",
  55458=>"11111011",
  55459=>"11111111",
  55460=>"00000000",
  55461=>"00000001",
  55462=>"00000010",
  55463=>"00000011",
  55464=>"11111101",
  55465=>"00000100",
  55466=>"00000000",
  55467=>"00000000",
  55468=>"00000011",
  55469=>"11111111",
  55470=>"11111111",
  55471=>"00000011",
  55472=>"11111110",
  55473=>"00000100",
  55474=>"11111110",
  55475=>"11111101",
  55476=>"00000001",
  55477=>"11111110",
  55478=>"11111101",
  55479=>"00000001",
  55480=>"00000001",
  55481=>"00000011",
  55482=>"00000001",
  55483=>"11111111",
  55484=>"11111101",
  55485=>"00000001",
  55486=>"11111111",
  55487=>"00000000",
  55488=>"00000111",
  55489=>"11111111",
  55490=>"00000010",
  55491=>"00000000",
  55492=>"00000001",
  55493=>"11111111",
  55494=>"11111111",
  55495=>"00000010",
  55496=>"00000010",
  55497=>"00000101",
  55498=>"11111110",
  55499=>"00000000",
  55500=>"11111100",
  55501=>"00000001",
  55502=>"00000000",
  55503=>"11111111",
  55504=>"00000000",
  55505=>"00000100",
  55506=>"00000000",
  55507=>"11111110",
  55508=>"11111110",
  55509=>"00000010",
  55510=>"00000100",
  55511=>"11111111",
  55512=>"11111111",
  55513=>"11111111",
  55514=>"00000001",
  55515=>"11111111",
  55516=>"11111110",
  55517=>"00000001",
  55518=>"00000011",
  55519=>"11111111",
  55520=>"11111101",
  55521=>"00000000",
  55522=>"00000010",
  55523=>"00000100",
  55524=>"11111110",
  55525=>"11111110",
  55526=>"00000011",
  55527=>"00000001",
  55528=>"11111111",
  55529=>"11111100",
  55530=>"11111111",
  55531=>"11111111",
  55532=>"00000011",
  55533=>"00000001",
  55534=>"00000000",
  55535=>"00000000",
  55536=>"00000000",
  55537=>"00000111",
  55538=>"00000010",
  55539=>"00000010",
  55540=>"00000001",
  55541=>"00000001",
  55542=>"00000010",
  55543=>"00000100",
  55544=>"00000000",
  55545=>"11111111",
  55546=>"11111100",
  55547=>"00000000",
  55548=>"00000011",
  55549=>"11111101",
  55550=>"00000001",
  55551=>"11111101",
  55552=>"00000001",
  55553=>"11111111",
  55554=>"11111101",
  55555=>"00000001",
  55556=>"00000010",
  55557=>"00000010",
  55558=>"00000001",
  55559=>"11111100",
  55560=>"11111110",
  55561=>"11111110",
  55562=>"00000000",
  55563=>"11111110",
  55564=>"00000011",
  55565=>"00000010",
  55566=>"00000001",
  55567=>"00000000",
  55568=>"00000011",
  55569=>"11111111",
  55570=>"11111110",
  55571=>"00000011",
  55572=>"00000001",
  55573=>"11111101",
  55574=>"11111111",
  55575=>"11111101",
  55576=>"11111110",
  55577=>"00000011",
  55578=>"00000000",
  55579=>"11111111",
  55580=>"11111100",
  55581=>"11111101",
  55582=>"00000000",
  55583=>"00000010",
  55584=>"00000011",
  55585=>"11111111",
  55586=>"00000001",
  55587=>"00000011",
  55588=>"11111101",
  55589=>"11111111",
  55590=>"00000100",
  55591=>"11111111",
  55592=>"00000000",
  55593=>"00000000",
  55594=>"00000000",
  55595=>"00000000",
  55596=>"11111110",
  55597=>"11111111",
  55598=>"11111101",
  55599=>"11111101",
  55600=>"00000001",
  55601=>"11111110",
  55602=>"11111111",
  55603=>"00000011",
  55604=>"11111111",
  55605=>"11111101",
  55606=>"00000010",
  55607=>"00000010",
  55608=>"00000010",
  55609=>"11111110",
  55610=>"11111111",
  55611=>"00000011",
  55612=>"00000001",
  55613=>"00000001",
  55614=>"00000000",
  55615=>"00000001",
  55616=>"11111110",
  55617=>"00000100",
  55618=>"11111111",
  55619=>"11111111",
  55620=>"00000011",
  55621=>"11111101",
  55622=>"00000101",
  55623=>"00000001",
  55624=>"00000001",
  55625=>"00000100",
  55626=>"11111110",
  55627=>"00000001",
  55628=>"00000101",
  55629=>"11111111",
  55630=>"00000000",
  55631=>"11111111",
  55632=>"00000010",
  55633=>"00000000",
  55634=>"00000000",
  55635=>"11111101",
  55636=>"11111101",
  55637=>"11111111",
  55638=>"11111111",
  55639=>"00000100",
  55640=>"00000001",
  55641=>"00000010",
  55642=>"00000100",
  55643=>"11111110",
  55644=>"11111110",
  55645=>"00000001",
  55646=>"11111101",
  55647=>"11111111",
  55648=>"00000010",
  55649=>"00000010",
  55650=>"00000001",
  55651=>"00000010",
  55652=>"00000001",
  55653=>"00000001",
  55654=>"00000100",
  55655=>"11111101",
  55656=>"11111111",
  55657=>"00000011",
  55658=>"00000000",
  55659=>"11111101",
  55660=>"11111110",
  55661=>"11111111",
  55662=>"11111101",
  55663=>"00000011",
  55664=>"11111111",
  55665=>"00000000",
  55666=>"11111111",
  55667=>"00000000",
  55668=>"00000011",
  55669=>"11111110",
  55670=>"11111110",
  55671=>"00000010",
  55672=>"11111110",
  55673=>"00000011",
  55674=>"11111111",
  55675=>"11111111",
  55676=>"00000100",
  55677=>"11111111",
  55678=>"00000010",
  55679=>"00000010",
  55680=>"00000000",
  55681=>"00000011",
  55682=>"00000011",
  55683=>"11111111",
  55684=>"00000000",
  55685=>"00000000",
  55686=>"00000001",
  55687=>"00000001",
  55688=>"11111110",
  55689=>"11111100",
  55690=>"11111101",
  55691=>"00000000",
  55692=>"00000001",
  55693=>"11111110",
  55694=>"00000000",
  55695=>"00000001",
  55696=>"00000001",
  55697=>"00000010",
  55698=>"11111111",
  55699=>"00000001",
  55700=>"11111111",
  55701=>"00000001",
  55702=>"11111110",
  55703=>"00000001",
  55704=>"11111101",
  55705=>"00000010",
  55706=>"11111101",
  55707=>"11111101",
  55708=>"11111101",
  55709=>"00000001",
  55710=>"11111101",
  55711=>"00000100",
  55712=>"00000001",
  55713=>"00000011",
  55714=>"11111101",
  55715=>"11111101",
  55716=>"00000000",
  55717=>"00000001",
  55718=>"00000101",
  55719=>"00000001",
  55720=>"00000010",
  55721=>"00000100",
  55722=>"11111110",
  55723=>"11111101",
  55724=>"11111101",
  55725=>"00000001",
  55726=>"00000000",
  55727=>"00000010",
  55728=>"11111110",
  55729=>"00000000",
  55730=>"00000000",
  55731=>"00000001",
  55732=>"11111110",
  55733=>"00001000",
  55734=>"11111110",
  55735=>"00000000",
  55736=>"00000001",
  55737=>"11111110",
  55738=>"00000000",
  55739=>"00000001",
  55740=>"11111111",
  55741=>"00000010",
  55742=>"11111111",
  55743=>"00000011",
  55744=>"00000000",
  55745=>"00000001",
  55746=>"00000010",
  55747=>"00000001",
  55748=>"11111110",
  55749=>"00000100",
  55750=>"00000001",
  55751=>"00000010",
  55752=>"11111111",
  55753=>"00000001",
  55754=>"00000011",
  55755=>"00000010",
  55756=>"11111110",
  55757=>"00000010",
  55758=>"00000000",
  55759=>"00000001",
  55760=>"00000000",
  55761=>"11111101",
  55762=>"11111111",
  55763=>"00000010",
  55764=>"11111101",
  55765=>"00000000",
  55766=>"11111101",
  55767=>"00000001",
  55768=>"00000010",
  55769=>"00000001",
  55770=>"11111111",
  55771=>"11111100",
  55772=>"11111101",
  55773=>"00000101",
  55774=>"11111110",
  55775=>"00000011",
  55776=>"11111111",
  55777=>"00000010",
  55778=>"11111110",
  55779=>"00000010",
  55780=>"00000001",
  55781=>"00000001",
  55782=>"11111110",
  55783=>"11111111",
  55784=>"11111111",
  55785=>"11111101",
  55786=>"00000010",
  55787=>"00000000",
  55788=>"00000101",
  55789=>"11111111",
  55790=>"00000000",
  55791=>"00000010",
  55792=>"00000000",
  55793=>"00000011",
  55794=>"11111110",
  55795=>"00000000",
  55796=>"00000000",
  55797=>"11111110",
  55798=>"11111101",
  55799=>"11111111",
  55800=>"00000001",
  55801=>"00000011",
  55802=>"00000001",
  55803=>"00000010",
  55804=>"00000001",
  55805=>"00000011",
  55806=>"11111111",
  55807=>"11111110",
  55808=>"00000001",
  55809=>"00000001",
  55810=>"11111110",
  55811=>"11111110",
  55812=>"00000001",
  55813=>"11111111",
  55814=>"11111111",
  55815=>"00000010",
  55816=>"11111111",
  55817=>"11111111",
  55818=>"00000010",
  55819=>"11111111",
  55820=>"00000100",
  55821=>"11111110",
  55822=>"00000000",
  55823=>"11111110",
  55824=>"11111110",
  55825=>"00000011",
  55826=>"00000010",
  55827=>"00000010",
  55828=>"11111101",
  55829=>"11111110",
  55830=>"11111110",
  55831=>"00000011",
  55832=>"00000010",
  55833=>"00000000",
  55834=>"00000010",
  55835=>"00000000",
  55836=>"00000000",
  55837=>"11111111",
  55838=>"00000000",
  55839=>"11111100",
  55840=>"11111011",
  55841=>"00000000",
  55842=>"11111110",
  55843=>"00000001",
  55844=>"00000010",
  55845=>"00000000",
  55846=>"00000010",
  55847=>"11111110",
  55848=>"11111110",
  55849=>"11111110",
  55850=>"00000010",
  55851=>"00000010",
  55852=>"00000000",
  55853=>"11111110",
  55854=>"11111111",
  55855=>"00000001",
  55856=>"11111101",
  55857=>"11111110",
  55858=>"00000000",
  55859=>"11111110",
  55860=>"00000000",
  55861=>"00000001",
  55862=>"11111110",
  55863=>"11111110",
  55864=>"11111111",
  55865=>"00000010",
  55866=>"00000000",
  55867=>"00000010",
  55868=>"00000000",
  55869=>"00000110",
  55870=>"11111101",
  55871=>"11111111",
  55872=>"00000000",
  55873=>"11111111",
  55874=>"00000001",
  55875=>"11111111",
  55876=>"11111100",
  55877=>"11111111",
  55878=>"00000000",
  55879=>"11111100",
  55880=>"00000010",
  55881=>"11111110",
  55882=>"11111101",
  55883=>"11111110",
  55884=>"11111110",
  55885=>"11111111",
  55886=>"11111101",
  55887=>"00000001",
  55888=>"00000001",
  55889=>"00000000",
  55890=>"00000000",
  55891=>"11111101",
  55892=>"00000000",
  55893=>"00000000",
  55894=>"11111111",
  55895=>"00000001",
  55896=>"00000000",
  55897=>"00000010",
  55898=>"00000001",
  55899=>"00000010",
  55900=>"00000001",
  55901=>"00000010",
  55902=>"11111101",
  55903=>"00000000",
  55904=>"11111110",
  55905=>"11111100",
  55906=>"00000010",
  55907=>"11111100",
  55908=>"00000000",
  55909=>"00000001",
  55910=>"11111110",
  55911=>"11111110",
  55912=>"11111111",
  55913=>"11111110",
  55914=>"00000000",
  55915=>"00000010",
  55916=>"00000001",
  55917=>"00000001",
  55918=>"11111110",
  55919=>"00000000",
  55920=>"11111101",
  55921=>"00000010",
  55922=>"00000000",
  55923=>"11111111",
  55924=>"11111111",
  55925=>"11111101",
  55926=>"11111110",
  55927=>"00000010",
  55928=>"11111101",
  55929=>"11111110",
  55930=>"00000001",
  55931=>"00000101",
  55932=>"00000010",
  55933=>"00000001",
  55934=>"11111101",
  55935=>"11111101",
  55936=>"00000011",
  55937=>"11111110",
  55938=>"11111111",
  55939=>"11111110",
  55940=>"00000000",
  55941=>"11111111",
  55942=>"00000010",
  55943=>"11111110",
  55944=>"00000001",
  55945=>"11111101",
  55946=>"11111101",
  55947=>"00000001",
  55948=>"00000001",
  55949=>"00000001",
  55950=>"11111110",
  55951=>"00000010",
  55952=>"11111111",
  55953=>"11111101",
  55954=>"00000001",
  55955=>"00000001",
  55956=>"11111111",
  55957=>"00000001",
  55958=>"00000011",
  55959=>"11111110",
  55960=>"00000010",
  55961=>"11111101",
  55962=>"00000000",
  55963=>"00000001",
  55964=>"11111101",
  55965=>"00000001",
  55966=>"00000100",
  55967=>"00000011",
  55968=>"00000011",
  55969=>"11111110",
  55970=>"11111111",
  55971=>"00000000",
  55972=>"00000010",
  55973=>"00000011",
  55974=>"00000010",
  55975=>"00000000",
  55976=>"00000001",
  55977=>"00000001",
  55978=>"11111110",
  55979=>"00000000",
  55980=>"11111110",
  55981=>"00000001",
  55982=>"00000000",
  55983=>"11111111",
  55984=>"11111100",
  55985=>"00000111",
  55986=>"00000010",
  55987=>"00000000",
  55988=>"00000000",
  55989=>"11111111",
  55990=>"00000010",
  55991=>"00000001",
  55992=>"00000001",
  55993=>"11111111",
  55994=>"00000000",
  55995=>"00000010",
  55996=>"11111101",
  55997=>"11111110",
  55998=>"00000000",
  55999=>"11111101",
  56000=>"00000001",
  56001=>"11111101",
  56002=>"00000000",
  56003=>"11111110",
  56004=>"00000010",
  56005=>"00000000",
  56006=>"00000101",
  56007=>"00000011",
  56008=>"11111110",
  56009=>"11111110",
  56010=>"11111111",
  56011=>"11111110",
  56012=>"11111101",
  56013=>"00000010",
  56014=>"00000010",
  56015=>"11111110",
  56016=>"00000010",
  56017=>"00000010",
  56018=>"00000000",
  56019=>"00000000",
  56020=>"11111101",
  56021=>"11111111",
  56022=>"11111110",
  56023=>"00000100",
  56024=>"00000011",
  56025=>"00000000",
  56026=>"00000001",
  56027=>"00000010",
  56028=>"00000010",
  56029=>"00000000",
  56030=>"00000011",
  56031=>"11111110",
  56032=>"00000001",
  56033=>"00000000",
  56034=>"00000100",
  56035=>"11111111",
  56036=>"11111100",
  56037=>"00000001",
  56038=>"00000000",
  56039=>"11111101",
  56040=>"00000100",
  56041=>"00000010",
  56042=>"00000001",
  56043=>"11111101",
  56044=>"00000010",
  56045=>"11111111",
  56046=>"11111101",
  56047=>"11111111",
  56048=>"11111101",
  56049=>"00000010",
  56050=>"11111101",
  56051=>"11111111",
  56052=>"11111110",
  56053=>"11111110",
  56054=>"11111111",
  56055=>"00000001",
  56056=>"11111111",
  56057=>"00000001",
  56058=>"00000010",
  56059=>"00000000",
  56060=>"00000000",
  56061=>"00000011",
  56062=>"00000011",
  56063=>"11111101",
  56064=>"11111101",
  56065=>"00000010",
  56066=>"00000000",
  56067=>"11111110",
  56068=>"11111111",
  56069=>"11111101",
  56070=>"00000000",
  56071=>"11111111",
  56072=>"00000001",
  56073=>"11111110",
  56074=>"00000000",
  56075=>"00000011",
  56076=>"00000001",
  56077=>"00000001",
  56078=>"11111101",
  56079=>"00000010",
  56080=>"00000000",
  56081=>"11111110",
  56082=>"11111100",
  56083=>"00000011",
  56084=>"11111111",
  56085=>"00000000",
  56086=>"00000010",
  56087=>"11111101",
  56088=>"00000001",
  56089=>"00000000",
  56090=>"11111111",
  56091=>"00000001",
  56092=>"11111110",
  56093=>"00000011",
  56094=>"00000010",
  56095=>"00000000",
  56096=>"11111110",
  56097=>"11111111",
  56098=>"00000100",
  56099=>"00000001",
  56100=>"11111111",
  56101=>"00000000",
  56102=>"11111101",
  56103=>"11111110",
  56104=>"00000010",
  56105=>"00000011",
  56106=>"00000010",
  56107=>"11111111",
  56108=>"11111111",
  56109=>"00000010",
  56110=>"11111101",
  56111=>"00000010",
  56112=>"00000001",
  56113=>"11111101",
  56114=>"00000011",
  56115=>"11111111",
  56116=>"11111111",
  56117=>"00000000",
  56118=>"00000010",
  56119=>"00000000",
  56120=>"11111101",
  56121=>"11111111",
  56122=>"11111111",
  56123=>"11111101",
  56124=>"00000011",
  56125=>"11111110",
  56126=>"11111101",
  56127=>"11111110",
  56128=>"00000011",
  56129=>"00000011",
  56130=>"00000011",
  56131=>"00000101",
  56132=>"00000000",
  56133=>"00000010",
  56134=>"11111101",
  56135=>"11111110",
  56136=>"11111101",
  56137=>"00000011",
  56138=>"00000000",
  56139=>"00000011",
  56140=>"00000001",
  56141=>"00000000",
  56142=>"00000000",
  56143=>"11111100",
  56144=>"00000010",
  56145=>"00000000",
  56146=>"00000010",
  56147=>"11111100",
  56148=>"00000011",
  56149=>"00000001",
  56150=>"00000001",
  56151=>"11111101",
  56152=>"00000101",
  56153=>"11111101",
  56154=>"11111111",
  56155=>"00000101",
  56156=>"11111111",
  56157=>"11111110",
  56158=>"11111101",
  56159=>"00000001",
  56160=>"11111111",
  56161=>"11111101",
  56162=>"00000000",
  56163=>"00000011",
  56164=>"11111100",
  56165=>"00000010",
  56166=>"00000000",
  56167=>"11111111",
  56168=>"00000001",
  56169=>"00000100",
  56170=>"00000000",
  56171=>"00000100",
  56172=>"00000010",
  56173=>"11111100",
  56174=>"00000111",
  56175=>"11111110",
  56176=>"00000011",
  56177=>"00000001",
  56178=>"11111111",
  56179=>"11111110",
  56180=>"11111111",
  56181=>"11111101",
  56182=>"11111111",
  56183=>"11111111",
  56184=>"11111101",
  56185=>"00000001",
  56186=>"11111110",
  56187=>"00000000",
  56188=>"00000001",
  56189=>"11111110",
  56190=>"11111101",
  56191=>"00000000",
  56192=>"11111111",
  56193=>"00000010",
  56194=>"00000011",
  56195=>"11111110",
  56196=>"00000000",
  56197=>"00000011",
  56198=>"00000011",
  56199=>"11111110",
  56200=>"00000001",
  56201=>"11111110",
  56202=>"11111110",
  56203=>"11111111",
  56204=>"11111110",
  56205=>"11111110",
  56206=>"00000010",
  56207=>"00000001",
  56208=>"00000011",
  56209=>"11111101",
  56210=>"00000101",
  56211=>"11111111",
  56212=>"11111110",
  56213=>"11111110",
  56214=>"00000000",
  56215=>"00000000",
  56216=>"11111110",
  56217=>"00000000",
  56218=>"00000001",
  56219=>"00000000",
  56220=>"00000100",
  56221=>"00000010",
  56222=>"11111101",
  56223=>"11111110",
  56224=>"11111111",
  56225=>"00000001",
  56226=>"00000000",
  56227=>"00000001",
  56228=>"00000001",
  56229=>"00000000",
  56230=>"00000100",
  56231=>"11111111",
  56232=>"00000000",
  56233=>"11111110",
  56234=>"00000010",
  56235=>"00000001",
  56236=>"11111101",
  56237=>"00000001",
  56238=>"11111110",
  56239=>"11111110",
  56240=>"00000001",
  56241=>"11111111",
  56242=>"00000010",
  56243=>"11111101",
  56244=>"00000010",
  56245=>"11111110",
  56246=>"00000000",
  56247=>"00000001",
  56248=>"00000010",
  56249=>"11111101",
  56250=>"00000000",
  56251=>"00000010",
  56252=>"11111110",
  56253=>"00000000",
  56254=>"11111101",
  56255=>"00000100",
  56256=>"00000000",
  56257=>"00000001",
  56258=>"11111111",
  56259=>"00000100",
  56260=>"11111110",
  56261=>"11111110",
  56262=>"00000000",
  56263=>"00000001",
  56264=>"11111110",
  56265=>"11111111",
  56266=>"00000001",
  56267=>"11111111",
  56268=>"11111101",
  56269=>"00000001",
  56270=>"00000010",
  56271=>"00000011",
  56272=>"11111110",
  56273=>"00000000",
  56274=>"00000011",
  56275=>"00000100",
  56276=>"00000000",
  56277=>"11111110",
  56278=>"00000100",
  56279=>"11111100",
  56280=>"00000000",
  56281=>"11111111",
  56282=>"00000011",
  56283=>"00000000",
  56284=>"00000001",
  56285=>"11111101",
  56286=>"00000000",
  56287=>"00000010",
  56288=>"00000000",
  56289=>"00000010",
  56290=>"11111111",
  56291=>"00000010",
  56292=>"11111110",
  56293=>"00000000",
  56294=>"00000010",
  56295=>"00000000",
  56296=>"11111110",
  56297=>"11111110",
  56298=>"11111110",
  56299=>"11111100",
  56300=>"00000011",
  56301=>"00000011",
  56302=>"11111100",
  56303=>"11111101",
  56304=>"11111111",
  56305=>"00000011",
  56306=>"11111101",
  56307=>"00000010",
  56308=>"11111110",
  56309=>"11111100",
  56310=>"11111101",
  56311=>"00000001",
  56312=>"00000000",
  56313=>"00000010",
  56314=>"11111101",
  56315=>"11111111",
  56316=>"00000010",
  56317=>"00001000",
  56318=>"00000001",
  56319=>"00000001",
  56320=>"00000001",
  56321=>"00000010",
  56322=>"11111111",
  56323=>"11111101",
  56324=>"11111111",
  56325=>"11111101",
  56326=>"00000000",
  56327=>"00000001",
  56328=>"11111111",
  56329=>"00000001",
  56330=>"00000011",
  56331=>"11111110",
  56332=>"00000000",
  56333=>"11111100",
  56334=>"11111110",
  56335=>"11111101",
  56336=>"00000101",
  56337=>"00000001",
  56338=>"00000110",
  56339=>"11111101",
  56340=>"11111110",
  56341=>"00000010",
  56342=>"00000010",
  56343=>"11111101",
  56344=>"00000010",
  56345=>"11111100",
  56346=>"11111111",
  56347=>"00000010",
  56348=>"11111101",
  56349=>"11111110",
  56350=>"00000011",
  56351=>"11111100",
  56352=>"11111101",
  56353=>"11111101",
  56354=>"11111101",
  56355=>"00000001",
  56356=>"11111110",
  56357=>"00000100",
  56358=>"00000000",
  56359=>"11111110",
  56360=>"11111110",
  56361=>"00000000",
  56362=>"00000000",
  56363=>"11111101",
  56364=>"00000001",
  56365=>"00000001",
  56366=>"11111110",
  56367=>"00000000",
  56368=>"11111111",
  56369=>"11111100",
  56370=>"00000010",
  56371=>"00000001",
  56372=>"00000011",
  56373=>"11111111",
  56374=>"00000001",
  56375=>"00000010",
  56376=>"11111111",
  56377=>"11111111",
  56378=>"00000010",
  56379=>"11111111",
  56380=>"11111111",
  56381=>"11111110",
  56382=>"00000000",
  56383=>"11111111",
  56384=>"11111101",
  56385=>"00000000",
  56386=>"11111110",
  56387=>"11111111",
  56388=>"11111111",
  56389=>"11111100",
  56390=>"00000011",
  56391=>"00000000",
  56392=>"00000000",
  56393=>"11111101",
  56394=>"00000001",
  56395=>"11111110",
  56396=>"11111100",
  56397=>"00000001",
  56398=>"00000000",
  56399=>"11111110",
  56400=>"11111101",
  56401=>"11111111",
  56402=>"00000011",
  56403=>"00000101",
  56404=>"00000001",
  56405=>"00000010",
  56406=>"00000000",
  56407=>"11111110",
  56408=>"00000010",
  56409=>"00000010",
  56410=>"00000001",
  56411=>"11111111",
  56412=>"00000011",
  56413=>"11111111",
  56414=>"00000011",
  56415=>"00000001",
  56416=>"11111101",
  56417=>"11111110",
  56418=>"11111111",
  56419=>"11111111",
  56420=>"11111111",
  56421=>"11111101",
  56422=>"11111101",
  56423=>"00000010",
  56424=>"11111110",
  56425=>"00000010",
  56426=>"11111101",
  56427=>"11111111",
  56428=>"00000100",
  56429=>"00000100",
  56430=>"11111111",
  56431=>"00000001",
  56432=>"11111111",
  56433=>"11111111",
  56434=>"00000000",
  56435=>"11111100",
  56436=>"11111110",
  56437=>"00000000",
  56438=>"11111110",
  56439=>"11111110",
  56440=>"11111100",
  56441=>"11111101",
  56442=>"11111111",
  56443=>"00000001",
  56444=>"11111110",
  56445=>"00000000",
  56446=>"00000000",
  56447=>"11111110",
  56448=>"00000000",
  56449=>"11111100",
  56450=>"00000011",
  56451=>"11111110",
  56452=>"11111101",
  56453=>"00000001",
  56454=>"11111110",
  56455=>"11111101",
  56456=>"00000010",
  56457=>"11111110",
  56458=>"00000010",
  56459=>"00000001",
  56460=>"11111110",
  56461=>"00000000",
  56462=>"11111101",
  56463=>"00000000",
  56464=>"00000100",
  56465=>"00000100",
  56466=>"00000001",
  56467=>"11111101",
  56468=>"00000001",
  56469=>"00000100",
  56470=>"11111101",
  56471=>"00000100",
  56472=>"00000101",
  56473=>"00000000",
  56474=>"11111101",
  56475=>"11111111",
  56476=>"11111110",
  56477=>"00000010",
  56478=>"00000010",
  56479=>"00000000",
  56480=>"00000011",
  56481=>"00000000",
  56482=>"11111101",
  56483=>"00000011",
  56484=>"00000000",
  56485=>"11111110",
  56486=>"00000001",
  56487=>"11111101",
  56488=>"00000000",
  56489=>"11111110",
  56490=>"00000010",
  56491=>"11111110",
  56492=>"00000000",
  56493=>"11111101",
  56494=>"00000000",
  56495=>"11111110",
  56496=>"00000011",
  56497=>"11111110",
  56498=>"11111110",
  56499=>"11111111",
  56500=>"00000001",
  56501=>"00000001",
  56502=>"00000101",
  56503=>"00000000",
  56504=>"11111101",
  56505=>"11111110",
  56506=>"00000000",
  56507=>"00000010",
  56508=>"11111101",
  56509=>"00000000",
  56510=>"00000000",
  56511=>"00000011",
  56512=>"11111110",
  56513=>"00000000",
  56514=>"00000010",
  56515=>"00000001",
  56516=>"00000010",
  56517=>"11111101",
  56518=>"11111111",
  56519=>"00000000",
  56520=>"11111111",
  56521=>"00000101",
  56522=>"00000001",
  56523=>"11111100",
  56524=>"00000101",
  56525=>"00000000",
  56526=>"11111111",
  56527=>"00000011",
  56528=>"00000100",
  56529=>"00000000",
  56530=>"11111111",
  56531=>"11111111",
  56532=>"11111110",
  56533=>"11111111",
  56534=>"00000100",
  56535=>"00000000",
  56536=>"11111111",
  56537=>"11111111",
  56538=>"00000000",
  56539=>"00000000",
  56540=>"00000011",
  56541=>"11111100",
  56542=>"11111111",
  56543=>"11111101",
  56544=>"00000001",
  56545=>"11111110",
  56546=>"11111100",
  56547=>"00000000",
  56548=>"11111111",
  56549=>"11111101",
  56550=>"00000000",
  56551=>"11111101",
  56552=>"11111110",
  56553=>"11111101",
  56554=>"11111110",
  56555=>"11111101",
  56556=>"00000001",
  56557=>"11111111",
  56558=>"00000100",
  56559=>"00000000",
  56560=>"11111100",
  56561=>"11111101",
  56562=>"00000011",
  56563=>"11111111",
  56564=>"11111111",
  56565=>"11111111",
  56566=>"00000001",
  56567=>"00000100",
  56568=>"00000110",
  56569=>"11111111",
  56570=>"11111110",
  56571=>"00000001",
  56572=>"00000000",
  56573=>"00000010",
  56574=>"11111100",
  56575=>"11111111",
  56576=>"11111101",
  56577=>"11111101",
  56578=>"00000100",
  56579=>"00000000",
  56580=>"11111111",
  56581=>"11111111",
  56582=>"00000001",
  56583=>"11111111",
  56584=>"00000000",
  56585=>"00000101",
  56586=>"00000000",
  56587=>"11111111",
  56588=>"11111110",
  56589=>"11111111",
  56590=>"00000010",
  56591=>"11111111",
  56592=>"11111111",
  56593=>"00000010",
  56594=>"00000010",
  56595=>"11111111",
  56596=>"11111111",
  56597=>"00000001",
  56598=>"11111110",
  56599=>"11111111",
  56600=>"00000010",
  56601=>"00000000",
  56602=>"11111111",
  56603=>"00000000",
  56604=>"11111111",
  56605=>"11111110",
  56606=>"00000001",
  56607=>"11111111",
  56608=>"11111111",
  56609=>"00000001",
  56610=>"11111101",
  56611=>"00000010",
  56612=>"11111110",
  56613=>"00000011",
  56614=>"11111101",
  56615=>"00000001",
  56616=>"00000010",
  56617=>"00000001",
  56618=>"11111101",
  56619=>"00000010",
  56620=>"00000011",
  56621=>"11111101",
  56622=>"11111101",
  56623=>"00000000",
  56624=>"00000011",
  56625=>"11111101",
  56626=>"00000000",
  56627=>"11111111",
  56628=>"00000001",
  56629=>"00000101",
  56630=>"00000001",
  56631=>"00000010",
  56632=>"00000000",
  56633=>"11111101",
  56634=>"11111110",
  56635=>"00000011",
  56636=>"00000000",
  56637=>"11111110",
  56638=>"11111111",
  56639=>"11111101",
  56640=>"00000010",
  56641=>"11111110",
  56642=>"00000010",
  56643=>"11111101",
  56644=>"11111101",
  56645=>"00000001",
  56646=>"00000100",
  56647=>"00000000",
  56648=>"11111110",
  56649=>"11111110",
  56650=>"11111110",
  56651=>"11111111",
  56652=>"11111101",
  56653=>"00000000",
  56654=>"00000011",
  56655=>"11111100",
  56656=>"00000010",
  56657=>"00000010",
  56658=>"00000001",
  56659=>"11111111",
  56660=>"00000001",
  56661=>"11111111",
  56662=>"11111110",
  56663=>"11111101",
  56664=>"00000001",
  56665=>"00000000",
  56666=>"00000100",
  56667=>"11111110",
  56668=>"00000000",
  56669=>"11111110",
  56670=>"11111110",
  56671=>"11111111",
  56672=>"00000000",
  56673=>"00000110",
  56674=>"00000000",
  56675=>"00000000",
  56676=>"00000001",
  56677=>"11111111",
  56678=>"11111101",
  56679=>"11111111",
  56680=>"11111111",
  56681=>"00000000",
  56682=>"00000001",
  56683=>"00000000",
  56684=>"11111100",
  56685=>"00000000",
  56686=>"00000000",
  56687=>"11111100",
  56688=>"11111111",
  56689=>"11111110",
  56690=>"00000001",
  56691=>"00000010",
  56692=>"11111111",
  56693=>"00000011",
  56694=>"11111101",
  56695=>"11111101",
  56696=>"11111110",
  56697=>"11111110",
  56698=>"11111110",
  56699=>"00000011",
  56700=>"00000000",
  56701=>"00000100",
  56702=>"11111110",
  56703=>"00000011",
  56704=>"00000010",
  56705=>"00000010",
  56706=>"00000000",
  56707=>"11111111",
  56708=>"11111110",
  56709=>"00000010",
  56710=>"00000010",
  56711=>"00000000",
  56712=>"00000000",
  56713=>"11111111",
  56714=>"11111110",
  56715=>"11111111",
  56716=>"00000001",
  56717=>"00000010",
  56718=>"11111111",
  56719=>"11111111",
  56720=>"11111110",
  56721=>"00000011",
  56722=>"11111110",
  56723=>"00000011",
  56724=>"00000000",
  56725=>"00000000",
  56726=>"00000010",
  56727=>"00000010",
  56728=>"11111110",
  56729=>"11111111",
  56730=>"00000001",
  56731=>"00000001",
  56732=>"00000010",
  56733=>"00000011",
  56734=>"00000001",
  56735=>"00000000",
  56736=>"00000010",
  56737=>"11111110",
  56738=>"00000001",
  56739=>"00000011",
  56740=>"00000010",
  56741=>"00000010",
  56742=>"11111111",
  56743=>"00000011",
  56744=>"00000011",
  56745=>"00000010",
  56746=>"11111111",
  56747=>"00000001",
  56748=>"00000001",
  56749=>"00000001",
  56750=>"00000010",
  56751=>"00000001",
  56752=>"00000011",
  56753=>"11111100",
  56754=>"00000000",
  56755=>"11111111",
  56756=>"11111101",
  56757=>"11111110",
  56758=>"11111111",
  56759=>"11111111",
  56760=>"00000001",
  56761=>"11111110",
  56762=>"11111111",
  56763=>"11111111",
  56764=>"11111110",
  56765=>"00000001",
  56766=>"00000010",
  56767=>"00000001",
  56768=>"11111101",
  56769=>"00000001",
  56770=>"11111111",
  56771=>"00000100",
  56772=>"11111110",
  56773=>"11111101",
  56774=>"00000001",
  56775=>"11111101",
  56776=>"00000100",
  56777=>"11111101",
  56778=>"00000010",
  56779=>"00000000",
  56780=>"00000010",
  56781=>"00000001",
  56782=>"11111111",
  56783=>"00000000",
  56784=>"00000000",
  56785=>"00000001",
  56786=>"00000101",
  56787=>"00000101",
  56788=>"11111110",
  56789=>"11111111",
  56790=>"00000000",
  56791=>"00000010",
  56792=>"00000001",
  56793=>"00000010",
  56794=>"11111111",
  56795=>"00000011",
  56796=>"00000000",
  56797=>"11111110",
  56798=>"00000000",
  56799=>"00000010",
  56800=>"00000011",
  56801=>"00000010",
  56802=>"11111111",
  56803=>"11111111",
  56804=>"00000011",
  56805=>"11111111",
  56806=>"11111111",
  56807=>"00000001",
  56808=>"11111110",
  56809=>"11111101",
  56810=>"00000000",
  56811=>"11111101",
  56812=>"00000001",
  56813=>"00000010",
  56814=>"00000001",
  56815=>"11111111",
  56816=>"00000001",
  56817=>"00000011",
  56818=>"11111110",
  56819=>"00000001",
  56820=>"11111101",
  56821=>"00000001",
  56822=>"00000001",
  56823=>"00000001",
  56824=>"00000000",
  56825=>"00000001",
  56826=>"11111110",
  56827=>"11111111",
  56828=>"11111101",
  56829=>"00000001",
  56830=>"00000001",
  56831=>"11111101",
  56832=>"00000001",
  56833=>"11111101",
  56834=>"00000001",
  56835=>"00000010",
  56836=>"11111110",
  56837=>"00000001",
  56838=>"00000000",
  56839=>"00000000",
  56840=>"00000000",
  56841=>"00000001",
  56842=>"00000001",
  56843=>"00000001",
  56844=>"00000011",
  56845=>"11111110",
  56846=>"00000101",
  56847=>"11111100",
  56848=>"00000100",
  56849=>"11111110",
  56850=>"00000011",
  56851=>"00000100",
  56852=>"00000011",
  56853=>"00000000",
  56854=>"00000000",
  56855=>"00000000",
  56856=>"00000010",
  56857=>"00000011",
  56858=>"00000000",
  56859=>"00000001",
  56860=>"00000001",
  56861=>"11111111",
  56862=>"00000000",
  56863=>"00000000",
  56864=>"11111111",
  56865=>"11111110",
  56866=>"11111111",
  56867=>"00000010",
  56868=>"00000010",
  56869=>"11111101",
  56870=>"11111111",
  56871=>"00000100",
  56872=>"00000001",
  56873=>"00000110",
  56874=>"11111111",
  56875=>"00000010",
  56876=>"11111101",
  56877=>"11111111",
  56878=>"00000000",
  56879=>"11111111",
  56880=>"00000000",
  56881=>"00000000",
  56882=>"11111101",
  56883=>"00000001",
  56884=>"11111101",
  56885=>"00000000",
  56886=>"11111111",
  56887=>"00000001",
  56888=>"11111111",
  56889=>"00000001",
  56890=>"11111101",
  56891=>"11111111",
  56892=>"11111110",
  56893=>"00000111",
  56894=>"00000001",
  56895=>"00000010",
  56896=>"11111110",
  56897=>"11111110",
  56898=>"11111101",
  56899=>"11111100",
  56900=>"11111110",
  56901=>"00000000",
  56902=>"00000010",
  56903=>"11111101",
  56904=>"11111111",
  56905=>"11111111",
  56906=>"00000001",
  56907=>"00000100",
  56908=>"00000001",
  56909=>"11111111",
  56910=>"00000011",
  56911=>"00000001",
  56912=>"00000011",
  56913=>"00000100",
  56914=>"11111111",
  56915=>"11111101",
  56916=>"11111111",
  56917=>"00000010",
  56918=>"00000010",
  56919=>"00000101",
  56920=>"11111111",
  56921=>"00000011",
  56922=>"11111101",
  56923=>"11111111",
  56924=>"00000000",
  56925=>"00000010",
  56926=>"11111101",
  56927=>"00000001",
  56928=>"11111110",
  56929=>"11111110",
  56930=>"00000000",
  56931=>"00000011",
  56932=>"00000001",
  56933=>"00000010",
  56934=>"00000010",
  56935=>"11111100",
  56936=>"11111110",
  56937=>"11111111",
  56938=>"00000001",
  56939=>"11111110",
  56940=>"00000011",
  56941=>"00000000",
  56942=>"11111100",
  56943=>"00000011",
  56944=>"11111110",
  56945=>"00000001",
  56946=>"00000011",
  56947=>"00000000",
  56948=>"11111111",
  56949=>"00000000",
  56950=>"00000010",
  56951=>"00000001",
  56952=>"11111110",
  56953=>"00000000",
  56954=>"11111110",
  56955=>"00000011",
  56956=>"00000000",
  56957=>"11111111",
  56958=>"00000101",
  56959=>"00000001",
  56960=>"11111110",
  56961=>"00000001",
  56962=>"11111101",
  56963=>"11111011",
  56964=>"00000001",
  56965=>"00000001",
  56966=>"11111101",
  56967=>"00000001",
  56968=>"11111110",
  56969=>"00000001",
  56970=>"11111110",
  56971=>"11111101",
  56972=>"11111111",
  56973=>"11111101",
  56974=>"11111101",
  56975=>"00000001",
  56976=>"00000000",
  56977=>"11111100",
  56978=>"00000000",
  56979=>"00000001",
  56980=>"00000001",
  56981=>"11111100",
  56982=>"00000010",
  56983=>"00000100",
  56984=>"00000101",
  56985=>"00000101",
  56986=>"00000001",
  56987=>"11111110",
  56988=>"11111011",
  56989=>"00000000",
  56990=>"00000011",
  56991=>"00000011",
  56992=>"11111110",
  56993=>"11111111",
  56994=>"00000011",
  56995=>"00000010",
  56996=>"11111101",
  56997=>"00000001",
  56998=>"11111111",
  56999=>"00000001",
  57000=>"00000000",
  57001=>"00000010",
  57002=>"00000101",
  57003=>"00000011",
  57004=>"00000001",
  57005=>"00000010",
  57006=>"00000000",
  57007=>"00000000",
  57008=>"00000001",
  57009=>"11111101",
  57010=>"11111111",
  57011=>"11111111",
  57012=>"11111110",
  57013=>"11111100",
  57014=>"00000000",
  57015=>"00000000",
  57016=>"00000010",
  57017=>"11111111",
  57018=>"11111101",
  57019=>"11111110",
  57020=>"00000011",
  57021=>"11111100",
  57022=>"00000001",
  57023=>"11111111",
  57024=>"11111110",
  57025=>"11111111",
  57026=>"11111101",
  57027=>"11111111",
  57028=>"11111110",
  57029=>"11111111",
  57030=>"00000001",
  57031=>"00000011",
  57032=>"11111101",
  57033=>"00000001",
  57034=>"00000001",
  57035=>"11111100",
  57036=>"00000101",
  57037=>"11111111",
  57038=>"00000000",
  57039=>"11111111",
  57040=>"00000000",
  57041=>"11111101",
  57042=>"00000011",
  57043=>"00000000",
  57044=>"11111110",
  57045=>"11111110",
  57046=>"00000000",
  57047=>"00001001",
  57048=>"00000001",
  57049=>"11111111",
  57050=>"11111110",
  57051=>"00000000",
  57052=>"00000001",
  57053=>"00000010",
  57054=>"00000001",
  57055=>"00000010",
  57056=>"11111110",
  57057=>"00000010",
  57058=>"11111110",
  57059=>"00000000",
  57060=>"00000000",
  57061=>"11111101",
  57062=>"00000000",
  57063=>"00000110",
  57064=>"00000010",
  57065=>"11111111",
  57066=>"00000011",
  57067=>"11111110",
  57068=>"00000010",
  57069=>"11111110",
  57070=>"00000001",
  57071=>"00000011",
  57072=>"11111111",
  57073=>"11111111",
  57074=>"11111110",
  57075=>"00000000",
  57076=>"00000001",
  57077=>"00000010",
  57078=>"00000000",
  57079=>"11111110",
  57080=>"11111100",
  57081=>"00000001",
  57082=>"00000010",
  57083=>"00000010",
  57084=>"00000000",
  57085=>"00000000",
  57086=>"00000000",
  57087=>"00000001",
  57088=>"00000001",
  57089=>"00000010",
  57090=>"00000000",
  57091=>"00000011",
  57092=>"00000001",
  57093=>"11111110",
  57094=>"00000000",
  57095=>"11111110",
  57096=>"11111111",
  57097=>"11111111",
  57098=>"00000000",
  57099=>"11111111",
  57100=>"00000010",
  57101=>"00000100",
  57102=>"00000101",
  57103=>"11111110",
  57104=>"11111100",
  57105=>"11111101",
  57106=>"00000001",
  57107=>"00000000",
  57108=>"00000101",
  57109=>"11111110",
  57110=>"00000010",
  57111=>"11111110",
  57112=>"00000001",
  57113=>"00000100",
  57114=>"00000100",
  57115=>"11111101",
  57116=>"00000000",
  57117=>"11111111",
  57118=>"11111100",
  57119=>"00000010",
  57120=>"11111110",
  57121=>"00000001",
  57122=>"00000001",
  57123=>"11111101",
  57124=>"00000001",
  57125=>"11111111",
  57126=>"00000000",
  57127=>"11111110",
  57128=>"00000001",
  57129=>"00000010",
  57130=>"00000010",
  57131=>"11111111",
  57132=>"11111111",
  57133=>"00000000",
  57134=>"00000001",
  57135=>"00000001",
  57136=>"00000010",
  57137=>"11111111",
  57138=>"11111110",
  57139=>"00000000",
  57140=>"00000000",
  57141=>"00000000",
  57142=>"00000000",
  57143=>"11111100",
  57144=>"11111101",
  57145=>"00000000",
  57146=>"00000001",
  57147=>"00000011",
  57148=>"11111101",
  57149=>"00000000",
  57150=>"00000000",
  57151=>"11111110",
  57152=>"11111111",
  57153=>"11111101",
  57154=>"11111110",
  57155=>"11111110",
  57156=>"00000000",
  57157=>"00000010",
  57158=>"11111111",
  57159=>"11111101",
  57160=>"11111111",
  57161=>"11111101",
  57162=>"00000000",
  57163=>"00000011",
  57164=>"00000000",
  57165=>"11111110",
  57166=>"00000001",
  57167=>"11111111",
  57168=>"00000000",
  57169=>"11111101",
  57170=>"11111101",
  57171=>"11111101",
  57172=>"00000001",
  57173=>"00000101",
  57174=>"00000000",
  57175=>"00000001",
  57176=>"00000001",
  57177=>"11111110",
  57178=>"00000010",
  57179=>"11111110",
  57180=>"11111100",
  57181=>"11111100",
  57182=>"00000000",
  57183=>"11111111",
  57184=>"11111110",
  57185=>"00000001",
  57186=>"00000000",
  57187=>"00000011",
  57188=>"00000000",
  57189=>"11111110",
  57190=>"00000010",
  57191=>"11111110",
  57192=>"11111110",
  57193=>"00000000",
  57194=>"11111101",
  57195=>"00000010",
  57196=>"00000001",
  57197=>"00000011",
  57198=>"11111101",
  57199=>"11111111",
  57200=>"00000010",
  57201=>"11111111",
  57202=>"00000001",
  57203=>"00000001",
  57204=>"00000100",
  57205=>"11111111",
  57206=>"11111111",
  57207=>"11111111",
  57208=>"11111110",
  57209=>"00000001",
  57210=>"00000010",
  57211=>"00000000",
  57212=>"00000001",
  57213=>"11111110",
  57214=>"11111100",
  57215=>"00000100",
  57216=>"11111101",
  57217=>"11111111",
  57218=>"00000000",
  57219=>"00000000",
  57220=>"00000010",
  57221=>"11111110",
  57222=>"00000000",
  57223=>"00000100",
  57224=>"00000011",
  57225=>"00000000",
  57226=>"00000010",
  57227=>"00000000",
  57228=>"00000000",
  57229=>"11111110",
  57230=>"11111101",
  57231=>"11111110",
  57232=>"11111111",
  57233=>"00000001",
  57234=>"11111111",
  57235=>"00000000",
  57236=>"11111101",
  57237=>"00000000",
  57238=>"00000000",
  57239=>"11111111",
  57240=>"00000011",
  57241=>"11111111",
  57242=>"11111101",
  57243=>"11111110",
  57244=>"11111111",
  57245=>"11111101",
  57246=>"11111110",
  57247=>"11111111",
  57248=>"00000010",
  57249=>"11111101",
  57250=>"11111011",
  57251=>"00000000",
  57252=>"00000000",
  57253=>"00000001",
  57254=>"11111110",
  57255=>"00000000",
  57256=>"11111111",
  57257=>"11111111",
  57258=>"11111111",
  57259=>"00000010",
  57260=>"11111111",
  57261=>"11111110",
  57262=>"00000011",
  57263=>"00000011",
  57264=>"11111101",
  57265=>"11111111",
  57266=>"11111110",
  57267=>"11111101",
  57268=>"00000000",
  57269=>"11111100",
  57270=>"00000001",
  57271=>"11111110",
  57272=>"11111111",
  57273=>"00000010",
  57274=>"11111111",
  57275=>"00000000",
  57276=>"00000010",
  57277=>"00000100",
  57278=>"11111101",
  57279=>"00000001",
  57280=>"00000000",
  57281=>"11111110",
  57282=>"11111111",
  57283=>"00000000",
  57284=>"00000010",
  57285=>"00000010",
  57286=>"00000110",
  57287=>"11111111",
  57288=>"11111101",
  57289=>"11111110",
  57290=>"11111110",
  57291=>"00000000",
  57292=>"00000000",
  57293=>"11111110",
  57294=>"11111111",
  57295=>"00000000",
  57296=>"00000001",
  57297=>"00000010",
  57298=>"11111100",
  57299=>"11111110",
  57300=>"00000010",
  57301=>"00000011",
  57302=>"11111110",
  57303=>"11111110",
  57304=>"00000001",
  57305=>"00000100",
  57306=>"00000001",
  57307=>"00000000",
  57308=>"11111111",
  57309=>"00000010",
  57310=>"11111111",
  57311=>"11111011",
  57312=>"11111110",
  57313=>"00000000",
  57314=>"00000000",
  57315=>"11111110",
  57316=>"11111111",
  57317=>"11111111",
  57318=>"11111111",
  57319=>"00000000",
  57320=>"00000001",
  57321=>"00000010",
  57322=>"00000000",
  57323=>"11111101",
  57324=>"00000100",
  57325=>"00000001",
  57326=>"11111101",
  57327=>"00000000",
  57328=>"00000011",
  57329=>"11111101",
  57330=>"00000100",
  57331=>"00000000",
  57332=>"00000010",
  57333=>"11111101",
  57334=>"00000100",
  57335=>"00000010",
  57336=>"11111111",
  57337=>"00000000",
  57338=>"11111110",
  57339=>"00000010",
  57340=>"00000000",
  57341=>"00000010",
  57342=>"11111101",
  57343=>"00000001",
  57344=>"11111111",
  57345=>"00000010",
  57346=>"11111110",
  57347=>"00000000",
  57348=>"00000110",
  57349=>"00000110",
  57350=>"11111110",
  57351=>"00000010",
  57352=>"00000000",
  57353=>"11111110",
  57354=>"11111101",
  57355=>"00000000",
  57356=>"11111101",
  57357=>"11111111",
  57358=>"11111101",
  57359=>"00000010",
  57360=>"11111110",
  57361=>"11111111",
  57362=>"00000000",
  57363=>"11111101",
  57364=>"11111110",
  57365=>"11111110",
  57366=>"00000000",
  57367=>"00000001",
  57368=>"00000011",
  57369=>"00000010",
  57370=>"00000001",
  57371=>"00000011",
  57372=>"00000000",
  57373=>"00000010",
  57374=>"00000001",
  57375=>"00000001",
  57376=>"11111110",
  57377=>"00000011",
  57378=>"00000000",
  57379=>"11111110",
  57380=>"00000000",
  57381=>"00000011",
  57382=>"00000100",
  57383=>"00000011",
  57384=>"11111010",
  57385=>"00000110",
  57386=>"11111110",
  57387=>"00000000",
  57388=>"11111100",
  57389=>"00000001",
  57390=>"11111101",
  57391=>"11111111",
  57392=>"00000001",
  57393=>"00000000",
  57394=>"00000000",
  57395=>"00000101",
  57396=>"00000001",
  57397=>"11111111",
  57398=>"00000001",
  57399=>"00000000",
  57400=>"11111101",
  57401=>"00000010",
  57402=>"11111110",
  57403=>"00000001",
  57404=>"11111110",
  57405=>"00000010",
  57406=>"00000000",
  57407=>"11111110",
  57408=>"00000001",
  57409=>"00000010",
  57410=>"00000100",
  57411=>"00000011",
  57412=>"11111111",
  57413=>"00000001",
  57414=>"00000100",
  57415=>"11111111",
  57416=>"00000000",
  57417=>"11111110",
  57418=>"00000000",
  57419=>"00000010",
  57420=>"00000011",
  57421=>"00000010",
  57422=>"11111110",
  57423=>"00000010",
  57424=>"11111111",
  57425=>"00000001",
  57426=>"00000001",
  57427=>"11111111",
  57428=>"00000001",
  57429=>"11111101",
  57430=>"00000100",
  57431=>"00000011",
  57432=>"00000001",
  57433=>"11111100",
  57434=>"00000000",
  57435=>"00000100",
  57436=>"11111101",
  57437=>"11111111",
  57438=>"11111110",
  57439=>"11111111",
  57440=>"11111111",
  57441=>"00000011",
  57442=>"00000000",
  57443=>"00000000",
  57444=>"00000000",
  57445=>"11111100",
  57446=>"11111110",
  57447=>"00000101",
  57448=>"11111101",
  57449=>"11111011",
  57450=>"00000101",
  57451=>"11111110",
  57452=>"00000011",
  57453=>"00000010",
  57454=>"00000010",
  57455=>"11111101",
  57456=>"11111110",
  57457=>"11111110",
  57458=>"11111110",
  57459=>"00000010",
  57460=>"00000001",
  57461=>"11111111",
  57462=>"00000010",
  57463=>"11111101",
  57464=>"11111111",
  57465=>"00000001",
  57466=>"11111110",
  57467=>"00000000",
  57468=>"00000001",
  57469=>"11111111",
  57470=>"00000010",
  57471=>"11111110",
  57472=>"00000101",
  57473=>"11111101",
  57474=>"00000001",
  57475=>"11111111",
  57476=>"11111110",
  57477=>"00000100",
  57478=>"11111111",
  57479=>"00000001",
  57480=>"00000011",
  57481=>"11111101",
  57482=>"00000001",
  57483=>"00000001",
  57484=>"00000010",
  57485=>"11111111",
  57486=>"11111101",
  57487=>"00000100",
  57488=>"11111110",
  57489=>"00000010",
  57490=>"00000010",
  57491=>"00000010",
  57492=>"00000100",
  57493=>"00000011",
  57494=>"11111110",
  57495=>"11111111",
  57496=>"00000000",
  57497=>"11111101",
  57498=>"00000011",
  57499=>"00000000",
  57500=>"11111111",
  57501=>"00000011",
  57502=>"00000000",
  57503=>"11111111",
  57504=>"11111110",
  57505=>"00000000",
  57506=>"00000010",
  57507=>"00000011",
  57508=>"11111110",
  57509=>"11111100",
  57510=>"11111110",
  57511=>"11111101",
  57512=>"11111110",
  57513=>"00000100",
  57514=>"00000010",
  57515=>"00000011",
  57516=>"11111111",
  57517=>"11111101",
  57518=>"00000100",
  57519=>"00000001",
  57520=>"00000001",
  57521=>"00000011",
  57522=>"11111101",
  57523=>"00000000",
  57524=>"00000001",
  57525=>"00000000",
  57526=>"11111100",
  57527=>"11111100",
  57528=>"00000010",
  57529=>"00000010",
  57530=>"00000000",
  57531=>"00000000",
  57532=>"00000011",
  57533=>"11111110",
  57534=>"11111110",
  57535=>"00000100",
  57536=>"00000000",
  57537=>"00000010",
  57538=>"11111110",
  57539=>"11111111",
  57540=>"11111110",
  57541=>"11111111",
  57542=>"00000001",
  57543=>"11111111",
  57544=>"11111101",
  57545=>"00000010",
  57546=>"11111111",
  57547=>"00000011",
  57548=>"00000011",
  57549=>"11111110",
  57550=>"11111111",
  57551=>"00000001",
  57552=>"00000100",
  57553=>"00000001",
  57554=>"11111110",
  57555=>"11111110",
  57556=>"00000010",
  57557=>"11111110",
  57558=>"00000001",
  57559=>"11111111",
  57560=>"11111101",
  57561=>"00000000",
  57562=>"11111110",
  57563=>"00000001",
  57564=>"11111111",
  57565=>"11111111",
  57566=>"11111110",
  57567=>"00000010",
  57568=>"11111110",
  57569=>"00000011",
  57570=>"11111110",
  57571=>"00000001",
  57572=>"11111110",
  57573=>"00000100",
  57574=>"00000001",
  57575=>"00000000",
  57576=>"00000010",
  57577=>"00000000",
  57578=>"11111110",
  57579=>"11111111",
  57580=>"11111110",
  57581=>"00000000",
  57582=>"00000010",
  57583=>"11111111",
  57584=>"00000001",
  57585=>"00000001",
  57586=>"00000100",
  57587=>"11111111",
  57588=>"11111110",
  57589=>"00000000",
  57590=>"00000011",
  57591=>"11111101",
  57592=>"11111111",
  57593=>"00000010",
  57594=>"00000010",
  57595=>"00000010",
  57596=>"11111111",
  57597=>"11111110",
  57598=>"00000010",
  57599=>"11111111",
  57600=>"11111111",
  57601=>"00000101",
  57602=>"11111100",
  57603=>"00000001",
  57604=>"00000001",
  57605=>"00000010",
  57606=>"11111100",
  57607=>"11111101",
  57608=>"11111110",
  57609=>"00000011",
  57610=>"11111110",
  57611=>"11111101",
  57612=>"00000000",
  57613=>"11111111",
  57614=>"00000000",
  57615=>"00000010",
  57616=>"11111110",
  57617=>"11111111",
  57618=>"11111110",
  57619=>"11111010",
  57620=>"00000000",
  57621=>"00000011",
  57622=>"11111111",
  57623=>"11111100",
  57624=>"00000001",
  57625=>"00000000",
  57626=>"00000011",
  57627=>"11111110",
  57628=>"11111111",
  57629=>"00000000",
  57630=>"00000101",
  57631=>"00000011",
  57632=>"11111110",
  57633=>"11111110",
  57634=>"11111111",
  57635=>"00000010",
  57636=>"00000100",
  57637=>"00000010",
  57638=>"11111111",
  57639=>"00000000",
  57640=>"11111111",
  57641=>"11111111",
  57642=>"11111110",
  57643=>"11111101",
  57644=>"00000010",
  57645=>"00000011",
  57646=>"00000100",
  57647=>"11111011",
  57648=>"11111101",
  57649=>"11111111",
  57650=>"11111111",
  57651=>"00000001",
  57652=>"11111111",
  57653=>"00000010",
  57654=>"00000001",
  57655=>"11111110",
  57656=>"00000001",
  57657=>"00000000",
  57658=>"11111111",
  57659=>"00000001",
  57660=>"00000010",
  57661=>"11111110",
  57662=>"11111111",
  57663=>"11111110",
  57664=>"11111111",
  57665=>"11111011",
  57666=>"11111101",
  57667=>"11111111",
  57668=>"00000010",
  57669=>"11111101",
  57670=>"11111011",
  57671=>"00000001",
  57672=>"00000001",
  57673=>"00000000",
  57674=>"11111111",
  57675=>"00000000",
  57676=>"00000010",
  57677=>"11111111",
  57678=>"00000010",
  57679=>"00000010",
  57680=>"00000010",
  57681=>"00000100",
  57682=>"11111111",
  57683=>"00000001",
  57684=>"00000000",
  57685=>"00000011",
  57686=>"00000001",
  57687=>"11111111",
  57688=>"11111110",
  57689=>"00000000",
  57690=>"00000101",
  57691=>"00000000",
  57692=>"00000010",
  57693=>"00000000",
  57694=>"00000001",
  57695=>"00000001",
  57696=>"00000010",
  57697=>"00000011",
  57698=>"11111110",
  57699=>"11111110",
  57700=>"00000000",
  57701=>"11111111",
  57702=>"00000100",
  57703=>"11111111",
  57704=>"11111110",
  57705=>"11111110",
  57706=>"11111101",
  57707=>"00000011",
  57708=>"00000001",
  57709=>"00000000",
  57710=>"11111111",
  57711=>"00000000",
  57712=>"11111111",
  57713=>"11111111",
  57714=>"00000000",
  57715=>"11111110",
  57716=>"11111110",
  57717=>"11111111",
  57718=>"00000001",
  57719=>"00000001",
  57720=>"11111111",
  57721=>"00000000",
  57722=>"00000110",
  57723=>"00000100",
  57724=>"00000010",
  57725=>"00000010",
  57726=>"00000001",
  57727=>"00000001",
  57728=>"11111100",
  57729=>"00000011",
  57730=>"00000011",
  57731=>"00000010",
  57732=>"11111101",
  57733=>"00000011",
  57734=>"00000000",
  57735=>"00000000",
  57736=>"11111110",
  57737=>"00000000",
  57738=>"00000001",
  57739=>"00000011",
  57740=>"11111110",
  57741=>"00000010",
  57742=>"00000000",
  57743=>"00000010",
  57744=>"11111111",
  57745=>"11111111",
  57746=>"11111111",
  57747=>"11111110",
  57748=>"00000100",
  57749=>"11111110",
  57750=>"11111101",
  57751=>"11111101",
  57752=>"00000011",
  57753=>"00000011",
  57754=>"00000011",
  57755=>"00000010",
  57756=>"00000000",
  57757=>"00000001",
  57758=>"11111111",
  57759=>"11111111",
  57760=>"00000001",
  57761=>"11111110",
  57762=>"00000001",
  57763=>"00000011",
  57764=>"00000011",
  57765=>"00000010",
  57766=>"00000010",
  57767=>"00000101",
  57768=>"11111111",
  57769=>"00000000",
  57770=>"00000100",
  57771=>"00000000",
  57772=>"00000001",
  57773=>"11111101",
  57774=>"00000010",
  57775=>"00000011",
  57776=>"00000011",
  57777=>"11111111",
  57778=>"11111110",
  57779=>"11111111",
  57780=>"00000000",
  57781=>"11111101",
  57782=>"11111111",
  57783=>"00000000",
  57784=>"11111010",
  57785=>"11111111",
  57786=>"00000100",
  57787=>"00000000",
  57788=>"00000001",
  57789=>"11111110",
  57790=>"11111101",
  57791=>"11111101",
  57792=>"11111110",
  57793=>"00000001",
  57794=>"00000011",
  57795=>"11111101",
  57796=>"11111110",
  57797=>"00000001",
  57798=>"11111101",
  57799=>"00000010",
  57800=>"00000100",
  57801=>"00000010",
  57802=>"00000010",
  57803=>"11111111",
  57804=>"00000001",
  57805=>"00000000",
  57806=>"11111110",
  57807=>"00000010",
  57808=>"11111101",
  57809=>"11111110",
  57810=>"00000101",
  57811=>"11111110",
  57812=>"00000010",
  57813=>"11111100",
  57814=>"00000011",
  57815=>"00000010",
  57816=>"11111101",
  57817=>"00000100",
  57818=>"11111111",
  57819=>"00000011",
  57820=>"00000001",
  57821=>"00000001",
  57822=>"00000011",
  57823=>"11111111",
  57824=>"11111011",
  57825=>"11111111",
  57826=>"00000001",
  57827=>"11111111",
  57828=>"00000001",
  57829=>"00000001",
  57830=>"11111110",
  57831=>"00000011",
  57832=>"11111110",
  57833=>"00000000",
  57834=>"11111101",
  57835=>"11111110",
  57836=>"11111011",
  57837=>"00000001",
  57838=>"11111111",
  57839=>"11111110",
  57840=>"00000010",
  57841=>"00000011",
  57842=>"11111101",
  57843=>"00000010",
  57844=>"11111110",
  57845=>"11111111",
  57846=>"00000010",
  57847=>"11111101",
  57848=>"00000011",
  57849=>"00000011",
  57850=>"00000100",
  57851=>"00000011",
  57852=>"00000001",
  57853=>"00000101",
  57854=>"11111100",
  57855=>"00000000",
  57856=>"11111111",
  57857=>"00000000",
  57858=>"00000000",
  57859=>"11111101",
  57860=>"00000001",
  57861=>"11111101",
  57862=>"00000111",
  57863=>"11111100",
  57864=>"11111100",
  57865=>"11111110",
  57866=>"00000000",
  57867=>"11111111",
  57868=>"00000010",
  57869=>"00000010",
  57870=>"11111100",
  57871=>"00000011",
  57872=>"11111111",
  57873=>"11111101",
  57874=>"11111110",
  57875=>"00000001",
  57876=>"00000001",
  57877=>"00000000",
  57878=>"11111111",
  57879=>"11111101",
  57880=>"00000010",
  57881=>"00000000",
  57882=>"00000001",
  57883=>"00000000",
  57884=>"00000000",
  57885=>"11111111",
  57886=>"00000010",
  57887=>"00000011",
  57888=>"00000011",
  57889=>"11111101",
  57890=>"11111101",
  57891=>"00000010",
  57892=>"11111110",
  57893=>"00000010",
  57894=>"00000000",
  57895=>"11111110",
  57896=>"11111101",
  57897=>"11111110",
  57898=>"00000001",
  57899=>"00000011",
  57900=>"00000101",
  57901=>"00000100",
  57902=>"11111100",
  57903=>"00000010",
  57904=>"00000011",
  57905=>"11111110",
  57906=>"11111110",
  57907=>"11111111",
  57908=>"11111101",
  57909=>"00000100",
  57910=>"00000010",
  57911=>"00000010",
  57912=>"00000100",
  57913=>"00000011",
  57914=>"11111110",
  57915=>"11111110",
  57916=>"11111110",
  57917=>"00000011",
  57918=>"11111101",
  57919=>"11111100",
  57920=>"00000100",
  57921=>"11111110",
  57922=>"00000011",
  57923=>"00000000",
  57924=>"11111100",
  57925=>"11111111",
  57926=>"11111101",
  57927=>"11111100",
  57928=>"00000001",
  57929=>"00000011",
  57930=>"00000101",
  57931=>"00000000",
  57932=>"00000001",
  57933=>"00000011",
  57934=>"11111101",
  57935=>"00000000",
  57936=>"00000000",
  57937=>"11111110",
  57938=>"00000000",
  57939=>"00000000",
  57940=>"00000001",
  57941=>"11111100",
  57942=>"11111110",
  57943=>"11111110",
  57944=>"00000100",
  57945=>"11111101",
  57946=>"00000001",
  57947=>"11111101",
  57948=>"11111110",
  57949=>"00000011",
  57950=>"11111011",
  57951=>"00000000",
  57952=>"00000011",
  57953=>"00000001",
  57954=>"00000000",
  57955=>"11111101",
  57956=>"11111110",
  57957=>"00000000",
  57958=>"11111101",
  57959=>"00000100",
  57960=>"00000000",
  57961=>"00000011",
  57962=>"00000000",
  57963=>"11111111",
  57964=>"00000100",
  57965=>"00000010",
  57966=>"11111110",
  57967=>"11111110",
  57968=>"00000001",
  57969=>"00000011",
  57970=>"00000010",
  57971=>"00000100",
  57972=>"00000000",
  57973=>"11111101",
  57974=>"11111111",
  57975=>"00000010",
  57976=>"11111110",
  57977=>"00000011",
  57978=>"00000010",
  57979=>"00000010",
  57980=>"00000010",
  57981=>"00000011",
  57982=>"00000011",
  57983=>"11111111",
  57984=>"00000010",
  57985=>"00000001",
  57986=>"00000000",
  57987=>"00000001",
  57988=>"11111101",
  57989=>"00000010",
  57990=>"00000001",
  57991=>"11111111",
  57992=>"00000001",
  57993=>"11111101",
  57994=>"11111111",
  57995=>"00000010",
  57996=>"11111101",
  57997=>"11111110",
  57998=>"00000110",
  57999=>"11111110",
  58000=>"00000100",
  58001=>"00000001",
  58002=>"00000010",
  58003=>"00000000",
  58004=>"00000011",
  58005=>"00000101",
  58006=>"11111101",
  58007=>"11111110",
  58008=>"00000000",
  58009=>"00000010",
  58010=>"00000100",
  58011=>"11111110",
  58012=>"00000100",
  58013=>"00000011",
  58014=>"00000000",
  58015=>"11111101",
  58016=>"00000010",
  58017=>"11111110",
  58018=>"11111101",
  58019=>"00000101",
  58020=>"00000100",
  58021=>"00000011",
  58022=>"11111111",
  58023=>"00000000",
  58024=>"00000010",
  58025=>"00000000",
  58026=>"11111101",
  58027=>"00000100",
  58028=>"00000001",
  58029=>"11111111",
  58030=>"11111111",
  58031=>"00000000",
  58032=>"00000010",
  58033=>"00000010",
  58034=>"00000100",
  58035=>"00000010",
  58036=>"11111111",
  58037=>"11111101",
  58038=>"11111111",
  58039=>"11111101",
  58040=>"00000011",
  58041=>"11111101",
  58042=>"11111110",
  58043=>"11111111",
  58044=>"00000110",
  58045=>"00000100",
  58046=>"00000000",
  58047=>"00000001",
  58048=>"00000011",
  58049=>"00000010",
  58050=>"00000000",
  58051=>"00000001",
  58052=>"00000000",
  58053=>"00000000",
  58054=>"11111111",
  58055=>"11111101",
  58056=>"00000000",
  58057=>"00000100",
  58058=>"11111111",
  58059=>"11111111",
  58060=>"00000010",
  58061=>"11111111",
  58062=>"00000001",
  58063=>"00000001",
  58064=>"11111111",
  58065=>"00000001",
  58066=>"11111111",
  58067=>"00000010",
  58068=>"11111110",
  58069=>"00000001",
  58070=>"00000001",
  58071=>"11111100",
  58072=>"00000000",
  58073=>"11111100",
  58074=>"00000010",
  58075=>"00000001",
  58076=>"00000010",
  58077=>"00000001",
  58078=>"00000011",
  58079=>"00000100",
  58080=>"00000001",
  58081=>"11111111",
  58082=>"11111110",
  58083=>"00000011",
  58084=>"11111101",
  58085=>"11111111",
  58086=>"11111100",
  58087=>"00000001",
  58088=>"00000011",
  58089=>"11111110",
  58090=>"00000010",
  58091=>"11111110",
  58092=>"00000010",
  58093=>"11111101",
  58094=>"11111111",
  58095=>"11111100",
  58096=>"00000100",
  58097=>"11111101",
  58098=>"00000100",
  58099=>"11111111",
  58100=>"00000001",
  58101=>"00000001",
  58102=>"00000011",
  58103=>"11111101",
  58104=>"00000111",
  58105=>"00000010",
  58106=>"00000000",
  58107=>"00000100",
  58108=>"00000000",
  58109=>"11111111",
  58110=>"11111110",
  58111=>"00000011",
  58112=>"00000011",
  58113=>"11111100",
  58114=>"00000000",
  58115=>"11111101",
  58116=>"11111101",
  58117=>"00000011",
  58118=>"00000000",
  58119=>"00000010",
  58120=>"11111101",
  58121=>"00000000",
  58122=>"11111101",
  58123=>"00000010",
  58124=>"00000001",
  58125=>"00000010",
  58126=>"00000101",
  58127=>"11111110",
  58128=>"00000101",
  58129=>"00000010",
  58130=>"00000011",
  58131=>"00000001",
  58132=>"00000001",
  58133=>"00000001",
  58134=>"00000001",
  58135=>"00000011",
  58136=>"11111101",
  58137=>"00000000",
  58138=>"11111111",
  58139=>"00000001",
  58140=>"00000011",
  58141=>"00000010",
  58142=>"00000001",
  58143=>"00000010",
  58144=>"00000001",
  58145=>"11111101",
  58146=>"00000001",
  58147=>"00000001",
  58148=>"00000001",
  58149=>"11111111",
  58150=>"11111110",
  58151=>"00000011",
  58152=>"00000011",
  58153=>"00000010",
  58154=>"00000010",
  58155=>"11111110",
  58156=>"11111111",
  58157=>"00000010",
  58158=>"00000000",
  58159=>"11111110",
  58160=>"00000100",
  58161=>"11111110",
  58162=>"00000000",
  58163=>"11111100",
  58164=>"00000000",
  58165=>"00000010",
  58166=>"00000001",
  58167=>"00000100",
  58168=>"00000101",
  58169=>"00000010",
  58170=>"11111111",
  58171=>"11111110",
  58172=>"00000000",
  58173=>"00000011",
  58174=>"11111111",
  58175=>"00000000",
  58176=>"11111111",
  58177=>"00001000",
  58178=>"00000001",
  58179=>"00000001",
  58180=>"00000000",
  58181=>"00000010",
  58182=>"00000000",
  58183=>"11111100",
  58184=>"11111011",
  58185=>"11111111",
  58186=>"11111111",
  58187=>"11111111",
  58188=>"00000010",
  58189=>"00000110",
  58190=>"00000010",
  58191=>"00000001",
  58192=>"00000010",
  58193=>"00000010",
  58194=>"00000010",
  58195=>"00000001",
  58196=>"00000000",
  58197=>"00000001",
  58198=>"11111101",
  58199=>"00000001",
  58200=>"00000000",
  58201=>"00000001",
  58202=>"00000101",
  58203=>"00000100",
  58204=>"00000000",
  58205=>"00000011",
  58206=>"11111111",
  58207=>"11111101",
  58208=>"00000100",
  58209=>"11111111",
  58210=>"00000001",
  58211=>"11111110",
  58212=>"00000010",
  58213=>"00000000",
  58214=>"00000000",
  58215=>"11111101",
  58216=>"00000000",
  58217=>"00000010",
  58218=>"00000001",
  58219=>"00000001",
  58220=>"00000001",
  58221=>"00000011",
  58222=>"11111100",
  58223=>"00000000",
  58224=>"00000001",
  58225=>"00000100",
  58226=>"11111110",
  58227=>"00000001",
  58228=>"11111110",
  58229=>"11111101",
  58230=>"00000000",
  58231=>"00000001",
  58232=>"00000101",
  58233=>"00000001",
  58234=>"00000000",
  58235=>"11111111",
  58236=>"11111111",
  58237=>"00000010",
  58238=>"00000000",
  58239=>"00000001",
  58240=>"11111101",
  58241=>"11111101",
  58242=>"00000011",
  58243=>"00000011",
  58244=>"00000001",
  58245=>"00000001",
  58246=>"11111101",
  58247=>"11111110",
  58248=>"11111111",
  58249=>"00000001",
  58250=>"11111101",
  58251=>"11111111",
  58252=>"11111101",
  58253=>"11111101",
  58254=>"11111011",
  58255=>"00000000",
  58256=>"00000011",
  58257=>"11111110",
  58258=>"11111111",
  58259=>"11111101",
  58260=>"00000000",
  58261=>"00000101",
  58262=>"00000000",
  58263=>"00000001",
  58264=>"00000000",
  58265=>"11111101",
  58266=>"00000100",
  58267=>"11111111",
  58268=>"00000001",
  58269=>"11111111",
  58270=>"00000001",
  58271=>"00000011",
  58272=>"00000010",
  58273=>"00000001",
  58274=>"00000100",
  58275=>"11111111",
  58276=>"00000011",
  58277=>"00000011",
  58278=>"00000001",
  58279=>"11111101",
  58280=>"00000010",
  58281=>"00000100",
  58282=>"00000001",
  58283=>"00000011",
  58284=>"00000010",
  58285=>"00000011",
  58286=>"11111111",
  58287=>"00000010",
  58288=>"00000000",
  58289=>"11111111",
  58290=>"00000101",
  58291=>"00000001",
  58292=>"00000000",
  58293=>"00000000",
  58294=>"11111110",
  58295=>"11111111",
  58296=>"00000001",
  58297=>"11111110",
  58298=>"11111111",
  58299=>"00000000",
  58300=>"11111111",
  58301=>"00000010",
  58302=>"00000001",
  58303=>"11111101",
  58304=>"11111101",
  58305=>"11111111",
  58306=>"00000011",
  58307=>"00000000",
  58308=>"11111111",
  58309=>"11111110",
  58310=>"00000000",
  58311=>"11111101",
  58312=>"11111101",
  58313=>"00000000",
  58314=>"00000100",
  58315=>"11111101",
  58316=>"11111101",
  58317=>"11111101",
  58318=>"11111110",
  58319=>"00000000",
  58320=>"11111111",
  58321=>"00000010",
  58322=>"00000100",
  58323=>"11111110",
  58324=>"00000001",
  58325=>"11111111",
  58326=>"11111101",
  58327=>"11111100",
  58328=>"11111110",
  58329=>"00000000",
  58330=>"00000001",
  58331=>"00000001",
  58332=>"11111100",
  58333=>"11111111",
  58334=>"00000001",
  58335=>"00000000",
  58336=>"00000101",
  58337=>"11111110",
  58338=>"00000001",
  58339=>"11111110",
  58340=>"00000000",
  58341=>"11111110",
  58342=>"11111110",
  58343=>"00000001",
  58344=>"11111111",
  58345=>"11111110",
  58346=>"00000001",
  58347=>"00000010",
  58348=>"11111110",
  58349=>"00000011",
  58350=>"00000010",
  58351=>"00000101",
  58352=>"00000011",
  58353=>"00000011",
  58354=>"11111101",
  58355=>"00000000",
  58356=>"11111110",
  58357=>"11111110",
  58358=>"00000001",
  58359=>"00000001",
  58360=>"00000000",
  58361=>"11111111",
  58362=>"11111111",
  58363=>"00000001",
  58364=>"00000111",
  58365=>"00000101",
  58366=>"00000010",
  58367=>"00000010",
  58368=>"11111101",
  58369=>"00000001",
  58370=>"00000101",
  58371=>"00000000",
  58372=>"00000011",
  58373=>"11111110",
  58374=>"11111110",
  58375=>"00000000",
  58376=>"11111110",
  58377=>"11111100",
  58378=>"11111110",
  58379=>"00000000",
  58380=>"00000011",
  58381=>"11111110",
  58382=>"00000000",
  58383=>"11111111",
  58384=>"00000011",
  58385=>"00000100",
  58386=>"00000011",
  58387=>"11111110",
  58388=>"00000110",
  58389=>"00000010",
  58390=>"00000000",
  58391=>"11111111",
  58392=>"00000010",
  58393=>"00000000",
  58394=>"00000010",
  58395=>"00000010",
  58396=>"11111111",
  58397=>"00000010",
  58398=>"00000000",
  58399=>"00000000",
  58400=>"11111111",
  58401=>"11111111",
  58402=>"11111101",
  58403=>"00000000",
  58404=>"00000010",
  58405=>"00000000",
  58406=>"00000010",
  58407=>"11111101",
  58408=>"11111110",
  58409=>"11111100",
  58410=>"00000010",
  58411=>"11111111",
  58412=>"11111101",
  58413=>"11111111",
  58414=>"00000001",
  58415=>"11111101",
  58416=>"11111111",
  58417=>"00000000",
  58418=>"11111110",
  58419=>"11111101",
  58420=>"11111101",
  58421=>"00000001",
  58422=>"00000000",
  58423=>"00000001",
  58424=>"11111111",
  58425=>"11111111",
  58426=>"00000000",
  58427=>"00000100",
  58428=>"11111101",
  58429=>"11111110",
  58430=>"11111110",
  58431=>"00000010",
  58432=>"00000001",
  58433=>"11111110",
  58434=>"11111110",
  58435=>"11111111",
  58436=>"11111111",
  58437=>"11111110",
  58438=>"00000000",
  58439=>"00000010",
  58440=>"11111110",
  58441=>"00000000",
  58442=>"00000001",
  58443=>"11111111",
  58444=>"11111101",
  58445=>"00000000",
  58446=>"11111111",
  58447=>"11111111",
  58448=>"00000011",
  58449=>"00000001",
  58450=>"11111111",
  58451=>"11111101",
  58452=>"11111110",
  58453=>"11111101",
  58454=>"00000010",
  58455=>"00000001",
  58456=>"00000000",
  58457=>"00000010",
  58458=>"11111111",
  58459=>"00000101",
  58460=>"00000010",
  58461=>"11111111",
  58462=>"00000011",
  58463=>"00000011",
  58464=>"00000010",
  58465=>"00000010",
  58466=>"00000011",
  58467=>"00000010",
  58468=>"11111110",
  58469=>"11111111",
  58470=>"11111111",
  58471=>"11111111",
  58472=>"11111110",
  58473=>"11111110",
  58474=>"00000001",
  58475=>"11111110",
  58476=>"00000010",
  58477=>"11111111",
  58478=>"11111110",
  58479=>"00000001",
  58480=>"00000011",
  58481=>"00000100",
  58482=>"00000010",
  58483=>"11111110",
  58484=>"00000011",
  58485=>"00000001",
  58486=>"00000001",
  58487=>"11111111",
  58488=>"11111110",
  58489=>"00000000",
  58490=>"11111111",
  58491=>"00000011",
  58492=>"00000001",
  58493=>"00000010",
  58494=>"11111111",
  58495=>"11111110",
  58496=>"00000100",
  58497=>"11111111",
  58498=>"11111110",
  58499=>"11111101",
  58500=>"00000001",
  58501=>"00000001",
  58502=>"00000000",
  58503=>"00000000",
  58504=>"11111110",
  58505=>"11111111",
  58506=>"00000010",
  58507=>"00000010",
  58508=>"00000011",
  58509=>"11111110",
  58510=>"11111111",
  58511=>"00000001",
  58512=>"11111110",
  58513=>"11111111",
  58514=>"11111110",
  58515=>"11111101",
  58516=>"00000011",
  58517=>"11111100",
  58518=>"00000001",
  58519=>"11111101",
  58520=>"11111111",
  58521=>"00000010",
  58522=>"00000011",
  58523=>"11111110",
  58524=>"00000010",
  58525=>"11111110",
  58526=>"00000001",
  58527=>"00000000",
  58528=>"00000001",
  58529=>"00000011",
  58530=>"00000100",
  58531=>"00000000",
  58532=>"00000001",
  58533=>"11111110",
  58534=>"00000000",
  58535=>"00000000",
  58536=>"00000011",
  58537=>"00000000",
  58538=>"00000000",
  58539=>"00000001",
  58540=>"00000010",
  58541=>"00000011",
  58542=>"11111111",
  58543=>"11111101",
  58544=>"11111110",
  58545=>"00000000",
  58546=>"00000000",
  58547=>"11111101",
  58548=>"00000000",
  58549=>"00000001",
  58550=>"11111101",
  58551=>"11111101",
  58552=>"11111110",
  58553=>"11111101",
  58554=>"11111110",
  58555=>"00000000",
  58556=>"11111111",
  58557=>"00000010",
  58558=>"00000011",
  58559=>"11111101",
  58560=>"00000000",
  58561=>"00000001",
  58562=>"00000100",
  58563=>"11111110",
  58564=>"00000010",
  58565=>"11111110",
  58566=>"00000001",
  58567=>"00000001",
  58568=>"00000000",
  58569=>"11111111",
  58570=>"00000000",
  58571=>"11111111",
  58572=>"00000000",
  58573=>"00000010",
  58574=>"00000000",
  58575=>"00000000",
  58576=>"11111111",
  58577=>"00000001",
  58578=>"00000000",
  58579=>"00000011",
  58580=>"11111111",
  58581=>"00000001",
  58582=>"11111100",
  58583=>"00000010",
  58584=>"00000000",
  58585=>"11111111",
  58586=>"11111111",
  58587=>"11111101",
  58588=>"11111101",
  58589=>"11111101",
  58590=>"11111101",
  58591=>"00000011",
  58592=>"00000010",
  58593=>"00000010",
  58594=>"00000011",
  58595=>"00000000",
  58596=>"11111101",
  58597=>"00000010",
  58598=>"00000001",
  58599=>"00000001",
  58600=>"11111101",
  58601=>"00000011",
  58602=>"11111110",
  58603=>"11111111",
  58604=>"00000001",
  58605=>"00000001",
  58606=>"00000010",
  58607=>"11111110",
  58608=>"00000001",
  58609=>"00000000",
  58610=>"11111111",
  58611=>"00000010",
  58612=>"00000010",
  58613=>"11111101",
  58614=>"00000010",
  58615=>"00000000",
  58616=>"11111111",
  58617=>"11111110",
  58618=>"11111111",
  58619=>"11111111",
  58620=>"11111110",
  58621=>"00000001",
  58622=>"11111100",
  58623=>"11111110",
  58624=>"11111111",
  58625=>"00000001",
  58626=>"00000010",
  58627=>"00000000",
  58628=>"00000000",
  58629=>"11111110",
  58630=>"11111110",
  58631=>"00000010",
  58632=>"11111111",
  58633=>"11111110",
  58634=>"00000001",
  58635=>"11111111",
  58636=>"11111110",
  58637=>"00000010",
  58638=>"11111110",
  58639=>"00000000",
  58640=>"11111101",
  58641=>"11111110",
  58642=>"00000001",
  58643=>"11111100",
  58644=>"11111111",
  58645=>"00000000",
  58646=>"00000010",
  58647=>"00000000",
  58648=>"00000001",
  58649=>"11111110",
  58650=>"11111101",
  58651=>"11111101",
  58652=>"00000001",
  58653=>"11111110",
  58654=>"11111110",
  58655=>"11111111",
  58656=>"00000011",
  58657=>"11111110",
  58658=>"00000010",
  58659=>"11111111",
  58660=>"11111111",
  58661=>"11111101",
  58662=>"11111110",
  58663=>"00000001",
  58664=>"11111111",
  58665=>"11111101",
  58666=>"00000010",
  58667=>"00000001",
  58668=>"00000001",
  58669=>"00000010",
  58670=>"11111111",
  58671=>"11111101",
  58672=>"11111110",
  58673=>"00000100",
  58674=>"11111110",
  58675=>"11111111",
  58676=>"00000000",
  58677=>"00000010",
  58678=>"00000100",
  58679=>"11111111",
  58680=>"11111101",
  58681=>"00000011",
  58682=>"11111110",
  58683=>"00000001",
  58684=>"11111101",
  58685=>"00000000",
  58686=>"11111111",
  58687=>"11111101",
  58688=>"00000000",
  58689=>"11111101",
  58690=>"00000000",
  58691=>"00000101",
  58692=>"11111111",
  58693=>"00000010",
  58694=>"00000001",
  58695=>"00000101",
  58696=>"00000100",
  58697=>"11111111",
  58698=>"00000000",
  58699=>"00000001",
  58700=>"00000000",
  58701=>"00000011",
  58702=>"00000010",
  58703=>"00000001",
  58704=>"00000010",
  58705=>"00000001",
  58706=>"00000001",
  58707=>"11111110",
  58708=>"00000001",
  58709=>"00000011",
  58710=>"00000011",
  58711=>"00000001",
  58712=>"00000001",
  58713=>"00000010",
  58714=>"00000001",
  58715=>"00000011",
  58716=>"11111110",
  58717=>"00000100",
  58718=>"00000001",
  58719=>"00000001",
  58720=>"11111110",
  58721=>"00000000",
  58722=>"00000010",
  58723=>"00000001",
  58724=>"11111111",
  58725=>"00000000",
  58726=>"11111111",
  58727=>"11111110",
  58728=>"11111101",
  58729=>"11111101",
  58730=>"00000011",
  58731=>"11111111",
  58732=>"00000010",
  58733=>"00000001",
  58734=>"11111101",
  58735=>"00000010",
  58736=>"00000000",
  58737=>"11111101",
  58738=>"11111111",
  58739=>"11111111",
  58740=>"00000010",
  58741=>"00000110",
  58742=>"11111101",
  58743=>"00000010",
  58744=>"00000010",
  58745=>"00000000",
  58746=>"00000101",
  58747=>"11111101",
  58748=>"00000010",
  58749=>"00000000",
  58750=>"00000010",
  58751=>"00000011",
  58752=>"11111110",
  58753=>"00000000",
  58754=>"11111111",
  58755=>"00000001",
  58756=>"11111110",
  58757=>"00000010",
  58758=>"00000001",
  58759=>"11111110",
  58760=>"00000010",
  58761=>"00000010",
  58762=>"00000001",
  58763=>"00000010",
  58764=>"00000000",
  58765=>"00000001",
  58766=>"00000001",
  58767=>"11111101",
  58768=>"00000001",
  58769=>"00000100",
  58770=>"00000000",
  58771=>"00000001",
  58772=>"00000011",
  58773=>"00000000",
  58774=>"00000000",
  58775=>"00000000",
  58776=>"11111100",
  58777=>"11111101",
  58778=>"00000100",
  58779=>"00000010",
  58780=>"00000001",
  58781=>"00000011",
  58782=>"00000010",
  58783=>"00000001",
  58784=>"00000000",
  58785=>"11111110",
  58786=>"00000000",
  58787=>"00000100",
  58788=>"11111110",
  58789=>"11111110",
  58790=>"11111101",
  58791=>"11111110",
  58792=>"00000010",
  58793=>"00000010",
  58794=>"00000110",
  58795=>"00000000",
  58796=>"00000000",
  58797=>"00000000",
  58798=>"11111111",
  58799=>"11111111",
  58800=>"11111111",
  58801=>"00000011",
  58802=>"00000010",
  58803=>"11111111",
  58804=>"11111111",
  58805=>"00000000",
  58806=>"11111101",
  58807=>"00000010",
  58808=>"00000001",
  58809=>"11111110",
  58810=>"11111110",
  58811=>"11111110",
  58812=>"00000010",
  58813=>"11111100",
  58814=>"11111101",
  58815=>"11111111",
  58816=>"11111111",
  58817=>"00000000",
  58818=>"11111110",
  58819=>"00000001",
  58820=>"00000000",
  58821=>"11111111",
  58822=>"00000000",
  58823=>"11111111",
  58824=>"11111100",
  58825=>"11111111",
  58826=>"00000000",
  58827=>"00000000",
  58828=>"00000001",
  58829=>"00000011",
  58830=>"00000010",
  58831=>"00000000",
  58832=>"00000010",
  58833=>"00000010",
  58834=>"00000011",
  58835=>"11111101",
  58836=>"11111110",
  58837=>"00000100",
  58838=>"00000000",
  58839=>"00000001",
  58840=>"11111110",
  58841=>"00000011",
  58842=>"00000001",
  58843=>"00000010",
  58844=>"11111110",
  58845=>"00000011",
  58846=>"11111111",
  58847=>"11111110",
  58848=>"00000001",
  58849=>"00000000",
  58850=>"00000010",
  58851=>"00000010",
  58852=>"00000001",
  58853=>"11111111",
  58854=>"11111111",
  58855=>"00000001",
  58856=>"00000000",
  58857=>"00000010",
  58858=>"11111111",
  58859=>"00000100",
  58860=>"00000011",
  58861=>"00000000",
  58862=>"00000010",
  58863=>"11111111",
  58864=>"00000010",
  58865=>"00000001",
  58866=>"00000001",
  58867=>"11111110",
  58868=>"00000000",
  58869=>"11111110",
  58870=>"00000011",
  58871=>"00000010",
  58872=>"11111110",
  58873=>"00000000",
  58874=>"00000001",
  58875=>"11111111",
  58876=>"00000000",
  58877=>"00000001",
  58878=>"00000000",
  58879=>"11111101",
  58880=>"11111111",
  58881=>"11111111",
  58882=>"00000010",
  58883=>"11111111",
  58884=>"00000000",
  58885=>"11111101",
  58886=>"00000011",
  58887=>"11111111",
  58888=>"11111101",
  58889=>"00000001",
  58890=>"00000001",
  58891=>"00000001",
  58892=>"00000000",
  58893=>"00000001",
  58894=>"00000000",
  58895=>"00000000",
  58896=>"11111111",
  58897=>"11111101",
  58898=>"00000000",
  58899=>"11111101",
  58900=>"11111111",
  58901=>"00000000",
  58902=>"00000010",
  58903=>"00000000",
  58904=>"11111110",
  58905=>"11111111",
  58906=>"00000010",
  58907=>"00000011",
  58908=>"00000000",
  58909=>"11111110",
  58910=>"00000010",
  58911=>"00000101",
  58912=>"00000001",
  58913=>"00000100",
  58914=>"00000011",
  58915=>"11111110",
  58916=>"11111101",
  58917=>"00000010",
  58918=>"11111111",
  58919=>"11111101",
  58920=>"11111111",
  58921=>"11111110",
  58922=>"00000001",
  58923=>"00000001",
  58924=>"00000010",
  58925=>"11111110",
  58926=>"11111111",
  58927=>"00000010",
  58928=>"11111111",
  58929=>"00000100",
  58930=>"11111101",
  58931=>"00000001",
  58932=>"11111111",
  58933=>"00000001",
  58934=>"11111110",
  58935=>"00000001",
  58936=>"11111111",
  58937=>"00000011",
  58938=>"00000000",
  58939=>"00000010",
  58940=>"11111110",
  58941=>"11111111",
  58942=>"00000001",
  58943=>"00000010",
  58944=>"11111110",
  58945=>"00000001",
  58946=>"11111110",
  58947=>"11111110",
  58948=>"00000000",
  58949=>"00000000",
  58950=>"11111110",
  58951=>"00000011",
  58952=>"00000000",
  58953=>"11111110",
  58954=>"00000010",
  58955=>"11111110",
  58956=>"00000000",
  58957=>"11111110",
  58958=>"00000100",
  58959=>"00000010",
  58960=>"11111110",
  58961=>"11111110",
  58962=>"00000000",
  58963=>"00000000",
  58964=>"00000001",
  58965=>"00000010",
  58966=>"11111111",
  58967=>"11111110",
  58968=>"00000001",
  58969=>"00000000",
  58970=>"11111110",
  58971=>"11111100",
  58972=>"11111110",
  58973=>"00000001",
  58974=>"00000101",
  58975=>"00000000",
  58976=>"11111110",
  58977=>"11111101",
  58978=>"00000000",
  58979=>"00000011",
  58980=>"00000000",
  58981=>"00000011",
  58982=>"00000001",
  58983=>"11111101",
  58984=>"11111110",
  58985=>"00000001",
  58986=>"11111110",
  58987=>"00000000",
  58988=>"00000010",
  58989=>"11111110",
  58990=>"00000001",
  58991=>"00000100",
  58992=>"11111110",
  58993=>"11111100",
  58994=>"11111111",
  58995=>"11111110",
  58996=>"00000010",
  58997=>"00000000",
  58998=>"00000001",
  58999=>"00000000",
  59000=>"11111110",
  59001=>"00000000",
  59002=>"00000000",
  59003=>"11111110",
  59004=>"11111101",
  59005=>"11111111",
  59006=>"00000001",
  59007=>"11111111",
  59008=>"11111111",
  59009=>"11111111",
  59010=>"11111110",
  59011=>"11111100",
  59012=>"00000010",
  59013=>"11111101",
  59014=>"11111110",
  59015=>"00000001",
  59016=>"00000011",
  59017=>"11111101",
  59018=>"11111111",
  59019=>"00000000",
  59020=>"11111111",
  59021=>"00000001",
  59022=>"11111101",
  59023=>"11111111",
  59024=>"00000000",
  59025=>"00000000",
  59026=>"00000000",
  59027=>"00000000",
  59028=>"11111111",
  59029=>"00000010",
  59030=>"11111100",
  59031=>"00000000",
  59032=>"11111110",
  59033=>"00000000",
  59034=>"00000001",
  59035=>"11111111",
  59036=>"11111101",
  59037=>"11111111",
  59038=>"00000010",
  59039=>"00000000",
  59040=>"00000010",
  59041=>"11111101",
  59042=>"00000001",
  59043=>"11111111",
  59044=>"11111101",
  59045=>"00000001",
  59046=>"00000011",
  59047=>"00000010",
  59048=>"00000010",
  59049=>"11111101",
  59050=>"11111110",
  59051=>"11111110",
  59052=>"00000100",
  59053=>"00000001",
  59054=>"00000010",
  59055=>"00000001",
  59056=>"11111101",
  59057=>"11111111",
  59058=>"11111111",
  59059=>"11111110",
  59060=>"11111110",
  59061=>"11111110",
  59062=>"11111111",
  59063=>"11111111",
  59064=>"00000001",
  59065=>"11111111",
  59066=>"00000010",
  59067=>"00000010",
  59068=>"00000001",
  59069=>"11111111",
  59070=>"11111111",
  59071=>"00000001",
  59072=>"00000001",
  59073=>"11111101",
  59074=>"11111100",
  59075=>"00000001",
  59076=>"00000001",
  59077=>"00000100",
  59078=>"00000000",
  59079=>"00000100",
  59080=>"11111111",
  59081=>"00000001",
  59082=>"11111101",
  59083=>"11111101",
  59084=>"11111111",
  59085=>"00000100",
  59086=>"00000001",
  59087=>"00000010",
  59088=>"11111111",
  59089=>"00000010",
  59090=>"00000001",
  59091=>"00000000",
  59092=>"00000001",
  59093=>"11111110",
  59094=>"11111110",
  59095=>"00000010",
  59096=>"11111110",
  59097=>"00000010",
  59098=>"00000000",
  59099=>"11111110",
  59100=>"00000001",
  59101=>"00000010",
  59102=>"00000001",
  59103=>"11111101",
  59104=>"11111101",
  59105=>"00000001",
  59106=>"00000010",
  59107=>"00000100",
  59108=>"00000011",
  59109=>"00000000",
  59110=>"00000001",
  59111=>"00000100",
  59112=>"11111110",
  59113=>"00000001",
  59114=>"00000100",
  59115=>"00000010",
  59116=>"00000000",
  59117=>"00000000",
  59118=>"11111110",
  59119=>"11111101",
  59120=>"11111111",
  59121=>"00000001",
  59122=>"00000000",
  59123=>"11111110",
  59124=>"11111101",
  59125=>"00000001",
  59126=>"00000001",
  59127=>"11111111",
  59128=>"00000000",
  59129=>"11111110",
  59130=>"00000000",
  59131=>"11111100",
  59132=>"11111110",
  59133=>"11111111",
  59134=>"11111110",
  59135=>"11111110",
  59136=>"11111110",
  59137=>"00000110",
  59138=>"00000010",
  59139=>"11111101",
  59140=>"11111111",
  59141=>"00000010",
  59142=>"11111101",
  59143=>"00000001",
  59144=>"00000010",
  59145=>"11111101",
  59146=>"11111111",
  59147=>"11111110",
  59148=>"00000001",
  59149=>"11111111",
  59150=>"11111110",
  59151=>"00000010",
  59152=>"11111110",
  59153=>"00000100",
  59154=>"00000010",
  59155=>"11111110",
  59156=>"00000001",
  59157=>"00000100",
  59158=>"00000001",
  59159=>"00000010",
  59160=>"00000001",
  59161=>"11111101",
  59162=>"11111100",
  59163=>"00000100",
  59164=>"00000001",
  59165=>"11111101",
  59166=>"00000101",
  59167=>"11111100",
  59168=>"11111101",
  59169=>"00000010",
  59170=>"11111101",
  59171=>"11111111",
  59172=>"00000000",
  59173=>"11111101",
  59174=>"00000110",
  59175=>"00000101",
  59176=>"11111101",
  59177=>"11111110",
  59178=>"11111111",
  59179=>"00000010",
  59180=>"00000000",
  59181=>"11111111",
  59182=>"00000011",
  59183=>"00000010",
  59184=>"11111101",
  59185=>"00000000",
  59186=>"11111101",
  59187=>"00000001",
  59188=>"11111111",
  59189=>"00000010",
  59190=>"00000000",
  59191=>"11111101",
  59192=>"11111100",
  59193=>"00000001",
  59194=>"00000010",
  59195=>"00000110",
  59196=>"00000010",
  59197=>"00000001",
  59198=>"00000101",
  59199=>"00000000",
  59200=>"00000010",
  59201=>"00000001",
  59202=>"11111101",
  59203=>"11111110",
  59204=>"00000101",
  59205=>"11111101",
  59206=>"00000000",
  59207=>"11111111",
  59208=>"11111111",
  59209=>"00000000",
  59210=>"00000100",
  59211=>"11111100",
  59212=>"00000010",
  59213=>"00000010",
  59214=>"00000001",
  59215=>"00000100",
  59216=>"11111111",
  59217=>"00000011",
  59218=>"00000000",
  59219=>"00000010",
  59220=>"00000001",
  59221=>"11111110",
  59222=>"00000001",
  59223=>"00000000",
  59224=>"00000001",
  59225=>"00000010",
  59226=>"11111110",
  59227=>"11111111",
  59228=>"00000011",
  59229=>"11111110",
  59230=>"11111110",
  59231=>"00000000",
  59232=>"11111101",
  59233=>"11111111",
  59234=>"11111101",
  59235=>"11111101",
  59236=>"00000001",
  59237=>"00000001",
  59238=>"11111110",
  59239=>"00000011",
  59240=>"11111101",
  59241=>"11111101",
  59242=>"00000101",
  59243=>"00000011",
  59244=>"00000000",
  59245=>"00000011",
  59246=>"00000010",
  59247=>"00000010",
  59248=>"00000011",
  59249=>"11111111",
  59250=>"00000000",
  59251=>"11111111",
  59252=>"00000000",
  59253=>"11111111",
  59254=>"11111101",
  59255=>"11111111",
  59256=>"11111101",
  59257=>"00000001",
  59258=>"00000010",
  59259=>"00000010",
  59260=>"00000010",
  59261=>"00000011",
  59262=>"00000000",
  59263=>"00000011",
  59264=>"00000000",
  59265=>"11111111",
  59266=>"00000001",
  59267=>"00000011",
  59268=>"11111101",
  59269=>"11111110",
  59270=>"00000001",
  59271=>"11111101",
  59272=>"11111101",
  59273=>"00000001",
  59274=>"00000011",
  59275=>"00000010",
  59276=>"00000010",
  59277=>"00000001",
  59278=>"00000101",
  59279=>"00000000",
  59280=>"11111111",
  59281=>"00000001",
  59282=>"00000100",
  59283=>"00000010",
  59284=>"00000010",
  59285=>"11111110",
  59286=>"11111111",
  59287=>"00000100",
  59288=>"00000001",
  59289=>"11111101",
  59290=>"00000010",
  59291=>"11111111",
  59292=>"11111111",
  59293=>"11111111",
  59294=>"11111111",
  59295=>"00000000",
  59296=>"00000011",
  59297=>"11111110",
  59298=>"11111110",
  59299=>"00000010",
  59300=>"11111110",
  59301=>"11111110",
  59302=>"00000101",
  59303=>"11111111",
  59304=>"11111110",
  59305=>"00000011",
  59306=>"11111110",
  59307=>"00000010",
  59308=>"00000001",
  59309=>"00000010",
  59310=>"11111111",
  59311=>"11111110",
  59312=>"11111111",
  59313=>"11111111",
  59314=>"11111110",
  59315=>"11111110",
  59316=>"00000001",
  59317=>"00000001",
  59318=>"11111111",
  59319=>"11111101",
  59320=>"00000001",
  59321=>"11111110",
  59322=>"00000001",
  59323=>"00000000",
  59324=>"11111111",
  59325=>"00000010",
  59326=>"11111110",
  59327=>"11111111",
  59328=>"11111110",
  59329=>"11111111",
  59330=>"11111110",
  59331=>"11111111",
  59332=>"00000001",
  59333=>"11111110",
  59334=>"00000011",
  59335=>"00000001",
  59336=>"11111110",
  59337=>"00000011",
  59338=>"00000010",
  59339=>"11111101",
  59340=>"00000010",
  59341=>"11111100",
  59342=>"11111110",
  59343=>"11111111",
  59344=>"11111111",
  59345=>"00000000",
  59346=>"00000001",
  59347=>"00000010",
  59348=>"11111110",
  59349=>"00000111",
  59350=>"11111101",
  59351=>"00000000",
  59352=>"11111101",
  59353=>"00000010",
  59354=>"11111111",
  59355=>"11111111",
  59356=>"00000011",
  59357=>"00000010",
  59358=>"00000001",
  59359=>"00000010",
  59360=>"11111101",
  59361=>"11111110",
  59362=>"11111111",
  59363=>"00000001",
  59364=>"11111111",
  59365=>"11111110",
  59366=>"00000000",
  59367=>"00000000",
  59368=>"11111110",
  59369=>"11111110",
  59370=>"00000000",
  59371=>"11111101",
  59372=>"11111110",
  59373=>"00000010",
  59374=>"11111111",
  59375=>"00000010",
  59376=>"11111111",
  59377=>"11111101",
  59378=>"00000000",
  59379=>"11111111",
  59380=>"11111101",
  59381=>"00000010",
  59382=>"11111101",
  59383=>"11111100",
  59384=>"00000010",
  59385=>"00000000",
  59386=>"00000011",
  59387=>"00000000",
  59388=>"11111100",
  59389=>"11111111",
  59390=>"00000010",
  59391=>"11111101",
  59392=>"00000000",
  59393=>"00000010",
  59394=>"00000010",
  59395=>"00000001",
  59396=>"11111101",
  59397=>"11111101",
  59398=>"11111111",
  59399=>"11111110",
  59400=>"11111111",
  59401=>"00000101",
  59402=>"11111110",
  59403=>"00000100",
  59404=>"00000011",
  59405=>"00000000",
  59406=>"00000001",
  59407=>"11111110",
  59408=>"00000101",
  59409=>"11111101",
  59410=>"00000000",
  59411=>"00000001",
  59412=>"11111101",
  59413=>"00000001",
  59414=>"00000100",
  59415=>"00000010",
  59416=>"11111101",
  59417=>"11111110",
  59418=>"11111110",
  59419=>"11111110",
  59420=>"00000010",
  59421=>"00000001",
  59422=>"11111110",
  59423=>"11111110",
  59424=>"00000010",
  59425=>"00000100",
  59426=>"11111101",
  59427=>"00000000",
  59428=>"11111110",
  59429=>"00000000",
  59430=>"00000100",
  59431=>"00000010",
  59432=>"00000010",
  59433=>"11111101",
  59434=>"11111111",
  59435=>"11111111",
  59436=>"00000001",
  59437=>"00000011",
  59438=>"00000001",
  59439=>"00000000",
  59440=>"11111110",
  59441=>"11111101",
  59442=>"11111110",
  59443=>"11111101",
  59444=>"00000001",
  59445=>"11111101",
  59446=>"00000010",
  59447=>"00000101",
  59448=>"00000000",
  59449=>"11111110",
  59450=>"11111101",
  59451=>"11111111",
  59452=>"00000010",
  59453=>"11111111",
  59454=>"00000001",
  59455=>"11111110",
  59456=>"11111110",
  59457=>"11111110",
  59458=>"11111111",
  59459=>"00000000",
  59460=>"00000011",
  59461=>"00000010",
  59462=>"11111110",
  59463=>"11111110",
  59464=>"00000101",
  59465=>"00000011",
  59466=>"00000001",
  59467=>"00000001",
  59468=>"00000110",
  59469=>"11111110",
  59470=>"11111111",
  59471=>"00000010",
  59472=>"11111111",
  59473=>"00000001",
  59474=>"00000100",
  59475=>"11111101",
  59476=>"00000010",
  59477=>"00000011",
  59478=>"11111101",
  59479=>"00000000",
  59480=>"00000010",
  59481=>"11111111",
  59482=>"00000001",
  59483=>"00000001",
  59484=>"00000000",
  59485=>"00000001",
  59486=>"11111101",
  59487=>"11111101",
  59488=>"00000001",
  59489=>"11111100",
  59490=>"11111111",
  59491=>"11111111",
  59492=>"00000010",
  59493=>"00000010",
  59494=>"00000010",
  59495=>"00000001",
  59496=>"00000000",
  59497=>"00000000",
  59498=>"11111111",
  59499=>"11111110",
  59500=>"00000000",
  59501=>"00000010",
  59502=>"11111111",
  59503=>"11111101",
  59504=>"00000001",
  59505=>"11111101",
  59506=>"11111111",
  59507=>"11111111",
  59508=>"00000010",
  59509=>"11111111",
  59510=>"00000101",
  59511=>"00000011",
  59512=>"00000010",
  59513=>"00000010",
  59514=>"11111110",
  59515=>"11111111",
  59516=>"00000001",
  59517=>"11111111",
  59518=>"00000000",
  59519=>"00000000",
  59520=>"00000001",
  59521=>"00000010",
  59522=>"00000001",
  59523=>"00000000",
  59524=>"00000001",
  59525=>"00000000",
  59526=>"11111111",
  59527=>"11111111",
  59528=>"11111110",
  59529=>"11111101",
  59530=>"00000010",
  59531=>"00000001",
  59532=>"00000010",
  59533=>"00000001",
  59534=>"11111101",
  59535=>"11111111",
  59536=>"00000010",
  59537=>"11111110",
  59538=>"00000011",
  59539=>"00000000",
  59540=>"00000001",
  59541=>"00000000",
  59542=>"11111110",
  59543=>"11111110",
  59544=>"00000010",
  59545=>"00000001",
  59546=>"00000010",
  59547=>"11111111",
  59548=>"11111110",
  59549=>"11111101",
  59550=>"00000010",
  59551=>"00000000",
  59552=>"11111110",
  59553=>"00000000",
  59554=>"00000010",
  59555=>"00000010",
  59556=>"11111111",
  59557=>"11111111",
  59558=>"11111110",
  59559=>"00000000",
  59560=>"11111111",
  59561=>"11111101",
  59562=>"00000010",
  59563=>"11111111",
  59564=>"00000011",
  59565=>"00000000",
  59566=>"00000010",
  59567=>"00000001",
  59568=>"00000010",
  59569=>"00000000",
  59570=>"11111110",
  59571=>"00000000",
  59572=>"00000000",
  59573=>"00000011",
  59574=>"00000001",
  59575=>"11111111",
  59576=>"11111111",
  59577=>"00000000",
  59578=>"00000100",
  59579=>"11111110",
  59580=>"00000001",
  59581=>"00000000",
  59582=>"00000001",
  59583=>"00000010",
  59584=>"11111110",
  59585=>"00000001",
  59586=>"00000010",
  59587=>"00000000",
  59588=>"11111101",
  59589=>"11111110",
  59590=>"11111101",
  59591=>"11111110",
  59592=>"00000001",
  59593=>"00000010",
  59594=>"00000000",
  59595=>"11111100",
  59596=>"11111101",
  59597=>"00000000",
  59598=>"00000010",
  59599=>"00000010",
  59600=>"11111110",
  59601=>"00000101",
  59602=>"00000000",
  59603=>"00000011",
  59604=>"00000000",
  59605=>"11111111",
  59606=>"11111111",
  59607=>"00000011",
  59608=>"11111101",
  59609=>"11111110",
  59610=>"00000010",
  59611=>"00000001",
  59612=>"00000000",
  59613=>"11111111",
  59614=>"00000111",
  59615=>"00000001",
  59616=>"11111110",
  59617=>"00000000",
  59618=>"11111111",
  59619=>"11111111",
  59620=>"00000001",
  59621=>"11111111",
  59622=>"00000000",
  59623=>"11111110",
  59624=>"11111101",
  59625=>"11111110",
  59626=>"11111111",
  59627=>"11111110",
  59628=>"00000001",
  59629=>"11111110",
  59630=>"11111101",
  59631=>"00000010",
  59632=>"11111101",
  59633=>"00000001",
  59634=>"00000000",
  59635=>"00000001",
  59636=>"11111101",
  59637=>"11111101",
  59638=>"11111110",
  59639=>"11111110",
  59640=>"11111101",
  59641=>"11111110",
  59642=>"00000101",
  59643=>"00000010",
  59644=>"00000001",
  59645=>"00000000",
  59646=>"00000100",
  59647=>"00000001",
  59648=>"11111111",
  59649=>"11111110",
  59650=>"11111110",
  59651=>"11111111",
  59652=>"00000001",
  59653=>"00000001",
  59654=>"11111111",
  59655=>"00000000",
  59656=>"11111101",
  59657=>"00000010",
  59658=>"00000011",
  59659=>"00000000",
  59660=>"11111110",
  59661=>"11111101",
  59662=>"00000001",
  59663=>"00000010",
  59664=>"00000010",
  59665=>"11111110",
  59666=>"11111100",
  59667=>"00000010",
  59668=>"11111110",
  59669=>"11111111",
  59670=>"00000010",
  59671=>"00000000",
  59672=>"11111111",
  59673=>"00000001",
  59674=>"00000000",
  59675=>"11111110",
  59676=>"11111110",
  59677=>"11111110",
  59678=>"11111101",
  59679=>"00000011",
  59680=>"00000000",
  59681=>"11111111",
  59682=>"11111101",
  59683=>"11111101",
  59684=>"11111011",
  59685=>"11111111",
  59686=>"00000001",
  59687=>"11111100",
  59688=>"00000000",
  59689=>"00000001",
  59690=>"00000000",
  59691=>"00000000",
  59692=>"00000001",
  59693=>"11111110",
  59694=>"00000010",
  59695=>"00000000",
  59696=>"00000000",
  59697=>"00000011",
  59698=>"11111110",
  59699=>"00000011",
  59700=>"11111110",
  59701=>"11111101",
  59702=>"11111110",
  59703=>"00000001",
  59704=>"00000010",
  59705=>"00000000",
  59706=>"00000010",
  59707=>"11111101",
  59708=>"00000010",
  59709=>"00000010",
  59710=>"11111101",
  59711=>"11111110",
  59712=>"11111110",
  59713=>"00000000",
  59714=>"11111110",
  59715=>"11111110",
  59716=>"00000000",
  59717=>"11111101",
  59718=>"11111111",
  59719=>"11111101",
  59720=>"00000100",
  59721=>"00000001",
  59722=>"00000000",
  59723=>"00000000",
  59724=>"11111101",
  59725=>"00000001",
  59726=>"11111101",
  59727=>"11111111",
  59728=>"00000011",
  59729=>"11111110",
  59730=>"11111110",
  59731=>"00000110",
  59732=>"00000000",
  59733=>"11111111",
  59734=>"00000000",
  59735=>"00000000",
  59736=>"00000010",
  59737=>"00000001",
  59738=>"00000000",
  59739=>"00000010",
  59740=>"00000000",
  59741=>"00000001",
  59742=>"00000011",
  59743=>"00000100",
  59744=>"00000001",
  59745=>"11111101",
  59746=>"11111101",
  59747=>"00000000",
  59748=>"11111110",
  59749=>"11111110",
  59750=>"00000000",
  59751=>"00000011",
  59752=>"11111110",
  59753=>"11111110",
  59754=>"00000000",
  59755=>"11111101",
  59756=>"00000001",
  59757=>"00000000",
  59758=>"00000100",
  59759=>"11111111",
  59760=>"00000010",
  59761=>"00000001",
  59762=>"00000000",
  59763=>"11111111",
  59764=>"00000000",
  59765=>"11111101",
  59766=>"00000001",
  59767=>"11111111",
  59768=>"00000010",
  59769=>"00000000",
  59770=>"00000010",
  59771=>"00000000",
  59772=>"11111101",
  59773=>"00000101",
  59774=>"00000001",
  59775=>"11111101",
  59776=>"11111101",
  59777=>"11111110",
  59778=>"11111111",
  59779=>"11111111",
  59780=>"00000001",
  59781=>"00000001",
  59782=>"11111110",
  59783=>"00000000",
  59784=>"00000010",
  59785=>"00000011",
  59786=>"00000101",
  59787=>"00000010",
  59788=>"00000000",
  59789=>"00000001",
  59790=>"11111111",
  59791=>"11111111",
  59792=>"00000000",
  59793=>"00000011",
  59794=>"00000101",
  59795=>"00000001",
  59796=>"11111100",
  59797=>"00000001",
  59798=>"11111101",
  59799=>"11111101",
  59800=>"11111110",
  59801=>"11111110",
  59802=>"00000000",
  59803=>"00000000",
  59804=>"00000011",
  59805=>"00000100",
  59806=>"00000000",
  59807=>"11111110",
  59808=>"11111111",
  59809=>"00000010",
  59810=>"00000000",
  59811=>"00000010",
  59812=>"00000010",
  59813=>"00000000",
  59814=>"00000100",
  59815=>"00000000",
  59816=>"11111111",
  59817=>"00000010",
  59818=>"00000010",
  59819=>"00000010",
  59820=>"11111111",
  59821=>"00000010",
  59822=>"11111110",
  59823=>"00000010",
  59824=>"00000010",
  59825=>"11111110",
  59826=>"00000001",
  59827=>"00000010",
  59828=>"11111101",
  59829=>"00000010",
  59830=>"00000100",
  59831=>"00000000",
  59832=>"00000010",
  59833=>"00000000",
  59834=>"00000010",
  59835=>"00000001",
  59836=>"00000000",
  59837=>"00000001",
  59838=>"00000001",
  59839=>"00000101",
  59840=>"00000000",
  59841=>"11111101",
  59842=>"00000010",
  59843=>"11111110",
  59844=>"00000010",
  59845=>"11111111",
  59846=>"00000001",
  59847=>"11111110",
  59848=>"11111110",
  59849=>"00000011",
  59850=>"11111110",
  59851=>"00000010",
  59852=>"11111111",
  59853=>"00000001",
  59854=>"00000000",
  59855=>"11111110",
  59856=>"11111101",
  59857=>"11111111",
  59858=>"11111101",
  59859=>"11111101",
  59860=>"11111101",
  59861=>"11111100",
  59862=>"00000000",
  59863=>"00000001",
  59864=>"00000001",
  59865=>"00000000",
  59866=>"00000000",
  59867=>"11111110",
  59868=>"11111101",
  59869=>"11111111",
  59870=>"11111101",
  59871=>"11111111",
  59872=>"00000000",
  59873=>"00000001",
  59874=>"00000010",
  59875=>"00000000",
  59876=>"00000000",
  59877=>"00000001",
  59878=>"00000010",
  59879=>"00000001",
  59880=>"11111110",
  59881=>"11111111",
  59882=>"11111111",
  59883=>"00000000",
  59884=>"00000101",
  59885=>"11111100",
  59886=>"00000001",
  59887=>"00000101",
  59888=>"11111111",
  59889=>"00000011",
  59890=>"11111110",
  59891=>"11111111",
  59892=>"11111100",
  59893=>"00000001",
  59894=>"11111101",
  59895=>"00000000",
  59896=>"00000000",
  59897=>"00000010",
  59898=>"00000001",
  59899=>"11111111",
  59900=>"11111111",
  59901=>"00000001",
  59902=>"11111101",
  59903=>"00000011",
  59904=>"00000001",
  59905=>"00000001",
  59906=>"11111111",
  59907=>"11111110",
  59908=>"00000000",
  59909=>"11111110",
  59910=>"11111101",
  59911=>"00000110",
  59912=>"11111111",
  59913=>"00000011",
  59914=>"00000000",
  59915=>"11111111",
  59916=>"11111111",
  59917=>"00000001",
  59918=>"11111111",
  59919=>"00000011",
  59920=>"00000010",
  59921=>"00000000",
  59922=>"11111110",
  59923=>"11111110",
  59924=>"11111110",
  59925=>"00000000",
  59926=>"11111110",
  59927=>"00000001",
  59928=>"11111101",
  59929=>"00000110",
  59930=>"11111101",
  59931=>"11111110",
  59932=>"00000001",
  59933=>"11111110",
  59934=>"11111110",
  59935=>"11111111",
  59936=>"00000010",
  59937=>"00000001",
  59938=>"00000010",
  59939=>"11111111",
  59940=>"00000001",
  59941=>"11111110",
  59942=>"11111111",
  59943=>"11111111",
  59944=>"00000000",
  59945=>"00000010",
  59946=>"00000001",
  59947=>"11111110",
  59948=>"11111111",
  59949=>"11111101",
  59950=>"11111110",
  59951=>"00000001",
  59952=>"00000001",
  59953=>"11111110",
  59954=>"11111111",
  59955=>"11111110",
  59956=>"00000000",
  59957=>"00000001",
  59958=>"00000100",
  59959=>"00000010",
  59960=>"11111111",
  59961=>"00000011",
  59962=>"11111110",
  59963=>"11111111",
  59964=>"11111101",
  59965=>"11111111",
  59966=>"00000010",
  59967=>"11111101",
  59968=>"11111101",
  59969=>"00000100",
  59970=>"00000000",
  59971=>"11111101",
  59972=>"00000100",
  59973=>"00000010",
  59974=>"11111110",
  59975=>"00000000",
  59976=>"00000010",
  59977=>"11111111",
  59978=>"00000001",
  59979=>"11111111",
  59980=>"00000010",
  59981=>"00000010",
  59982=>"11111101",
  59983=>"00000000",
  59984=>"11111111",
  59985=>"00000001",
  59986=>"00000010",
  59987=>"11111101",
  59988=>"11111101",
  59989=>"00000000",
  59990=>"00000010",
  59991=>"11111111",
  59992=>"11111111",
  59993=>"11111110",
  59994=>"00000001",
  59995=>"00000100",
  59996=>"00000011",
  59997=>"00000000",
  59998=>"00000100",
  59999=>"00000101",
  60000=>"11111111",
  60001=>"11111111",
  60002=>"11111110",
  60003=>"11111110",
  60004=>"11111110",
  60005=>"11111110",
  60006=>"00000010",
  60007=>"11111101",
  60008=>"00000011",
  60009=>"00000001",
  60010=>"00000000",
  60011=>"00000001",
  60012=>"00000001",
  60013=>"00000011",
  60014=>"00000010",
  60015=>"00000001",
  60016=>"11111110",
  60017=>"00000000",
  60018=>"11111101",
  60019=>"11111111",
  60020=>"11111110",
  60021=>"11111101",
  60022=>"00000001",
  60023=>"00000001",
  60024=>"11111111",
  60025=>"00000000",
  60026=>"11111111",
  60027=>"11111101",
  60028=>"11111110",
  60029=>"11111101",
  60030=>"11111100",
  60031=>"00000000",
  60032=>"11111111",
  60033=>"11111110",
  60034=>"00000011",
  60035=>"11111111",
  60036=>"00000001",
  60037=>"00000001",
  60038=>"00000000",
  60039=>"00000000",
  60040=>"11111111",
  60041=>"11111111",
  60042=>"11111101",
  60043=>"11111101",
  60044=>"00000011",
  60045=>"11111101",
  60046=>"11111101",
  60047=>"11111110",
  60048=>"00000001",
  60049=>"00000010",
  60050=>"00000000",
  60051=>"00000011",
  60052=>"11111101",
  60053=>"11111111",
  60054=>"00000011",
  60055=>"00000000",
  60056=>"11111110",
  60057=>"11111110",
  60058=>"00000101",
  60059=>"11111111",
  60060=>"11111111",
  60061=>"00000001",
  60062=>"00000101",
  60063=>"00000001",
  60064=>"11111110",
  60065=>"00000001",
  60066=>"11111110",
  60067=>"00000000",
  60068=>"00000001",
  60069=>"11111101",
  60070=>"11111111",
  60071=>"11111100",
  60072=>"11111110",
  60073=>"00000001",
  60074=>"11111101",
  60075=>"11111111",
  60076=>"00000001",
  60077=>"11111110",
  60078=>"11111110",
  60079=>"11111110",
  60080=>"11111110",
  60081=>"00000011",
  60082=>"11111111",
  60083=>"11111111",
  60084=>"11111110",
  60085=>"11111101",
  60086=>"00000010",
  60087=>"11111111",
  60088=>"11111110",
  60089=>"00000001",
  60090=>"00000010",
  60091=>"00000001",
  60092=>"00000001",
  60093=>"11111111",
  60094=>"00000001",
  60095=>"00000000",
  60096=>"11111111",
  60097=>"00000000",
  60098=>"11111101",
  60099=>"11111101",
  60100=>"00000001",
  60101=>"00000100",
  60102=>"11111100",
  60103=>"00000010",
  60104=>"11111111",
  60105=>"11111101",
  60106=>"11111100",
  60107=>"00000001",
  60108=>"11111110",
  60109=>"11111111",
  60110=>"11111101",
  60111=>"00000000",
  60112=>"11111110",
  60113=>"11111110",
  60114=>"00000001",
  60115=>"00000010",
  60116=>"11111111",
  60117=>"00000001",
  60118=>"00000010",
  60119=>"00000000",
  60120=>"00000100",
  60121=>"00000000",
  60122=>"00000001",
  60123=>"11111101",
  60124=>"11111110",
  60125=>"00000001",
  60126=>"00000001",
  60127=>"00000000",
  60128=>"00000001",
  60129=>"11111101",
  60130=>"00000011",
  60131=>"11111101",
  60132=>"00000011",
  60133=>"00000001",
  60134=>"11111101",
  60135=>"11111110",
  60136=>"00000000",
  60137=>"11111101",
  60138=>"11111101",
  60139=>"00000011",
  60140=>"11111111",
  60141=>"11111110",
  60142=>"11111111",
  60143=>"00000001",
  60144=>"00000000",
  60145=>"11111111",
  60146=>"11111110",
  60147=>"11111110",
  60148=>"11111101",
  60149=>"11111101",
  60150=>"00000010",
  60151=>"00000010",
  60152=>"11111111",
  60153=>"11111110",
  60154=>"00000001",
  60155=>"00000001",
  60156=>"11111110",
  60157=>"11111110",
  60158=>"11111111",
  60159=>"00000010",
  60160=>"11111111",
  60161=>"11111101",
  60162=>"00000000",
  60163=>"00000000",
  60164=>"00000000",
  60165=>"00000001",
  60166=>"00000000",
  60167=>"11111111",
  60168=>"00000011",
  60169=>"00000001",
  60170=>"11111110",
  60171=>"00000000",
  60172=>"00000011",
  60173=>"00000000",
  60174=>"00000010",
  60175=>"00000010",
  60176=>"00000001",
  60177=>"11111101",
  60178=>"00000000",
  60179=>"00000100",
  60180=>"11111101",
  60181=>"00000000",
  60182=>"00000001",
  60183=>"00000001",
  60184=>"00000011",
  60185=>"11111101",
  60186=>"00000000",
  60187=>"11111100",
  60188=>"00000010",
  60189=>"11111100",
  60190=>"11111111",
  60191=>"11111101",
  60192=>"11111101",
  60193=>"11111111",
  60194=>"00000001",
  60195=>"00000001",
  60196=>"11111110",
  60197=>"11111110",
  60198=>"11111101",
  60199=>"11111110",
  60200=>"00000001",
  60201=>"11111111",
  60202=>"11111111",
  60203=>"00000001",
  60204=>"00000011",
  60205=>"00000000",
  60206=>"11111111",
  60207=>"00000010",
  60208=>"00000000",
  60209=>"11111101",
  60210=>"00000010",
  60211=>"00000000",
  60212=>"00000001",
  60213=>"11111110",
  60214=>"00000000",
  60215=>"11111110",
  60216=>"11111111",
  60217=>"11111110",
  60218=>"00000000",
  60219=>"11111110",
  60220=>"11111111",
  60221=>"11111111",
  60222=>"00000000",
  60223=>"11111110",
  60224=>"11111111",
  60225=>"00000001",
  60226=>"11111101",
  60227=>"00000001",
  60228=>"00000001",
  60229=>"11111110",
  60230=>"11111101",
  60231=>"00000001",
  60232=>"00000010",
  60233=>"00000001",
  60234=>"00000000",
  60235=>"00000000",
  60236=>"11111110",
  60237=>"11111101",
  60238=>"11111110",
  60239=>"00000011",
  60240=>"11111101",
  60241=>"11111101",
  60242=>"11111111",
  60243=>"00000001",
  60244=>"11111110",
  60245=>"11111101",
  60246=>"11111111",
  60247=>"00000001",
  60248=>"11111110",
  60249=>"11111101",
  60250=>"11111101",
  60251=>"11111111",
  60252=>"11111110",
  60253=>"11111110",
  60254=>"00000000",
  60255=>"00000001",
  60256=>"11111110",
  60257=>"00000101",
  60258=>"00000001",
  60259=>"11111110",
  60260=>"00000011",
  60261=>"00000001",
  60262=>"00000011",
  60263=>"11111111",
  60264=>"00000000",
  60265=>"00000010",
  60266=>"00000001",
  60267=>"00000000",
  60268=>"00000001",
  60269=>"11111011",
  60270=>"00000000",
  60271=>"00000001",
  60272=>"11111100",
  60273=>"00000010",
  60274=>"00000000",
  60275=>"11111111",
  60276=>"00000011",
  60277=>"00000010",
  60278=>"11111110",
  60279=>"00000010",
  60280=>"00000011",
  60281=>"00000000",
  60282=>"11111111",
  60283=>"11111101",
  60284=>"00000101",
  60285=>"00000011",
  60286=>"00000111",
  60287=>"11111110",
  60288=>"00000001",
  60289=>"00000100",
  60290=>"00000000",
  60291=>"11111111",
  60292=>"11111111",
  60293=>"11111111",
  60294=>"00000100",
  60295=>"00000010",
  60296=>"11111100",
  60297=>"00000001",
  60298=>"11111110",
  60299=>"00000001",
  60300=>"00000000",
  60301=>"00000010",
  60302=>"00000000",
  60303=>"00000011",
  60304=>"11111110",
  60305=>"00000001",
  60306=>"11111110",
  60307=>"11111101",
  60308=>"00000001",
  60309=>"00000000",
  60310=>"00000010",
  60311=>"00000010",
  60312=>"11111101",
  60313=>"11111111",
  60314=>"00000010",
  60315=>"11111101",
  60316=>"11111110",
  60317=>"00000010",
  60318=>"11111110",
  60319=>"11111101",
  60320=>"11111111",
  60321=>"00000010",
  60322=>"00000000",
  60323=>"00000010",
  60324=>"11111110",
  60325=>"00000000",
  60326=>"00000011",
  60327=>"11111110",
  60328=>"11111110",
  60329=>"00000001",
  60330=>"00000001",
  60331=>"11111101",
  60332=>"00000000",
  60333=>"11111101",
  60334=>"00000010",
  60335=>"00000000",
  60336=>"00000001",
  60337=>"11111110",
  60338=>"00000100",
  60339=>"00000001",
  60340=>"00000010",
  60341=>"00000100",
  60342=>"11111111",
  60343=>"11111101",
  60344=>"11111101",
  60345=>"11111110",
  60346=>"11111110",
  60347=>"11111111",
  60348=>"11111110",
  60349=>"11111110",
  60350=>"11111111",
  60351=>"00000001",
  60352=>"11111101",
  60353=>"00000011",
  60354=>"11111111",
  60355=>"11111110",
  60356=>"00000000",
  60357=>"11111101",
  60358=>"11111111",
  60359=>"00000001",
  60360=>"00000001",
  60361=>"11111101",
  60362=>"00000001",
  60363=>"11111111",
  60364=>"11111110",
  60365=>"00000010",
  60366=>"11111101",
  60367=>"11111101",
  60368=>"11111101",
  60369=>"00000001",
  60370=>"00000000",
  60371=>"00000011",
  60372=>"00000000",
  60373=>"11111101",
  60374=>"00000001",
  60375=>"00000001",
  60376=>"11111111",
  60377=>"11111101",
  60378=>"00000011",
  60379=>"00000000",
  60380=>"11111111",
  60381=>"11111110",
  60382=>"11111101",
  60383=>"00000010",
  60384=>"11111110",
  60385=>"00000000",
  60386=>"00000001",
  60387=>"00000010",
  60388=>"00000001",
  60389=>"11111110",
  60390=>"11111111",
  60391=>"00000000",
  60392=>"11111111",
  60393=>"11111111",
  60394=>"00000010",
  60395=>"11111111",
  60396=>"11111110",
  60397=>"11111101",
  60398=>"11111111",
  60399=>"00000000",
  60400=>"00000001",
  60401=>"11111101",
  60402=>"11111110",
  60403=>"11111111",
  60404=>"11111111",
  60405=>"11111111",
  60406=>"00000010",
  60407=>"11111111",
  60408=>"11111101",
  60409=>"00000010",
  60410=>"11111110",
  60411=>"11111111",
  60412=>"11111110",
  60413=>"11111111",
  60414=>"00000010",
  60415=>"00000001",
  60416=>"00000010",
  60417=>"00000011",
  60418=>"11111111",
  60419=>"11111111",
  60420=>"00000001",
  60421=>"00000011",
  60422=>"00000011",
  60423=>"11111101",
  60424=>"00000000",
  60425=>"00000010",
  60426=>"00000001",
  60427=>"00000000",
  60428=>"00000100",
  60429=>"00000010",
  60430=>"00000000",
  60431=>"00000011",
  60432=>"00000000",
  60433=>"11111100",
  60434=>"11111110",
  60435=>"00000001",
  60436=>"11111101",
  60437=>"11111110",
  60438=>"11111110",
  60439=>"11111111",
  60440=>"11111100",
  60441=>"00000011",
  60442=>"00000011",
  60443=>"00000000",
  60444=>"00000011",
  60445=>"00000010",
  60446=>"00000011",
  60447=>"00000010",
  60448=>"11111111",
  60449=>"11111111",
  60450=>"11111101",
  60451=>"00000001",
  60452=>"11111111",
  60453=>"11111110",
  60454=>"00000000",
  60455=>"00000010",
  60456=>"11111100",
  60457=>"00000001",
  60458=>"11111111",
  60459=>"00000101",
  60460=>"00000011",
  60461=>"11111111",
  60462=>"00000000",
  60463=>"11111101",
  60464=>"11111111",
  60465=>"00000011",
  60466=>"00000001",
  60467=>"11111110",
  60468=>"11111110",
  60469=>"11111110",
  60470=>"00000000",
  60471=>"11111110",
  60472=>"11111100",
  60473=>"11111110",
  60474=>"00000000",
  60475=>"00000001",
  60476=>"00000010",
  60477=>"11111111",
  60478=>"00000000",
  60479=>"00000100",
  60480=>"00000001",
  60481=>"00000001",
  60482=>"11111110",
  60483=>"00000011",
  60484=>"00000001",
  60485=>"00000100",
  60486=>"00000100",
  60487=>"00000010",
  60488=>"11111110",
  60489=>"00000011",
  60490=>"00000001",
  60491=>"00000011",
  60492=>"11111110",
  60493=>"00000000",
  60494=>"00000010",
  60495=>"00000000",
  60496=>"11111111",
  60497=>"00000010",
  60498=>"00000110",
  60499=>"11111110",
  60500=>"00000011",
  60501=>"11111111",
  60502=>"11111111",
  60503=>"00000100",
  60504=>"00000000",
  60505=>"11111011",
  60506=>"00000100",
  60507=>"11111100",
  60508=>"00000000",
  60509=>"11111111",
  60510=>"00000100",
  60511=>"00001000",
  60512=>"11111101",
  60513=>"11111101",
  60514=>"00000011",
  60515=>"11111101",
  60516=>"11111101",
  60517=>"11111111",
  60518=>"00000011",
  60519=>"11111111",
  60520=>"00000000",
  60521=>"00000001",
  60522=>"00000100",
  60523=>"11111111",
  60524=>"00000100",
  60525=>"00000001",
  60526=>"00000000",
  60527=>"00000011",
  60528=>"11111111",
  60529=>"11111101",
  60530=>"11111110",
  60531=>"11111101",
  60532=>"11111111",
  60533=>"00000011",
  60534=>"11111100",
  60535=>"00000001",
  60536=>"00000101",
  60537=>"11111111",
  60538=>"00000001",
  60539=>"11111110",
  60540=>"00000010",
  60541=>"00000001",
  60542=>"11111110",
  60543=>"00000011",
  60544=>"11111100",
  60545=>"11111110",
  60546=>"00000010",
  60547=>"11111110",
  60548=>"00000001",
  60549=>"00000011",
  60550=>"00000000",
  60551=>"00000010",
  60552=>"00000000",
  60553=>"11111101",
  60554=>"00000000",
  60555=>"11111101",
  60556=>"00000010",
  60557=>"00000010",
  60558=>"11111111",
  60559=>"00000000",
  60560=>"00000000",
  60561=>"00000001",
  60562=>"11111111",
  60563=>"11111101",
  60564=>"11111111",
  60565=>"00000000",
  60566=>"00000011",
  60567=>"00000000",
  60568=>"00000010",
  60569=>"00000011",
  60570=>"00000011",
  60571=>"00000000",
  60572=>"00000001",
  60573=>"11111100",
  60574=>"11111111",
  60575=>"00000000",
  60576=>"11111110",
  60577=>"00000000",
  60578=>"00000001",
  60579=>"00000010",
  60580=>"11111111",
  60581=>"11111101",
  60582=>"00000101",
  60583=>"11111101",
  60584=>"11111111",
  60585=>"11111101",
  60586=>"11111111",
  60587=>"11111100",
  60588=>"00000000",
  60589=>"00000000",
  60590=>"11111110",
  60591=>"00000000",
  60592=>"11111101",
  60593=>"00000010",
  60594=>"11111101",
  60595=>"00000010",
  60596=>"11111110",
  60597=>"11111101",
  60598=>"00000000",
  60599=>"11111100",
  60600=>"00000011",
  60601=>"11111100",
  60602=>"00000010",
  60603=>"11111110",
  60604=>"00000000",
  60605=>"11111110",
  60606=>"00000011",
  60607=>"11111111",
  60608=>"11111110",
  60609=>"00000001",
  60610=>"00000011",
  60611=>"00000001",
  60612=>"00000001",
  60613=>"00000000",
  60614=>"00000010",
  60615=>"00000101",
  60616=>"00000001",
  60617=>"11111101",
  60618=>"00000011",
  60619=>"00000001",
  60620=>"00000010",
  60621=>"11111111",
  60622=>"11111111",
  60623=>"00000100",
  60624=>"00000100",
  60625=>"00000000",
  60626=>"00000000",
  60627=>"11111101",
  60628=>"00000010",
  60629=>"00000010",
  60630=>"00000000",
  60631=>"00000010",
  60632=>"00000001",
  60633=>"00000100",
  60634=>"11111110",
  60635=>"00000000",
  60636=>"11111011",
  60637=>"00000111",
  60638=>"11111100",
  60639=>"00000010",
  60640=>"00000000",
  60641=>"11111101",
  60642=>"11111101",
  60643=>"11111100",
  60644=>"00000000",
  60645=>"00000101",
  60646=>"11111011",
  60647=>"11111101",
  60648=>"11111110",
  60649=>"00000000",
  60650=>"11111110",
  60651=>"00000011",
  60652=>"11111110",
  60653=>"00000001",
  60654=>"00000010",
  60655=>"11111110",
  60656=>"00000001",
  60657=>"11111111",
  60658=>"11111110",
  60659=>"11111111",
  60660=>"11111110",
  60661=>"00000010",
  60662=>"00000010",
  60663=>"00000001",
  60664=>"00000000",
  60665=>"00000100",
  60666=>"00000001",
  60667=>"00000001",
  60668=>"00000001",
  60669=>"00000010",
  60670=>"00000101",
  60671=>"11111111",
  60672=>"00000001",
  60673=>"11111110",
  60674=>"00000000",
  60675=>"11111110",
  60676=>"11111110",
  60677=>"00000010",
  60678=>"11111101",
  60679=>"11111111",
  60680=>"00000001",
  60681=>"00000000",
  60682=>"11111110",
  60683=>"00000010",
  60684=>"11111111",
  60685=>"11111111",
  60686=>"00000101",
  60687=>"00000000",
  60688=>"00000001",
  60689=>"00000000",
  60690=>"00000000",
  60691=>"00000001",
  60692=>"00000011",
  60693=>"00000000",
  60694=>"11111110",
  60695=>"00000000",
  60696=>"11111111",
  60697=>"00000010",
  60698=>"11111101",
  60699=>"11111111",
  60700=>"11111101",
  60701=>"11111110",
  60702=>"00000010",
  60703=>"00000011",
  60704=>"11111110",
  60705=>"11111111",
  60706=>"00000010",
  60707=>"11111111",
  60708=>"00000100",
  60709=>"11111101",
  60710=>"00000001",
  60711=>"00000001",
  60712=>"11111111",
  60713=>"00000001",
  60714=>"00000010",
  60715=>"00000000",
  60716=>"11111110",
  60717=>"00000000",
  60718=>"00000101",
  60719=>"00000011",
  60720=>"00000001",
  60721=>"00000011",
  60722=>"11111111",
  60723=>"00000010",
  60724=>"11111110",
  60725=>"00000010",
  60726=>"11111100",
  60727=>"11111111",
  60728=>"11111111",
  60729=>"11111110",
  60730=>"00000001",
  60731=>"00000011",
  60732=>"00000000",
  60733=>"00000000",
  60734=>"00000000",
  60735=>"11111111",
  60736=>"00000010",
  60737=>"11111110",
  60738=>"00000001",
  60739=>"00000010",
  60740=>"00000010",
  60741=>"11111110",
  60742=>"00000001",
  60743=>"11111110",
  60744=>"11111110",
  60745=>"11111100",
  60746=>"00000011",
  60747=>"11111111",
  60748=>"00000001",
  60749=>"00000011",
  60750=>"00000011",
  60751=>"00000010",
  60752=>"11111111",
  60753=>"11111110",
  60754=>"11111110",
  60755=>"00000001",
  60756=>"00000001",
  60757=>"11111111",
  60758=>"11111101",
  60759=>"11111111",
  60760=>"00000001",
  60761=>"00000010",
  60762=>"00000001",
  60763=>"00000100",
  60764=>"11111110",
  60765=>"11111110",
  60766=>"00000000",
  60767=>"11111110",
  60768=>"00000001",
  60769=>"11111110",
  60770=>"11111101",
  60771=>"11111110",
  60772=>"11111111",
  60773=>"00000001",
  60774=>"00000001",
  60775=>"00000010",
  60776=>"00000001",
  60777=>"11111111",
  60778=>"00000010",
  60779=>"00000001",
  60780=>"11111101",
  60781=>"00000001",
  60782=>"00000011",
  60783=>"00000010",
  60784=>"11111110",
  60785=>"11111100",
  60786=>"11111110",
  60787=>"00000011",
  60788=>"00000000",
  60789=>"00000000",
  60790=>"11111101",
  60791=>"11111111",
  60792=>"11111101",
  60793=>"00000001",
  60794=>"11111101",
  60795=>"00000000",
  60796=>"11111101",
  60797=>"00000001",
  60798=>"00000010",
  60799=>"00000011",
  60800=>"11111111",
  60801=>"00000010",
  60802=>"11111111",
  60803=>"00000011",
  60804=>"11111111",
  60805=>"00000010",
  60806=>"00000000",
  60807=>"00000011",
  60808=>"11111110",
  60809=>"11111111",
  60810=>"11111110",
  60811=>"00000001",
  60812=>"11111111",
  60813=>"00000011",
  60814=>"11111110",
  60815=>"00000100",
  60816=>"11111101",
  60817=>"11111111",
  60818=>"00000001",
  60819=>"11111111",
  60820=>"00000101",
  60821=>"00000001",
  60822=>"00000000",
  60823=>"00000011",
  60824=>"00000001",
  60825=>"00000010",
  60826=>"00000001",
  60827=>"11111111",
  60828=>"00000011",
  60829=>"11111101",
  60830=>"11111110",
  60831=>"11111111",
  60832=>"00000010",
  60833=>"00000000",
  60834=>"00000000",
  60835=>"11111110",
  60836=>"11111111",
  60837=>"00000011",
  60838=>"11111101",
  60839=>"00000011",
  60840=>"11111111",
  60841=>"11111110",
  60842=>"00000000",
  60843=>"00000010",
  60844=>"11111111",
  60845=>"00000010",
  60846=>"11111110",
  60847=>"11111110",
  60848=>"00000011",
  60849=>"00000010",
  60850=>"00000010",
  60851=>"11111110",
  60852=>"00000001",
  60853=>"11111110",
  60854=>"11111101",
  60855=>"00000011",
  60856=>"00000011",
  60857=>"00000000",
  60858=>"00000000",
  60859=>"00000011",
  60860=>"00000001",
  60861=>"00000001",
  60862=>"11111111",
  60863=>"00000000",
  60864=>"11111100",
  60865=>"00000101",
  60866=>"00000101",
  60867=>"11111111",
  60868=>"00000001",
  60869=>"00000010",
  60870=>"00000000",
  60871=>"11111101",
  60872=>"11111110",
  60873=>"00000000",
  60874=>"00000011",
  60875=>"00000000",
  60876=>"00000010",
  60877=>"11111110",
  60878=>"00000010",
  60879=>"00000010",
  60880=>"11111111",
  60881=>"00000000",
  60882=>"11111101",
  60883=>"00000001",
  60884=>"00000100",
  60885=>"11111111",
  60886=>"00000001",
  60887=>"00000100",
  60888=>"00000010",
  60889=>"11111100",
  60890=>"00000010",
  60891=>"11111101",
  60892=>"00000011",
  60893=>"11111111",
  60894=>"00000010",
  60895=>"00000001",
  60896=>"11111110",
  60897=>"00000001",
  60898=>"11111111",
  60899=>"00000011",
  60900=>"00000001",
  60901=>"00000000",
  60902=>"11111101",
  60903=>"00000001",
  60904=>"11111111",
  60905=>"00000100",
  60906=>"11111111",
  60907=>"11111100",
  60908=>"11111101",
  60909=>"11111100",
  60910=>"00000010",
  60911=>"00000000",
  60912=>"00000010",
  60913=>"11111100",
  60914=>"11111110",
  60915=>"00000000",
  60916=>"11111110",
  60917=>"00000010",
  60918=>"00000011",
  60919=>"00000011",
  60920=>"00000011",
  60921=>"11111111",
  60922=>"11111101",
  60923=>"11111111",
  60924=>"00000010",
  60925=>"00000010",
  60926=>"11111110",
  60927=>"00000010",
  60928=>"00000000",
  60929=>"00000011",
  60930=>"00000100",
  60931=>"11111100",
  60932=>"11111101",
  60933=>"00000011",
  60934=>"00000100",
  60935=>"00000000",
  60936=>"00000011",
  60937=>"00000000",
  60938=>"00000001",
  60939=>"11111101",
  60940=>"11111110",
  60941=>"00000001",
  60942=>"11111110",
  60943=>"00000111",
  60944=>"00000000",
  60945=>"00000000",
  60946=>"00000000",
  60947=>"00000000",
  60948=>"00000010",
  60949=>"11111101",
  60950=>"11111111",
  60951=>"11111111",
  60952=>"00000000",
  60953=>"11111111",
  60954=>"11111101",
  60955=>"11111111",
  60956=>"00000000",
  60957=>"11111110",
  60958=>"11111111",
  60959=>"00000101",
  60960=>"00000010",
  60961=>"11111111",
  60962=>"11111101",
  60963=>"11111100",
  60964=>"11111100",
  60965=>"11111101",
  60966=>"00000010",
  60967=>"00000001",
  60968=>"00000000",
  60969=>"11111110",
  60970=>"00000100",
  60971=>"11111111",
  60972=>"00000010",
  60973=>"11111111",
  60974=>"11111111",
  60975=>"11111111",
  60976=>"00000100",
  60977=>"11111101",
  60978=>"11111110",
  60979=>"11111111",
  60980=>"11111110",
  60981=>"00000011",
  60982=>"00000001",
  60983=>"00000001",
  60984=>"11111110",
  60985=>"00000010",
  60986=>"00000100",
  60987=>"11111111",
  60988=>"11111111",
  60989=>"11111111",
  60990=>"00000000",
  60991=>"11111101",
  60992=>"00000001",
  60993=>"11111111",
  60994=>"11111110",
  60995=>"00000001",
  60996=>"00000001",
  60997=>"00000010",
  60998=>"11111111",
  60999=>"00000010",
  61000=>"11111110",
  61001=>"11111111",
  61002=>"00000000",
  61003=>"11111111",
  61004=>"00000000",
  61005=>"00000011",
  61006=>"11111111",
  61007=>"00000000",
  61008=>"00000011",
  61009=>"00000001",
  61010=>"00000010",
  61011=>"11111110",
  61012=>"11111110",
  61013=>"00000010",
  61014=>"00000010",
  61015=>"11111101",
  61016=>"00000011",
  61017=>"00000000",
  61018=>"00000011",
  61019=>"11111110",
  61020=>"00000111",
  61021=>"11111110",
  61022=>"00000001",
  61023=>"11111111",
  61024=>"11111111",
  61025=>"00000010",
  61026=>"00000110",
  61027=>"11111100",
  61028=>"00000000",
  61029=>"11111111",
  61030=>"00000010",
  61031=>"00000100",
  61032=>"00000000",
  61033=>"11111110",
  61034=>"11111110",
  61035=>"00000110",
  61036=>"11111110",
  61037=>"00000001",
  61038=>"11111111",
  61039=>"00000011",
  61040=>"11111101",
  61041=>"11111110",
  61042=>"11111101",
  61043=>"00000001",
  61044=>"11111110",
  61045=>"00000010",
  61046=>"00000001",
  61047=>"00000010",
  61048=>"00000011",
  61049=>"11111111",
  61050=>"11111101",
  61051=>"00000001",
  61052=>"00000000",
  61053=>"11111111",
  61054=>"00000110",
  61055=>"00000011",
  61056=>"11111110",
  61057=>"00000010",
  61058=>"00000001",
  61059=>"00000110",
  61060=>"11111100",
  61061=>"00000100",
  61062=>"00000010",
  61063=>"11111111",
  61064=>"11111110",
  61065=>"00000110",
  61066=>"11111111",
  61067=>"11111110",
  61068=>"11111111",
  61069=>"00000001",
  61070=>"11111101",
  61071=>"00000001",
  61072=>"00000100",
  61073=>"11111111",
  61074=>"11111100",
  61075=>"11111101",
  61076=>"00000010",
  61077=>"00000010",
  61078=>"00000010",
  61079=>"11111101",
  61080=>"11111100",
  61081=>"11111110",
  61082=>"00000001",
  61083=>"00000000",
  61084=>"11111111",
  61085=>"00000010",
  61086=>"11111111",
  61087=>"00000001",
  61088=>"00000000",
  61089=>"11111111",
  61090=>"11111111",
  61091=>"00000001",
  61092=>"11111110",
  61093=>"11111110",
  61094=>"11111100",
  61095=>"11111110",
  61096=>"11111101",
  61097=>"11111110",
  61098=>"00000001",
  61099=>"00000011",
  61100=>"11111101",
  61101=>"00000010",
  61102=>"11111111",
  61103=>"00000100",
  61104=>"00000111",
  61105=>"00000000",
  61106=>"00000010",
  61107=>"00000001",
  61108=>"11111110",
  61109=>"00000100",
  61110=>"11111110",
  61111=>"11111101",
  61112=>"00000011",
  61113=>"11111110",
  61114=>"00000000",
  61115=>"11111111",
  61116=>"00000101",
  61117=>"00000011",
  61118=>"11111101",
  61119=>"00000000",
  61120=>"11111110",
  61121=>"00000011",
  61122=>"11111110",
  61123=>"11111110",
  61124=>"00000010",
  61125=>"11111101",
  61126=>"00000001",
  61127=>"11111110",
  61128=>"11111111",
  61129=>"00000000",
  61130=>"00000010",
  61131=>"11111111",
  61132=>"11111110",
  61133=>"11111100",
  61134=>"11111111",
  61135=>"11111100",
  61136=>"00000000",
  61137=>"11111110",
  61138=>"00000011",
  61139=>"00000101",
  61140=>"11111110",
  61141=>"11111101",
  61142=>"00000001",
  61143=>"11111101",
  61144=>"11111110",
  61145=>"11111111",
  61146=>"00000000",
  61147=>"11111101",
  61148=>"00000011",
  61149=>"00000001",
  61150=>"00000010",
  61151=>"00000001",
  61152=>"11111101",
  61153=>"00000001",
  61154=>"11111111",
  61155=>"11111101",
  61156=>"00000011",
  61157=>"11111110",
  61158=>"11111101",
  61159=>"00000000",
  61160=>"00000010",
  61161=>"00000011",
  61162=>"00000101",
  61163=>"00000000",
  61164=>"11111101",
  61165=>"11111111",
  61166=>"00000000",
  61167=>"11111111",
  61168=>"00000000",
  61169=>"00000000",
  61170=>"11111101",
  61171=>"00000010",
  61172=>"00000101",
  61173=>"00000101",
  61174=>"00000001",
  61175=>"00000011",
  61176=>"00000101",
  61177=>"11111111",
  61178=>"11111110",
  61179=>"00000110",
  61180=>"00000010",
  61181=>"00000001",
  61182=>"11111111",
  61183=>"11111110",
  61184=>"00000000",
  61185=>"11111111",
  61186=>"11111110",
  61187=>"00000000",
  61188=>"00000000",
  61189=>"00000000",
  61190=>"11111101",
  61191=>"11111110",
  61192=>"00000011",
  61193=>"00000100",
  61194=>"00000100",
  61195=>"00000000",
  61196=>"11111110",
  61197=>"00000000",
  61198=>"11111110",
  61199=>"00000010",
  61200=>"11111110",
  61201=>"11111111",
  61202=>"00000001",
  61203=>"00000010",
  61204=>"11111101",
  61205=>"11111110",
  61206=>"00000010",
  61207=>"11111101",
  61208=>"00000001",
  61209=>"00000011",
  61210=>"00000101",
  61211=>"00000010",
  61212=>"00000010",
  61213=>"11111101",
  61214=>"00000111",
  61215=>"11111111",
  61216=>"11111111",
  61217=>"11111101",
  61218=>"11111110",
  61219=>"11111111",
  61220=>"00000010",
  61221=>"11111100",
  61222=>"00000000",
  61223=>"00000000",
  61224=>"11111011",
  61225=>"00000000",
  61226=>"11111100",
  61227=>"11111111",
  61228=>"11111101",
  61229=>"11111111",
  61230=>"11111111",
  61231=>"11111110",
  61232=>"00000000",
  61233=>"00000000",
  61234=>"00000010",
  61235=>"00000001",
  61236=>"11111110",
  61237=>"00000000",
  61238=>"00000000",
  61239=>"00000100",
  61240=>"00000000",
  61241=>"00000001",
  61242=>"00000000",
  61243=>"11111100",
  61244=>"00000001",
  61245=>"00000000",
  61246=>"00000001",
  61247=>"11111110",
  61248=>"11111101",
  61249=>"00000010",
  61250=>"00000010",
  61251=>"11111110",
  61252=>"00000001",
  61253=>"11111100",
  61254=>"00000100",
  61255=>"00000000",
  61256=>"00000011",
  61257=>"00000000",
  61258=>"11111110",
  61259=>"00000001",
  61260=>"00000011",
  61261=>"00000000",
  61262=>"11111100",
  61263=>"00000001",
  61264=>"00000100",
  61265=>"11111101",
  61266=>"11111101",
  61267=>"11111100",
  61268=>"00000011",
  61269=>"00000010",
  61270=>"00000011",
  61271=>"11111110",
  61272=>"11111110",
  61273=>"11111111",
  61274=>"11111111",
  61275=>"11111101",
  61276=>"00000000",
  61277=>"00000101",
  61278=>"11111110",
  61279=>"11111101",
  61280=>"00000010",
  61281=>"00000011",
  61282=>"11111111",
  61283=>"11111110",
  61284=>"00000011",
  61285=>"00000100",
  61286=>"00000011",
  61287=>"11111110",
  61288=>"00000000",
  61289=>"11111100",
  61290=>"11111111",
  61291=>"00000010",
  61292=>"11111110",
  61293=>"00000001",
  61294=>"11111100",
  61295=>"11111110",
  61296=>"00000000",
  61297=>"11111111",
  61298=>"11111111",
  61299=>"00000100",
  61300=>"00000100",
  61301=>"11111111",
  61302=>"11111101",
  61303=>"11111111",
  61304=>"00000011",
  61305=>"11111111",
  61306=>"00000000",
  61307=>"00000000",
  61308=>"11111101",
  61309=>"00000001",
  61310=>"11111110",
  61311=>"00000000",
  61312=>"00000000",
  61313=>"00000011",
  61314=>"00000101",
  61315=>"11111111",
  61316=>"00000001",
  61317=>"00000010",
  61318=>"00000010",
  61319=>"11111111",
  61320=>"00000110",
  61321=>"11111110",
  61322=>"00000011",
  61323=>"11111110",
  61324=>"00000000",
  61325=>"11111101",
  61326=>"11111111",
  61327=>"00000100",
  61328=>"11111110",
  61329=>"00000010",
  61330=>"00000101",
  61331=>"11111110",
  61332=>"00000100",
  61333=>"00000111",
  61334=>"00000000",
  61335=>"00000001",
  61336=>"11111110",
  61337=>"11111101",
  61338=>"11111101",
  61339=>"00000001",
  61340=>"00000010",
  61341=>"00000010",
  61342=>"11111101",
  61343=>"11111111",
  61344=>"11111111",
  61345=>"11111111",
  61346=>"00000111",
  61347=>"00000010",
  61348=>"00000011",
  61349=>"00000001",
  61350=>"00000001",
  61351=>"00000011",
  61352=>"11111101",
  61353=>"11111110",
  61354=>"00000010",
  61355=>"00000001",
  61356=>"00000000",
  61357=>"11111110",
  61358=>"11111111",
  61359=>"00000001",
  61360=>"00000000",
  61361=>"11111110",
  61362=>"00000001",
  61363=>"00000001",
  61364=>"11111111",
  61365=>"00000010",
  61366=>"11111111",
  61367=>"11111111",
  61368=>"00000000",
  61369=>"11111111",
  61370=>"11111111",
  61371=>"11111110",
  61372=>"00000011",
  61373=>"00000001",
  61374=>"00000001",
  61375=>"11111110",
  61376=>"00000110",
  61377=>"00000000",
  61378=>"11111110",
  61379=>"00000010",
  61380=>"11111111",
  61381=>"00000000",
  61382=>"00000010",
  61383=>"00000000",
  61384=>"00000001",
  61385=>"11111111",
  61386=>"00000100",
  61387=>"00000010",
  61388=>"11111111",
  61389=>"11111111",
  61390=>"11111111",
  61391=>"00000000",
  61392=>"00000010",
  61393=>"11111101",
  61394=>"00000100",
  61395=>"11111110",
  61396=>"11111111",
  61397=>"11111110",
  61398=>"00000000",
  61399=>"00000011",
  61400=>"00000001",
  61401=>"11111011",
  61402=>"11111110",
  61403=>"00000001",
  61404=>"00000001",
  61405=>"00000010",
  61406=>"00000011",
  61407=>"00000000",
  61408=>"11111111",
  61409=>"11111110",
  61410=>"11111111",
  61411=>"00000000",
  61412=>"00000001",
  61413=>"00000100",
  61414=>"00000001",
  61415=>"11111111",
  61416=>"00000000",
  61417=>"00000011",
  61418=>"11111111",
  61419=>"00000011",
  61420=>"00000000",
  61421=>"00000010",
  61422=>"00000011",
  61423=>"11111101",
  61424=>"00000001",
  61425=>"00000001",
  61426=>"11111101",
  61427=>"11111101",
  61428=>"00000001",
  61429=>"00000110",
  61430=>"00000001",
  61431=>"00000010",
  61432=>"00000010",
  61433=>"00000011",
  61434=>"11111110",
  61435=>"11111110",
  61436=>"00000011",
  61437=>"11111100",
  61438=>"11111101",
  61439=>"00000101",
  61440=>"11111111",
  61441=>"00000000",
  61442=>"11111111",
  61443=>"00000100",
  61444=>"00000000",
  61445=>"00000001",
  61446=>"11111101",
  61447=>"00000010",
  61448=>"00000000",
  61449=>"11111111",
  61450=>"00000000",
  61451=>"00000010",
  61452=>"11111101",
  61453=>"11111101",
  61454=>"00000110",
  61455=>"00000000",
  61456=>"00000001",
  61457=>"11111101",
  61458=>"11111101",
  61459=>"00000101",
  61460=>"00000010",
  61461=>"00000010",
  61462=>"11111101",
  61463=>"00000000",
  61464=>"00000110",
  61465=>"00000000",
  61466=>"11111111",
  61467=>"11111111",
  61468=>"00000000",
  61469=>"11111111",
  61470=>"11111110",
  61471=>"00000011",
  61472=>"00000101",
  61473=>"00000010",
  61474=>"00000001",
  61475=>"11111111",
  61476=>"11111110",
  61477=>"11111011",
  61478=>"11111101",
  61479=>"00000000",
  61480=>"11111110",
  61481=>"11111111",
  61482=>"00000001",
  61483=>"00000000",
  61484=>"00000000",
  61485=>"11111111",
  61486=>"11111111",
  61487=>"11111111",
  61488=>"11111111",
  61489=>"00000000",
  61490=>"00000110",
  61491=>"11111110",
  61492=>"00000000",
  61493=>"11111110",
  61494=>"11111110",
  61495=>"11111111",
  61496=>"00000010",
  61497=>"11111110",
  61498=>"00000011",
  61499=>"11111110",
  61500=>"00000000",
  61501=>"11111110",
  61502=>"11111110",
  61503=>"00000000",
  61504=>"00000011",
  61505=>"11111101",
  61506=>"00000001",
  61507=>"11111110",
  61508=>"11111110",
  61509=>"11111110",
  61510=>"00000001",
  61511=>"00000100",
  61512=>"00000100",
  61513=>"11111111",
  61514=>"00000000",
  61515=>"11111110",
  61516=>"00000000",
  61517=>"00000010",
  61518=>"00000001",
  61519=>"11111101",
  61520=>"11111111",
  61521=>"00000000",
  61522=>"11111111",
  61523=>"00000011",
  61524=>"00000001",
  61525=>"00000000",
  61526=>"00000010",
  61527=>"11111111",
  61528=>"00000001",
  61529=>"00000001",
  61530=>"00000011",
  61531=>"00000000",
  61532=>"11111101",
  61533=>"11111110",
  61534=>"11111100",
  61535=>"11111011",
  61536=>"11111110",
  61537=>"11111100",
  61538=>"11111101",
  61539=>"00000001",
  61540=>"11111101",
  61541=>"11111101",
  61542=>"00000101",
  61543=>"00000000",
  61544=>"00000000",
  61545=>"00000000",
  61546=>"00000001",
  61547=>"11111101",
  61548=>"00000010",
  61549=>"00000000",
  61550=>"11111110",
  61551=>"11111101",
  61552=>"11111101",
  61553=>"00000000",
  61554=>"00000001",
  61555=>"00000100",
  61556=>"11111110",
  61557=>"00000001",
  61558=>"11111110",
  61559=>"11111101",
  61560=>"11111111",
  61561=>"11111101",
  61562=>"00000011",
  61563=>"11111111",
  61564=>"11111101",
  61565=>"00000000",
  61566=>"11111111",
  61567=>"11111111",
  61568=>"00000000",
  61569=>"00000001",
  61570=>"00000100",
  61571=>"00000001",
  61572=>"00000011",
  61573=>"00000000",
  61574=>"00000000",
  61575=>"00000000",
  61576=>"00000010",
  61577=>"11111110",
  61578=>"00000001",
  61579=>"00000001",
  61580=>"00000101",
  61581=>"00000010",
  61582=>"00000011",
  61583=>"00000010",
  61584=>"11111111",
  61585=>"11111110",
  61586=>"00000000",
  61587=>"00000001",
  61588=>"11111110",
  61589=>"00000100",
  61590=>"00000010",
  61591=>"00000000",
  61592=>"00000010",
  61593=>"11111111",
  61594=>"11111110",
  61595=>"00000101",
  61596=>"11111110",
  61597=>"00000001",
  61598=>"11111101",
  61599=>"00000100",
  61600=>"00000000",
  61601=>"00000000",
  61602=>"00000000",
  61603=>"11111111",
  61604=>"00000000",
  61605=>"11111101",
  61606=>"00000001",
  61607=>"11111100",
  61608=>"11111110",
  61609=>"11111110",
  61610=>"00000001",
  61611=>"00000100",
  61612=>"00000100",
  61613=>"00000001",
  61614=>"00000011",
  61615=>"11111111",
  61616=>"00000010",
  61617=>"11111101",
  61618=>"11111111",
  61619=>"11111110",
  61620=>"00000101",
  61621=>"00000011",
  61622=>"00000011",
  61623=>"00000110",
  61624=>"11111110",
  61625=>"11111110",
  61626=>"00000000",
  61627=>"00000001",
  61628=>"00000010",
  61629=>"00000010",
  61630=>"11111111",
  61631=>"00000000",
  61632=>"11111111",
  61633=>"11111110",
  61634=>"00000010",
  61635=>"00000100",
  61636=>"11111110",
  61637=>"00000010",
  61638=>"00000101",
  61639=>"11111111",
  61640=>"00000001",
  61641=>"11111111",
  61642=>"00000000",
  61643=>"00000010",
  61644=>"11111100",
  61645=>"11111110",
  61646=>"11111111",
  61647=>"00000010",
  61648=>"11111110",
  61649=>"11111111",
  61650=>"11111110",
  61651=>"11111101",
  61652=>"11111111",
  61653=>"00000100",
  61654=>"11111101",
  61655=>"00000100",
  61656=>"11111110",
  61657=>"00000010",
  61658=>"11111111",
  61659=>"00000110",
  61660=>"00000000",
  61661=>"00000001",
  61662=>"11111111",
  61663=>"11111110",
  61664=>"00000110",
  61665=>"11111111",
  61666=>"00000011",
  61667=>"11111110",
  61668=>"00000111",
  61669=>"00000001",
  61670=>"00000011",
  61671=>"00000011",
  61672=>"11111111",
  61673=>"11111100",
  61674=>"00000010",
  61675=>"11111111",
  61676=>"11111101",
  61677=>"00000011",
  61678=>"00000000",
  61679=>"11111111",
  61680=>"11111110",
  61681=>"11111111",
  61682=>"00000000",
  61683=>"00000001",
  61684=>"00000000",
  61685=>"00000000",
  61686=>"00000000",
  61687=>"00000001",
  61688=>"11111111",
  61689=>"00000100",
  61690=>"00000000",
  61691=>"00000001",
  61692=>"00000101",
  61693=>"00000010",
  61694=>"00000010",
  61695=>"00000011",
  61696=>"11111101",
  61697=>"00000001",
  61698=>"00000100",
  61699=>"00000000",
  61700=>"00000001",
  61701=>"00000001",
  61702=>"00000100",
  61703=>"11111101",
  61704=>"00000001",
  61705=>"00000000",
  61706=>"11111111",
  61707=>"00000010",
  61708=>"11111111",
  61709=>"00000001",
  61710=>"11111110",
  61711=>"00000011",
  61712=>"11111111",
  61713=>"00000000",
  61714=>"00000000",
  61715=>"00000011",
  61716=>"11111101",
  61717=>"11111110",
  61718=>"11111111",
  61719=>"00000000",
  61720=>"00000010",
  61721=>"11111101",
  61722=>"11111111",
  61723=>"00000001",
  61724=>"00000110",
  61725=>"11111110",
  61726=>"00000000",
  61727=>"11111101",
  61728=>"11111110",
  61729=>"00000001",
  61730=>"11111110",
  61731=>"00000001",
  61732=>"00000000",
  61733=>"11111111",
  61734=>"00000000",
  61735=>"00000011",
  61736=>"00000100",
  61737=>"11111111",
  61738=>"00000000",
  61739=>"00000000",
  61740=>"11111101",
  61741=>"00000000",
  61742=>"11111101",
  61743=>"00000000",
  61744=>"11111111",
  61745=>"11111111",
  61746=>"11111110",
  61747=>"00000000",
  61748=>"00000010",
  61749=>"00000001",
  61750=>"11111100",
  61751=>"00000001",
  61752=>"00000011",
  61753=>"11111111",
  61754=>"00000000",
  61755=>"00000001",
  61756=>"00000001",
  61757=>"00000000",
  61758=>"00000100",
  61759=>"00000010",
  61760=>"00000010",
  61761=>"11111110",
  61762=>"00000010",
  61763=>"11111111",
  61764=>"00000000",
  61765=>"00000000",
  61766=>"11111100",
  61767=>"00000000",
  61768=>"00000010",
  61769=>"00000010",
  61770=>"00000100",
  61771=>"00000010",
  61772=>"11111111",
  61773=>"11111110",
  61774=>"11111111",
  61775=>"00000010",
  61776=>"00000010",
  61777=>"00000001",
  61778=>"11111111",
  61779=>"11111110",
  61780=>"11111111",
  61781=>"11111111",
  61782=>"11111101",
  61783=>"11111110",
  61784=>"00000001",
  61785=>"00000000",
  61786=>"11111101",
  61787=>"11111111",
  61788=>"00000001",
  61789=>"00000011",
  61790=>"11111110",
  61791=>"00000001",
  61792=>"11111110",
  61793=>"11111100",
  61794=>"00000100",
  61795=>"00000011",
  61796=>"00000001",
  61797=>"00000010",
  61798=>"11111101",
  61799=>"00000000",
  61800=>"00000001",
  61801=>"11111110",
  61802=>"00000000",
  61803=>"11111101",
  61804=>"11111110",
  61805=>"00000100",
  61806=>"00000010",
  61807=>"00000100",
  61808=>"00000001",
  61809=>"11111111",
  61810=>"00000001",
  61811=>"11111110",
  61812=>"00000001",
  61813=>"11111110",
  61814=>"11111111",
  61815=>"00000000",
  61816=>"00000100",
  61817=>"00000001",
  61818=>"11111101",
  61819=>"00000001",
  61820=>"11111111",
  61821=>"11111110",
  61822=>"11111110",
  61823=>"00000001",
  61824=>"00000001",
  61825=>"00000100",
  61826=>"11111111",
  61827=>"11111111",
  61828=>"00000101",
  61829=>"00000010",
  61830=>"00000011",
  61831=>"00000001",
  61832=>"11111110",
  61833=>"11111101",
  61834=>"00000000",
  61835=>"00000000",
  61836=>"11111110",
  61837=>"00000001",
  61838=>"11111110",
  61839=>"00000001",
  61840=>"00000011",
  61841=>"00000001",
  61842=>"00000010",
  61843=>"00000011",
  61844=>"00000010",
  61845=>"11111111",
  61846=>"11111111",
  61847=>"00000001",
  61848=>"00000010",
  61849=>"00000000",
  61850=>"11111111",
  61851=>"11111110",
  61852=>"00000010",
  61853=>"00000000",
  61854=>"11111110",
  61855=>"11111111",
  61856=>"00000000",
  61857=>"00000001",
  61858=>"00000001",
  61859=>"11111110",
  61860=>"00000000",
  61861=>"00000001",
  61862=>"00000001",
  61863=>"00000001",
  61864=>"00000101",
  61865=>"11111111",
  61866=>"11111011",
  61867=>"11111101",
  61868=>"11111101",
  61869=>"00000001",
  61870=>"00000110",
  61871=>"11111110",
  61872=>"00000001",
  61873=>"00000011",
  61874=>"00000011",
  61875=>"00000011",
  61876=>"11111110",
  61877=>"11111101",
  61878=>"00000000",
  61879=>"11111101",
  61880=>"00000000",
  61881=>"11111110",
  61882=>"11111111",
  61883=>"11111111",
  61884=>"00000001",
  61885=>"11111110",
  61886=>"00000010",
  61887=>"11111110",
  61888=>"11111101",
  61889=>"11111111",
  61890=>"00000000",
  61891=>"11111110",
  61892=>"11111101",
  61893=>"11111110",
  61894=>"11111110",
  61895=>"11111110",
  61896=>"00000000",
  61897=>"11111101",
  61898=>"11111110",
  61899=>"00000010",
  61900=>"00000000",
  61901=>"11111110",
  61902=>"00000000",
  61903=>"00000010",
  61904=>"11111101",
  61905=>"00000001",
  61906=>"11111111",
  61907=>"11111110",
  61908=>"00000000",
  61909=>"11111111",
  61910=>"11111110",
  61911=>"11111110",
  61912=>"11111111",
  61913=>"00000000",
  61914=>"00000000",
  61915=>"00000100",
  61916=>"11111101",
  61917=>"11111101",
  61918=>"11111101",
  61919=>"11111100",
  61920=>"00000001",
  61921=>"00000001",
  61922=>"00000001",
  61923=>"00000001",
  61924=>"00000001",
  61925=>"00000001",
  61926=>"00000111",
  61927=>"00000000",
  61928=>"00000010",
  61929=>"11111110",
  61930=>"11111111",
  61931=>"00000000",
  61932=>"11111111",
  61933=>"11111010",
  61934=>"11111101",
  61935=>"00000001",
  61936=>"00000001",
  61937=>"00000010",
  61938=>"00000001",
  61939=>"00000001",
  61940=>"11111111",
  61941=>"11111110",
  61942=>"11111111",
  61943=>"00000010",
  61944=>"00000001",
  61945=>"00000100",
  61946=>"00000010",
  61947=>"00000001",
  61948=>"11111110",
  61949=>"11111110",
  61950=>"00000101",
  61951=>"00000001",
  61952=>"00000000",
  61953=>"11111111",
  61954=>"00000000",
  61955=>"00000000",
  61956=>"11111110",
  61957=>"00000000",
  61958=>"00000101",
  61959=>"11111100",
  61960=>"00000011",
  61961=>"11111110",
  61962=>"00000000",
  61963=>"11111111",
  61964=>"11111101",
  61965=>"00000000",
  61966=>"00000011",
  61967=>"00000000",
  61968=>"11111101",
  61969=>"00000100",
  61970=>"00000000",
  61971=>"00000000",
  61972=>"00000010",
  61973=>"00000010",
  61974=>"00000001",
  61975=>"00000000",
  61976=>"00000001",
  61977=>"00000001",
  61978=>"11111111",
  61979=>"00000001",
  61980=>"00000010",
  61981=>"00000000",
  61982=>"00000001",
  61983=>"11111110",
  61984=>"00000101",
  61985=>"11111110",
  61986=>"00000001",
  61987=>"00000010",
  61988=>"00000010",
  61989=>"00000100",
  61990=>"00000010",
  61991=>"00000011",
  61992=>"00000100",
  61993=>"00000001",
  61994=>"00000010",
  61995=>"11111100",
  61996=>"11111111",
  61997=>"00000001",
  61998=>"00000100",
  61999=>"00000001",
  62000=>"00000000",
  62001=>"11111100",
  62002=>"11111110",
  62003=>"00000000",
  62004=>"00000110",
  62005=>"00000011",
  62006=>"11111101",
  62007=>"00000001",
  62008=>"00000000",
  62009=>"00000000",
  62010=>"11111111",
  62011=>"11111111",
  62012=>"00000001",
  62013=>"11111100",
  62014=>"00000010",
  62015=>"00000000",
  62016=>"11111101",
  62017=>"11111110",
  62018=>"11111110",
  62019=>"11111101",
  62020=>"00000010",
  62021=>"11111110",
  62022=>"00000010",
  62023=>"00000001",
  62024=>"00000100",
  62025=>"00000001",
  62026=>"00000001",
  62027=>"11111101",
  62028=>"00000000",
  62029=>"00000010",
  62030=>"00000000",
  62031=>"11111110",
  62032=>"00000010",
  62033=>"00000010",
  62034=>"00000000",
  62035=>"00000001",
  62036=>"00000010",
  62037=>"00000001",
  62038=>"11111111",
  62039=>"11111111",
  62040=>"11111110",
  62041=>"00000110",
  62042=>"00000010",
  62043=>"11111101",
  62044=>"11111101",
  62045=>"11111111",
  62046=>"00000000",
  62047=>"11111101",
  62048=>"00000010",
  62049=>"00000000",
  62050=>"11111110",
  62051=>"00000000",
  62052=>"00000100",
  62053=>"11111100",
  62054=>"11111111",
  62055=>"11111111",
  62056=>"00000001",
  62057=>"11111111",
  62058=>"00000010",
  62059=>"11111110",
  62060=>"00000001",
  62061=>"11111111",
  62062=>"11111111",
  62063=>"00000011",
  62064=>"00000000",
  62065=>"00000001",
  62066=>"11111111",
  62067=>"11111110",
  62068=>"11111111",
  62069=>"00000110",
  62070=>"00000000",
  62071=>"00000000",
  62072=>"00000010",
  62073=>"00000000",
  62074=>"00000000",
  62075=>"00000100",
  62076=>"00000000",
  62077=>"11111110",
  62078=>"11111011",
  62079=>"11111111",
  62080=>"00000001",
  62081=>"00000010",
  62082=>"11111100",
  62083=>"00000010",
  62084=>"00000010",
  62085=>"11111111",
  62086=>"00000000",
  62087=>"11111111",
  62088=>"00000001",
  62089=>"11111110",
  62090=>"00000000",
  62091=>"00000000",
  62092=>"00000001",
  62093=>"00000000",
  62094=>"11111111",
  62095=>"11111100",
  62096=>"11111111",
  62097=>"00000001",
  62098=>"11111101",
  62099=>"00000001",
  62100=>"00000001",
  62101=>"00000010",
  62102=>"11111110",
  62103=>"00000011",
  62104=>"11111100",
  62105=>"00000011",
  62106=>"00000001",
  62107=>"00000001",
  62108=>"11111101",
  62109=>"00000011",
  62110=>"11111100",
  62111=>"00000001",
  62112=>"00000000",
  62113=>"11111110",
  62114=>"00000010",
  62115=>"11111101",
  62116=>"00000000",
  62117=>"00000001",
  62118=>"11111111",
  62119=>"11111111",
  62120=>"11111110",
  62121=>"00000100",
  62122=>"00000001",
  62123=>"00000001",
  62124=>"00000000",
  62125=>"11111100",
  62126=>"00000011",
  62127=>"00000000",
  62128=>"00000001",
  62129=>"11111111",
  62130=>"11111111",
  62131=>"00000010",
  62132=>"00000100",
  62133=>"00000010",
  62134=>"00000000",
  62135=>"11111101",
  62136=>"00000001",
  62137=>"11111101",
  62138=>"00000001",
  62139=>"00000010",
  62140=>"00000010",
  62141=>"00000001",
  62142=>"11111111",
  62143=>"00000000",
  62144=>"11111101",
  62145=>"00000011",
  62146=>"00000000",
  62147=>"00000100",
  62148=>"00000010",
  62149=>"00000001",
  62150=>"00000010",
  62151=>"11111101",
  62152=>"00000001",
  62153=>"00000010",
  62154=>"00000011",
  62155=>"11111110",
  62156=>"00000000",
  62157=>"00000011",
  62158=>"00000001",
  62159=>"00000010",
  62160=>"11111110",
  62161=>"11111111",
  62162=>"11111110",
  62163=>"11111101",
  62164=>"00000011",
  62165=>"11111111",
  62166=>"11111110",
  62167=>"00000001",
  62168=>"00000000",
  62169=>"00000001",
  62170=>"11111110",
  62171=>"00000001",
  62172=>"00000010",
  62173=>"00000001",
  62174=>"00000010",
  62175=>"00000001",
  62176=>"00000000",
  62177=>"11111111",
  62178=>"00000001",
  62179=>"11111110",
  62180=>"11111110",
  62181=>"00000001",
  62182=>"00000000",
  62183=>"00000001",
  62184=>"11111110",
  62185=>"00000000",
  62186=>"11111100",
  62187=>"11111100",
  62188=>"00000000",
  62189=>"00000010",
  62190=>"00000001",
  62191=>"00000001",
  62192=>"11111100",
  62193=>"00000000",
  62194=>"00000100",
  62195=>"00000010",
  62196=>"11111110",
  62197=>"11111011",
  62198=>"11111110",
  62199=>"00000010",
  62200=>"00000010",
  62201=>"00000001",
  62202=>"11111110",
  62203=>"00000001",
  62204=>"11111101",
  62205=>"00000011",
  62206=>"00000001",
  62207=>"00000000",
  62208=>"11111101",
  62209=>"11111111",
  62210=>"00000000",
  62211=>"00000001",
  62212=>"00000101",
  62213=>"00000001",
  62214=>"00000000",
  62215=>"11111110",
  62216=>"11111110",
  62217=>"11111111",
  62218=>"11111110",
  62219=>"00000000",
  62220=>"11111101",
  62221=>"00000011",
  62222=>"00000011",
  62223=>"11111110",
  62224=>"00000000",
  62225=>"11111110",
  62226=>"11111101",
  62227=>"00000001",
  62228=>"00000000",
  62229=>"11111111",
  62230=>"11111110",
  62231=>"00000000",
  62232=>"00000011",
  62233=>"00000001",
  62234=>"11111111",
  62235=>"00000010",
  62236=>"00000000",
  62237=>"00000011",
  62238=>"00000001",
  62239=>"00000011",
  62240=>"11111110",
  62241=>"00000100",
  62242=>"11111111",
  62243=>"11111110",
  62244=>"00000000",
  62245=>"00000000",
  62246=>"11111110",
  62247=>"00000000",
  62248=>"00000011",
  62249=>"00000001",
  62250=>"11111110",
  62251=>"11111111",
  62252=>"11111111",
  62253=>"00000010",
  62254=>"11111110",
  62255=>"00000010",
  62256=>"11111111",
  62257=>"11111110",
  62258=>"00000000",
  62259=>"00000000",
  62260=>"00000001",
  62261=>"00000111",
  62262=>"00000011",
  62263=>"11111111",
  62264=>"11111111",
  62265=>"11111101",
  62266=>"00000000",
  62267=>"11111101",
  62268=>"00000001",
  62269=>"00000001",
  62270=>"11111101",
  62271=>"11111101",
  62272=>"11111111",
  62273=>"11111110",
  62274=>"11111101",
  62275=>"00000010",
  62276=>"11111111",
  62277=>"00000001",
  62278=>"11111110",
  62279=>"00000010",
  62280=>"11111110",
  62281=>"00000001",
  62282=>"11111101",
  62283=>"11111111",
  62284=>"00000001",
  62285=>"11111110",
  62286=>"00000000",
  62287=>"00000010",
  62288=>"00000001",
  62289=>"00000010",
  62290=>"00000000",
  62291=>"11111111",
  62292=>"00000001",
  62293=>"11111111",
  62294=>"00000001",
  62295=>"00000000",
  62296=>"11111110",
  62297=>"11111110",
  62298=>"00000001",
  62299=>"11111110",
  62300=>"00000100",
  62301=>"00000001",
  62302=>"00000000",
  62303=>"11111111",
  62304=>"11111111",
  62305=>"11111111",
  62306=>"00000111",
  62307=>"11111101",
  62308=>"00000100",
  62309=>"11111110",
  62310=>"11111111",
  62311=>"11111111",
  62312=>"00000101",
  62313=>"11111110",
  62314=>"00000000",
  62315=>"11111111",
  62316=>"00000000",
  62317=>"00000001",
  62318=>"11111101",
  62319=>"11111101",
  62320=>"00000010",
  62321=>"11111111",
  62322=>"00000000",
  62323=>"00000010",
  62324=>"00000001",
  62325=>"11111110",
  62326=>"00000000",
  62327=>"11111101",
  62328=>"11111101",
  62329=>"00000010",
  62330=>"11111101",
  62331=>"11111100",
  62332=>"11111111",
  62333=>"00000010",
  62334=>"11111110",
  62335=>"00000010",
  62336=>"00000010",
  62337=>"11111101",
  62338=>"11111111",
  62339=>"00000010",
  62340=>"00000000",
  62341=>"00000000",
  62342=>"00000010",
  62343=>"11111110",
  62344=>"11111111",
  62345=>"11111111",
  62346=>"00000001",
  62347=>"11111101",
  62348=>"00000001",
  62349=>"00000010",
  62350=>"11111110",
  62351=>"11111111",
  62352=>"11111110",
  62353=>"00000001",
  62354=>"11111100",
  62355=>"00000100",
  62356=>"00000011",
  62357=>"11111110",
  62358=>"00000110",
  62359=>"00000010",
  62360=>"00000110",
  62361=>"11111111",
  62362=>"00000011",
  62363=>"11111110",
  62364=>"00000001",
  62365=>"11111110",
  62366=>"00000100",
  62367=>"00000000",
  62368=>"11111111",
  62369=>"00000000",
  62370=>"11111110",
  62371=>"00000001",
  62372=>"00000010",
  62373=>"00000001",
  62374=>"11111110",
  62375=>"00000000",
  62376=>"00000101",
  62377=>"00000011",
  62378=>"00000011",
  62379=>"00000000",
  62380=>"00000001",
  62381=>"00000010",
  62382=>"00000001",
  62383=>"11111110",
  62384=>"00000000",
  62385=>"00000100",
  62386=>"11111100",
  62387=>"11111110",
  62388=>"11111101",
  62389=>"11111110",
  62390=>"11111110",
  62391=>"11111100",
  62392=>"11111111",
  62393=>"11111110",
  62394=>"00000000",
  62395=>"00000011",
  62396=>"11111111",
  62397=>"11111101",
  62398=>"11111111",
  62399=>"00000001",
  62400=>"11111111",
  62401=>"00000011",
  62402=>"00000001",
  62403=>"00000000",
  62404=>"00000000",
  62405=>"00000100",
  62406=>"11111100",
  62407=>"11111111",
  62408=>"00000101",
  62409=>"00000100",
  62410=>"00000000",
  62411=>"00000101",
  62412=>"00000001",
  62413=>"00000010",
  62414=>"00000010",
  62415=>"11111100",
  62416=>"00000000",
  62417=>"00000010",
  62418=>"11111101",
  62419=>"00000001",
  62420=>"00000010",
  62421=>"11111111",
  62422=>"00000110",
  62423=>"11111101",
  62424=>"00000001",
  62425=>"11111111",
  62426=>"11111101",
  62427=>"00000110",
  62428=>"00000001",
  62429=>"11111111",
  62430=>"00000010",
  62431=>"11111101",
  62432=>"00000000",
  62433=>"00000001",
  62434=>"00000000",
  62435=>"00000001",
  62436=>"00000001",
  62437=>"00000001",
  62438=>"00000011",
  62439=>"11111101",
  62440=>"00000000",
  62441=>"00000001",
  62442=>"11111101",
  62443=>"00000011",
  62444=>"11111111",
  62445=>"00000001",
  62446=>"00000000",
  62447=>"00000010",
  62448=>"00000011",
  62449=>"11111101",
  62450=>"00000000",
  62451=>"11111111",
  62452=>"00000010",
  62453=>"00000000",
  62454=>"00000001",
  62455=>"11111101",
  62456=>"00000100",
  62457=>"00000010",
  62458=>"11111110",
  62459=>"11111111",
  62460=>"11111011",
  62461=>"00000010",
  62462=>"11111110",
  62463=>"00000001",
  62464=>"00000000",
  62465=>"00000001",
  62466=>"11111110",
  62467=>"00000010",
  62468=>"11111111",
  62469=>"00000000",
  62470=>"11111110",
  62471=>"00000001",
  62472=>"00000111",
  62473=>"11111110",
  62474=>"00000001",
  62475=>"11111110",
  62476=>"00000010",
  62477=>"00000000",
  62478=>"11111101",
  62479=>"00000001",
  62480=>"11111111",
  62481=>"00000011",
  62482=>"11111110",
  62483=>"11111110",
  62484=>"11111111",
  62485=>"00000010",
  62486=>"11111111",
  62487=>"00000011",
  62488=>"00000000",
  62489=>"00000001",
  62490=>"11111101",
  62491=>"00000001",
  62492=>"00000001",
  62493=>"11111111",
  62494=>"11111110",
  62495=>"11111110",
  62496=>"11111110",
  62497=>"11111111",
  62498=>"00000010",
  62499=>"00000000",
  62500=>"00000001",
  62501=>"00000001",
  62502=>"11111101",
  62503=>"00000010",
  62504=>"00000001",
  62505=>"00000011",
  62506=>"00000011",
  62507=>"00000001",
  62508=>"11111101",
  62509=>"00000010",
  62510=>"11111111",
  62511=>"00000001",
  62512=>"00000001",
  62513=>"00000000",
  62514=>"00000101",
  62515=>"11111100",
  62516=>"11111110",
  62517=>"11111111",
  62518=>"00000010",
  62519=>"00000001",
  62520=>"00000011",
  62521=>"11111110",
  62522=>"00000001",
  62523=>"11111111",
  62524=>"00000000",
  62525=>"00000011",
  62526=>"00000100",
  62527=>"11111111",
  62528=>"11111111",
  62529=>"11111111",
  62530=>"00000010",
  62531=>"00000010",
  62532=>"11111110",
  62533=>"11111110",
  62534=>"11111111",
  62535=>"00000011",
  62536=>"00000011",
  62537=>"11111111",
  62538=>"00000001",
  62539=>"11111110",
  62540=>"11111101",
  62541=>"00000100",
  62542=>"00000011",
  62543=>"00000011",
  62544=>"00000000",
  62545=>"00000010",
  62546=>"00000010",
  62547=>"00000001",
  62548=>"11111110",
  62549=>"00000010",
  62550=>"00000000",
  62551=>"11111110",
  62552=>"00000010",
  62553=>"11111101",
  62554=>"00000010",
  62555=>"11111110",
  62556=>"00000001",
  62557=>"11111111",
  62558=>"00000010",
  62559=>"11111101",
  62560=>"00000000",
  62561=>"00000100",
  62562=>"11111110",
  62563=>"00000011",
  62564=>"00000010",
  62565=>"00000010",
  62566=>"00000100",
  62567=>"00000011",
  62568=>"00000010",
  62569=>"11111111",
  62570=>"00000011",
  62571=>"11111101",
  62572=>"11111110",
  62573=>"00000010",
  62574=>"11111110",
  62575=>"00000010",
  62576=>"00000000",
  62577=>"00000010",
  62578=>"00000000",
  62579=>"00000010",
  62580=>"00000010",
  62581=>"11111100",
  62582=>"00000010",
  62583=>"00000001",
  62584=>"11111111",
  62585=>"00000000",
  62586=>"11111101",
  62587=>"00000100",
  62588=>"00000000",
  62589=>"00000011",
  62590=>"11111110",
  62591=>"11111110",
  62592=>"00000000",
  62593=>"00000000",
  62594=>"00000010",
  62595=>"00000010",
  62596=>"00000101",
  62597=>"00000000",
  62598=>"11111111",
  62599=>"00000011",
  62600=>"00000110",
  62601=>"11111110",
  62602=>"00000110",
  62603=>"11111111",
  62604=>"11111110",
  62605=>"11111110",
  62606=>"11111110",
  62607=>"00000001",
  62608=>"00000011",
  62609=>"00000001",
  62610=>"00000000",
  62611=>"00000001",
  62612=>"00000000",
  62613=>"11111111",
  62614=>"11111111",
  62615=>"00000001",
  62616=>"00000000",
  62617=>"00000000",
  62618=>"00000000",
  62619=>"11111110",
  62620=>"00000000",
  62621=>"00000001",
  62622=>"11111111",
  62623=>"00000001",
  62624=>"00000001",
  62625=>"11111110",
  62626=>"00000000",
  62627=>"00000011",
  62628=>"00000001",
  62629=>"00000011",
  62630=>"00000000",
  62631=>"00000001",
  62632=>"11111110",
  62633=>"00000001",
  62634=>"00000001",
  62635=>"11111111",
  62636=>"00000000",
  62637=>"00000010",
  62638=>"11111110",
  62639=>"00000000",
  62640=>"11111111",
  62641=>"00000000",
  62642=>"11111110",
  62643=>"00000100",
  62644=>"00000001",
  62645=>"00000011",
  62646=>"00000000",
  62647=>"11111111",
  62648=>"11111110",
  62649=>"11111101",
  62650=>"00000001",
  62651=>"00000010",
  62652=>"00000001",
  62653=>"00000010",
  62654=>"00000001",
  62655=>"11111111",
  62656=>"11111101",
  62657=>"00000011",
  62658=>"11111110",
  62659=>"00000001",
  62660=>"00000010",
  62661=>"00000001",
  62662=>"11111110",
  62663=>"00000001",
  62664=>"11111110",
  62665=>"11111110",
  62666=>"11111110",
  62667=>"00000100",
  62668=>"11111100",
  62669=>"11111111",
  62670=>"11111111",
  62671=>"00000000",
  62672=>"00000010",
  62673=>"00000000",
  62674=>"00000000",
  62675=>"00000010",
  62676=>"00000000",
  62677=>"00000010",
  62678=>"11111101",
  62679=>"00000001",
  62680=>"00000110",
  62681=>"00000001",
  62682=>"00000000",
  62683=>"00000000",
  62684=>"00000100",
  62685=>"11111101",
  62686=>"11111110",
  62687=>"00000010",
  62688=>"11111101",
  62689=>"11111111",
  62690=>"00000000",
  62691=>"00000001",
  62692=>"11111110",
  62693=>"00000100",
  62694=>"00000000",
  62695=>"00000000",
  62696=>"11111110",
  62697=>"00000010",
  62698=>"00000000",
  62699=>"11111111",
  62700=>"11111110",
  62701=>"00000011",
  62702=>"00000010",
  62703=>"00000011",
  62704=>"11111111",
  62705=>"00000000",
  62706=>"00000001",
  62707=>"00000010",
  62708=>"11111110",
  62709=>"00000001",
  62710=>"11111111",
  62711=>"11111101",
  62712=>"11111111",
  62713=>"11111101",
  62714=>"00000010",
  62715=>"11111111",
  62716=>"11111100",
  62717=>"00000010",
  62718=>"11111101",
  62719=>"11111111",
  62720=>"11111111",
  62721=>"00000001",
  62722=>"00000001",
  62723=>"11111111",
  62724=>"00000001",
  62725=>"00000000",
  62726=>"00000010",
  62727=>"00000010",
  62728=>"11111111",
  62729=>"00000110",
  62730=>"11111101",
  62731=>"11111111",
  62732=>"00000001",
  62733=>"00000011",
  62734=>"11111111",
  62735=>"00000001",
  62736=>"11111111",
  62737=>"00000010",
  62738=>"00000000",
  62739=>"11111111",
  62740=>"00000010",
  62741=>"11111110",
  62742=>"00000001",
  62743=>"11111111",
  62744=>"11111110",
  62745=>"00000000",
  62746=>"00000001",
  62747=>"11111111",
  62748=>"11111101",
  62749=>"00000001",
  62750=>"11111111",
  62751=>"11111111",
  62752=>"11111110",
  62753=>"11111111",
  62754=>"00000010",
  62755=>"00000001",
  62756=>"00000100",
  62757=>"11111111",
  62758=>"11111111",
  62759=>"11111101",
  62760=>"11111111",
  62761=>"00000000",
  62762=>"00000001",
  62763=>"00000011",
  62764=>"00000001",
  62765=>"00000010",
  62766=>"00000011",
  62767=>"00000010",
  62768=>"00000010",
  62769=>"00000001",
  62770=>"11111100",
  62771=>"00000000",
  62772=>"00000011",
  62773=>"00000000",
  62774=>"00000010",
  62775=>"11111110",
  62776=>"00000011",
  62777=>"00000010",
  62778=>"00000000",
  62779=>"11111101",
  62780=>"11111111",
  62781=>"00000011",
  62782=>"00000001",
  62783=>"00000001",
  62784=>"11111110",
  62785=>"11111111",
  62786=>"11111110",
  62787=>"00000011",
  62788=>"00000001",
  62789=>"00000100",
  62790=>"11111100",
  62791=>"11111101",
  62792=>"11111101",
  62793=>"00000001",
  62794=>"00000101",
  62795=>"00000000",
  62796=>"11111111",
  62797=>"00000010",
  62798=>"11111110",
  62799=>"11111110",
  62800=>"11111111",
  62801=>"11111111",
  62802=>"00000011",
  62803=>"11111110",
  62804=>"00000101",
  62805=>"00000011",
  62806=>"00000000",
  62807=>"00000010",
  62808=>"11111111",
  62809=>"00000010",
  62810=>"11111101",
  62811=>"00000001",
  62812=>"00000010",
  62813=>"00000001",
  62814=>"11111111",
  62815=>"00000010",
  62816=>"00000011",
  62817=>"11111111",
  62818=>"00000010",
  62819=>"00000000",
  62820=>"11111110",
  62821=>"00000011",
  62822=>"11111110",
  62823=>"11111111",
  62824=>"00000000",
  62825=>"00000000",
  62826=>"00000001",
  62827=>"00000011",
  62828=>"00000000",
  62829=>"00000101",
  62830=>"11111101",
  62831=>"00000011",
  62832=>"11111111",
  62833=>"00000001",
  62834=>"11111110",
  62835=>"11111110",
  62836=>"00000001",
  62837=>"00000001",
  62838=>"11111101",
  62839=>"11111110",
  62840=>"00000000",
  62841=>"11111101",
  62842=>"00000011",
  62843=>"11111101",
  62844=>"00000001",
  62845=>"11111110",
  62846=>"00000011",
  62847=>"00000001",
  62848=>"00000010",
  62849=>"00000010",
  62850=>"11111110",
  62851=>"00000010",
  62852=>"00000000",
  62853=>"00000000",
  62854=>"11111101",
  62855=>"00000100",
  62856=>"11111110",
  62857=>"00000011",
  62858=>"00000010",
  62859=>"00000001",
  62860=>"00000010",
  62861=>"00000010",
  62862=>"00000010",
  62863=>"11111110",
  62864=>"00000010",
  62865=>"00000001",
  62866=>"11111110",
  62867=>"11111111",
  62868=>"11111111",
  62869=>"11111110",
  62870=>"00000000",
  62871=>"00000100",
  62872=>"11111111",
  62873=>"00000000",
  62874=>"11111110",
  62875=>"11111101",
  62876=>"00000001",
  62877=>"11111101",
  62878=>"00000001",
  62879=>"11111110",
  62880=>"00000000",
  62881=>"00000010",
  62882=>"11111110",
  62883=>"11111110",
  62884=>"11111111",
  62885=>"11111111",
  62886=>"11111110",
  62887=>"00000000",
  62888=>"00000010",
  62889=>"11111101",
  62890=>"11111110",
  62891=>"00000001",
  62892=>"00000100",
  62893=>"00000001",
  62894=>"00000010",
  62895=>"00000010",
  62896=>"11111111",
  62897=>"00000011",
  62898=>"11111110",
  62899=>"00000011",
  62900=>"11111101",
  62901=>"00000000",
  62902=>"00000010",
  62903=>"00000000",
  62904=>"11111101",
  62905=>"00000101",
  62906=>"00000000",
  62907=>"00000011",
  62908=>"00000011",
  62909=>"11111100",
  62910=>"11111110",
  62911=>"00000010",
  62912=>"00000110",
  62913=>"11111110",
  62914=>"00000011",
  62915=>"11111100",
  62916=>"00000001",
  62917=>"11111110",
  62918=>"00000001",
  62919=>"11111110",
  62920=>"11111111",
  62921=>"00000010",
  62922=>"11111110",
  62923=>"11111111",
  62924=>"00000010",
  62925=>"00000001",
  62926=>"00000011",
  62927=>"11111101",
  62928=>"00000001",
  62929=>"11111111",
  62930=>"11111100",
  62931=>"00000000",
  62932=>"00000100",
  62933=>"00000010",
  62934=>"11111101",
  62935=>"11111101",
  62936=>"00000010",
  62937=>"11111111",
  62938=>"00000011",
  62939=>"00000001",
  62940=>"00000001",
  62941=>"11111110",
  62942=>"00000000",
  62943=>"11111110",
  62944=>"11111111",
  62945=>"11111111",
  62946=>"11111111",
  62947=>"00000010",
  62948=>"00000001",
  62949=>"11111101",
  62950=>"11111110",
  62951=>"00000010",
  62952=>"00000011",
  62953=>"11111111",
  62954=>"00000101",
  62955=>"00000001",
  62956=>"00000001",
  62957=>"00000101",
  62958=>"00000010",
  62959=>"11111111",
  62960=>"11111110",
  62961=>"00000001",
  62962=>"11111101",
  62963=>"11111101",
  62964=>"00000010",
  62965=>"11111110",
  62966=>"11111110",
  62967=>"11111111",
  62968=>"00000000",
  62969=>"11111110",
  62970=>"11111111",
  62971=>"00000011",
  62972=>"11111110",
  62973=>"00000000",
  62974=>"11111110",
  62975=>"00000001",
  62976=>"00000010",
  62977=>"11111111",
  62978=>"11111110",
  62979=>"00000000",
  62980=>"11111111",
  62981=>"00000010",
  62982=>"00000100",
  62983=>"11111110",
  62984=>"00000011",
  62985=>"00000010",
  62986=>"00000011",
  62987=>"00000010",
  62988=>"00000010",
  62989=>"00000010",
  62990=>"11111110",
  62991=>"00000011",
  62992=>"00000000",
  62993=>"11111110",
  62994=>"00000010",
  62995=>"11111100",
  62996=>"11111111",
  62997=>"11111110",
  62998=>"00000000",
  62999=>"00000000",
  63000=>"11111110",
  63001=>"11111111",
  63002=>"00000000",
  63003=>"11111111",
  63004=>"11111110",
  63005=>"00000001",
  63006=>"00000000",
  63007=>"00000101",
  63008=>"11111111",
  63009=>"00000001",
  63010=>"11111101",
  63011=>"11111111",
  63012=>"00000001",
  63013=>"11111100",
  63014=>"00000010",
  63015=>"00000000",
  63016=>"00000100",
  63017=>"00000001",
  63018=>"11111101",
  63019=>"00000011",
  63020=>"11111111",
  63021=>"11111110",
  63022=>"00000001",
  63023=>"00000011",
  63024=>"00000001",
  63025=>"00000010",
  63026=>"00000011",
  63027=>"00000000",
  63028=>"00000001",
  63029=>"11111111",
  63030=>"11111110",
  63031=>"00000011",
  63032=>"00000100",
  63033=>"00000010",
  63034=>"00000000",
  63035=>"11111101",
  63036=>"00000000",
  63037=>"00000000",
  63038=>"11111101",
  63039=>"00000001",
  63040=>"11111111",
  63041=>"11111110",
  63042=>"00000011",
  63043=>"00000010",
  63044=>"00000000",
  63045=>"00000101",
  63046=>"00000101",
  63047=>"00000000",
  63048=>"00000000",
  63049=>"00000011",
  63050=>"11111101",
  63051=>"00000010",
  63052=>"11111110",
  63053=>"00000110",
  63054=>"00000100",
  63055=>"00000001",
  63056=>"00000000",
  63057=>"00000000",
  63058=>"11111110",
  63059=>"11111110",
  63060=>"11111101",
  63061=>"11111111",
  63062=>"11111111",
  63063=>"11111101",
  63064=>"11111110",
  63065=>"00000000",
  63066=>"11111111",
  63067=>"00000011",
  63068=>"11111111",
  63069=>"11111111",
  63070=>"11111110",
  63071=>"11111111",
  63072=>"11111111",
  63073=>"11111111",
  63074=>"11111111",
  63075=>"00000011",
  63076=>"11111101",
  63077=>"11111101",
  63078=>"00000100",
  63079=>"00000000",
  63080=>"11111111",
  63081=>"11111100",
  63082=>"00000000",
  63083=>"00000000",
  63084=>"00000010",
  63085=>"11111111",
  63086=>"00000011",
  63087=>"11111111",
  63088=>"00000010",
  63089=>"11111101",
  63090=>"00000001",
  63091=>"11111111",
  63092=>"00000000",
  63093=>"00000011",
  63094=>"11111111",
  63095=>"00000000",
  63096=>"11111111",
  63097=>"11111111",
  63098=>"11111111",
  63099=>"00000000",
  63100=>"00000001",
  63101=>"00000010",
  63102=>"11111101",
  63103=>"00000010",
  63104=>"00000011",
  63105=>"11111111",
  63106=>"00000000",
  63107=>"00000101",
  63108=>"00000001",
  63109=>"11111111",
  63110=>"11111111",
  63111=>"11111111",
  63112=>"00000000",
  63113=>"00000011",
  63114=>"00000010",
  63115=>"11111111",
  63116=>"11111110",
  63117=>"00000001",
  63118=>"00000010",
  63119=>"11111110",
  63120=>"00000000",
  63121=>"11111101",
  63122=>"11111101",
  63123=>"11111110",
  63124=>"00000000",
  63125=>"00000000",
  63126=>"00000000",
  63127=>"11111100",
  63128=>"11111111",
  63129=>"11111100",
  63130=>"00000001",
  63131=>"11111111",
  63132=>"00000001",
  63133=>"11111110",
  63134=>"11111101",
  63135=>"00000001",
  63136=>"00000000",
  63137=>"00000001",
  63138=>"11111111",
  63139=>"00000001",
  63140=>"11111110",
  63141=>"00000010",
  63142=>"00000001",
  63143=>"00000000",
  63144=>"00000011",
  63145=>"11111101",
  63146=>"00000001",
  63147=>"00000001",
  63148=>"00000011",
  63149=>"11111111",
  63150=>"00000100",
  63151=>"00000000",
  63152=>"00000000",
  63153=>"11111101",
  63154=>"00000000",
  63155=>"11111111",
  63156=>"00000000",
  63157=>"11111110",
  63158=>"11111111",
  63159=>"11111110",
  63160=>"11111110",
  63161=>"11111110",
  63162=>"11111111",
  63163=>"00000001",
  63164=>"11111111",
  63165=>"11111111",
  63166=>"11111110",
  63167=>"00000011",
  63168=>"00000011",
  63169=>"00000001",
  63170=>"11111110",
  63171=>"11111101",
  63172=>"11111111",
  63173=>"00000010",
  63174=>"00000000",
  63175=>"11111101",
  63176=>"00000011",
  63177=>"11111111",
  63178=>"00000100",
  63179=>"00000010",
  63180=>"00000001",
  63181=>"00000010",
  63182=>"11111110",
  63183=>"11111101",
  63184=>"00000011",
  63185=>"00000001",
  63186=>"11111111",
  63187=>"11111111",
  63188=>"00000100",
  63189=>"00000001",
  63190=>"00000001",
  63191=>"00000001",
  63192=>"11111101",
  63193=>"00000001",
  63194=>"00000000",
  63195=>"11111110",
  63196=>"11111110",
  63197=>"00000010",
  63198=>"11111110",
  63199=>"11111110",
  63200=>"00000000",
  63201=>"11111111",
  63202=>"11111111",
  63203=>"00000011",
  63204=>"11111101",
  63205=>"00000010",
  63206=>"11111110",
  63207=>"00000001",
  63208=>"11111101",
  63209=>"00000011",
  63210=>"00000000",
  63211=>"00000000",
  63212=>"00000001",
  63213=>"00000010",
  63214=>"00000000",
  63215=>"00000000",
  63216=>"11111111",
  63217=>"11111101",
  63218=>"11111101",
  63219=>"11111101",
  63220=>"00000011",
  63221=>"00000000",
  63222=>"00000001",
  63223=>"00000010",
  63224=>"00000001",
  63225=>"11111111",
  63226=>"11111110",
  63227=>"00000001",
  63228=>"11111110",
  63229=>"11111101",
  63230=>"11111111",
  63231=>"00000001",
  63232=>"11111111",
  63233=>"11111111",
  63234=>"00000000",
  63235=>"11111111",
  63236=>"11111111",
  63237=>"00000001",
  63238=>"11111111",
  63239=>"11111111",
  63240=>"00000000",
  63241=>"11111110",
  63242=>"11111110",
  63243=>"11111110",
  63244=>"00000010",
  63245=>"00000010",
  63246=>"11111110",
  63247=>"11111110",
  63248=>"00000010",
  63249=>"11111110",
  63250=>"11111111",
  63251=>"00000001",
  63252=>"00000010",
  63253=>"11111101",
  63254=>"11111110",
  63255=>"11111111",
  63256=>"11111111",
  63257=>"11111110",
  63258=>"11111100",
  63259=>"00000010",
  63260=>"00000000",
  63261=>"11111110",
  63262=>"11111111",
  63263=>"00000001",
  63264=>"00000011",
  63265=>"00000010",
  63266=>"11111111",
  63267=>"00000011",
  63268=>"11111111",
  63269=>"11111111",
  63270=>"11111110",
  63271=>"00000010",
  63272=>"00000000",
  63273=>"11111110",
  63274=>"11111101",
  63275=>"00000000",
  63276=>"11111101",
  63277=>"11111111",
  63278=>"00000010",
  63279=>"00000011",
  63280=>"11111110",
  63281=>"00000011",
  63282=>"11111110",
  63283=>"00000110",
  63284=>"00000100",
  63285=>"00000000",
  63286=>"11111111",
  63287=>"11111111",
  63288=>"00000100",
  63289=>"00000000",
  63290=>"00000010",
  63291=>"00000000",
  63292=>"00000000",
  63293=>"00000011",
  63294=>"11111110",
  63295=>"11111110",
  63296=>"00000010",
  63297=>"11111111",
  63298=>"11111110",
  63299=>"00000101",
  63300=>"00000011",
  63301=>"11111111",
  63302=>"00000000",
  63303=>"00000011",
  63304=>"00000100",
  63305=>"00000010",
  63306=>"11111110",
  63307=>"00000011",
  63308=>"11111101",
  63309=>"00000010",
  63310=>"00000010",
  63311=>"11111110",
  63312=>"00000010",
  63313=>"11111110",
  63314=>"11111111",
  63315=>"00000001",
  63316=>"00000010",
  63317=>"00000000",
  63318=>"11111110",
  63319=>"00000010",
  63320=>"00000001",
  63321=>"00000100",
  63322=>"11111101",
  63323=>"00000000",
  63324=>"00000010",
  63325=>"11111111",
  63326=>"00000001",
  63327=>"00000000",
  63328=>"00000010",
  63329=>"00000010",
  63330=>"11111111",
  63331=>"00000001",
  63332=>"00000000",
  63333=>"11111111",
  63334=>"11111111",
  63335=>"11111111",
  63336=>"11111101",
  63337=>"11111110",
  63338=>"11111111",
  63339=>"11111110",
  63340=>"11111110",
  63341=>"11111101",
  63342=>"11111111",
  63343=>"00000011",
  63344=>"11111111",
  63345=>"00000000",
  63346=>"00000000",
  63347=>"11111110",
  63348=>"11111110",
  63349=>"00000010",
  63350=>"00000011",
  63351=>"00000011",
  63352=>"00000010",
  63353=>"11111101",
  63354=>"11111111",
  63355=>"00000000",
  63356=>"11111110",
  63357=>"11111110",
  63358=>"00000010",
  63359=>"11111100",
  63360=>"11111110",
  63361=>"11111110",
  63362=>"00000001",
  63363=>"00000001",
  63364=>"00000001",
  63365=>"11111101",
  63366=>"00000011",
  63367=>"00000001",
  63368=>"00000000",
  63369=>"00000000",
  63370=>"00000010",
  63371=>"11111111",
  63372=>"00000001",
  63373=>"11111110",
  63374=>"00000000",
  63375=>"11111101",
  63376=>"00000001",
  63377=>"11111101",
  63378=>"11111110",
  63379=>"00000001",
  63380=>"00000010",
  63381=>"11111111",
  63382=>"00000000",
  63383=>"00000000",
  63384=>"11111111",
  63385=>"11111110",
  63386=>"00000010",
  63387=>"00000000",
  63388=>"11111101",
  63389=>"00000001",
  63390=>"00000000",
  63391=>"11111111",
  63392=>"11111110",
  63393=>"11111111",
  63394=>"00000001",
  63395=>"00000010",
  63396=>"00000000",
  63397=>"00000010",
  63398=>"11111111",
  63399=>"00000010",
  63400=>"11111110",
  63401=>"11111101",
  63402=>"11111110",
  63403=>"00000011",
  63404=>"11111101",
  63405=>"00000100",
  63406=>"00000010",
  63407=>"00000010",
  63408=>"00000101",
  63409=>"11111111",
  63410=>"00000000",
  63411=>"00000001",
  63412=>"11111111",
  63413=>"11111110",
  63414=>"11111110",
  63415=>"11111111",
  63416=>"11111111",
  63417=>"00000010",
  63418=>"00000010",
  63419=>"00000001",
  63420=>"00000001",
  63421=>"00000000",
  63422=>"00000010",
  63423=>"00000011",
  63424=>"00000011",
  63425=>"00000001",
  63426=>"00000000",
  63427=>"11111101",
  63428=>"00000000",
  63429=>"11111110",
  63430=>"00000011",
  63431=>"00000010",
  63432=>"11111110",
  63433=>"11111111",
  63434=>"00000001",
  63435=>"11111111",
  63436=>"11111110",
  63437=>"00000001",
  63438=>"00000011",
  63439=>"11111111",
  63440=>"00000010",
  63441=>"00000000",
  63442=>"00000100",
  63443=>"00000000",
  63444=>"00000001",
  63445=>"11111101",
  63446=>"00000001",
  63447=>"00000101",
  63448=>"00000011",
  63449=>"00000001",
  63450=>"00000000",
  63451=>"11111111",
  63452=>"11111110",
  63453=>"11111111",
  63454=>"00000001",
  63455=>"00000010",
  63456=>"11111101",
  63457=>"11111101",
  63458=>"11111101",
  63459=>"00000000",
  63460=>"11111110",
  63461=>"11111101",
  63462=>"11111101",
  63463=>"11111110",
  63464=>"11111111",
  63465=>"00000010",
  63466=>"11111111",
  63467=>"00000001",
  63468=>"11111111",
  63469=>"11111111",
  63470=>"00000011",
  63471=>"11111111",
  63472=>"00000001",
  63473=>"00000011",
  63474=>"00000000",
  63475=>"00000001",
  63476=>"00000011",
  63477=>"00000001",
  63478=>"00000000",
  63479=>"00000011",
  63480=>"00000101",
  63481=>"00000011",
  63482=>"11111111",
  63483=>"11111110",
  63484=>"11111110",
  63485=>"00000000",
  63486=>"11111111",
  63487=>"00000001",
  63488=>"00000000",
  63489=>"00000000",
  63490=>"00000000",
  63491=>"00000000",
  63492=>"00000000",
  63493=>"00000000",
  63494=>"00000000",
  63495=>"00000000",
  63496=>"00000000",
  63497=>"00000000",
  63498=>"00000000",
  63499=>"00000000",
  63500=>"00000000",
  63501=>"00000000",
  63502=>"00000000",
  63503=>"00000000",
  63504=>"00000000",
  63505=>"00000000",
  63506=>"00000000",
  63507=>"00000000",
  63508=>"00000000",
  63509=>"00000000",
  63510=>"00000000",
  63511=>"00000000",
  63512=>"00000000",
  63513=>"00000000",
  63514=>"00000000",
  63515=>"00000000",
  63516=>"00000000",
  63517=>"00000000",
  63518=>"00000000",
  63519=>"00000000",
  63520=>"00000000",
  63521=>"00000000",
  63522=>"00000000",
  63523=>"00000000",
  63524=>"00000000",
  63525=>"00000000",
  63526=>"00000000",
  63527=>"00000000",
  63528=>"00000000",
  63529=>"00000000",
  63530=>"00000000",
  63531=>"00000000",
  63532=>"00000000",
  63533=>"00000000",
  63534=>"00000000",
  63535=>"00000000",
  63536=>"00000000",
  63537=>"00000000",
  63538=>"00000000",
  63539=>"00000000",
  63540=>"00000000",
  63541=>"00000000",
  63542=>"00000000",
  63543=>"00000000",
  63544=>"00000000",
  63545=>"00000000",
  63546=>"00000000",
  63547=>"00000000",
  63548=>"00000000",
  63549=>"00000000",
  63550=>"00000000",
  63551=>"00000000",
  63552=>"00000000",
  63553=>"00000000",
  63554=>"00000000",
  63555=>"00000000",
  63556=>"00000000",
  63557=>"00000000",
  63558=>"00000000",
  63559=>"00000000",
  63560=>"00000000",
  63561=>"00000000",
  63562=>"00000000",
  63563=>"00000000",
  63564=>"00000000",
  63565=>"00000000",
  63566=>"00000000",
  63567=>"00000000",
  63568=>"00000000",
  63569=>"00000000",
  63570=>"00000000",
  63571=>"00000000",
  63572=>"00000000",
  63573=>"00000000",
  63574=>"00000000",
  63575=>"00000000",
  63576=>"00000000",
  63577=>"00000000",
  63578=>"00000000",
  63579=>"00000000",
  63580=>"00000000",
  63581=>"00000000",
  63582=>"00000000",
  63583=>"00000000",
  63584=>"00000000",
  63585=>"00000000",
  63586=>"00000000",
  63587=>"00000000",
  63588=>"00000000",
  63589=>"00000000",
  63590=>"00000000",
  63591=>"00000000",
  63592=>"00000000",
  63593=>"00000000",
  63594=>"00000000",
  63595=>"00000000",
  63596=>"00000000",
  63597=>"00000000",
  63598=>"00000000",
  63599=>"00000000",
  63600=>"00000000",
  63601=>"00000000",
  63602=>"00000000",
  63603=>"00000000",
  63604=>"00000000",
  63605=>"00000000",
  63606=>"00000000",
  63607=>"00000000",
  63608=>"00000000",
  63609=>"00000000",
  63610=>"00000000",
  63611=>"00000000",
  63612=>"00000000",
  63613=>"00000000",
  63614=>"00000000",
  63615=>"00000000",
  63616=>"00000000",
  63617=>"00000000",
  63618=>"00000000",
  63619=>"00000000",
  63620=>"00000000",
  63621=>"00000000",
  63622=>"00000000",
  63623=>"00000000",
  63624=>"00000000",
  63625=>"00000000",
  63626=>"00000000",
  63627=>"00000000",
  63628=>"00000000",
  63629=>"00000000",
  63630=>"00000000",
  63631=>"00000000",
  63632=>"00000000",
  63633=>"00000000",
  63634=>"00000000",
  63635=>"00000000",
  63636=>"00000000",
  63637=>"00000000",
  63638=>"00000000",
  63639=>"00000000",
  63640=>"00000000",
  63641=>"00000000",
  63642=>"00000000",
  63643=>"00000000",
  63644=>"00000000",
  63645=>"00000000",
  63646=>"00000000",
  63647=>"00000000",
  63648=>"00000000",
  63649=>"00000000",
  63650=>"00000000",
  63651=>"00000000",
  63652=>"00000000",
  63653=>"00000000",
  63654=>"00000000",
  63655=>"00000000",
  63656=>"00000000",
  63657=>"00000000",
  63658=>"00000000",
  63659=>"00000000",
  63660=>"00000000",
  63661=>"00000000",
  63662=>"00000000",
  63663=>"00000000",
  63664=>"00000000",
  63665=>"00000000",
  63666=>"00000000",
  63667=>"00000000",
  63668=>"00000000",
  63669=>"00000000",
  63670=>"00000000",
  63671=>"00000000",
  63672=>"00000000",
  63673=>"00000000",
  63674=>"00000000",
  63675=>"00000000",
  63676=>"00000000",
  63677=>"00000000",
  63678=>"00000000",
  63679=>"00000000",
  63680=>"00000000",
  63681=>"00000000",
  63682=>"00000000",
  63683=>"00000000",
  63684=>"00000000",
  63685=>"00000000",
  63686=>"00000000",
  63687=>"00000000",
  63688=>"00000000",
  63689=>"00000000",
  63690=>"00000000",
  63691=>"00000000",
  63692=>"00000000",
  63693=>"00000000",
  63694=>"00000000",
  63695=>"00000000",
  63696=>"00000000",
  63697=>"00000000",
  63698=>"00000000",
  63699=>"00000000",
  63700=>"00000000",
  63701=>"00000000",
  63702=>"00000000",
  63703=>"00000000",
  63704=>"00000000",
  63705=>"00000000",
  63706=>"00000000",
  63707=>"00000000",
  63708=>"00000000",
  63709=>"00000000",
  63710=>"00000000",
  63711=>"00000000",
  63712=>"00000000",
  63713=>"00000000",
  63714=>"00000000",
  63715=>"00000000",
  63716=>"00000000",
  63717=>"00000000",
  63718=>"00000000",
  63719=>"00000000",
  63720=>"00000000",
  63721=>"00000000",
  63722=>"00000000",
  63723=>"00000000",
  63724=>"00000000",
  63725=>"00000000",
  63726=>"00000000",
  63727=>"00000000",
  63728=>"00000000",
  63729=>"00000000",
  63730=>"00000000",
  63731=>"00000000",
  63732=>"00000000",
  63733=>"00000000",
  63734=>"00000000",
  63735=>"00000000",
  63736=>"00000000",
  63737=>"00000000",
  63738=>"00000000",
  63739=>"00000000",
  63740=>"00000000",
  63741=>"00000000",
  63742=>"00000000",
  63743=>"00000000",
  63744=>"00000000",
  63745=>"00000000",
  63746=>"00000000",
  63747=>"00000000",
  63748=>"00000000",
  63749=>"00000000",
  63750=>"00000000",
  63751=>"00000000",
  63752=>"00000000",
  63753=>"00000000",
  63754=>"00000000",
  63755=>"00000000",
  63756=>"00000000",
  63757=>"00000000",
  63758=>"00000000",
  63759=>"00000000",
  63760=>"00000000",
  63761=>"00000000",
  63762=>"00000000",
  63763=>"00000000",
  63764=>"00000000",
  63765=>"00000000",
  63766=>"00000000",
  63767=>"00000000",
  63768=>"00000000",
  63769=>"00000000",
  63770=>"00000000",
  63771=>"00000000",
  63772=>"00000000",
  63773=>"00000000",
  63774=>"00000000",
  63775=>"00000000",
  63776=>"00000000",
  63777=>"00000000",
  63778=>"00000000",
  63779=>"00000000",
  63780=>"00000000",
  63781=>"00000000",
  63782=>"00000000",
  63783=>"00000000",
  63784=>"00000000",
  63785=>"00000000",
  63786=>"00000000",
  63787=>"00000000",
  63788=>"00000000",
  63789=>"00000000",
  63790=>"00000000",
  63791=>"00000000",
  63792=>"00000000",
  63793=>"00000000",
  63794=>"00000000",
  63795=>"00000000",
  63796=>"00000000",
  63797=>"00000000",
  63798=>"00000000",
  63799=>"00000000",
  63800=>"00000000",
  63801=>"00000000",
  63802=>"00000000",
  63803=>"00000000",
  63804=>"00000000",
  63805=>"00000000",
  63806=>"00000000",
  63807=>"00000000",
  63808=>"00000000",
  63809=>"00000000",
  63810=>"00000000",
  63811=>"00000000",
  63812=>"00000000",
  63813=>"00000000",
  63814=>"00000000",
  63815=>"00000000",
  63816=>"00000000",
  63817=>"00000000",
  63818=>"00000000",
  63819=>"00000000",
  63820=>"00000000",
  63821=>"00000000",
  63822=>"00000000",
  63823=>"00000000",
  63824=>"00000000",
  63825=>"00000000",
  63826=>"00000000",
  63827=>"00000000",
  63828=>"00000000",
  63829=>"00000000",
  63830=>"00000000",
  63831=>"00000000",
  63832=>"00000000",
  63833=>"00000000",
  63834=>"00000000",
  63835=>"00000000",
  63836=>"00000000",
  63837=>"00000000",
  63838=>"00000000",
  63839=>"00000000",
  63840=>"00000000",
  63841=>"00000000",
  63842=>"00000000",
  63843=>"00000000",
  63844=>"00000000",
  63845=>"00000000",
  63846=>"00000000",
  63847=>"00000000",
  63848=>"00000000",
  63849=>"00000000",
  63850=>"00000000",
  63851=>"00000000",
  63852=>"00000000",
  63853=>"00000000",
  63854=>"00000000",
  63855=>"00000000",
  63856=>"00000000",
  63857=>"00000000",
  63858=>"00000000",
  63859=>"00000000",
  63860=>"00000000",
  63861=>"00000000",
  63862=>"00000000",
  63863=>"00000000",
  63864=>"00000000",
  63865=>"00000000",
  63866=>"00000000",
  63867=>"00000000",
  63868=>"00000000",
  63869=>"00000000",
  63870=>"00000000",
  63871=>"00000000",
  63872=>"00000000",
  63873=>"00000000",
  63874=>"00000000",
  63875=>"00000000",
  63876=>"00000000",
  63877=>"00000000",
  63878=>"00000000",
  63879=>"00000000",
  63880=>"00000000",
  63881=>"00000000",
  63882=>"00000000",
  63883=>"00000000",
  63884=>"00000000",
  63885=>"00000000",
  63886=>"00000000",
  63887=>"00000000",
  63888=>"00000000",
  63889=>"00000000",
  63890=>"00000000",
  63891=>"00000000",
  63892=>"00000000",
  63893=>"00000000",
  63894=>"00000000",
  63895=>"00000000",
  63896=>"00000000",
  63897=>"00000000",
  63898=>"00000000",
  63899=>"00000000",
  63900=>"00000000",
  63901=>"00000000",
  63902=>"00000000",
  63903=>"00000000",
  63904=>"00000000",
  63905=>"00000000",
  63906=>"00000000",
  63907=>"00000000",
  63908=>"00000000",
  63909=>"00000000",
  63910=>"00000000",
  63911=>"00000000",
  63912=>"00000000",
  63913=>"00000000",
  63914=>"00000000",
  63915=>"00000000",
  63916=>"00000000",
  63917=>"00000000",
  63918=>"00000000",
  63919=>"00000000",
  63920=>"00000000",
  63921=>"00000000",
  63922=>"00000000",
  63923=>"00000000",
  63924=>"00000000",
  63925=>"00000000",
  63926=>"00000000",
  63927=>"00000000",
  63928=>"00000000",
  63929=>"00000000",
  63930=>"00000000",
  63931=>"00000000",
  63932=>"00000000",
  63933=>"00000000",
  63934=>"00000000",
  63935=>"00000000",
  63936=>"00000000",
  63937=>"00000000",
  63938=>"00000000",
  63939=>"00000000",
  63940=>"00000000",
  63941=>"00000000",
  63942=>"00000000",
  63943=>"00000000",
  63944=>"00000000",
  63945=>"00000000",
  63946=>"00000000",
  63947=>"00000000",
  63948=>"00000000",
  63949=>"00000000",
  63950=>"00000000",
  63951=>"00000000",
  63952=>"00000000",
  63953=>"00000000",
  63954=>"00000000",
  63955=>"00000000",
  63956=>"00000000",
  63957=>"00000000",
  63958=>"00000000",
  63959=>"00000000",
  63960=>"00000000",
  63961=>"00000000",
  63962=>"00000000",
  63963=>"00000000",
  63964=>"00000000",
  63965=>"00000000",
  63966=>"00000000",
  63967=>"00000000",
  63968=>"00000000",
  63969=>"00000000",
  63970=>"00000000",
  63971=>"00000000",
  63972=>"00000000",
  63973=>"00000000",
  63974=>"00000000",
  63975=>"00000000",
  63976=>"00000000",
  63977=>"00000000",
  63978=>"00000000",
  63979=>"00000000",
  63980=>"00000000",
  63981=>"00000000",
  63982=>"00000000",
  63983=>"00000000",
  63984=>"00000000",
  63985=>"00000000",
  63986=>"00000000",
  63987=>"00000000",
  63988=>"00000000",
  63989=>"00000000",
  63990=>"00000000",
  63991=>"00000000",
  63992=>"00000000",
  63993=>"00000000",
  63994=>"00000000",
  63995=>"00000000",
  63996=>"00000000",
  63997=>"00000000",
  63998=>"00000000",
  63999=>"00000000",
  64000=>"00000000",
  64001=>"00000000",
  64002=>"00000000",
  64003=>"00000000",
  64004=>"00000000",
  64005=>"00000000",
  64006=>"00000000",
  64007=>"00000000",
  64008=>"00000000",
  64009=>"00000000",
  64010=>"00000000",
  64011=>"00000000",
  64012=>"00000000",
  64013=>"00000000",
  64014=>"00000000",
  64015=>"00000000",
  64016=>"00000000",
  64017=>"00000000",
  64018=>"00000000",
  64019=>"00000000",
  64020=>"00000000",
  64021=>"00000000",
  64022=>"00000000",
  64023=>"00000000",
  64024=>"00000000",
  64025=>"00000000",
  64026=>"00000000",
  64027=>"00000000",
  64028=>"00000000",
  64029=>"00000000",
  64030=>"00000000",
  64031=>"00000000",
  64032=>"00000000",
  64033=>"00000000",
  64034=>"00000000",
  64035=>"00000000",
  64036=>"00000000",
  64037=>"00000000",
  64038=>"00000000",
  64039=>"00000000",
  64040=>"00000000",
  64041=>"00000000",
  64042=>"00000000",
  64043=>"00000000",
  64044=>"00000000",
  64045=>"00000000",
  64046=>"00000000",
  64047=>"00000000",
  64048=>"00000000",
  64049=>"00000000",
  64050=>"00000000",
  64051=>"00000000",
  64052=>"00000000",
  64053=>"00000000",
  64054=>"00000000",
  64055=>"00000000",
  64056=>"00000000",
  64057=>"00000000",
  64058=>"00000000",
  64059=>"00000000",
  64060=>"00000000",
  64061=>"00000000",
  64062=>"00000000",
  64063=>"00000000",
  64064=>"00000000",
  64065=>"00000000",
  64066=>"00000000",
  64067=>"00000000",
  64068=>"00000000",
  64069=>"00000000",
  64070=>"00000000",
  64071=>"00000000",
  64072=>"00000000",
  64073=>"00000000",
  64074=>"00000000",
  64075=>"00000000",
  64076=>"00000000",
  64077=>"00000000",
  64078=>"00000000",
  64079=>"00000000",
  64080=>"00000000",
  64081=>"00000000",
  64082=>"00000000",
  64083=>"00000000",
  64084=>"00000000",
  64085=>"00000000",
  64086=>"00000000",
  64087=>"00000000",
  64088=>"00000000",
  64089=>"00000000",
  64090=>"00000000",
  64091=>"00000000",
  64092=>"00000000",
  64093=>"00000000",
  64094=>"00000000",
  64095=>"00000000",
  64096=>"00000000",
  64097=>"00000000",
  64098=>"00000000",
  64099=>"00000000",
  64100=>"00000000",
  64101=>"00000000",
  64102=>"00000000",
  64103=>"00000000",
  64104=>"00000000",
  64105=>"00000000",
  64106=>"00000000",
  64107=>"00000000",
  64108=>"00000000",
  64109=>"00000000",
  64110=>"00000000",
  64111=>"00000000",
  64112=>"00000000",
  64113=>"00000000",
  64114=>"00000000",
  64115=>"00000000",
  64116=>"00000000",
  64117=>"00000000",
  64118=>"00000000",
  64119=>"00000000",
  64120=>"00000000",
  64121=>"00000000",
  64122=>"00000000",
  64123=>"00000000",
  64124=>"00000000",
  64125=>"00000000",
  64126=>"00000000",
  64127=>"00000000",
  64128=>"00000000",
  64129=>"00000000",
  64130=>"00000000",
  64131=>"00000000",
  64132=>"00000000",
  64133=>"00000000",
  64134=>"00000000",
  64135=>"00000000",
  64136=>"00000000",
  64137=>"00000000",
  64138=>"00000000",
  64139=>"00000000",
  64140=>"00000000",
  64141=>"00000000",
  64142=>"00000000",
  64143=>"00000000",
  64144=>"00000000",
  64145=>"00000000",
  64146=>"00000000",
  64147=>"00000000",
  64148=>"00000000",
  64149=>"00000000",
  64150=>"00000000",
  64151=>"00000000",
  64152=>"00000000",
  64153=>"00000000",
  64154=>"00000000",
  64155=>"00000000",
  64156=>"00000000",
  64157=>"00000000",
  64158=>"00000000",
  64159=>"00000000",
  64160=>"00000000",
  64161=>"00000000",
  64162=>"00000000",
  64163=>"00000000",
  64164=>"00000000",
  64165=>"00000000",
  64166=>"00000000",
  64167=>"00000000",
  64168=>"00000000",
  64169=>"00000000",
  64170=>"00000000",
  64171=>"00000000",
  64172=>"00000000",
  64173=>"00000000",
  64174=>"00000000",
  64175=>"00000000",
  64176=>"00000000",
  64177=>"00000000",
  64178=>"00000000",
  64179=>"00000000",
  64180=>"00000000",
  64181=>"00000000",
  64182=>"00000000",
  64183=>"00000000",
  64184=>"00000000",
  64185=>"00000000",
  64186=>"00000000",
  64187=>"00000000",
  64188=>"00000000",
  64189=>"00000000",
  64190=>"00000000",
  64191=>"00000000",
  64192=>"00000000",
  64193=>"00000000",
  64194=>"00000000",
  64195=>"00000000",
  64196=>"00000000",
  64197=>"00000000",
  64198=>"00000000",
  64199=>"00000000",
  64200=>"00000000",
  64201=>"00000000",
  64202=>"00000000",
  64203=>"00000000",
  64204=>"00000000",
  64205=>"00000000",
  64206=>"00000000",
  64207=>"00000000",
  64208=>"00000000",
  64209=>"00000000",
  64210=>"00000000",
  64211=>"00000000",
  64212=>"00000000",
  64213=>"00000000",
  64214=>"00000000",
  64215=>"00000000",
  64216=>"00000000",
  64217=>"00000000",
  64218=>"00000000",
  64219=>"00000000",
  64220=>"00000000",
  64221=>"00000000",
  64222=>"00000000",
  64223=>"00000000",
  64224=>"00000000",
  64225=>"00000000",
  64226=>"00000000",
  64227=>"00000000",
  64228=>"00000000",
  64229=>"00000000",
  64230=>"00000000",
  64231=>"00000000",
  64232=>"00000000",
  64233=>"00000000",
  64234=>"00000000",
  64235=>"00000000",
  64236=>"00000000",
  64237=>"00000000",
  64238=>"00000000",
  64239=>"00000000",
  64240=>"00000000",
  64241=>"00000000",
  64242=>"00000000",
  64243=>"00000000",
  64244=>"00000000",
  64245=>"00000000",
  64246=>"00000000",
  64247=>"00000000",
  64248=>"00000000",
  64249=>"00000000",
  64250=>"00000000",
  64251=>"00000000",
  64252=>"00000000",
  64253=>"00000000",
  64254=>"00000000",
  64255=>"00000000",
  64256=>"00000000",
  64257=>"00000000",
  64258=>"00000000",
  64259=>"00000000",
  64260=>"00000000",
  64261=>"00000000",
  64262=>"00000000",
  64263=>"00000000",
  64264=>"00000000",
  64265=>"00000000",
  64266=>"00000000",
  64267=>"00000000",
  64268=>"00000000",
  64269=>"00000000",
  64270=>"00000000",
  64271=>"00000000",
  64272=>"00000000",
  64273=>"00000000",
  64274=>"00000000",
  64275=>"00000000",
  64276=>"00000000",
  64277=>"00000000",
  64278=>"00000000",
  64279=>"00000000",
  64280=>"00000000",
  64281=>"00000000",
  64282=>"00000000",
  64283=>"00000000",
  64284=>"00000000",
  64285=>"00000000",
  64286=>"00000000",
  64287=>"00000000",
  64288=>"00000000",
  64289=>"00000000",
  64290=>"00000000",
  64291=>"00000000",
  64292=>"00000000",
  64293=>"00000000",
  64294=>"00000000",
  64295=>"00000000",
  64296=>"00000000",
  64297=>"00000000",
  64298=>"00000000",
  64299=>"00000000",
  64300=>"00000000",
  64301=>"00000000",
  64302=>"00000000",
  64303=>"00000000",
  64304=>"00000000",
  64305=>"00000000",
  64306=>"00000000",
  64307=>"00000000",
  64308=>"00000000",
  64309=>"00000000",
  64310=>"00000000",
  64311=>"00000000",
  64312=>"00000000",
  64313=>"00000000",
  64314=>"00000000",
  64315=>"00000000",
  64316=>"00000000",
  64317=>"00000000",
  64318=>"00000000",
  64319=>"00000000",
  64320=>"00000000",
  64321=>"00000000",
  64322=>"00000000",
  64323=>"00000000",
  64324=>"00000000",
  64325=>"00000000",
  64326=>"00000000",
  64327=>"00000000",
  64328=>"00000000",
  64329=>"00000000",
  64330=>"00000000",
  64331=>"00000000",
  64332=>"00000000",
  64333=>"00000000",
  64334=>"00000000",
  64335=>"00000000",
  64336=>"00000000",
  64337=>"00000000",
  64338=>"00000000",
  64339=>"00000000",
  64340=>"00000000",
  64341=>"00000000",
  64342=>"00000000",
  64343=>"00000000",
  64344=>"00000000",
  64345=>"00000000",
  64346=>"00000000",
  64347=>"00000000",
  64348=>"00000000",
  64349=>"00000000",
  64350=>"00000000",
  64351=>"00000000",
  64352=>"00000000",
  64353=>"00000000",
  64354=>"00000000",
  64355=>"00000000",
  64356=>"00000000",
  64357=>"00000000",
  64358=>"00000000",
  64359=>"00000000",
  64360=>"00000000",
  64361=>"00000000",
  64362=>"00000000",
  64363=>"00000000",
  64364=>"00000000",
  64365=>"00000000",
  64366=>"00000000",
  64367=>"00000000",
  64368=>"00000000",
  64369=>"00000000",
  64370=>"00000000",
  64371=>"00000000",
  64372=>"00000000",
  64373=>"00000000",
  64374=>"00000000",
  64375=>"00000000",
  64376=>"00000000",
  64377=>"00000000",
  64378=>"00000000",
  64379=>"00000000",
  64380=>"00000000",
  64381=>"00000000",
  64382=>"00000000",
  64383=>"00000000",
  64384=>"00000000",
  64385=>"00000000",
  64386=>"00000000",
  64387=>"00000000",
  64388=>"00000000",
  64389=>"00000000",
  64390=>"00000000",
  64391=>"00000000",
  64392=>"00000000",
  64393=>"00000000",
  64394=>"00000000",
  64395=>"00000000",
  64396=>"00000000",
  64397=>"00000000",
  64398=>"00000000",
  64399=>"00000000",
  64400=>"00000000",
  64401=>"00000000",
  64402=>"00000000",
  64403=>"00000000",
  64404=>"00000000",
  64405=>"00000000",
  64406=>"00000000",
  64407=>"00000000",
  64408=>"00000000",
  64409=>"00000000",
  64410=>"00000000",
  64411=>"00000000",
  64412=>"00000000",
  64413=>"00000000",
  64414=>"00000000",
  64415=>"00000000",
  64416=>"00000000",
  64417=>"00000000",
  64418=>"00000000",
  64419=>"00000000",
  64420=>"00000000",
  64421=>"00000000",
  64422=>"00000000",
  64423=>"00000000",
  64424=>"00000000",
  64425=>"00000000",
  64426=>"00000000",
  64427=>"00000000",
  64428=>"00000000",
  64429=>"00000000",
  64430=>"00000000",
  64431=>"00000000",
  64432=>"00000000",
  64433=>"00000000",
  64434=>"00000000",
  64435=>"00000000",
  64436=>"00000000",
  64437=>"00000000",
  64438=>"00000000",
  64439=>"00000000",
  64440=>"00000000",
  64441=>"00000000",
  64442=>"00000000",
  64443=>"00000000",
  64444=>"00000000",
  64445=>"00000000",
  64446=>"00000000",
  64447=>"00000000",
  64448=>"00000000",
  64449=>"00000000",
  64450=>"00000000",
  64451=>"00000000",
  64452=>"00000000",
  64453=>"00000000",
  64454=>"00000000",
  64455=>"00000000",
  64456=>"00000000",
  64457=>"00000000",
  64458=>"00000000",
  64459=>"00000000",
  64460=>"00000000",
  64461=>"00000000",
  64462=>"00000000",
  64463=>"00000000",
  64464=>"00000000",
  64465=>"00000000",
  64466=>"00000000",
  64467=>"00000000",
  64468=>"00000000",
  64469=>"00000000",
  64470=>"00000000",
  64471=>"00000000",
  64472=>"00000000",
  64473=>"00000000",
  64474=>"00000000",
  64475=>"00000000",
  64476=>"00000000",
  64477=>"00000000",
  64478=>"00000000",
  64479=>"00000000",
  64480=>"00000000",
  64481=>"00000000",
  64482=>"00000000",
  64483=>"00000000",
  64484=>"00000000",
  64485=>"00000000",
  64486=>"00000000",
  64487=>"00000000",
  64488=>"00000000",
  64489=>"00000000",
  64490=>"00000000",
  64491=>"00000000",
  64492=>"00000000",
  64493=>"00000000",
  64494=>"00000000",
  64495=>"00000000",
  64496=>"00000000",
  64497=>"00000000",
  64498=>"00000000",
  64499=>"00000000",
  64500=>"00000000",
  64501=>"00000000",
  64502=>"00000000",
  64503=>"00000000",
  64504=>"00000000",
  64505=>"00000000",
  64506=>"00000000",
  64507=>"00000000",
  64508=>"00000000",
  64509=>"00000000",
  64510=>"00000000",
  64511=>"00000000");

  BEGIN
  weight <= ROM_content(to_integer(address));
END RTL;